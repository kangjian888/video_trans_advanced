

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CvmaYyJzAT4gGJRlCkE1yXt5Lv9gJbr2gC0wBzixkhI3TupXRLTg9s4Z9WVWp43QDkUuM3VRZjAj
RVnqESt3JA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hHyS2uxRkJ6sHR79RwG8dxYfMwySDoNzo0ZpVSoiAp/93R212I5J1LxM+7EujDw/cO/x9djlyxbz
erzC6/tIqQ2nS2hUZANmmER9YkiA1RlXlIqDOWo8pOFHNj1c4jf7Zdq7OJMDPvKF+fLgmk5Lu9Y0
15oIyfQw7L+gXpW1qEU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Cfhh7YIOGyVJiZpd5j8xa2ugbHZdDDpkNcw6vvVCCgnGCfzlen3wlGk0omzzJqyVapnfg0aPFCVf
eH/noQVGu1bQkowx0JKcNE5x1v5DKH//UNI+lq09SNF0WKlMcTAGlNSUzO8kgVv9uNbKUHDXodcD
5iGh6bHMhVPSu1QKpTfJlIMd2CMz0JfDQiVbfTaAGKvrQhaqVte7pYpnqiXM7povPwt/ntWHBH4s
XSF4J4eDVLMuQmQNy3vrqFdEUqmQFtLWgNRpG2fwo19Y2lRzT3ux5SiA0Iv55uR6x7AG21x8BZlD
JC102ufirdrREfWUzlClY8zmr+TUHpTF/SgPMw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UWceDgHVHZAg17Yudaw03bncVn75AJ6y0RYlYeqdZU3kMG9E1W6q5REaQAI7sMZSrC2g0zavsx4w
utskoq80P2avoebtdvBfjr/nBCQqUN3AvM3GSk85froboZgk4fCQ8UtEj2Qk7ob+ox/md7d9P9dw
2YULi+eG04dUc1g45wwF0ZoZdARk7Ml+fXMnm7zxmvqVieAEsVq6ETZN/P0pwvIpAakLTayKriGC
qcrb1S28bOuV+Na/FX9rxN6hM5aK7vSdFqja5GGs32r9UVRIkX6i7uqS9pWQDR0Qa31W3z6wrRrT
+2wzEwNMDKYuWVIM1FQo/Tp0NKa1Y+kyjahSGA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tLsJPLnIUk5FSxPTGLkNhAFldHrP7oFH8h39nfqyEmnC/AmGzR3fePfCEcee3I4TYySABpWhyXIf
m1jGiCuHfIpFkF2EJqjWmBev0bD33cbw1av2xtJRFa5gaQjxChO9URfjedFvCQWWwjlxejc9nD0N
O0V2XUDQxd573YmSBuByzshlxt3bujEd6Xeeb8N8NI8c2ZsfY4693LGdb3k6gtY9ZEoo4XuYVt6n
S2tNFVJTfQjyBEXbuCPqpwGf6bPdy2SKvTE/s4rSIVTO08J6bXDaEOBUGg13XVoJJqrayiJRVuQL
LhoiPzgOqS6ude1uUaMHE/SN9X/vt/6uOsOl2w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jgk19ieS+ZYiySHKvgAHMus0OAx0HPJ59p64LMaYK8CyW0wSM8LIn++sFz9tsOBdLj2gb8IKpSVr
SOX9XXXM2pQFSME7x8q0m+EPg9m1+ghIpW4bU/w4zVq4NBjYydZCI0Hpy+X3op0a3+eENVEw5SoK
4R/zOL7aV/2nZ//wkaw=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
L/BPRr/PHH5da1O06dKRr5ST8eskM6lzR1UPuTvZQ6RCsFEjTD1HgyqjW7/ypnIq7V5TYDC553+Y
rJnEENzDc6RSpzenrYxw7NrURpUedIWlCc/PEf5Zq9gu1ESkpND7t98rc+uiAz7zsn/pHD/K50NR
q9l/gcWkOCgArmADo1Lw9usrfZ8ECIPKY2kLxeTYbh4fsrCpPQsQUk4NxX3N1Q0h3RRUCdHSFc0O
lvGip/vd24OK8zXDMaQv4fPmgToFQMUvLrJXErEUeRlkpxkcX6g6Zu4RMWwwmkNIfZHpc5K8Q3RL
MMc5rARUSXbNbpf28H3iyAMZ0y+EgI0CrKwooA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967856)
`protect data_block
QCm4HuQKiYy3DVHsH65D6Aj9OL3RtWCCXGwahQ37x8ObWwLS5rgEIP+a8OTS0lZU+UJWkzITZQfF
WIUzBu096DKRrTIiKaceWHrTRneNTzXfw5TZPQQguRfJIVTocvUXcaAGiyS/K6F48tezM5qi2JLl
CS6awmxqjObHRrONz+OkLBhxLXLi0K8/LY/H1mCYPXt/fzMxwk8p+dlp767kXFiq9yeXh2y4MTPw
P1bhg+JjRsGmdpVcetIoTEVANIjExCPoNV2f7ZstvPFT8HK80wG9kTNocsrhN1gsXbN3btGH7I3o
iYxcgJ8GvohWXsEfm4N4TVvc7S+xpUjHfZ7v/7mwwoOMR+pWTNn3SXuJFs4W4WW1iNGmedoaL5PU
79Xqbfpbi72A0rZ1/36Z07fS/VqnzWb7oUnk825oGxyC5trHrTgdoM7yqu8xJz8fx20gDfJ1gjFC
Odk9eylzFp0OZnYtzKvUw9NnvUfcLKuGpOksdZJ8w36n3sWwIZdtSht7kCPhxEcicDZ9M8ivRnEh
F+yX5kLHjuOdJv93SbqnGUXHurnl2t2IB/h/ukVIizxwR6AyYF05X+gz7FoXwPGnoaSkfbvypCoN
4XiObqUYyt7/1cMF9VD+diTFBXjFrSPRySBZppW9/hSGJeefUFGXSvfCtInoKFVG2LdeOUCdLRzV
zUtaw7VhFDYruj4CLKkR0MJCkG7sQDna+5oSTYfzz3ujC9bsbYsuxziXWeUOZtooG29F7X8czKK2
72D+F0ZavFnIrNLLquIdrK601My8hPAe3ho/4ZoOovB9YFfBBdwYD1Qx1YUzuGxMHBzyNno/h8Wk
79zG1uV6wikxfVb6J+gMJi+CDHjtbJlXSszzN6QAKS28z+bltZvYLbf6C3lRKQ/cXoMZ5BLEnmF4
5iGo6SUPg+w6ohOudjHofPLKrrBErz1DazqyuuxVziqQZ1GMEbzD9H7Hzy90RY+I/adLqjTgsuho
eF2FoO2KVJSGiWMymkb82hBSrq30cyuz4z7or9pd7jgDp+bc+z8vICFvAYctYn0v1XJGrnWKHJv6
2gcCF6k7SRz7HTkuZyDuhPKg5lyRWr1SBdD8B9DKO0EzVeLEq643zrTWRkVwiGNlO8S6dRlSyM7C
jtiVKi2T/fsJEqmzyCi238tZfBmGNZ7BH8MKfrK8kdt1I2zV6r9P7vNcHFTs+W1SIgeblGsnwhF/
ILlBVms/G8DWDPw/gT0Cl8qFkCU0HERdY9v1iE/nvg9UkjIjCWx+L3A4ENKGSwos9mAPPTdAsj/t
0dMC0zG90eqFxYx9jGN4ohRhuj8BWCUXn45tViIaC0r4HFq/ZP1q88FcEsBlL0PB5maZlpmih5J3
efcAMYpfrfRkLBGvylxtgytKGRmSch6mupT3Jv6gegdkZBiloYm/bQUvWecMLDRB320IDVSKw1tu
79ucz0w4HabBaIP/aeIQNBAfF4b4nuV/dflSm/te6f8sF8yTxRBjie4cTKSRTrcEF3NGZZC4i3UQ
rCKIphMF6Rtp3R9ZF0JXYfcC4mhEoWxZz+9z2nsnlJfqJsw5w1fdr7NRyHzv04Nd6OqD+6GLDbt5
lX+9jYf0D2/SW6mOkFoofm/A5qzm87WJeIN4jI9lABFOaXObZpfr7tbUbjQo2gUOtmcDuudxepTe
QHOfYbPQ49Ny+uBro4xPOoLlgePgwkZGIP1w3sI3GE/k36boEDZIpvLHr//064MjN3mFMjzbfXpW
pvqSz7dEt0mGDT4Qu1hysNFR6bkN+oW/fjlYuvrXaX5rIF0JZ7g1ReToEjisPRH2JmIZG6hHwsK5
A6sdpsazED2BjQd/sh9FN1mH5erjVn5liBzCX9BeO9tj3mAVVZvap5rEKOkIGpFQ3ertLk43e5i9
WwCsuCrtLgrynYREOZRvGXQQVCTTtNDHlqFebW9QN/zfBnFO6SR+xQulQQWrJDcQFZtndY1jnwOo
0smoi07GZpy2tJ1nR/twrtUa42TkLW5E+eMVj8ySxNEUx/N8lju/C+NtdrCDhR7CIL4TX/1qxaoa
/rz/6/OxM8lAqhnigMFvOSPopU1MKJ20qz7deMqP36vNwS7OqMFy3Cdp7d35hNJjH3QTOuK+TrUu
lr9at7W+DYucx7TQA+Wlh3REaoBxeV4KboeRs4msmLsq1M169QfdQ1/G+ieWv7F6/Fm/ZRay93Bf
FPqCNbXv+GT2aZ7s8p1SM5N78itspAAUf2OaPLEzuYmu+q8dBKfYv5lFsmd5qfZLM4CzWrwnC22Z
cWK2V//27dc3qOsSKJaSvLkciqoEsH/dog02iEHs9UHoxPTMO/gxUs1g0Bd0Tpo3TqnUpr7tUFht
scO2vLpZWTgkF4IEfGnpNdA8c4SI3mmaVdsMhIqxqmWEeSqikos2SP/huRZzKwiMyyvdD4adxCgh
lO9ynaH0p8OvGUk8cIWvhxjt3teV1SrUqcAeA4A+LNyh9/336vUj4S2OcncUYxh13fTatswKuuiO
KmjpxdfMYkoE0GPtXiOaA7484LhB2GEyIxDf2/Sevxl7PjHQYp7ROnaZjbENCkczlQgvSrJyEBGJ
OebmsA9AUETl6QnsNmb6MvTnezZNLJ1niSMXB4Ux0utBW5/82fsU7PmoqNp1Io8mEy95FfFlVzFA
ND1MWK44st8UZNA/n1ZJXkgD/1OMX+nyfsGCZTKUOVIiKndpuSxJRGAtL6IPEtH7dv4Thd+UlpBK
EHbOwojfW+igXitsc9NnUGAyhSRHVGFJg7r+u9Ngjp4SlZBkxa7tWjPEUdqDOLHXoMqSvAKFIJU2
/cGmR5NgNN/RUrrAqJwe3joOKpxTMZgqXO254HDsUIHzgRbHU2ppFY6G6Yn5XM8PGbL+Y2+Mo6RA
DtAXAkl9EiJr3jMROyrmSJGRhvz/rfj1R6RmZHBW6YAAGqT7Z0DP87HRF9+zRBnGon/hphXrBMa8
aY+iqZmqcqCMQWf6WPH0SRU0BHWhtNkvL7oblqrih8aKroXVh1Miv3hE76cxCzNmM64E0IzIsFtl
LxXQICyPWxv61KSA6qdtAeuL9vOzGdlj/NNwGUr3FqL8E5DJdzBRNYeWXbRB7he+fRVGklEgtkn9
wNdeg9VH7qB3g2/WSfGOWD1JTRMPYXhmqPvv9nt3y84MNyqNN0vhHbKTY+tZdYVy6fC3YQvBub1Z
uCUFAwoUc5vg+TIm9MVETeHc1nYCpmn2VjiaPtxCQHoKkvzEjTMRQGBLqtThFnpaduPLBftx7en5
zWIGAfplxFduyXTyQTh4TeCdQ1fksVtZ/QdSqwoExcev5VeUZLXo9KntNboGoBaUISy/khY6Roa7
T534K5v+j97iOLEflaFUXAKe4CKdJ4beqGfjOt0dG01fm1Zrw8B7o+oqSFlmxyT8IJgScfDTen9r
IQdEqiomvwTu9Xvn7zphQSiVrW8dwCJ7YxccWzBgMJ535ybAXdVOenMWqMl3mPIjvdzdEXeF+hmc
uRbfUXbbE2V/f4Q0L/OLHOnEkMYj3Zr7E0sPTT+Y6wBDdQChUZUuvH8O7f9OkuMC5bq0qKq0aRKj
a9/f+EtSfn9ddlgJCF4tFX9lVZInA4Q7byPUiyWkZfHJXqY0CXJTY+SmZCSi7xUgWLLlp+1DtT1a
MZYBMha6jjGWP7hZYUCGabTpFd8I5Nqtcq4I5BTUDuoIBsgWReNjglC7ZDNDzLfI2lIcTog2NqQA
uqqQZsXBY1Q2vagBMhMNoHbkZzU3EdAI/KjLoUG0xDvEnCARYD3I8xKRe8IJVIw+FLJ7JNW/WhHd
lwQkSE8Ut24jvtNK5+pjfO6v7g7bG62SAP2gdKV5tfXo5zacDa6pp1erOoZe53qrX00C9wEOE9Ax
5/Q/zvc4tfMwGYrF4PHT02aXmFCycx2Xg2ZQ9Jl5RVLnAq/UIOkeyEmzLPkFQ6dGI9oKChwy5RJw
mdVZSyWRZzbgR42+KtnODjFvk4J7YQmrz8L8RIvE8Wtv/0RYrzWtfj8dRCnWu4fxh83XBqtNx9n/
fhx++KIq+nu73KyQPODrYE6uGyj5VWv6nVVqP5p4E5P/jqwl8RdLYkhmJmgLGfBG+TlVpXNF5YYM
AXwPOp7Smk3Y0yhqK/ph5GLDf2xlAUqA1apLzkxswtLFdSKaZANJh7FmbmLhsoLlm3m4qnd0I3st
8TSP7lFRD9FGOI8ScDySSq5Q8IZQD7hcR5Ah2KeHuP2iHYrfxT6ZZDokQy/nDy1+0XGKYAIhtpfW
Z1kKiXu5Dl4tmjz8iKGxnJgOi5frmyrIF40r70NsZAX7OqSpkCVgxRQ1vwEo1kefVc9QbiLSzZDm
mUPCpqVsnZKRuSgJTHnmOpuNSGZzWlloYGSbA1yF8qjfB8MopiC12JIt6YZ0OSCYb/0dmivL7R23
hP0npWeB+ChbdZIcuDBagYTaC7gJdAPb5qBkpLKiZnBEDKTHrcklAoR/a65fSntOPSQr6auWmtG2
sXl0dkmUZLJr51t2gWKa7oKSz+e2ZMHFeBL46tys4QchxMqkynhUQPouX3en9mqpOgxm6xrKHrRH
p/cEByaeFUXrXxbQcUyWQDcQv+cqzPowkbZiLzrGZw6AGiX2rsWfZcM+pfjMjo/yu0hpzErvoYSK
i7W4Bq/nhKvFPVZgLX4ramwIXvvUDQ72IU5a4UauN0cYhVCYP8l1kWPFwnAOuqaajUWKpez9wDh9
HclgWNm/Wfe5UDC2F6aMBd82pSxy6aqtmbLqV/dWU2UICRppdi83PzCJwHmAqL/MNpUv+RfQz3Sp
RP/JuDG8ErBteTWFQWLHj5A5s7InAkoySXQ8BMuTa53TWFvt9XzDGsR//oc0NXxOaYRoG6WmwLtC
RYhYhIazES0vG3Ij4I3TeghbmOnmmj8RWYYts2vFvty55VH7STkdfJMciYLKGxmKAhB/Jo7QtCXa
2tzvshwA/wVAjtcoobh23bjdb+upMR0Y7NoB2RPhU4/zIo22KmlmSiGlXps151YO/UrUk0ZS4d7w
/5VHRAlii0c6lKNAk2LGenELhs5Qg/muxjEOvqWbB1PVgMyy4XXC//Gi9TnjNRw7QoBMtVbCh2l0
u2QWz38PzX8EPMUmfGoEXNU9bqtxx3KVsSw2MLIdqFdYY4GqyyJKS4nEdKMcLVy3dhFi8wrW8Tel
kwaYvT4oWt1zzuJRY1W4y8utfO4fhyJnTWx90NQRQ5p/Gfjdxv69SWWp+7d99E/s0hQFcS0iSbyJ
6WlZ3erEFJX8TfWdv5B75BfR/+HgigJBq17UiaW/dlCtNDXZmel2GOgziQbCsDVFN0/2+uc2o+ja
UmV4nzkU0JMGrqRzlqdWfp6uPtHEYh8/xHcMlskbXgokEZw4hXajqgeGHLdQrvYd+HD41xyz89LM
qIu9MHpRpyuxOH9IxTo5ECdmbBLmQKlUWG0XoZLucQq17MXDO2GffsC1kCgnqbwwWEITMjLABelP
irnM1See+HdVFVVZkUcvu2Bo86M+BtTFyFrFHw5GICh2N0d4g5ZwLGUzidxUD07yni8Y8CzmlNAT
5q6Dhrnso16ttbQa043U48O8RZuG5locrZQ4yNmjJkay/T3lV66wEa2YaGf/Y260T8vCV6JCqn7O
XfYKpTRW91jN0fBAd08lfyLzY+Ld/SHwl/0jFyVOhDrdbTGa2cYJFz8dOe020CQJhazI4/3U7P2b
RzdhNt1LgaOxB5EfcB70xDDlaDiXwWAbNWgDLUYI5GzyXzKlKHRHIclWYXfyHXrRGyW642K3HRuU
ikyHZYBTrTh6DLG/cYXyz4tPiwmsUrOOebOysn9ehgfbwyGpzuO8et06BAY7p0I7L7HjbW9EfP2W
5VBrCQGO/ZMWuOdD9Flwya0vU6krwMENGQcxTzChJxd/aD8hO1lzTn0cyqTNYXZP8UnT99JD38cx
+odm3GU1zynMG837Ezun6lemjchyDFGhEpRpQKIyyxhwLiotDOBYH73zrwZs0p0gOACdljyoHNuR
ZKRDx57P8lCYycXh6BmwDfV6cKKhpiqlba/DyaScnbyBve4NTTxW/Vq5yIH+ppLQISJ8tDQIa3IX
ouncsuKZppkRpT45ER1Z9Ec7SIteM2GVs2qTpwZ2SVb3l5rJ2IuPjaAi9A9T88vpToP737/O8aMu
97y1ZXYT3e4XeFcq1POSPAiSLNAPxUZBOYtUqHo/doQ0korXIXSi+pyOoWQkrCh2rkBjOjGiaudr
I9vXyfV5TCAfKPJ7d1J834f+yiqN1YdC/lu/Mnavyr9bErlounstdVRRxzlpnOOVLp51E6WbxZx+
LslIpDLv6QhuamgO/K19CiEbpkG+UkVu/tUWTJlTnW+KebGRT9GgGlnUbRFTm20FQjfeJRyDreZC
Zaelz5nldQQhAyY+KzEqxeEzEi6a13kEuIsUm/8+uAEGm1YB65jkvjwkpUvffKInCl2az90ZcxBs
+I4U9iILgcJCv3Zmd1ModEygK/Lb0lc6RBl2TauvqNjcdpJQjsgBkWMypXSYh94I/hKTMRJ6Wgpf
cOnbySaWEtnWqL+zjP2wS+ahn/YrGVjTEvAOh7jmpOzLTusjkNew5YjnhIdudC0n/11r/5VHXw59
EBqWafjq/M71QybV9naKolQ0STDaWIV9/54Y/nlnlmGy7FgC4iQeEZigruhkcTp6WOJFtNoVZD3E
sn7k0tedXTcGI+OqU9M5hFSVpypYxez77OhIlpc3Egw5pu3j14XSZem4kcEQv3f4FRlk+05UXEE9
cEsCp4+PXyhWZZ2tVHALoIsujXRx+cWlqpn1idH5UdJw5uECG7UoNGYytupiXvjbrcJHjk1goCd/
b7B4eLLs+WeacHxgFOK5yJQUFAduzh+UBUARQrc7MSu1CzzJtpyivMhBjKIj+oaM/KUcBazPE4uo
Rt5i7yCLRc+uWSegCjgK8eQIzzWaoIHg2+epEH8f03zfAJ7nIMsgcGzCUQuEyqDk4BJRHe9RSs8K
lkT8fqLy3Xc11dbqwkqaZnaudAY2PF0JNRAwzwkLCNK4WZAAqFTNopJ0ZxMn3M+9RP9l5NUw4saW
MckL5d5V1a4uNzN/wIiZHM97DQy15AA66gzP0YUZOdhkzkanvKIiY+zQ/EySZ8ZkuWl6KZmv6ClT
KULMOBIQtBP2kpuufRA8FnfLyc5Douif95KKCtrZ0Bhyeju+NK2WQIi32Ui9uQjlcQqsBakQeM+J
zj7zpsO0Bz+c9E2kljdc8jpaaKzHcBxGAt60Yh1XblN0MFIWDolfIyy9J/kBWUU9dAbnUhEcYUSw
5tWZLmaDWiQdr11DZl+v6F4zvRjx3XyLMVxiaOzLbCVxwo0TLUM0bnTjdt0D0bu0h2DA5ymdORBd
iiIElFZ1JPEpEcSB+GzTuGodd29rwSGvOR3RW8XeajsPFsKPYyjet3WJcGIsg0nF4vxpxZS8oqUM
+1JJhDcVR9HPSa7rBD19Cn5ke9ocMFeES8csn9UiZyUIQebmX7B3HtEXLWEwUcAx3YRgDneCfN0R
lfR+xGCLVewhVKSXTVquy4bXCMDr+PVyNjsgvxErm7IqupUPtUx5nWhK5XlsmoOjDdKg8eDp8ubk
hJK86trRFFndquDKOOFUvEOoxvZvsOxf4EJEElYEVh1NfWB8PtnJeI+ncvmbX5a8H02aQmYY4VT1
VagHrOFwiFrPBxALb/nEG9eacOaerLsYDAb7Z33Yhngzh1q3LL8rNLxBZ7e23fvTkrAlSfEezqWr
1U66Pn1gJ7zXs2SVC+SStmPlAgB3WqPvqYvTtARi418qJhg5H7d7eLNgwok+WorVT41dEUOH5Wb7
qiXB68td0bB0/TtmuPrlJhS9xs9aaSL/Vn6ocdB4grQ2R29dSlt49NqEROm/pSdFS4gQmDMOa5NA
cBh1pGf0+wh50VzW6Ur6aKj249tPfPU3GocoxSPbaqThBj+jh9BsZ+9buJo+j42CggJwXijH7vR8
jxvjDuH1crl8sMGQZ1zuJdE3lz+97zwVWpc3ACzYVJ7ZSksNB03rGCh56/Up/sioExz1dcTRH8Fd
y8JXYA8l9LlL/GBMt+6f9wt6TjcgjwgXTow5C+ldRrsZz2yeiRx6+lLTbKY47tu6M8f7Q99047dK
ewULGJT+OuygojIb7Prl9R1SFnpVUoCiE6plUK6bqVAO8oQy+ZHqZ7UZibBlCJ0kEiEpVLJ5S/ZJ
mMY0cOp91i/nb3k9JfdXpCAR67D8ZDbQtICo8ctojCniOkJlxlEXXKJjPCMRV6Kd9ar7c0W234yC
k5Co9CtkoFaDshQaGQcV5d1HloNTJGrQbCfUbP+DF58/Wi7qdbQE1vQiIDYuz+/5jefPN3a3wS/C
riS1MtdkW3HyBdG3wuZHa45IGM7O9sh1/cak+hYAaDqXoNp6wEGNuKzg+BckAhPkGsPkwR5rr021
dkW65Ofy0w3SxZgRPrPUQlHARZS5rpRmFVjd/VmsLpdfephsy+JRucS1cKz9p5yx0rbKIwyy0x6x
rnP/3HR9UXsIHb9LLMTMdZaBIwlW+IiHIGngwdPiE32vecotC3MtXrM7G8sdX+ZINWiq3twlwPW/
xdWkvMk/ven2nYY66xNe+cTuDAimOfCP/rYnMGii27v4G7mi+QzZHSkDVixN5UyH7Etx9P2qD6BV
8XAVD1dgiAoNuolLcLdIIXqwVVVYopmGwC3vm1aM0blp2SruKqOp1TysYafb0c1oqgPbaBUFAkQM
vcite7tA2W2u7JhcfUF8DozTvglFwhzYD/UxR4Xhr4y7efnLKdGHz4tKj+XyBVVN08jsTZbbF86e
x3FWyge5kuU4Bz3AHWb7UWN3Q5uYOau7+f3OTPUWmaipLmiGMry00KpaIBUidG7mxSW6bgjx0nvS
onHV1+fITiLpVQAXnG/lK2OXqCANtYB7EBHOkUp3oARnyLOCplWCXWabS/yzo/BnCCtmCWiwSdvc
WkW4F09tWn/0/uhErHj93yNqFqEFHaS6yVMYG71cEBH3bfKQXueUbhnfKncLz9wksXeSLpaVHv6B
E96K0hT1co6C6CttSSktclf3Ag/nVlJDY3+tSuZU/MoIjn0NEgQhKw3wUMX8YFnqtUiu97X91bNc
LNRW9ehS6xvlwTroya8eUz9RpMX1RLvaFY+6XCxedrafOI5rKo6RF6Iayi43uZb736nWLVM1BYpY
0U/IuTW1FWz+WTPW6pPYA8muBM9hSOX0+IdDYXo9+A04BRew5g+m+Qg+RWQO38k6MLI+zVyDsBkN
AFe0Lj7wQXuMiCSJKw2M/shlPq9HPKFEvdVlKBKgRUsrnkvsGYLETRh63fXroA8Jl+/TEWpp+1QA
CsMnpDyshR2XLDMEZ/gdaaRp/u/DGwY+UY6SvqWlkxhB8UGmYwMeXfVW92bEzHh2U5GX6o2ISmqy
GD6chBvwYblCb3ART/q6J6s6Yz76s0jB5Gu1NEm8wgbLj9c7tzazJR75VwoSx9h3V7DWFDK6/FwN
3AeGZwu9vSFsVZ2VoHuKnxvUJbs09YUfR0l5S12i7xgDt/IOV7p2Lyb0QlRvUmVycvdByqflWsa5
usOdlbUe3HEfUPCvObyAh2j1955DuxGUWNNfjBgZucZ27lPO6SwDWJLzHEz4NqRUA5HXxz4mcp+n
3p9WCzh2Pt2rQ3/DcYYsB0U11tC2/kTh2+WPfM0vLcXH7QHsPOSuJLDrjSPudT9tV3gEKGOS3U6r
0k+rc2XVngu6FApUWjdYLHl6kkkI7y+tAgTGAOAx3XGY0rOGHAgvEZKX4lyfir5DPTVQnLN51Kb+
EAeu5bRPhcQpioa77FG0KDUgfH8aDnaFwc6kGIj1JUjqDjHF6z4epYOpmJrtxe1kwcqsP+l7/yVF
bqfI8RAZaZbHGnVLTtp/P/6O4usjIMwCy3PZYIXq6qyNorHoQxcq43RebBp2xbQ0xCdXe223p6mA
wRwI8l0GcnxWMTF0rb7VNWmm5zdP5sKnyWyMpXoXrdXScLet7HFtUSm0ZejH9uzRXNqkLUjtSS6u
8GBGcw8dknA4qdxOb4TrgewiLseAgGXd797/5uXoW8iIVqbD0kspHHiFevEkdMK89rm/FD/02RK5
+l79cJIp/p36MRHJv87CbbIGzZgY+ymw9JDp64V1evYYqG1AuHyXw5Hyjc5eu5jjdIoUWkxNa5oh
qSkQWFguGlc5UW70SGeb9ErV3eTrmg6tdw9Zbj//PPIJ8faUuVBxOAQ3btEtVWkpGaW1z2+R2XF2
EueTqxYR1eNjMcHpGGZFnYHF4qpV5pGUyIDh7hCcx9dV7v2GF2G2onceS6DtOBsuyf//8eUFleWH
cJa1aZ2iWMrAd5XzuRX4TgkRXJaKP4VX5oHpkQme5jsdUqvcjzQfJoiBqRl2Ur62nYcYK9iPsdeT
UFS4XTbwazUZ9exha/y42ncz44QyhdVrLtXfvSpY1OGw3dDs8gW7/EwwVo+SJrmJOw6QIQSZ/ul3
civWkM/gsEIIAlzYxLX9QZo1RbbjdlVbnKvETY37iddWBDZj/otPoxrn9QWAYw8CY9/U55/n+aJH
dpjwP9GwKOjd5ceEVDd7meb97ztnYTcoxarzzGObeHkf8dfqBoApm/ZMdtMgZRGKzX3dfr4+O8K0
LYDr/Oa/uTHZVdugCQbVXr8KcTa6O2Ich+EDNie+G8vysQA9LPwIQyQtqebBcZS4IMJF/SqritI4
GnJ0MqJaLvE/rwPdapQ1ludJ4J1w5w2eFqINjwPQCg0QmOKTbh1WO1RSiOq1raXFC08apRoDPu9K
EktSpUu73ieS8FSlf4L90zl6Cofu+ZEUvsGs/9cC3B1wfa8SMKBrimGimfwwaZbDxBNW5ADQKNSf
yMusfQ0aM72k0zd5fPgLLoPBdadY/n4BnzSoHKRhKTYlWMhJrA4ddhfnncjMEn0/SUEwJH9eviCT
fZg3NuF/McR1ulJCG02UV2ED+RckSQGRJ1XeV/PLa8l50QDckaXJK7cPuOdPA4A2G/UtP0zXGgco
Z842jHzUqC6GLw4G789LEqld88OyWitkPG1bWBF/4r5Pok3a5tcZgUQktWCa1x6BHP2kiTMVJ8/X
FaxT3kLRqryWxmgIkiSkzCPwlUxOXjrSlLmYj7VAxooUUiQj7I7QlEzT5re/yzM3K3SF7HSudan2
C4G5gBVPHToSiQozuhF76xHjnIZB/X1ZXX5tNQCaIlF1VcV4uVnXmC1gKIANH5bKwIjjKOWiDLaM
K5je23381QPBrk4fYzWefFOd54RAOscta0woD3Sp01z8s7AeW8Mvi/8uxqlpKUb9WhIMD+DbYix6
+16iUPZ2+LMOEuCnZsrbsJ2b9SYyUGUxa67JGgaJt0+k+Q12Afd2RmuT9PXoFgkptvli9toOxhAm
0AzUqnoAraMKrLBJokxq09JnPsGvAeOCKhkE1SFuT8ENQHgn/6ohy2LPDalHAUBzUu1sZbnqqLd3
FFPO5Mt7vcOiZtklEGH98h+dRr9f1K6vCAWJ9yLzbLRfiZDQdXoLy4ZFtamiqQI3VRSrNyhcUavd
EasPM5YxskX+riFcf36ZjsoNEFp9HhV+NDiPL1bvsRGp4ulD9jyjZHKJrk0oEQVKgLpfkaR+O5io
WoqbmxcgDOPTbiIoWb9tJLZN2Xn+9PEpOBGBTYIx5bpX4VQIHFGO5s9QgXkqisvLTnjagVkBu7cn
Y4dCppoLknQg8v0TAmlK838pb3maUI2VyRMeRmPrW49203i6UsNgBVs68/UgRIqF42qPGZ2ZH6Qf
Hs0oLDe5ycctS9WqZdgxnijY7Mm+hrk71rLdDvO9WOTIYLfd+ao1/yswq6TV82zi+d9b+uy/QcBT
/jKgXuFD2W4ozyIRKcIlwXJ2x8RGrxuVVJfe6y3KHMaeDveeI9+K5jN4XrykAPZoikTBU8Z5Z7WF
Lp0prHRfVn4pmn+itixJ9Cs6WVqUOD75Jd04FTv0O0r6A33lBvwmQ/5aHM370GJtUCfZFUo5HN5x
1ymwJaV2e5V3fvNKIvVfMw+sIqPXSGR8X5FSWrLR5KBJ4Oxx/O4fICIWWL+99ICTaOh7jW3ZTzWU
wSLN0PFKerSa8ahh8+lFSp8eYt/ZIqMI0m0RCnCFUuesF/y/U1kxcVfcMqWhiWTFM9Qd/0xVrHhV
SxTqFEho2c2prBfKbO9Qzmet3fvsQbDcMapnVgwiTEzfFYUrybSWsv2NmL59/M1+wipfkASpb1ag
S2UE4C0qQr0O/ohSpvJXVvT7Yl/U9rutvHiEbIjK5J6k+AWSkOIM0dubFdl0y3magHM25l6PU89B
LaSUEKlN3Bl8XL0qiDXmdZ1KyGgX33B/fEM+k/22UCRdkxHgLTkGC+XB4TWAO74LJTpUN0fpchNa
U5FwYQCZXWEf2Ty63Te+7mI3SwooISVVYvMHz00CjajDrXCiC/bIPEpukHyeIbmG4Ovx0Z+ys3KS
5YbB26EdrA+DbkopBmiQ6Rt3JBHs+orUz7HyuwhmNDEWHonMKiZuQDwleptV0Qz8UpjQm0IRzNVv
DlLT8AGPo9uyZjO8KUafwP4aRLTS7AWKo3233yqOXjCfWaylfR7mazVVS9qu02tRe14UjG9DsSG7
90TnJl7OYdvNL3X9hHsGdok0gQGh1GAsKcc4tA2pTnoRuIPnO11qn3ygR4Pda10YhW3yvqkyEw2w
CEI145EWPUZ1z1G7cRQtaVur6QkjJ/g8Tx86eiBmiqaRQ8PDXl3a3A+oJyXpYqEtpc+HYeBfeIUS
tBCyG3OQxwimMD9B77By2/KTjgqmf9gLcqOoAheX7lFPioc8sJIQKQYQFsYhhsgq3bgGkqlYgzXg
ItXKDv0Ga/ZcYG9WZ3zWLNBw4sOR9+JQqo3pXDW1PZYLOi/0/2LKuIXbY2hLlakdQ7JRsWApsX40
UVAAyaDjWunmcvN1yy8vPpR335v1d3NBxHCm9/d1hon2NjLeRaUaOZCA67GOOCqrUEKGEwjbStAo
DuZSBO0iLOtzYyHsjiO55wATgCD62Qo1mBn8wlcdGz2DhN2lnHl1ZlERPBeNjkotjMqMhkBqZTlx
GqQGqFOzNjbQ6PRkflobi6Y6voGhLmgQPP9InnhIdekJWRRkIj91XupvEnSYYJ4FBfCt5uHqNqSI
yAAwmUw1Vils7nDcQUw5yvEXPRK9oXdHtPG2ZeqWXlv33p8wupXUrN3Rrj7lq/nx2FtcMoc3A5aR
gpLPb/e8zwMmqyFbLyHhKvhG30MV6IC0h0o7KzupTyOY/yuwaiiGc6yO97c3bylxDId3yRmHk1Py
VRhm/GF1FrBAQ2tlzrk1k4eOEIUMrBsRsLrZfcV8cdlK4OmPuoDbENHIjRDjh7BJHV2/I8Q41gyw
5oMenCDldiIZ+63ffGudGcwDNtXdmObwyO8wplLwimB0+oiSuO3ZE9UMXwzSn/xQb6SOR6rlMs2E
xGKpd7U+eYl9I2H7mCJHXy6LI34Knk1JCKshjSKz4JayKE1eL42xb9bCwcNahEktWIVbQiBFZI7G
ptlafc2g7XspV9bjy89rX8cidDFziuEjN6xYuXSzKTgjDNRsXgAg1FdgkdBhi93z6Brrpi/Jj78Q
ZHgdx9n1ex5puMnYRufifBrhSZnZ1LCmaN8feafAPYGVL+7EADI+v9Z+Rs6EpphQE18hdZnya8Lj
8S3Stw3zbcF7Hdb7bJsTQWv9IHE+j+p6+Xkke/NyG+nbVcno3oJeyyYXMiT0mn3TjTE1Ql8e1jqI
ipffLN56QwEP3RmdzWWGI+IrSMNp552w/wS0nQ/CBQdTntVibiAtrfybRSbCczxn25O5xmqJeh1R
kol8NAY4rO+8EjQKTXq3brxLXrDd5qTMUdQtakyIKhVsmxl3HHH8NK+FGHBL/lk0aeDg2WHxaBRo
q2epHpjB1kTfQZPYSXKM+tB/bos7PD1FOfRdWmbRZQxg1EE5zwf9bAny0VwFKRmeoa29kIkvnAj0
SHyXKVHHMYdVDMCpf1NV8gqbvzMdwpPz5ujMzObUaffdOsYDNERimMn8pYaGQRYAgTGfe2Q3oe+/
fH8asHjMiIisTzC5C8IpldoIxoEFFWw1KInCM94kurxVmcElY+y7H7kKldGxAzhOSTNE+IQV2T88
3ycVhXjId+zKQ80jSwqaTyqWmBWOWvqLvONc6SGWVTKdZM9Hc1QGH3C6qJIL/n0hgq1wlKsNL1xK
iMSM0lOtoYKt2aE1m9HbgRZgWpKhisSY1VKamT+d/ZlIEWOg37k3snsMfw+zDGr0Ip/jMo/ZcdAV
onMagnyUMX6C6uQri9AtKnVeNm2PTBIBos3s/65YMuRmXaIYsl7Uk58Cb+OMOH+/eg2XhZfZUALQ
3BAAL3L3KG+0r5aYvX7s8NGIaZST6t2ChQAhRMWExOZwoP2n1v+wNNswT9RPVdhbYHObv5OHLCua
4FC5vdim+KEzC3aZcZghN5ja9kIhWO2UY8WjC9JKfC83HcoEZSRTTj1cg9tQdL1OlT3LuwZLRecT
+gZIuGfIZ0yKqbpb+iJRJoYhqV3/xmYgmbQyp7tXwfb8kih32CQm4+IGS/vgD3p03JiuvQZSSo+O
z9mOaAQSni/Cp4m31Z1QVfyrFVu/uGNPwtWHfljNaUFYez3hwnA3Yr5OJGTjFDN+FCLuV29WdyZ3
rzFZEMuVPya49BwbRzaU5QAUfIYdzao3qYG+p/Rshywe1TjCvc5Wt7KYS6sG0TvU+Qby/9/ApiiX
VobFDTxjVN7gZrqPo7gi/iYHHV9Nzc3tGyig9WDDVKYX36nsJKWz/T2ah0GANncrBQhsiF6ce5f5
TFpAR+kh3qFxBr+MjgeGu3ARtocvTRdNEUtdcTkjqMY/1rwYncl2tt5BpfSGiOevXQXSpgX3bcTm
67eRTqYXxlM+2PGiR1Q+7OWDfh58oJSKYC+sk8X779VmLTMVr3E1mWO4GlCp+41hp6LLxUVMT+Zk
ng03ns4LP5bfp27mnd56fM9FxqBlIDnV7VfBQ72zDufrhLxj8sRX9fZwp3ELF69n2Eg8z6bLjy9h
1XLNXGQn3MdFwKggGDHQxHKPWqx96cM6ZmljA1q54YJnbcsrcFhrFaKA8vnM98Ib3gKQBLcoQj1z
zBPQlSZHWWbxzFAMgADH/TT9ljvumURb2v0gpJio7QOuk60NtrmpX39y60GDperpfahVi32TOg2P
guxpb9dawUoT34Brv4VwKW/hwudPb5LGQFP5IGL9tdSj+YKma3qFMqpdK+fU2FaIKolVUp8LrGuz
cNbIxggVrMZ+jJqryy6U6q43mhQAGlcrrxY4S9IylcIno1KNjvwDY4ogqXwSZ3+eCPxwLdocODGS
mFzzlcJ32zLAWsqDEmBH/jv52Q07WoQv860qPMToFukot1E1rFQKjnKhDMZxryRyrzfi97gFD4zu
u0yCM72EsIhFYy5IUxnpiZmxdDUITkD14VdZ867QaJK9v/TLMeQYGNBHDtuYoMLasiCTQwUxlpVx
iLB2lzWm1CBa65c/Ibz6O40DZVZDlHtpl6j+R3mJIoTcxa2pHJzFQbQx/ElWGgCv0FzrTPpUdt5c
c8VWncN2Zj2hXVH1uiHVxhb0eFZBYg/IUGYf8P23yDNZ4ZreKAePGJDqAFXjOizyF20iQqys9WxK
hTaxMYsmQgjA7t6y5zagZaMMslccmTZn3hrJjgvibE+A+juX2fu7G0Ma7J7JIQaY8cOL8tLGC5Zp
tt5piSZ7lsPIScY6D8N6/ivYoqZMOQgQhy0pKV7r/kdyXJ2Duno9tJWM43y/k9wmBeKZSBJeq134
NV65sYFJw4MGND/PibqRq7SAwul/UDYkGzClYklJ20MqRrSfFA8EmbAbVM59nORqGq32S2eVdQTG
79mwtI8fFXKIZzHF2U9v7wJu2NDa77NO9M2KW5+p9xfQaAi8Gl1LKZfPVixhqmI/evDj9AzqEn9J
Hn8aIUlkecn59exJltWMdVkwv3s2EHF7FY/ftOrLkt1gX01vTGYrWlMqQ+/tFnZOWXr2j2pZQ0lT
ImIBQarW4dKDUd44cMe32ts/Nyq7bQ6Y6a1hf1a+k4Dp4Kce1cWF832NPO9OPpbrTdDqWE9c7YZI
8unJXTd+j9gGtER8slxBto/HiuHw9v9/e1n2AAa2l/AHKZxOuDze6BprKhZncfcmsZe1Z53Jo3HR
IXV1TPueaMNB3o6/K3uTkycP/vhOK+Xvl9rrmBzyOKXHA4XMzxJJMFYlMc3gG/YiJqYIby3rBewY
Gf3rN1Jblud0V2ZY+FKe/gO8Snsb5KrePVCylTaLuAEZdsOEhocqnX+fS8Nh8PsdLTBp2EFTA445
gFfzWknZTxRGkIfuF/bz4Z2RbbUF7HOn/1jWujh1eiTwdoPaSmQVUPrsuZjND9xXN5pcDfJfxKO5
Rvh151PssstUdpAXdXXBBeOnjJEm4FnOk1N+4CEBgf4G9xr2jCRDRpQYHwIi2cgFADY0vBt2LiLv
EipbOMNu9TKQKByoYNQZVIh/NUnn87SZpm9XXOuoB05HG7RgmKtssBrOV/inyuAABUpz3LXRsb5R
oT6+iM/76dnojA14hYtPvRuhWNPxN1Tqv2PEMHrHhLGrkDL9heKwDjIz/doi672k4EZpjEziBS+f
QGhA7rYjEfQ3rzRAw+bufNktqrKb38bor9bywOVkGvY6KaQPEtsNkOi6KEunU0NySrmGgdwBlU2X
QnxqeJgwNr5fapcV5+gQEC1LYfZCaQiStQzlc/ZJEGiz/774nzPAw24saazQO2dJrj7Wq6OtOpp6
/rzXxMmyAXzRQ7SZLRDsZD7reTNSxyuLCzigw6c5iGceBlCdG7kPAgn2hAT38sPxXAjytThCHqyr
D3P0391cWRS4DxxUY97INUifJhG/IyVG/6OK9otPPm2gzrCI6X3MGCxstlgkeyrqfC0z+yHYYnMM
ct8CHsUVlCUXKJDavMUm0aKLvjpMofswXqeHYzUk+QlkgQqvTAJSQter1ZMIZphna5nzEgt6mZlb
Vk0k6k/M98rV9td2FsniEmD0oMsmW4TBROAdJgSRgpH9Ml7ohJ7u9MO+lmEma+0hIHssS/cjn9bY
tBp7r3ge8Qkjw1X1Me5z5zc09ZFBz/63Sv9RUxnNw93AptDAdcVxpPLMsNQyTB9b6gbAecm67vjI
oNYvUw+Y+qmxx7nHnpfdXXo0X/XZHPg/2TQGg+/PhiIlli2Wl0wgf5EuoEYxpvriWZnX5E2Y2I1Z
/oXNrqCVMiVJUd0df3OliBO1z12KzsKMqq7Sex8ggPOKbKDnaF7M9/WwOL9fpuFG1RuosKhz+RIr
z60LbnD+KMImvpc9yDsUtUGtW4APAJh2UtI/D65m5lhuRi3uqE5SXKOCfax2GJYcxdMT/VpO3dWz
qpUwgSK75RLWfk7KxJC1lGTxNK61Rkg1LelAJrQHd3SKUcCh3U15j8ornbjTtOHe4tc6NeSZSoaj
SnlG4YoGSXC2F3oujuZZCFUiY3+/PP/JkK3WQlmPUFer+VC6QjgEp4rzTQOQw5IeHfrmWPmrFs2T
hRDDfd9K0fKCGjdIn2CYRpealHshMUDxOtIVKSIvRKJL2SPkt6/QIM8pUq07LQTk8oh1NDR5Am9E
IHZU9xOL7FCIcieIPaNeFsb5hQMyOH7y1yAIDfDjgYyaw4/yiDxcJJkwNkFvPOclqOuoFJRasS54
z1lBBNGkPS1Zud4z+BweqNFwx/8aP5timyt62/QHUGKEwb+vM6X7j3n16gxrol1eDh3nKC8gXIj6
o+dcp9gW/+IqxI4LvsVX7RWfru1RYlywNp0GKP2/slMKZyRVel1wVM9WZb7yygVr8XNK6wW2ceCI
A/8k+2DC1dJlGuWFeOaAQ8+PaoUC254MC/r7vV9xgHuqZyBTmKKxWvoIOwPcXmzv+QfLdRcl66nl
oVdljoHQxwO6GoZoNRnywq3i6N5TMEoTPCYyLwjnMdSabDx9CVNA/IwnXKdyNGsF15w7Zg9cDeRK
JdNMnlus4bP3qBQ6AxFV/qnc/HR0BeEosNqIfIgJnJRYzoqkmTweAqXrlY5UWesnjZ9eUhZTuYLR
araefsaWabpJfLarbEE2CmQZUw/Bbi66L+pAsaytGk01Qs9KiBpvTN/1PI/elaYgN+Xejc/ly/n5
pgQRzZuUCyMghRVAwF3wNiIpOaobpuKGcTPaM9ybC4067egsE+m5k4x9nA9M+kxoX6gahdDLPrkn
jaY5/Ab5VdQKKTq52+EsQIsIPA3qPfXnJCj/ri7Y0p6IUKzbYDzCzYXghL3rl8pFAO61U17dHue2
GyKAUHmIVgD84GBZ6OjgY/F9cN5EIWvlMB1qqAiquwqYVoLQqS688qI+4H2FUABrIyELGUYhlugH
8DI1yyZVYEUPr/5lPDs96j+qd6CPKeg3/5byKy5EPLh4vq/uQ3NbP1HezoDvbVEFtXGfI3Bv6Rb9
2Jqdkec+Tw0WLgmS61eDM9FR04d31EDXrULaL95g2pQ33IMIBaQZY254orrZcCqAhC4VieEsJEfO
MSG9iLvGodW1yFOqyWDylOr61TF0+zloFUZliTsz6elLF0Hqry4eKcCEriaVthZRRKDdvKtzW+p6
U1Xg9Lyjtie/54FS3NCcVfqME08EzlWGSZjpfd/ikBtqKLTTIaUqsy9F0jgKK6oWno9dDt0srYBi
oJSRFhLl3u54u2tnU8KsB6gejCgnr9Hfrp2r92LcGP5EwuL9XH4RPfVJlFcs/mpTQILpY1pPuSFs
mzTyv7u+KBRgyNBR9hcglkHvN6iX9KuqDb7rgu2lFstEZNGQSzWFN9DKThkTndPaW9/cAp7VCgGT
fsjYrhyKqgjni39ViWaUwpW3v4ygMOs8phNM2aHxEEpm3UMYY6LYQm+4Crf0vWJcgM34fRzX5Cyl
aVq0SrBJoJmL69H2wMlMJgetoxAzU77V04rO2qJW5P1sjtGF0ATj+pjrXWTOSMRpJKPFqm5G+ww+
37lLN/mA+fEOWGMWVpQCriicLu3PqllxHrDSgHBH017lcfDT+t6pApi3ld9kM2TgBSzIEjbFAFZd
cJbHMHyVfAqi4mxpipu66A904MeeZJULcrGJ4gQESziVxIEXqsafHMKfie045q7lQeJQcank/2Yt
8EBcJa0y9iVl0N29tA5FOIhnI0ZGkPZ5oZ3QVtBNV38kXWC1QC1R3HIstHKgznS8fSkmHu4pS1Nf
yHwfQDSIWkmZ0WXjXrT0ITANyV8th3mjahssA10b12IcnGAcf0iYXAlRr/Q53jvvWZYvArh7Oy5C
Jq5fa6FK96Pj2C7Yl2un6bHhfHl+pQUJgiL5FBH+MozvIYc9Bv7hSIqyCANgrpmcWmwrLrzrfi2Z
vL9397L6Xz7pBdxVZx0xkY88kfrXoBGWkjhFz0j2aBrkFVjMBwEyOJ2C1CEGU0CwiLp3TdbGDa3N
T3I+NdnthyVSLbzD0BwNjB5dvk49Cny7hMiArwkbbnkfzQTbf2/tTfW0h1Wa8Yz9wEOCSxx4VP1u
A3tW1F7KmMGy/mqsUwrOE6DcIk7duaaY+OQ0Lj3fcJrnl3CKUsHb8ERXCOXDFZxKuO5LF+J0dzXq
kzNVd7brPaeGxy7WaStNC2Z6CeJHpR4no5bWV+wiGB0Z/mvqMOH170Dlq1mOL1kCtnyJVQeappsm
b4P1wWmSkVKN+3eMZ34eDKCbwmowsnm1pDCc6cBEcMusW6yRmXB8AnqLWei2AWadABjOatCrDUcK
Bz746kCyOQSsdFgGdrhjWX1Q3wiH0JHrn3/8bB9LglYBzGOCaQ7Osy6Z0yuEE6u+2jfTOEPRE4uv
w6FvqOAIENUgouJH/Zhy+J9iqp+S0OVtQtPDrsEEsEqI3ZxvFGwR/8NSIa6gf/Lgn6qz8nTKsNWH
C4MwWPta+ZR7eGlRhIeMkzbMIWlltJnKtbG/2nTTLuK+if48H1y5RGjAfldpHKexEL9Qv+5wBxVL
br/Y2twnSBCMMh+SwRKEBNqqmYO2eKB9424cA+qIxx7Y8hUD99grbb475gS+P5NCAXJeoL0rnH3Y
309qmdoFXW7nCIVYPwfZTTITjH5eQbdC4/g9y9p0TQcjodclc/BQOhSWgwyxRyPRA8IhQD71CU/S
i3suSRHsNWYtpKc9kk/OocmU+fBfjd0OcQRl6bJRBKh0+XZOjZ7kQmMX0BWeIYtvjqCL9BqI9+Eh
ddIusyGBQrcErcnSzrR49lOC7pbxo5H417t4j7LeBKcO+/s4spJDmPm8P6c6LcwxCK8Iwph32j6k
Ihb6yyp2VUMqsUL8Y/Qw6AoL8K167cRII3OL2b3T1WkJpYbqHnmTiQxQ6K/dY3n1Aw4p7oBVxY6a
AE72di4k1sNdDyrdjFH/XYM2WhJSfx/P5Ex2U0z47EdwveVjtjXaCL9ALsBNkZriEyytzAktvh5j
XURX8t2AdE0/GKG3cWQbWoBcb80UOLgJX87ooTXlZuInN1PfQE1doOwv5eOfdtzeq+ZVQStl5qqu
FKCvyeX1aKTpjVZJaTAbyi2cSxEGL17p+fXToPxMw85dSxuo6JZ4qB1IHPr9B3Y66gtOEI/Dns3M
FFDsBqpXEM7ObkMYPZW+4Va5qh+14JE4Rfu7FNYTjMVNC47GlkLMpitYN+aJ/BPyN6E8Q0f7bQa9
LQK71xiZkiHgphsj8qy32Ks3ZFqZ1MkWsN24aT10rRP+oIxWiNwV3Ek0x5DU8KU4O1U9cScsiv1R
NChC5ahDFduRXKSuwDGz61ow2Rv1ZJS2WHdZoIyBxb06gDatWVY2J0Y5xG26SECFG1Pem6lXxlhF
5hdwKvpr0tw8tvD2ZCphQNxoLPgXnTMleYXLD4CYe7GcJZsdmu6bQtZEo8vRn3OH+i+8PI+BvFc/
b4D9GqOqhny6oy/p0rzjclRVXfhS+r3PYzBsl8rx1ZM4Aj58m4bfFQNV+mhGx2xIjt+WD1DBSIm6
axcw39Dju6sShfeAljRFSA8200frjs8AfwU/2gDaqtkv5saA7W5l3VCd9/qOsspAe9y66d3sO/ED
CK4Mzld0cx8oVldv754ywf1/5i+c72LRgnFGsTRsL7Z2aZPMNq+JiDONNzDaLnhaMCr+B/hhtcqF
YQzN4npaFav0uQRkXIXUpP/sbhUEfye4Fvjo9I4LHD3cZ6mhw/EcFvwS3owjvRzmWiR0mopY011c
nJqoI/87HmxfX2nR6dqRl0uX3LNy2zNVHbZQTzLsbydRcHQYHRy3IRuLXFO1WJUcp3+eLwtQ4dPj
aZLGYK8NSx4ezWQyZQbfyFBsOw/1XXJNxuGZ2AB30QJ1GzlsUfWXu27hzthNNMie9m6qsbWc7CxA
KORvTYNNZWcFPAJPZNie4uIBOoCmfY3eDU5mfL8KBMDkiOqNjOBmiphUNAFihUTTnWCCj6olOXd8
7kqcyJ77OtmNT9zwfAIPyJlZP5qrCHV6pgKLqT2fjeRSl2l5X4CYN7BD6052KSkxzpgGrVM6xJFF
lbYkwXuFbqwW0PGc/CjWsivclEcQdfbq4dIw+m1MnjCZHNiq0wCpeotj+ese4Z5m0vMLbnYZ+lSE
8dEh+qCmgKnpHpr5bg6CnGbdbgw8avgFTo2mKJffS/LQyqZQVFcEAFr+u8kQKGmSKfWFndMQmVQ0
i30NEcmFsg8vDYXJvlaPc3GltNwoCRm+W5DLsIwt5oYfmCWl5beuvzwDfvx8hi6wl42OFEJQuQkN
IPd4jmGWUuST+dxQJJhxCjY9vSh4f+OSH3hC+vPmKjEJhER4AS6pUsl1FugHfZ48IuSBXDai5ePB
WPKlQA4nfz2OdHLm6BBQSemcFmjnAKh8BZtBBcRvEbLIo8ZSkiJg4DC2CVi9ZKgRMcHpTEEPXbCo
ZojjuBvFTcVWYpGdk9DrEF7gBSK6RSuCs33PCRBRdDIWTX8Yp4lUJweYJfrlf27kRODuzstF4iCR
aX6YQ3Y/li57SaiMi0otkdpHuMOhfmws4NicGyuR2wOGvYkzhCQG5w4AVzBrhXMfeGusiJPfhmg9
oSgm1diV6tQctegnUiesn9pKzJK7gi1VZigOPhAsUo/vXW56nVzoOvN+HYai3hmuOUZ0um6fQg80
bc6rcLCw+YcSUh6orBf+alSFnomZ8LO2l1lFe8XcyolXPTEGw4RjSToWKlxIkOzYDFr7ykmr9XEG
xbvP8632cF7UNKH0B5JcZaF4BIRBZwkCLdie+Hi8RxJvkqd5qn2sQvfs5p+cSMLpCav4fctsF19l
FpcoQZxJtAPE5Zc+E5MEI4Kp17YseFDP/IKP/PKcdZEDuyD+vwXKykQOZKyDuD1Urv1c2Us+jJWd
cemZZ6UIuaLIFQlTRC6SZ1KYbDVJsTlr1CAOQqKjq1oz2ogInU8G08oJ71ggN7zx5kM2U5WexSYy
QTdD98ZREc9Ot77esJPQzXUCyIQe2IqBmMMQvywKBRIFvuXlt0AD/bkcJ4R8VnY7g8szsNzod37Y
6foJPI5QuaI92KdvTtPmd1m5yoFz7LdwzWZJ/LnEbwv/E8N6wNzCVSn8FAXI3KswpA348x0Ti/F1
2V68hKG4nl6VfcytsF1GEXT0uOHrdvZFhbqwZp8NLJoj/PSDaElSIvuUqSBPW6tva56JAk/lN22O
1S0nhjHlWrwggCiIVGQ3W8S2KVRzqhaOJD7ax1alj9JevPghvr2ZmtMoKu9VFE1pK7oTobkR5QtQ
6BX8+fJszIRrdRMxzIObSP+GFZT0VKyVrPP+Ry1N+zAK8n51Ttio1EGl/mwvkgCEFTWaWG8D/M/b
r23Nbi16dfNo+mWghUOKlhvVZCFlxp+2Ms8ewvnXexV8O/gB3xgdi2dd3pvmwVRQFvLGhIxpOpwD
OujmafiOk/GrK+y34ApzdYLBluTNoahLbdgetotgkcc7Z8vNR1sSFZNU+A4L7m9sCOV/UY0chPTu
9lC+CQgFX77Jr5lcP5n6Rul8W6w3F5PAkRTNIEnM/EtJyUsP4StWVVWGFDQ4fg8reX3S1tF77LQT
bC/jHjJCSi4oqShvM1mg8MJBrprtA79CoTl1EW04j+jJxW/XeAXkxNQcdaeskiT/mMsr5Kln/G8q
4gH67Bgmk4CJPWvinVcn850QhG5AcLFpdrbrK0MwgWcxqONUjY/ukyc9mMGO4nRoZSNiuWq79TDp
THE2sBaCFkM2BR1wEf7Jbymh659lhAopE3HlX5IdjBycUxkrIWgvISKx8RxbFRCpwDUK491UYQHb
js9KIxaBF/0VxcKlzulZQ4e+/PJsZThkXQM9AOU83M9B/bRMayRNsqKZ3gUzKq0SJ+pzRaZMPzjc
5w70+RSQCrw96ErtVe+v4GCsWSt/nNFkaS2UeXn1E5c7sWUitpmCUyfdbBs44hm41wPNgM4gM5GO
/VB3m6J+GKzeupUUs4jhs94k9PJ307ePKY/JMPCo0gmmGUtBx1/DBxz6OvfUSeiIo/yZLaSdrNmt
veJZ3CVvOY3YYn4lEIGZMeMUxhRfRHiv2OpCVq1x5VSZ+G80m6mjaZ+Y7PoxrdLWEiDnQJLF8iHR
25oAHTPIIEmFeJO6GEM4FcNC02rvK8hEpVJF5U21+rHsBI0V7rBzcOjVEwFV4v7HSt1OUN+VfiQv
xbDjD08b84T4SxZ4XOM26KjyXcJaE2wnohS2WkAJddv24QAIG5DrGuT3j5RD1AGa6EBeG1lHdk0k
QEdFRPL4h9hAB4BsRqdI4auM9WORgHNddB+QrmR2hxmcN/BuW5YWtliNesrrlw1CJSbxQ43H/5yA
7BWq+z/P3jQOmFTNMgDtfQjtC//dGezIIH5GLaQkLj3DzmcSw+qAZ09JHBMzv+nyZMa9YtDSr9xo
u410BzUennWGYWGU8QyFUgVhtiT3TVgkvSIkUqhFfq5OOq7Dx4DMX11WJwpEak535C24t9AO4F+M
zyBryeCTnof97G610dloCzaM4K7/VV1a5UqQ6KzGMO41CV9DSR96Toe5u2e0FGFheaO/5ccPLkbs
BamEaLAP+dULZ4XXZzHDDmYvQ8UN/jan2E8gWQ7NXDLBIUc8svwFmKUAeHL3uLhvOua9HClsUNFS
4anDH5R0Z57nymO/ZJeYX6gBxmO7Q5YAannl6xCG3YC2SzKRp0pzWteoecboX0YEYziqLWv8HkRn
WQRvaYQ7dGa3bSWAnaCLyY2BCMCfwolCjyAlsJHQxewPHPPeLKX2rQ/9OBwOcsd95lfEcPhG5bs5
CP4NGhhgqMIFQMcYilrdu/xweULaiAOIfsYpaf4LJoR44SxelNe1zDQQO3OrgsZykXbcbMs8O9vn
3O8Hasr42w3rE3aa1FCdJj58sYcTpq+uYxZSxvVayjkzG4aWnH4p7Y+pKOGgTTicoH+QM3YCEJFP
r5xvszxRRgYl2p6RC8clk4JjQsSU8hyyi5xTQ0V9jUgS0TkUSMttwn9+GcNJAGnT/P0NXFT7YHCe
0fwAh9xmy8Xuplt88iGQmCszUUyxy49J0/6N2bcgshC6WfNJngUWbEzz/lO5gSQO/6Ncp72XeOXs
5Oqz0oURd1DNGkUNAvuyrYuS58MSzEelwvAYzNC3FdsgSbw7jSsZLy1hc8p/ivYSZvarz09S+Dbl
AgZi/zRaNKM5zNSBNUrjeVZZi9u9Rbc+9Vk5Vl8fle/HYuuO/qQnpmywYYe+iXu1+yCLMy7+qUTR
D4w2S8ykwqJYXsLf65C2kIqqW3QAGCQZZ8g5n6Qxl5GFqK0qNbBBivyD5cETMoV2abTREdSJMUB2
Kg3NNeTFkFWiMgNoPZT0qXFkXZFaze6nMXy+kSHNJMOBapqFhE/B41mjyZQEPL3tgdM7KtaQnhAo
AWAOhVhSfBkP5/XdNZMUaNMz/1VRPR3+9AN4igTU2Jby0LRhz50f1o+FAiq6nnL7+gi5F9si5Bap
cS70ejRyNvSdLONq/TIx6tQOX4MKAwwK9kGz5OESCrHjRIIdc5l3hCLlB/29LZBrkcAq4xUr9x0m
8kGAmkGsDkX4zcbB5VEZRGN0QzwMqlwV7S/Zyejfhs1mZDXXDbPsH3NWRQOybCYvhScxFPCqul4h
veUjFS0ItR+CI28wdQHjEQAp49aB68IjFWmQfQlB+sSt5q6utoPer68Z0GiZCwUD8DvyPyMjxq5L
7PcY1ms6Z8DNs8g+UmhqKn8c6uuNDkR6emelcqR91xBavfjyW7SvO0TEONUZ2WZ/7DukwV26RtL/
m9XX/ZKkwj/96GHPhzfcr+93kJR7sFqw038T7ppTY36OMOMdF8UtNt/sahTjrou05xBIJjPC6r3b
flJgl+EjDt00ppbAEg8xIlirQtXL9MqclWkuIZCqDQG6/0VoYYR0TE3x8VxrFAl/lk+wkgghlR+A
+d/La6K0zrMcf3yQyN7Di1DbHAHpIf2DcnmIlUE/63TIQSKD3rNwsQ9p460eBh0+XBOOtwEd2Zkw
5mnIMEvIH5xvurdvmt85Wdc8f+Hd2fHLn/Yr9xiMtV+DfZCu6/Pd+ZkTe0lyExKWyA29hDPBlvf2
A4XAoJr38uUaJJ4KIkqBYyP7gg/j3cRl5X3VAEIPZP4v02nR7NaaSAhk5nc1WZB3QXUwwFIEr920
o0lSTMoJf2hN51fyCh1mNnQSFtkmwhwcngUn75EMbAHwULQV2A+PQTzb1F/RltRBuqVDk4rifVvQ
Xx4pM8rRzwHaViXl70ieTfwivvgVln7KUFsZz0oI9nx+KeWyUZqyyEIkHtdYAq7+JjEF0P+a3z2V
Zf4k9EKWI5lDcdDtHFrTfKLdWuPpwpZpbx8TxhP7qJOYZGVaFqMauIYk3q46yLB86Qeh1N/J8Tj0
wW6ftgBlvpESAOG2XzNOdkCM2zKnWkS9lV/0FoUFQIZqUVzvTA7gujDMPDV56R/pcpyISc5T9z+f
RD8lFyhKQnKBdJN6ni1pqfV2Kyvp9zlW5JIdpPN0C0yvnwS6SJwXmruCFifIQtG0CZbTCxrpGtYw
DiR6EzKHoK+490uyaspYVs7Rvv60K8sm4P7ChLXV5nQ6t9LmzZQHDnuArG4YRdyAT+g8dY9BSbUq
/2iG3cgO20v1IYXulwKdQ9dXjfxrLKnW0BUNGtrW+I8FTBtVeSToPxh8Xp1VPM/MWSBWj36h7AQy
ALtIB9Du1N6hJONnZrXjEubE0aqTzC0DnMURMbKDLwLQ9kULIa2D+0hdpbEhg53zcQxcICVN6yYL
N670nTfXL0AhISPEa+OfeEmSk+A1qtuhJOJqV/XeOR9N0zT7/4E/Was3M8CtWXgHy9PW+PpMfvAl
uOMbAANcnSSycJhxO364NvilwubsXKutSOAeB5hJJ/bcuPVPl1wcbU30o0jgP/73tlXo9y0CYNti
yuA8H/2jRhaAJUYFYZkIlbdc1JVI/0DF4zKtOwscfsj/oGwkpmC9wrz6QN3zskJxQTspw5U7UVz9
oehzHGBHw+CLgvZ1ls861smDi5FR8jenOYU+MSsvJwFvxQRBejiJ3BKFC0ogZGg9k4rbsYuB8dNu
8YVj5e1CANc1dTYi/1QkcYLRB3Q/SHremxEKlT3WXMggcysBqGBbMR+ikric3zSU06Kl6n2eQhT9
G74OmjPMYmjrPOun3jTA8uj3yyn/88wmao00stCW1t27OCtyw+5jV7LvtFO9MoDO+0OlBsl1wics
KNfD6SvwCwyOSdzIsOfywDMA3XRmcDkLUOuRATb3ZmTpDAViBZDu0QnkpIjQCQrweeLHZlo4+hj9
1d7CcOZz66a8sUlbZwT9Suf5HnwLs9JXVMsgQlhszjtaNEM165JL23bxDNOkRaJq3XwU/prYuimJ
+Vyr0YkD3IQpZ/H1zJyJRdSAZL99bUEFIQBpX7yUJUXxEyt+IriOsgm+Zf0IE1t9UauD7pr7widJ
1iZwdUNYo+tQCjYnMa7GGOnO0IWhHe47j7uNZE/ePTaacBjHrEkfLU+IGyh5bvax6OAb1Xg5oJp1
sTo9uwEAwj1MO94Z7Z/TEmVpdU8yzn39NI+pZH6VTHEvmjAuP3g5lbjaHszkg913tjU26KS1gGPJ
YV+qsZTKPqgNoyqS2oH0NkfmEtNu0lXMWboOm7tl6j3ER8O8KHrvP8iC5SzktVfOj5qFCs/gABi7
P0Nn4KPkqPs+CvMFIyZ3ITuOOum2rASxCgM7kgTRY+Yw57K4quIrttmLKlzXo03qd9hQqeJy8SLU
9OT0ncve8LCz+6a4rfxoMsD+lbk3JO76Yb3owLnthNNBSdg5pYmtErNyQ/EuWgqQshV/9lKNNKW/
OPUZ2cfSuiOwyfRxwyBPFMDfMg2aG3Rd/A0vbOiCwhWSB8kgGM8JNmLV8jiNZrTL8w69UU9BAOAs
w0e6V6c43cgGBghU8etMsDRcTXaGu1ubZZdxge11PX4Z0pYzVyJ+dBqbpweaP3hylucId4Wu1sFu
ieYkA0haaPfR5r96wahK3YWFTEsUBf7at3Rz/FzoczM1l9ddxrIhqKQ1mO0qm5z3jhLEWJ32UxAy
WHwaIZMKR678dws7hG/Lv6R7hT9ZBI/OMY68NtBNC9t3/xxfjrQfNgEOjsMn6slT1ItgIRKnk797
pbIRzGpTALTCeMFx6658mVHTLTUGTvAdZDI4c9nnb+Y909SLxyx+Bp/DxWhPL4PQ+vo0GeWEQ7Nq
GmP8t9smnjVaoX5aDJvpoVq/nFMZ38BXPAPWISUfhxcXbHydVTb/EQ3Wra3NPJxv1VQnRqoHUMU4
FASPI8tx6/ZtkEBPwyoE8CVzsPEZn4a86D3MkGFr8agD7d/EdYfQp2m9986iKJvCryG9rPeApjNl
javSjXUzF8vUjxjJ3dz+Gc5AChU8ZnDL4TZyllgiIH4YVf8nbcGTAyodRddvYyKfoEfD8hrJu54D
np4PH57n/H1Ws6RPWI7QYUctxGwt7VmMak3FFMsU2PhgfgUfzO1MXoes0tXDMc2IqlpoBLQUavOZ
VjMFDkW4JnqjkdtQrV8bXGw9YayW2YAaRomgrvYDAG04tF/+m5ldrat8zdlPPvme+rlpqHoIYNi4
gbYYOxDfX2kR2PtWoLqsluELNy9JHDwx97Z8oa/0F7VFD6eUTy8XFNy9Zl/Pu9+SuQnXz6S8coeC
JvdkO8EIgTx4jMBGGCkQ6u6oTfCxX1YgDSW+9I6ez/zyRNsK7i2PocBt7atQtnfspLaFjprJmCOo
Ej1Kndht096lf5y1kdXxx+NjjG0Y6zlSLcNKIZASbMK8q3V7Wfrbh5puPtW31+n7AtTL6PayXBKy
KhCmhd+JGtqGAT2DpnQNVY0KoUmt2BHrx3FjdY8+j55a3UcSWR9gpqXnm53BB21CyBSj4fcwJ7fp
k7mrP+0lJWWWqS+yh8ueGfJ24npFBmOgYGZUspl81fn4ymh6htOFdCqs5XAGd87hbxuL7NXdYmUx
Im6drHXiizokTWMTwhwcw7Mznz+CNF0ERA2JFZoUNB1stIzSoXVkQd7LUWxeKaR0uCSb5xCvoACp
P42YQV69cz78akiZq0/mo+3vP/BcSf2IUf6h6w0G1ZZJtwUgfb6XdPQb9DAPTkUZqNEyJgPyiSN/
riV1qmN2pc8Y13y+wh0F+nbvSauniWic6JQPAJNjUn4t/0nnxCc8FvLrmiuG5J1IoErlVH8sxQom
MMoxGjHjSThOPBkz8oPLSpYLcOxHd8tpsyhxPeRF05/dPJS+De4LFgdUL2oO753O8HleUNuMrOiD
s7XbFDRCFuuqnCZfORiT9JcwRI0p8cVx6P+iULMaeD75IfBwrD/k9mUxFI3l0RLK6h7cu8MUiVLU
Y/MUFLGrNw6rbWfdRkPCP4MNBymGrBEF9cwBvEUa5VHobcPrtJN27aORaNsyGI/yNIhw1an67xPi
IZa6obuB7qXy7JL6jRocGc+x5W2Xr7iSPzbblf7vuyQE4Di6VY6e8SsujJFgpk76rKccTOchtJPn
sEVFBlPqVmJxZk6EmErOOOAN6PwTvL/UTWKoAzJfxDInLWfmAlOyNqNi/x4IUFhFKN94SYuFu8kN
/ZMAYToIszispYVgY1FIRPY/r9g4ZYP8QBij6332sWKBW4Gmwor0i3JX8ilGIcnj2oYTIRlrp8k4
SDYgPCYLbmk26xswR+v0UlHuyNAM2H6uEgNuUmZjegUhAu/GMpYTQ3teeQnkScvWiO4/Ouz9bNfu
Z6oQ3lv45JHhPozF/igfLQs/R+iGxfnzk8G/jOctTfD/owoTPm7ERKfX2mWx/D7lSrqe7H9ChUIJ
uwVnhkg/taDtd0sfJe22H+tUxS0NMaK4eIA6gGgkiQcCsXKsFkvp5uT4aLC7Hy8IzrQd80q0qPIq
3tfnZ+xWNrb44NRD2k3bqGX0KosU0bSzUF2xmSmOPsUPaXXjyGEvvWPteJ9ImgwX02niSLCiDGtd
qPAxAFxigUe7nAf/i8yJVge1kMk5E2KUW/Nf4oQdkQJPAtoXN7ZWQ9KI9Zfiw7pjPfUyZXQ1PEyG
YtWN/xQJxJIlmF2kWsq7yjFYEM9affenYF2ul18z9jzS60wXaBRMnftqlr12BnDnUSOi4hzMd1ql
y9w1ubMkAnG76M+luU2ciUO6kCno+RkoCJSFCeL7RPaDaGF0KzJWZAhmO0JcrGosgfUWxtmfFNvW
fOaLmBZaVG0icOT/XwXNCYVvTscohUABQN13hOUStbXsfRGhayH7Rnzj+flr+rfW6LyxwlcJMyte
t3jQ6on/Mj8Km0ug5IJer+2A24VkNxXTGFHgsNLjFgRpiNru+ZnHgzOlfDEja6BdemXIZHrFs3x6
yYs/lxUw1RGw8kXxYdrgP+V11uau+PQ/WqO21rVwPEWo07dXm76nwAOcZcsdtUOJEaUkaJecjSn8
MxWpmbGQ7wLwwgW8MeQjW302iVOooDahIOKdaMhZvmUH7qvTq09d/Eup+v3AgETj9hpxnO8zw2BZ
yptdwuFyPmGMjYK3Y7+bpl4TdGPSyN3JsoHArC8oWTqI+UhyrRs4TbxHnjYBCkARz+VJs2vXH4Dh
bZVr2o0dprcAlBLfNR5OCjSYWnN5Fr4oVIUM63AJ6f0JrHqT+atvHrCMDgB/rvdvPxh7xWN4BdUO
K44mrKJUbl/ap8oNestnWcENMtJe+Aie5Vz1+s3w14HO/ApwK6x8n2yl1piYdaXivWJFzCYRaCXB
Q/alVzOrClyMRzgrcUiVkP3p7+AP4ajkx4NzLxExEAS62cyVIEbeSiqHrROsQokv5GiuXz2Fndwc
JLDUwoMMwCeEO1EOFux4fg/S6zG+iJzsUA1A5V6srkHVJ5opv6lBlrdXd11XlUn36eVWLxKiDvME
szSpbWUexeGoKHeFqGKp6VjDR90M6CGhdgm4x7oP7HDah7pIiStXHkBty5exyp2yUoG5ZeO9vx00
tJERCL8ev5kr0WTtzML9pjQy3tQyJRwVAutKa+KDGIOzWbWZiQePToRwDuoRRtQlCbAHZM3gJtLJ
H70LIv88OwMPTcU2obLFonJBB96ZGmNJaKpGn5WPl/h8mrDFs82w8IVi50GIuadP42yT3oLQs4mH
U0I+ax0Ydef3t11xatZK458elERU5v0UryIuKdzNdpe1Y3ApUYczOGa7nbgM61VWkoS4jQoLyLkN
VEDAe21/5YXqvlkfXm9a1COLretrGRos8U+74DW+3bhQ1FuaKoQ+BuWtjUxFxW1UVPtqkJcNuODA
hy/0JqCxyPHsbE8T4Hl9PXEJrJ7gdCnZ4J8LVTI3Lf4DzoIwMQk8fkrMLfU/5wijxm+IvopChtwd
/wujZzNyCeb/ziqd/ys+3QD+O06E8E0+WtqdcTW1Sd/T1vTvBq/vzBpRS2+DSgq3IF5pE0YLDOl3
RNa6xjO6XxpeNj49+7qPXWpJNGI9kx4s7ihgYGYotbxUdhI0j4AqC8ZeSppe9AKYuAStBkFco16H
LGgU1QzFoPliwkKYrVjuZNsJx/feE02AW+jan7Jxb/XK7i77qhE91c0wfY3yYkvSNz7KTJdldDga
jSNCMfqy3Ye8Gm9UNvtmR4ZnwiGWCw4sxrGPKXrZR2r/ApPA7Qect6FnHWrc0o6HpKlBcr8Q8OZ3
yDwCgqeMptTfn5myyQ3oWA/9lc+eMLr7gqPD0lu5gCnftRF6z7omsqZ/yOjn6XGyHmqlF4PneokE
85EvG99mgVtbQqpQr39rvM6yxeMQHG0YvJJn9RWdyH/wL7fdxwRdbKvGHesZnh6uJ68Cq1oGFMQ5
wek9e3bb42aWaEF+urClaZGUHxUEK67JrEcyhxXQ3h85BEkWcIQ1m8yWBfCZMMDfOonG8jfM3j/n
kkr+bC7jkOwqEibX4rm9tRd7K+l87ZAzL6dzLKlo0upN20yLkNorwlT6tBdlhiArCnVrk0qFnxlD
82zLbtXlro0BEsxONRXADMOx/rURTb4CdtSObw16c/LqOn1FmOdEalszY74T9bbKr4llJk9FAukv
Xv4JmbcwKYDta5RKepOTZGXrihrTzEy8NxInjNJhnCv6HpNmLf1ylgp2bE8zLyMO73JqPy04cpFs
1w2Q8/HiLxAve4KMFoysiLNrkWtO82kTh9kV5gX1kKOGASV9aypjokANZM+rmBMtejlvruiuAgVH
9KCekitqOY9nKxEYSMhgEttXHvvXEaYGIP/kVW6YPN8x0wJmyBmdVb47x3VqhRpgYtwFg8eE6HcO
/1Ij3gETBgpa/DCZHo2IDmntx6kGeoRjxZkchD5+hgZVf0hQ6A9feaZqF+/im7NEMoxCAX0RLA7u
uCPSlTJjiJCV0nR1QH2I9zBwokUyybMqRyBOPRjQ8RW8qz3CEpkmXx7UqGQpiosC6vUYXc4FBA9w
4WETS+/UGk/maPqp5IMFZYlpCb2Mpppmc4zZc2okJRbei88RIqE/tff6+XgKe6tORKR8g8Ga9mz7
J/E8QOixlE9KnyDhkIKk0ksxbjZNxnx/rBGN5iC5CRliJt0gVdVBSfe4GTgaqfEL0RpPstWj1jba
5mXU0bI5Ei5TLH58EjqZFpesXdSppHvwkUzHqC9VetezwhI6UhbZDvXvXRfKmMAt2ENg4NRHOBSY
59UaaA1X9jNBJnQP2EXnmqrSqlJxV58A8ytBsh27KRoeB+wItySk3d0MnVJD9RmC/mfnA2YLctvD
2uk+iBjOF88DK93Txi3f/vi8yU2QkuaTE5WSCQg7egZACR0YyAb8pdjfRdAZCW33XrLT2MsPIyHZ
T+55wMmcmTc6l+QcMZIsv3xzC0Tam/kf+aFWc9lo4X6nUGK1RvJuhIkFAijdtV9dBJBGEtYc9QsX
eR+gBXglYn3+OmM3mQD/8U//nHpvTvClEXxMnhAMG4FM6Bg7rm1W7GPy8Ljxt0OplrQFmzQQxlCE
qLCPBLJ+f6lAS0WYMcisl0AJ3w3Vn1ysz79iZFdmKwChsFf0lbjgsNP+FUX8x6zBO0YiS4ZcuF+K
fRKgd+bOsse4W+ksD7H537Lzj92OBDKN9rq4OOmwrpd2TIa1PPl0t+MKLzz3BZwuInrsTE+Rnd3k
DhWI7SKTSIlyBYGjxPVzJQoi1ysTz4V/kz/p5BUquvMZdGn3Nioqc4VjoHy6akZ/c0U37TC95xfA
Bsei9o0Jy2fnPiUQ0ut5Z6EyuyRtjkEYpE/WmxLJ1C00iOThkKM1Rn5LTINEMQpPAWWTEZfSnbrG
rLKXjGX8M9f0YXzXJSh6pqQgNH1NhOBt0cjZaB+vg1/dE5vwQsmE/QSMygHPOb3X5nxNlIVcyeuz
CkQ32CEEZ5oPDIrRPNjSrmVWJyia9+AaPzcd7WW3KvKZeNraEAS7JKGYnqEzaf1OURwLG8q2WtIR
l0GmmG9PWHvntPErEpW+RZhMjIuTr6A/BRsgalpygqaWOPPmCy6qJJuG1k1k/SVGWKCCYZ2gn9qb
zwcUpRhmATa1W7HwIer2LH3mkdkT6MqzX+043bTtRhkw8oys4Pe3A9qD+j7uNx7Yew6WflLTw+fR
xjo5T3CbcNOHgCedeAXgKRqD0nVqYF76ufP7TbYt4JDqiYwp5PdIxlbJPuqRPIpRGautosFKBtuW
pUkZT9OIU0DB5dTZgi1kzSAlFbRXOg9FcnMP4NjWHCeu7AI3KuTaUz4I6qBvMFAFUkj0AXX1L8d2
lw2Ahm9t5qtluN7AU/A12XmgVbAwHkOsNsgf4VregAhue3uHNqZ4pLwjxB41KqmX4RuCyn2uE1uo
W6yqW5VhsBkKixWn2uReCFBgO77fMRx6pASjICt5qLHmG6c11doJMQjDoF3kAs7hciB8tCvAZl/W
UYhwWLn0m3NdzfYHFeGZ//5gCZrcXM9tp5Eo000xrH1dJwZilqYsAWOBj2oyFb5hPCbiG0sJOwq5
pkMZNcA803mluwsJq5UaWE2E1dz3PoorSJp1CRBUVQT0NKdkz0p23ILZ/PcAqi2593sLFCVo04ic
FH0v1L1EX78+TWDf50LlYdqMaX41m7FMTx3/iDkIFvJMoR5Ncg7VDPHmw5w4zIn/avvTIWqUOMny
JGKZVS0VVHoETurZGsMQrQk+W3JE+RW0ydjBBfnHAulF2gollWHMWkSU3QlivsJqM7Tp5qbx+qkf
NgVfFxzR9TF6Y45jcTsg0xgdE4pPopMoTiqvJRnhBJZY0FeicnxB9Y3Qgv/RNdL50Eq4/2umvZdu
T8F6w0hiE52zE9u7q0VMtZteOAgUfzfzcScEqmO02XeF2yQkmhjHgruCO1lxwzlgRV1T9fUUPF2O
7/7R+ovan86wpFBrK2r5waMaCUyRS2tUqm0X4fT3Qlx47nd5hwVF/i7CslpWMIwvL3HXsDkzOcTM
nthpvr4CVeOLJKG/LiklL5mVXFtw/UOo3jPn1WUmTAqYJzMh7LEAz914XfzgNzQdqT8pLAsK7g/S
PcOSSzmNSsBOWBmOxyMh89f8tIth7qfidUfPuR2KXPPZwJKuY304GDqEdlj23xeV/toidnXXEcwT
zPZb+HTGQzuNT5FkwlIj1e3Spl8lPEupT+3hUg4lZ5pn1FzmAfyxw4R0mz3/PT6sEo4g1XDjdoIA
yLgDjEs7jBe0Ys7VI+N5QRBGqyjGpQsmY5I2AnPpLfprjt2PyGMnpCwDP/O5nwAXJtJcBMx5++jA
fRCAWIIcyW0Vb6+x58qu8FW7L4HtaFqof/AVpNPLr7iJnCBttZSlFA2EoSFWanb4fPpwjn57/NK8
3Xfn/Jg0cHRfJeqt29ABNjakWEZQoLbKbvxD0VNqEY0LtsCGcqmHjmelJSDVXQCF0RIn78Bi9/Sp
IWkOUCOjCJ1sqYjJmEkIJpjxF5zqB8BKWBjYYb4FiziYBrPFOGLh1RasIfvfRP2oNwxn45QhCDiE
TZqlkmy529n1zs7YA3LKNAoJJLR3JxSzjp6SR6iJAXcrAYHNxTWxM9OWfKRzJ+ymPvLWCRCJ+Yun
CWbwtYzSCQg+3Ri8aGmKfQ5LmOEnaJX2TygZcwTOPWd8L6qC98TVD+VYc6dnLG8guOqXP+27iwhA
2EXBHYYR7tXCj5iMNyJIHYsHipyCm4g2gxgoOnyFr5GCsCCzimgqeAEbcJpEw9U8AVv2gXpZd1FN
GODRHLogH6Nwa6EBA5j4hBnEFhrqjeXZRr7+Uh8p7cFmOBnHNaiVpuHlVqMi2pKero7t+jFAjJT4
SUOFYi07acAfe0EhRSDIDTibfTzL6+9kOVmReOopefetikr/Ipd61moGAFzoLCpcwLvTu8NQMR1p
Ivi2iDiJvFLCJKm067qWhApIqpWy/kJKkRK4Oc8nD/DzRXJ7zrd7fqRUdFGOWiQO1n20xgUZMCZW
VPE8CyfMUeuGVQUhJfyuNvfhKl4qr1rf5eEK5ERpBa9EXk+2InWMV5mQjVOTC8ykTRcrMhrJOSZK
wKySbIHIS3INlbijth0dvBL6dUIjRGlzUPyjwKxVioam89SXTa/TZr8lvZANK0Aga+1hnV3FTMIN
994NeGh1LSgqlEtgs74qUKXl4Wx4lru/LpXsdjF2nIBCYotjpWPHUgKxfbDCd0+7GEcwC7O+WJNI
Ecb7cnBrXn62QDyh8713O0HHVQev1l3ielCdIxDUmJ/yC61CXAvwsqZlr0sb+4Gka10svuB/UrKG
n42Mu+yoGcMR7+7eYKpHiLeyNsS8RAOVjBCTDmERE8fSTwwU9wbB4lCAJn5mkBkxPetnIX5PwHfG
B2NJFs3A6GoIJtVynrchpgoMjj8QgBwqBbY1uGcYU/0mu6XUZcTXtJyUvbSnePPgDN6NqJaljbXG
GxysA2I6Pa+68LURisQoqrTRSW5NFgqOi//ggvkyulERcW41amM4CM5Qn0dTmZbpQ/VnqFt9TSTo
QGCaa8U1y0cK+8julSvEBi0UpWBmL/L1/FQdNH2GNg7pC2sbkByyLDW44IxCZufoz1eqbbLqpWjw
PQba6Zk/Hg9K0CmOPT49dSNNXdiNVZJAQ1cWJYOhrf/6XhVFHD5u4wk9UTzS06cPcLkkSnHNRY3p
/kiYDcSf7982xmGefDDvW+ZFFNLHkM2G7+6xrzcAlg5HhsInggtkc4f7zrPRcW4FdEVmTg3LtbWP
CXyuqufREPcJEJZV6cAmJMFzdsDSbWQEy4Mh/DK/SrWGTb0NyavQmDtf5HynmqOtXoKcf7xCtQ3a
sJjwv8gtkLbucqnTZShUFF3WYCozqqffRlVgabYORVcZ8CQtYa+Mp8fX7e1Hw4BigZ/XNvdi2t7T
+rS3WLtOOO/uK39QsdpUtQXL3qM8RPLWTCxmeIhXJnr6/OtrTTp3bYlFXX3ER82PjP5GLvblNKpT
kNrLoevGFEk5WcNnO7LQq4NK5FGpzUTj4i/6dnNfKNOx6GfMObPgaduEkmH4oinjGXAteXPQZDLD
P1yoR8Qx2mMvi8V8zE+5F2OeSSJoVMG1/I7T47d6eSTz5mFO0qa7twnHtoZqu3HIvfwBuZx15GjR
zp86NCq9G25TO72g/JgZaal7UB8s8Uw48c8Nv+bM3Fzvgh11KaadyDmbNX5QnkPI4t9QXukSuKOo
fb2MoODy4xzzgMisA7XWm66kI77rpLbB5lL8uWfMsWo4vUn/8zmfqlqdyoRLlYS4w+dj408J43Xt
FO6btE4bXPUcokf2sO53n4ragFHlHQdXEmaBa97IPsPZMOtP/+sbQtmwsetu0a/CEaXRyI7zplUP
kAXyq+FzIU/4aQce+J3I0WC9AS96Lbs7xouF8f8etJ3j0k4gAdugSOITLSTS4PFvNdAMhSGPRoS8
8MCx3xbEYLVVLsNdYmZsqIPEfQwFnPFqXdbbucCYHINQMCcb9BchqxQfY152RrwIfd37/26Rpmx1
datWZMpQVhApdCGg8QFwKX2w1NBONmcJUogzbQopif6VzQIU/zqfvWDlWNkpzihNuoDAP5n0Cr1n
kZbuxymzB4lTqWJyI2qhHXegUdrt58+A/R5dF81LSAeG+vCc3gGHI8abg1y1+MPdDmtYTVsuCe4C
7Ul1ITrQYE8llCzohhfWSEW9LjbAzh0tpq6mtmqjgNKzXmpSVQocXz1j118RXiXy6W5eqNib9tPn
N9VNupEAMhxLdGhx67Bu9tXiJ4ZioxsWGPC5u/CleDp1SDjFxSp0JIWC2VD2aYs97lmtAXv7orcD
3bkwBxw3UDlcJsYyUVoM4XtIsqx/xqDgvuv3+4dU21iWkzc2VDMZvWnO4SznGpXqwuzcGZwvzSry
2iqnjSG8s74vBcPVHuqLxCC6D2gjx4PWauEvtihu30GxKZxq7MrCAAWROWBexMbCjiNwPpNfglkb
MV5Tcrj+UKlkqtTIA1nI8ualan+2aX50JTCNAAWbPu6qA9ui+1AukDYzVkhrcKaHWyRz+73LpBIn
FiPP3JfnwOVjkWpFI/VrUOcGSMBDMZwktdWXxCIinaKp1eVC5g+5+BXBnAnnKW8HKYJZgcOutwrL
GnQbjVBQGTrUGTULo6FXFtoEhXCPloKvKK42j6QekMwOdio0aTH5zsfqr6JmRiUykpJ9Wsq2R0wy
4Qjro5l+Frq+uxY4Q+qupyFOgqC9Z2Clq9JB+pBXWtjkfoCqIEa0lkS7UqQAREf5lQBqgiN0RWTx
HCk4H4hSrgRcTvCgH7BBL5ARVUcPUfxLryw0BRSFxzzUSEgCLf1hwOvdG+CWZfZxwG8FsIEhYzol
8zDuoRdAWMZXsZgzVcGMYw6hsZmEc1n0FumKjAK88sdsj7cYFokRwt5E2ihG+TmilPL8aVM4sUbv
/MR6+hLcPBpQ0I31csBGBNFavqDE07LB76jnWJ/e+u+njgzRFV+kBCgoM/x5rhmTs408TdGcpJ3T
ZFiJyGtEnvVlc8f3U27x7+ivIa/DAF6KVrDVDsBG0yjOhpdMOhC08mAYfQtv9ESibbRVYCDEC1I9
Fyo9399pWwAwmEYKYn/RqF42lOYfUR9kqzHSzTf82hsgWphsjdyIXwTTujH8G1PJC5R/EMd70YRs
/XK3uvfooXMekaQIyIk+T9k8nbmzxzkldsXcDLdCSi0JARv/0oeUos2h7y1trPA2RTXiCC21FE9X
EtmDM5YTlr1nBlkNnJQHX0WcgyND67oxQQGsNo+PzPvKlWUoPPC7oRKaRWiVpaHcbR9g//ddVRMc
ZlsPneD301BQzASOxHtozkJYUEnHGksblsHWeQUl/wQ6Q5s3CpV8Oj/qi2yLzmvyIgdP6wkw+9Y4
PXTzCy9li46CBgjNnYUJdxbWnN8U21W9ynTsfdN1qM5JRgehgCWcZMx4dlnxy/wglUbD/RxP47PC
+4R2O0xyJ46riQ8oftiXSkZLT8uzkr0mkgngNFmai1q5tTF0tbGC2IIFv8rjTKDzDDwLF+pXn4co
R0t7Vr/STzvQlkTvGefCNj/4kBbO2ZcjqeNI1REugISGevtbYLAXwe8QVeMdrN6YqCq6OJ5RGjZ0
DeKtsOyT3k4UYhlbB5NtH9ZrPNC9AgY/dxo9ZNe0MFNYWnAG55ubk8OyDf6cMZd9zhIDx4qxa4Fb
NAEUuMihrotJle0mmfDvPHXkrsu1CB6y99cKoikJXECVTz5l/2j3HCdRWmByCZ1tXQt+7T2A1LiD
gmcXyNYhCj/wUiJKQB7c2dn18H1tAfaLDiYKw+mH2YpQZt4O29OAlezYzXtWTHFSnCpjHkon48Rp
5nmItDYWbhYV8YKz1Nnr4MvEezhLnC06PXoVsb0DksU0HZ6GiTllHL0uvivI8AKmdmb7acpym0l4
pPTymyqdhbjoI9vaLl95o7xQCXAJSeR/zOwnkpSx5v6EFL1XnQhgPFm2c7MFcwoMOi+zfFcr/O9c
CVgAWSzsP9OIty0A9oUraqAbzQQbpNVHoNkuE8+00LS1rbPTATcVNx4r75PZSEkNKIzi6xDqMoZE
l70bEo+RPDVekmS0G+hQsJ6UqHKmxE/mUahqlOCLs9eGSP7H8zI/IRx0qsoSfbl+zPOzWtEGahFn
KyWTp7vhTci91T20EqVXLWAidmOwB22k6SRx0maapa32e18eySBfMzAp06GCbHNvcBFymtbHZciC
hD152DooBd+np2ti9QgWiLsbHIMF3US5YZAUINEcVhO1P8SCVI+4MtoKRg68qvIIsC/jqi+Byt4c
/ZrpjRwE3LumcYUa66c9e4Wg+hyvYc52ekn/GwfyS7an2L75ex0N3Mu3c0zDdO/ZIEK9d+SacyFb
BfXirhOdkjT7u+2LuRYDHrDa9Cxz+5x9bddWmXKgc3ex0wXPXuWuM9d6DUCSjgede5thlhxnH6Ne
EgUrYtCxwhWYScmOP8x1tJ3L6p2E0rA+xJz2auj9Zz/N+b0f5u6bw+UAIGO2S9DqWIcbVeyexhmw
IOehlIc3kJFpA9I2nwys2rBZ7h3HCUxLB4o38WjkclQ9rWwd/ARTkc7FYrcYV4mAYrAtjbHalDL1
eOzduIY0hqEIW2liqpf7iwJdbmXyIuH/xHlsWosOEI3PVcwMVd+Unmx31emSMsvwPAS/W6hqzha6
duC37/379/WCRNRPKYyBNQq6RsAUB6zRGP1ACzYy1WHvosBRp6le4Ucd85NZDc72UywT07cBVCSk
pk8IMc1HYfr1QDBLnUffMp9PTvk0Lp4Z2OEBZow9FzYdiSIlcQTGNEJm+kzW+Zf6/cBbY9GfIhQ3
cp3Z1w5sUCn516IIW7uzmw4ALXSXi6cDOCW/Sc3ag9qeuwyDc7aNEhFz532SW+4+SvB5a5OLpbq7
aV5yqCc1FImls8RY1Lsceg5LMCpU5rZ+mFq1WHOkrySWutclV4OeogIWZuAooNCEUvWP7CKVLxMa
yTL/gQYZlHXd3FmPMYkWzzvHgoij89/BYi+GEAISFoKxZRxrI7+DwJ+j7B0ek2jdzp3PdAkNkMWy
bO65JHZJ2pFvERK6jhz8J2Oj4te57IobJE0ChI3CBrW+DbHMOJkxkDgJ2149kkca4eDWOtGgVo2I
y7Kw1PyXxANVsf1opXGvMiPT02D7cb2Cu6vyxAFqGvtxwUoDc8LSorhKcb7Gat04jMi4mw6hzJRo
RcEn7NpyaHzMsh7dNBSQmGQ2VUU/G+xgZLY202FiUQwZACBQ+j6c/FjDhf4w/ppf1yWBQkAGpkwV
okqWtPouJlJvjuR3NkJHMyi4gu6g1A8Jlwv/XyDj6Ay98Zx5cvVtd3pbRSwKSQMtj8qpSzBp0PMa
qbU1+CmIRtEreJFCNJJGEkcCOkI7ysyCXM8+KWZS0cxzAaLo3RNeSHWxcQzbfcauMxyBdeOsnSZ0
oINhASntebLg/pdIdcnijONivOxlBRMsfuWpA5vuFEbhHAdZi0SwJwzB45xyY3hUrrJfYU2mhqXY
czeWkAKZ4fzox8K+z5e9/4Nxu3QFXMC3qfUZgre9zbbE3W1e5tL4z/mNQz20Nn2jy+gbyCXl/iVV
W2ytqTXRKiAyQs/OV7QVEmZyp63a3go9I3FnMTvm1IxyP7pREiCx7bZ1wIsNsP2i3qBtuo34N8XM
r3q+ADKh6v+qVAU/wdy+UJne01TP1sucxFR71f0ZMoqt6CBWtVkMLq0ScPZZ+FOpaVtYXwPr0eha
YNbXb0h3DX8Tv4HKxpofvOgn88b7ZO6djd2Or/Jpk3rkObQL58nn/mlQP0FyVAARnqleaaPPoimY
sneez3CFMae41XEmOtEw5xIictbueVK6L5ogaGGhTMWknTsTVBO1StVvIkcuYKcLjGY5IQGsoYds
54WDxr2qpA0UbrPS0ekbBBA5/G/Pitu9f9rC/nQD8SWcfLXUH8ykvFyyKUORngJ9RAe5xcp6y2Qt
5AvC7tBu2AvPS8aRu/lgwKM+u85N9jjDqayd9S0CXRLCrfyFt+thgk4ams89iPDvY9NZSi/GSSgm
f15tkZpev7CjFCSSTkvijRebocev22PojAmY0An+sRa2V05KYJPKdxuYJqBXRuf4n9KAL4U3VzAV
pghIrZvdfFxtz23GZTbQM3IvWWcR5VgCeBs3nDHfKJFw3n6iEIk5elz0ReFvQa57W8a4s9gvgupk
ZqUbjP68G/DZ7lpHhIEDFhmMHNZF2TZ7HML8w2fHgyalj5u9kzyWmsk6NL7iQ8M24u36SbkXyU3q
Z/a0e1tzFHIUmHYLzGboiu70q2unevO3NXQD6WaH9s/lmG7/Xgd0tQELDnIdfBD38Q+n8R4ZDd1R
YrnDh8tREXDBJVcJkvSk3U8/KexamYbtE7EEDjPEFPxEKZTQHCGd6ejs9fh2HA/3kLSJRneiftaU
/KwAuf2OkxuFYv2evlWelG+fmkbfS/CUf2zRolficEbvjspcfQZa5WGyDgpb3BYwLzrM1PyHZssc
aHWrTTdOxDexsqUcu3P8UP0xgivPCgGhfQiJSXXVwNqozj2WbM1lx8eHiFUeM+tQdXfrCl2adtcI
1dxqgHK7yICYG8jbw04XbmlQXgEqWP6uBm0E41xeJL2bHZgfYpJrdPGUWzGFjj/IEsHME1Culv6B
LIRzCDZDalWh8t/scoCWmmshXlcFr405GYvoZLjvKBBNooKB780n5D1P4xunJhGwGq3UD6qZ/Asi
/5NzQdi/ibbWjsYRyhrsfQf35PA75gsAd5wj5obRj0qXC/Yl8QBMvx2ux4QbgWkekldE4CH6JQ8q
s7E6NqJ0HazhQYbFuIGe4fctx09QWzox+3LwFTaelV3Qhc60H2hdrWEsN2zSaH/OreRE88jiULTH
xVfYB3y8JjJbZhBmc1k61ZyTLLcOwEkW5apqE8eV4ZpT2CqWfE7ExdgRq8JXJ91/hKDGChpSjSVy
pvrOyA/C2OH+4RB25kG7IW7hW1tjC6SWUchrUQfU7FjPwSh2aGg8I/2as2HwnWzat+9R/Md+XZ5o
jpO7pqIUl6DY3yaAvONpOOr5xFMy/G9iAEl4puh3Ro3gh8Ix/6fn1RSWPsPibwiMdWFhvjw1RdrI
nLT0vgMXo8CBTHjzQMNzsMum/pQnCRD7DtZvIgKIv33XuupVnENH/6kJMcrQ/AtUNobHWNP2xFCl
m9PbQ8TaZ5KyGIQHAc//L3lZGvEthvWDbvqjQV3WMnizuvnRa5GRHA8S7sqZq9wxIBxjtxclE3B/
SYoE/A4BYlYzyma9clED55BXLfEfAoLPxst2hqmDAkQSUXm1OfHkt7Cw/ztKsmaFgT2wDHARLYDw
cw0DSH321DSa3oHHbCHaDixr4ZZBpsbuDL9HIoxD5ygznslssXwL5LvaxLH0bhyysObEJKCOCXLX
51uIgTXtmahPaf5NbAnDJhC0Z5IBsvm7qtw3RBYClaprBrcwnJbmtY9BpxqphiPCPVXD1+BDtx5O
eDzLhYDgkvifa2VOlbD+ZuGVM9FuIp6SMrWVvn8EpsIfjKbzArafofTZb+1LlVkcS82LjbKbcqHz
nxL+LrZiyyr2XltjkVcCiLg1hJTYngsw+/WJ0hEJ7eP/CX2KhZSnODLTlJISs7oTiPWTcRq3YJel
H4SiMbZq5zZwHS7/BW2q8obSuICwLhwLAY4uUD+oM43/78nC4cXeiak4FqncNRiDSReOt8i94Fe1
tc/SnItJ9+w8ES4qC7ygzo5bclzRuO87zTXaXJ1s4ZbtqHMimp4nFDpSIvcZw0qYjTplrraNAt2L
DppNc5+Y4Gq7GcDRxVOsSp/V/hqMNcxjSgnB/tz/nfWO5iJznz2GCkkRIl4FXE6BNKunHF6S5QBc
r/CjLA/4KsRwr86K14D18ZSXFldJ4JG0lXtR550iGNY9riXJtoarQflV/eH/QYNVgphQOjUPDlrG
1W13f2YnjqVS9MkQ7SR16w5d+4prjrFCX0HGqg4eGV4pHjYneNCQ8t85KPVZ/7xZsBhkwIMJuv7i
GSsHND20IecgDz0MS4h++/W+183tkEZZqpXoN/mD/dBW4J/w7gp+LyL+umd7DbLhGIInPXiL9FYX
Ok5MFVAQGRe7auDIdJEIKpvc/adJPlNeWc7sYsPGyyXjo2hFvkj5Fds5elqJyPxOyN+Ny1NVoNhb
cjfeTJZIqTyccJySJkWaoIw7cS0lLq8IRCAR96/sxSoHpn/JK690s/ZI/NF824OMfKx+a4Kaa5L5
nfcxo+vvllYRpusejlgcMGUJr/9q2rd5qK3oeVYbrVLSQckX2/j763FCqi3Duvafi7uG09ZXK7GT
HF1ZcQZr5vtChrEMPXhNn9Cau5IYc6DSlUmeKHzuP3jlxY9rljFP44x19y947fH8OXd+7uldHJTq
cBEqlyjpqIKloX+leogjt9rSeoMLhx2p8UCNvk6AJ/MF4MZMBBI70sz+ZWy/mHj8jT2704P/U+cW
+qc+pyr2U+BD8M1wO669pWYcxn7r7bwtDJdlIij0d6S6kc48I24uAMLdJEUgM28a0FJidH1zuI8/
069GzA3MsngvRKsXk3JRSqD0S2GjMArMvi3usfVjAv4m3u5zLs8rRJGVShYI3TXjgLc9vc42z1zM
+PuM4UqlIXr89Jy05lHESwtTGymsxq+K8mDQQq2d64+Hy6LBejdfGzjOTJv1pSBY/CmcM1DRyrAb
44VAIb6rvu9QPwLFg9xfHBv4k43I1ZBkJsgyy0cId1jgQJp7DnGDgHmOv4Fag+jLuKgRiutGToHG
MxSQk1uyID1bNHIKTeDdDlVxeLCho7q0D9nbYiAtYoC9FyR9tQAQA73+b0P3Nax7vgNbtR7dQ2hM
AzhkayELAWaUpOK0Pwa1e8UPMVFMWcQJqKd+dxZXMEQC7SGcbSNTdCx/rrtlm5BIoXkLbgTJAS4G
ksSrmZcwTVYr1lOHvHUBI/HRml3EYZs//n8m02UcMf4rY0E1ueF+PaZVCDUBlGWYIAV7HthswpDl
cPiA6GcizuZvR2/UM1rf0c80v4gONa5HX9ptpzk8siQ63Qi19UkBQWSpOvN5rE9qlui+Sz05Qjzh
ELfgUGb66rCfCsTYBB+7OmPcJozw/X7pwnZHjOpF0F4j01nb1JjmhGZByxs/zAhnueYDt7An9UmD
SF+gj4N03CmcGVagf3xFljeFF8TkENnAN6+t5MmsXtmVPW6jbGlBpxcx9e87HMrtnndjgxi6OjPG
Ohh0Sdlqr22ky939Rap8wo8TVFpIDeLcbjIMslM303JV7b5aTArLcJfWFTs0zicg/oMx5NgUb1oX
X8AMGrt5FwXti3IS8Mey22oawWzl4bOfYL1hJJWrlhUOPPe7d+eIXQZNPquxuMIxq9vqmtqqAaLq
sLzkOCbdl6VO4db0zvT3KgeYzefRahxyuMe97wNVjIyHfejW5o4HYjmMmTAgZp1AMZVkNTXwA2xo
l7n2C4myzWA0S1T8u5fvMIbSlGyX8wwsquvmRmOsmLVAGGO2D0TtV3+YQdgwQSaFiW5C2VvMtV6L
s1Q5qgOzv7wELN9T2lyDcp+5E9vJzBwRLZZaQELzO+71G25+s/BnEpkNhakKhIXsqhTiQA0Td94o
rbJotGlOE/4P89f3NtR8sgSEuRatqpM1sbvXw4JvUFNdPxic9WjmhwWWJLyWYwW4/YW6xCRvscn4
9MpvbVhS+65ZeYy4EcgqjcDd+rDDJ8dI6OczGOzo+COqTmP+t4t+oa8Uu331K+iKOKk/3/X+oVxx
W5dYTNEa1NW7ObgOVvbfO8KivQT4sTSnLNoT78AsOEnjySDSG60/Bq4NSRpGIK1wDzONceD1++03
af76mQey9WXUrZ76ZZEnWD5cVulLEYdaw0V1aVYAyfRE7mAKc7QWutLiBLp4uTPOU0fthG7YFTJ9
HdCZYorVRWa8zisySDW9vZdt1gIMFkCGOVgVHmSBiVavmktRERrUV4fAYHj/2JsT4OvdDZoNanIF
rHiXIih9eRj5Ae4w2O6FOZ98oId2OFaKqJuBWbntsbCSJe51MeKQg47NTflh4Ua+ojmVk0rhyNn0
Due+piIWyFPLGcCDxjTQOyhw9E7ugjJ2tNfpOS4Ey0T4TkAD0e67TWbjeA2aN8jPV9hDCzQpQYQw
o3u/WvLSe5oD7dXpIUsXec5OBMs/YFLQ59vI0mQEqAd5zDY9GGaZkc2dDZr9xSHNHXy1fjPxgn4w
ry8uTi+2++9PD+F8N717PrWct9xF8EBfnqWe5RQ3Yr4SQMQU5ZEerq6j2IfgC7CVXFbW6iq/fnWz
ZIARRhJRkbA9h/U35O++qMITwxrkeMcJpw1sOUChFQ60yUO+0fxlJR9xsoxZi4L2+q6B7gvVP+hJ
swZr7Y8aQ+nOZu/TxQZryTep0Dt9AqF9WOXX+wck+J3UZEbJEpDQSANtk4arshbRMyQ+YWe3H0Fi
Acrw1LsLw5AgXlX1DlklE1/iAGBS85SrUlsWKgA8SxesH2ifoWkVvNar/Ewp2XqrL82EdFU8ufxU
NxBpWYzcJZgN0ZMr0UX/IOnJPXvaKOPpQAa9yKfTRMkRns1sq0y9XefhH6FsJw6QVYFzazN9ABU0
rS1IYJev+OQbI0OJPdXWAXo+lvrvjg/bqzcfRkLwBgKyT/pvLsTGbdSfPdodnTWyAymkLhEPG9rV
MDjJ4JHr6A1cQLkGX/KsrnCMM7yVlYvWvx/x+FwGnz3VkDXjPR+4mbLYdlpkLdCGhZz1ndrHMgov
KAXp7S0HyS4QNiXVIuf7xG/bCty4D8ED8fg2Wrv2HwwziCbG8d7Pe4nAy83c4A2PIV+9w+UwV8Ui
7kpmrP95fWPjsAPTeLsKBK+L2nA/W4zqgjr0SS/iZyzsuo9vngrnoe0+IlHNRKkad4WDAIoFcOJJ
otfazqqjD4ntaFA4MDP4K0DW7oL6tQIeQr3Ri3B+aATTyGKUKJLM5dqka33xdujytq+GpL2LBccp
j9yzdtRgy3+iPcOEVjyjIqDIrX7nIOdwgGszMoMOlpmIW07i3yc0KH2lqaXzVeuXCP/NTDP5NDO0
S4az/cQ72jxvtvqjEOuqvVCN84RsPOPX9bt9k8yeWqtLWTGxnCpQgaYRcDXJmlEhDio4asFtZmh4
Pi9O7FuEUvrg8TxGiwNIX6Hyd0CIZOPf6SQfzL6eT3/Sxa+pRlt04jQOYZDSq6tne2m76JbeQVt/
+8NJsDpmid1w4KtmvuAdIujBXoCg2uUQUbY2/ZGMaa3kSScu4iHg5bp59V35EDEH+QO2DRQxWLgN
uN9SbThJQ0pqVD1WqQrdAPu0rrvGl/fYnueV9EBe1aR1nsxH6lAbSE7/bHBxmHnHylau4qmvtY1b
wYym6zkUC/8bnpkN3OCBWgflTrOHGDBuahvXts6xYVazvM32dxETB5A5uymBFFgCplT8cxjPQ9p8
1BmkVzIa0AZN9kMzxCd+qGwn0Rdm1ssYrc+MOCIqCA3dxKhDOWeBidFJl4kIR+c51euHBOhGzugJ
YXA6BOOJbDJqYA3a0utus5VDitR6aWfURhTOFcgcoVVALgZ87RP1NuNz3b8jIwSZuIz74R+47Dk7
cihRdefD8KawkuWXKld6cnMN615wYJTQQ+0fhcA1ZB76RJMen440L0XdpMPaD9UveFjooQG7cMoQ
CIE9gLQIIoLAyUZ212MIZ1cnKquk7lx4TiUMCVAYKioYsWa8DPkTJ3YEh6TbIFCAkkDI0bmzopFh
oqwVCTX4AyQ0Gq8FmX6kYFHa7C0OWsGLnEo+XZlu5eoaHTnRACIf5+cTRd1yx1s9MQ1uvJJDVWDx
j+MVVP7FJvzlI2znOVXH/6O+OB8HGa0v1HK/TQz8XZI/4pCXIG+l7miovCkfpAUfFbybZHT/um3g
2uehEWUwnc8iRebwmII0Xp3DWLz7OXlBkTHuZXkmRhQbiZOK+W5qnT14arGagS68T1jD7LvqhCF/
qrlbkF1/LIKCFbwzTHU40ujRGNnWvMHuTaMfOot+b5Ib9Z6rNRzkomWuQA0l6LdfuTNiXXIYK8yr
BGyamOs0U1O1XNC5yKmXjNQlsZpokM4vNQeUlsUkbCfPNxPOl/5gQmHysRa7Ie/iPZjcWK/eaEJI
N9GQbivojIleHMo1CR4q+z9vV1XHqGze9OFkOaRWltRc9EqnhS2lmB/zQZvwUpstRpmaxGUH1cxr
r4vTO/qFi2jnibHSYx9H7a4wOqptTkLOfP18pjiasMn+XDLyIJw6tPGuPFpRwYwS0/ywbqVLQmPU
74fknIv9MHGk7ZHY3m23M/pokxF0dCK6WB6QpKTYYJEsOewdyPI1mzFrYvkxz+iYyrfifzTw+cAm
R/Oc4+u4ZKygGFqbXdslVGDDjNuxonwkflSeF6q4xXZMFuwdMV93PTv1RdmO37BYuCesb0J8UCj8
b782P2caksQVvWhy+4LKH7Nz5RcXVFnQcv9iSUD9vBpiC7TzFZj16BYBL7v24UPcjjnzbDAd3ify
SO53lhoho24ZNeNeJCwBF0VMbnWmq7wBjlHHIMRvy9LfKUpHlw0YB1R3oMGj/Lgq4spAX/Jdv+ud
anjUXNiuPxVuAAIR9Uk+oDIA0tAKPaNAMCdmbw8oKYBN6HSN8zTcnZsmGuDIymF3VAqK9Edlb9av
flQnL6Q/9g4RAS6O8mkuh9Z2qKzoGjA8U9AlcVGl+f2gkcchyefF7dk449SNEY8sTMF4x91vOIKr
Ny7LTDXtI4DcRBCVDMiY9+3KV5SNd8wA/NpuPHjME++20Vsmmap3LKqFhlUlHSwET43W2+fvUSrO
BLQSycllNa+PGQq6Er5tbIxuVkPNsuIYjaWbxXicEFD3b7aI6Rw3xUtskm0F1L++SBpezD8kVHfp
mty9u0Cy1nSyOLM9Q4/gyfZJJ0hKVHawXlPQGmNmSxYrcmX7Ci3lv4eH4U8sqQI2vp4/yzmHYtXe
sfPaA0JDTSAMO4sBqJfXLLG5D4l/SdOTeT98He74kwS98aSfpkhfPoVFO3zGRSrVmWU31SRxQQp4
TmCwIsPf3B4EnwcmZhkD7RbKsY9IeeazwSBMySHR324mfah/vFYEZIv46WSwxOpLf4/D5O+ZDznX
mdf1hGFbuKnUbPpjvMWh9/PxObpTzdAb2CPsaqGUqjkMH1R4f1xpzPWUutFj52jKTDWeG46c38KH
vRf0Djgul5YWtBj2nrkGW1X/2q/yOnfO7L6G70cPS1oDn5qaSFerX24vGM2NtM8M97h3tfFSKTel
pbFL5oG3p5cYShg1EmJMEa99VJyKhng4glJbZmU77T6HUITBd4VmD2beQ0TU/VnG8a+td6+rfzZj
R3I5zL/d2hHKxDFW+w3gA0VwRm27ztkeEvsrWqP9RjCHr4U4lGomq+GjgohmVmhjdqByO9hL7Yd7
CfOAREeB6ceGhAfcuOGLp81krgs2nHp/JhfV4AQM8mK4iVuyL+8lnwxKtDGwZYm0tjQYWloEmUG5
3Bc8oNHfFTkQBJeJ2gkcByZyblCV9m/53VBXTEXmWet4YSlNZyTQ3l/1riHhP/XAFafrEOmVXXVF
OO+YojuW5DMEcnHKDzu1JWAeSs1OJPjDgI9qmFnhIGHKH67igR3EBZQmE1GTmzJpWBIaEx/7cNp6
lVfWjmI8uAL5uUQOdmCWyCS8UNMBlRpfay4wfrIKdKFSicKVNnJQb67Tu9x3EndoUdUNfIxJWGZO
xTIOT7RvLogrcg1L876HxyhkJyzY38y+ye6tOk+M4dbMJOhJ+dAUfxC+LJrQE8ok7NAJX0u+VvSr
iuI0oKfW3UejTWEFmK3J8EcXIQEUnZweXN/5r8ypsa6vrb82X50PQJOq8XCxJ09o7vayPKFsLn3G
U3DLZUPOcoqtCKHQfxSIoWgD9G1iCpRQHRTFpV1eTzZgnDSiMZH2ljk42HBSaTRJuzYYj39epqm8
J+lZDFWnyAhxEce7PtwHo2E2f5DzugbulOURcj0q1LxqVqMYRvPQSc1wow8EVsWviCctyThRLpj4
EW4EgNZLPiMxGfWFitmICGav3meBduWZf7Q208zxM3bHfDmmIu3b/DXaavQs+UyX8CyDS4TIGHWW
e9ZVH4cQCr9NOqs9ZHjel/BfGsMJl25i44amqod1SdSZUNrK7+ndRYuw1gQLlwrjWhf8dal/+4iy
7k06EUNS5CEA9IhQdyA5hakHrEn37PEC+hNNZmymyVHjmoMIoDsRW0gvijJBTDxN2T/Dxc0J7jOS
7uTgQumhnXpVyOMGGqvK5NGXyd+ioEgUsBaR4DsVH0stEHjigzpBeg+9tzxS3uuyXiIfcp02qxR1
J+DzQgb9GHzM4Z7stIXR1woABRrc+Q/sWrvkjc1EtWHdXmwCIvj2Xn1U+sG/JwxtA/TObs41S28x
XvnUZQVyQXIPfYaD4uqAHihTC/W+hkhkBKu54UjmdMjrjOL9lYJ1KF/oAbU1G8s0SkaFLMtZfm88
JvYorcfFXByVSzODeXMs0a6M/VkCd1E1Zkcyou8WrA/S0wT/xaDwqQxsG4U7S99YKm1DV3vXgyHR
g4sUBTO8jxhfYDXHvSZtyz3ra0zWfSA59LXRu9ey1ZzN6Sg/ZnrqV64ZW5Z88fTybZjxAONxW3S6
jlvSw5n2MXeP5R7pGJwL07RWE9Ym8WfQ3FE37ftsvpbtsIix+Mhb3PH3fQPXgGZzhfTK2EL4nqVQ
M60hfLlKk3YPsV2FVDCIQ2USytlIdG7Ir+aNtLIudZEmX0GyTMLD6vJ5f4ZsgM9jDE6IOShtctz1
Crbt/RU9TNi6wjwGXw4GYIqdPZb9QdLF64zq0RqL6C7yww53qlNuZXwWRVjWs3dOmQXrMYosLjN/
4o5MuAkg+m+17iNCI7+14IhaHhlsrruEc3fpbUc6hVh74zMw4RROm8nFwJH/riF/SfpBOJd4Lsn1
lvfimuklbASuhTYhaKV9lGoVVnpSr2q/2D7xDRHWqgncQOdJWtD/pDsxmWnvx4QhrO4l9WNOuCPT
1kMYFojo1sGH2A8Fm4CMwM/5ouq3m9YKhVETfQPu0wnyHtAdwc/wGjfbvEMFnUmv04NMK+ROCkkh
Atji40mXJuhIG824xOZu3N+UeFYgPI0xNx8kPOqD3n2QJcMp9AFUn91vtxH3Fbl7zMMg/5vIhwJ1
bx+9KziMtI0wgCdmHsixSmst1iX8xbdgn9uo9/ijutN/92PDTMA4YJBOu/fJ6bmKBDWBEo5nJSdU
sESQ9YrfjF/fR+MLovOF0ps26W9ilfyeLohecg45dVWz9TS8d/EoSMQpV8oOucX+f3fKs8u/NuZn
z4RqSOw29H+k0YbYtd6ZNKgshmVo31fwVfh5AyBemSm++P4F3VVB00N1KpfIYCvTL6UhKDdY28CV
CeIJECWqGn8SM4tPbcE02cRiitwHut2sJg7toLfNGvdChrnJjBvjZOlIQuZEEAhheSgHxn5L1jMM
iOkWP7KNj1HtDSejRqK5fny5jvXUtvMWucTqFa6gvlRK+eiSIA56gVEA7mLbTjNfc9obgM1VxtbF
bWW9j6HY4HMK6FNkBX2kcRVTYxEQOJrUAXAtf1Z+fXOFrPx1B7qUtakLrpTytmX6LF7l4KOntB82
kOSFCHc67NkTieYZ5fyEpqUcckyDyo9ABT6CR+oqTI7OL4RmlvAEVflZuBA4RiAZIQfiKSf/7x/o
UdR6oNZ0aM4jcdU/QaS4FDz/ykn2QBNYXfSe3PHdSuUOwVtVimcbixDR30ru4SQuaNzXR4ecWDuG
YQAmFzdEFFDaZEn670es0ILXqDD613rRwWAf5xaU9O7HDo2n81tNYOlxUfpTO40OZ6CNlHxKkLFP
VE6Fhp+thXbm0aIouiOludXlsO5LhFtuBbh2vzFP+XlixGvOjRCGQ6BS6RAR9fe7dZe+9ZZRverB
tR+wO8gJya/X88FUkysDGfFPe5hlbuZLDi6wRxf3LT0RG+Q59f3CMIl1kkDtoJGWxYox1N+tEMTQ
J/p6VdPMwgOfnyObxdn4xHfmVl8MC6PQwGZasXBtJUAOASfOUAwHXy2o7Z+bX6kEpwdj/16uxs1R
VTYzUE46iJSdrcsFYnJFOFnoARdQqkXNnETA9JVUilmpebw53G38v00jFozGxXQHWWJ5rhjiYvRn
mxAIuBhEqQgdgCRi637vhqABC1sBRk24JejI4trF3DF3qSwrHCPVen3q5o/3AB6hN4zsVj0paTFW
V9p7/A4oYDYfLGp+VZ5MmNOr/9kvmQTg2UFn6EpeSyMd9iEXK58n76WjnwpUAoqZCC7qBQRpABas
PpLmeFXWWjHTErp8WavzciwJAvn+B7gPuRjRZepT2RVyVFRy91kDBDyz0dgXAxqhd6iGdT1TE5xj
88mBbiQGP+JIHb3Jz8Dz45wmA/mh/ifvp9bP8ivHVTy8/xNhrYvE1p3gu20fWOEsd/HHguHz2UZF
WCXPcY88Cnzhwgm3lqr3QEuo0F+A++iir/GsfZ9p9MpbZcerQFSdBuVxaCxTrtSkuTBwIWo320U7
Sds2/hcDLsJSditnw1XhN+fqBexk2gHSTzBalP0Zmfn592ltMGak6Tf2nYknpradcfa1ZMtBU2C+
t8NJAL6QaDtLjeVpouOyIuBOlNi5+k/3xOT40kB2QzzRrM54TmchHbtFepj7Nu0macC2JcK04eFK
m7qhm3Y/WSJF15+rdriusCbXWoZYcwe4P70yPL4Y6CclbsDH6+gmnZDKkNOQ1zNoWkdNcMB8AOwU
yKjVTHkTGPIZCJuQXwCg7ptCE3UggjysFm3e/JL5n4PBPwj/qwFyzWGKBI82Klwpnpjw9oDqqkTB
H8hD1VaQEaODy7WI5Ooqu5FmkVAcRpxWlc1eAxwcoQ7Zb8LrwuAGRN2HpTamfjggJj29EIbLF8PA
t4yF5S5otS64rCEBUJXc0JqjDtv/umnEkPpfS5Gm7eG5eno/K/C1iQP/UKH9Tfrrb9+bPs7BPpWs
iimufoeM9EoYUO5b9mIMFNap7O1jmr7zTwxSuLnGDnvoZqIb/Aq7nmE+ZlmiTTKgWZNDDkJPHFXt
Got0pGba8ob5bJ0IiihDvHmFGpWZW6YEdkS4+Ho5A+EwQWdPVKUsBeeCdW52C3e8my+SfpBTJax3
INlk5+Jb3Vvc/YMePMpDINJtZY+S7w/3I0a2OnjWYPP1qqGOgemHUQyD7OxoH085hjgcAzOLuwi+
B08GLg2lhgN4f469CWQbLy67K8i7QSp2CqfthnzXSaNdOnFJV2QjqCEt4jb/NUl1+rxgCfJ3y838
jZtkTPYDNGShhDMT5Q8CdwuWgMhFtkf5hzkRy2k+vJm0jUwXoO6CvOWrJA43Go/0b9vV5t5H179W
HI7ZfDQOtNwWbykKGp79PmHXrszANnqOXIqBMwJoMAHrHso6dbmxpQv/KD4vBH73ZFH0/YEk1lFl
aMs611a83BSm8WitJOpXgfz0AF5GWB+ylJGcR2O3r3TFs3GlwzDgd2VRNdcu9unljHoeI8UifHHE
RokjA7mx8m0SNU8MascPbs30QreqLihWz+1y3kAKsALGjDk9plZLxEeHDHAW/drZcjau0/Sik/wd
u0KcuQHDYMpdegS+yk5gGD9QYqeOM96JOFDYQCl9ZlK1uLGty/ZFPtjpgPJgjtc8STXSVWOATaxt
s4gbeejJLFOOm47oO3o39Kq2t54Nx7hi/SUGnZRrG0LRCzi2K/nbBQma80sywTWJmsmhgp2CUZr8
4RkKRapgDjdKvxtJ6C6GhNTiyTm2XkPsPE+/E5kLygH9JpUlyn9aSWe7EH+ABpQ8MUsv/CLvyVET
DsaviBCIkIAvrtIonXPVkXxCDWhbpXlwvbQ40I38s/F1WYHKNfWENK6e1BoVoziKFAGKE2O17HAb
veQyhWksTa+72u04YVS3XNVISSl2tP2kqHfSCugFKIXlUvMUJihisknTr5pUgXcIezCoOGUC3i8g
4mpvmqWUJ7rcezVT1UdEE0oWDwVXw5q7r9iQRnKm/JVma68Fx4C1vQu1bO6He+CB9h14r4AFRc4N
paI2+dNWhRUwa5r4HWsXNpW5rtr91le9WGfvTkqW4cjSQatJa0tkA3y3vhdKPV6ofjBPzT9R+CnP
L3/5HzNjKoyVgzMzscjm0IZJ1HvzehmZA7kP3ffO51JUA59kQUTf677ThHu+ZU6prqrbBmZaeQKP
t5JuNEqeJDDZbUWiiQTjGH+aDklbaPpK7Rm9a/Jn2m7zq8BGczCcrYH/WzNnq2xEsyXa+nWrCmn3
gt7B5xk8HOr2E/il8jyCvpQNRDeqhSz47jYpZW1spuyBAWYAsSg9rv5E1tMI6BPDmZCJoJ0UXcg/
M1t2yLtsWpvDy6m7xUGZRJNLd7fWHMOXRyaP1hzTokvgMirk0ORcEP4boR0885jbYMekzX5gLCW9
F3xn92G/zZLCcgIYDUTWMerXHW+yUno8ln+0Fa7FRPRgmwry0zesytdyFXUtu72k+JYtk/NEtRJD
DMuSsYZ1AVFM4UgzowccLH61cV4/sBuJHa+eMVAKDpHg7xA8724XI9CTooajK4vnbB6PMj2urNRr
snOFaJ/qIupl5fJnoguEkbTqjSVKRa9hLIwnbpNiU15B1peusisNi2SAwcd2+eP8vLuBMJse1AUK
W69zIJ/uZ7mo2kFxg0Z+TDJM0s5re4OqdgJ8fQF/5G1rbeeB1EOYWK63S68h2D2lgiBkehyDS1ym
UJm5FdokwYrO075XklmErfV978AzSk9S5HbFSgFfQHgVDthot2tKOKjNdef0AT9uIDTAmNGfUlSw
EeWgbYSq39ehf90B1UZC03GJXRI3uC+aCO9n8lIxzZVBAO2mDIzsBNhtcUAIx4M/XKTtfS4HMfgQ
5TS76Wmgyo91TMVqbaX2nKZ8930W8QVRwjcuTZ3OOQUU34FMwVXcInTg4ndIdl4s06b0jRtG3P8O
iRx/uXb0AW69b+Jq7bJHTgMp7h/ldw/sK7Ugl2VH+9dYpJ9j8pvZuU85akFp2pagXiv6119ULeAu
8eiKGDZTsxpJZLCAuhrPTzfByRn/ZPy80ixmGph5Eea+oRy5o3n37yuzzyS7v98bFcuzXojNkSPE
BQ6JolDeVyAPJV6MGoLV9+gJeTA9fw10D2sf6ogBd4O/ER/s+AY7D17DFyc7hyN9Ds4K9EU7aqRF
MdBC4OfVdRkFM/MU5YWUTXoKaiiRLSALm6k/zOfeILTvHYy57bgJqI0Na3e8mgKhcR1Ado35deKb
BJ24dWdHZhJ6gQfTyiTWtgoE2G5Zi/r1PxgnIqfx8i8HBxH0P0NsvlnyUbBRnME1uy8zfxbfO4/5
Ll+IhusD80qWmkFNni5URTO/8nPdLS5DXNzRf9URyI84Vst4CenUwRczK0vW7ik4242GNesIIiVW
j+oeR5DNuGpLNBzNMYW4YDTbjSjgjqwhwKOxhsVthJ7gAANSFub9D9EvV+5WRD5uHHgE6BLY3ovv
NviWdQCSFCsqesWoGvMBidPQxZRSgJEfWpZu6WkxjlRwkzPSFfdTyR7rnp2KDp9irTrEinvhlbzZ
9SpxPNrUAvuLeowmr38gl3gAMl9u+h17m+dcAVbrOmNbgV4JS3n8vCQZj8q3Z818XxhNXbiSd/M/
q3UCCzpGPRwv4ngimOTA0wvBeymdPVqQpY00otN4ohMIFuBiRDzSP1NzT2NUVahjXQHaBxcv8Qxy
ZVr4qb5fhnxyuRvTFKESIXjekhvTcRSoyDsi1K7umTbMlxE2d2BlEqqQUvRplW/wpa2z93AH5iOp
yqeR1m2gzv9wj0/At15Rd49TuyAzRJBLelnM0TRZ8inpqgH8LWCHlPCHMP8T+xD6fQWfVQjeSH6c
uML+pCzHOJwc78JIPwHQo/6Nc3Fdccj2lV6b+e3bfEh/tswgPqp2XhvDKcyvxBp71xG0V+JqJJBe
YWHpjj/aw4YeTQYV3olF5bsn1yEj2m6Ll0Cabx5to+mgHKI+kL8VuZf2swO0lfj64Zp66nJ/APmg
AqUMRgjtsic0F3iPzixriIzEMOgF9ZyLh7AKGX4Ve/zbGfE3etaRSLbTZ1mtyg2ZDNpY6er/0faM
eCY9asKqMHCfgWi3ZkpT0F3dvJitb8n+1WKtFGLHjkS7LMySOqPHXercugyAd0lN/Ou5ZHv0/GR0
cvEfwrhcZsEXGTGYAgw9UNiBHXMerQeDezYwbjanylaLF8f+BAIcHqrYa0A0paATV/002MmTvQQb
p5neFdZGF1gvc03/Yz36Hh5dcDBhlaGBzdlk2PsDa45r0GHoAY6bfu0n90T0RstQ5U7mAQJgYjB6
w/I/MqzWfkSAaa8CSC6n+xi7M2k6baLi2UAaC08vlzOuod2n4BtbPpWkoDv+Pt2q2i6wdR+fumeM
yyYccWLc7t07Rl8UmBzhAYHGJ1P6fopT75zI4oVhBzKdgHxXi7ttF9AXtxdGIGzs8s3FrARQ0W6K
i9HO4Kw3Kh09gwXHE7gAY9D2GC8XLGS0y2IzbCe6CpJwsNAyum8pJ3TOaf0Sz72TGd1PIeOgXVFa
cYBC12mQvFesuO27WxmQFV9hQ3TdO/37gH3qmrPyPBgQytTs6nT/mO/WrkjzAcxzQtoNadtAPW+F
HxqsTPyH3cZLzJsPonI+AEMjM/W7T9aWyuLMARIAGnLS6hA4OCqVgJdIyZRdvxnRmDjpV0RfFVy7
jjDw3sfX63kIbBg7yUVqvhb2ounCAS/D3D8U/Cc9+Lz/rpVaS/R9BbomKPycQ+NaGdkjWGNOuyOg
BXHvJChrcEyuHF0wxh61i1NQR7iGdBYWaKuDYJI5gmDStJab0m0l0ZvHK9tXXkIMusu4SJ36bqgr
sHDpbGqrWZ8O4nbxBlwgfCkrjOZ0Ymu5M577qdPRPG3gmL17bMo9mMzFnS26zye1gPOiz/omixM1
65xsl5fAZz/m/c1t80bIC0NBshH4c5qrJhmBBo0Q4b2NzCzoX+bFYKuQisi0e2c+rSi//3+0mFaO
qrn19opjQrlRXctbPFgfA1L9jZ2SO7nN6eU9ykP7/Fg9RF2p3uWlIGXCtrGNQENDEBJrda2gbQrc
hZznOcI9Cn0gAgGSmPqet4GpR5ExJ3ChChKDiskEQZN0zTZVT2Vikb0fXaUsA0uEETRLshFJsizm
WGk4qBaZZ80qd0CiFDbSQZLpXL/i9t7/j4CQ8DB3ArAbrcKhJE/tDnrKxflyBSLDDeQo5XzgFQpS
Ud2bMpDDdnKUnXHoPmhNkx+fR+29PgVc2e6jGqZE8YfJB27G7BwBpC3efnbWRLWxYv5JIIn9TMxX
ZyuIbI0WooOWwzDutcp9nyecnUoOf6he5gVDIDKY+lXZhE1wZnPqozvUgj8prr0X+McmQf4VnoyR
Os+3BnI9cNy9N0C1T6wKSDZhD25nYroZdT5OEecqRpVfn6qsxf7UI26/87AZs8Cj53lvQMwekRwO
LNc3j95pCYorbt8Yd+p0VX2TATbj1xf/7raMN5/rFKMRiYPEsAvjSL5UwzQPOBV03r54o3aKSr8R
uHb0RmmtxtZlP3qT+qs1IQWfKEwC3mOlnRbOKPgM5Z9k0OR1ZT5P1dH1vGt1vHnLUxTcZQjLRsMP
eQ1gWqATbCjZx0spmVHtnuBSZMQfWclQ3RDLl8VNxvv+T/DokrKraBibdRlqtyMnjF7TL78dCPOP
zd9Oo7K5RBfWpY1OWsT6PE9w4g2v1kzdOuPJxkmKUtyysFmq28WAx2+4ISD+FNe74DF4x0bFwXRg
+qvKV+Sh2oKOW8Z7T9f26AYC433Li3TalnjH7aFRjMrTHCdIlha6XraFwlOanBeeMpFL2UW5466r
husrGoRxaetCmcC3XZHK33q8i59/52h+tvIW0g2G+Y8SVLo6+D5HpXZqNhhUl7hQ+fkhESbuKLfZ
6i2c7RchoLCHqB6ibqtPOjWnbSncbBIBLx+kXKxfCn0f1PnnmG2lWpnrdiQgmwxrMmkZgGFuK4hw
ZUzwu6IFsJePMOsV0GWHcFacQDL1NFRzwByM07H3EwcNwE49yUsn81eoNhWM4W7kNEIPurBRFeA7
uCvwhui9Vn/7kw4PIX7ucSvFOm9eiGSqDySxyXU+Mw71WUWmHGKOuqgF57EqDZ7EaKhGPDxxYNoP
H7sujztqKhb1kJyO8mPd5KcQ9eJLoiCokAg3523/DB85T8/ju3aAhjTq/pxeJRMRgr/+++P2bj6B
qyhmr2xTvjICWucvoqnsbl/YHc1fo6k79AMSpeKnWhHjWBXPiepmWqAb/Y0Hm0O6WNKEYz8y7Ky0
XnkroE6jElLIyJuSJUjtkbGiAJ14nxlQC69dimXhUlmB2bp6ATRjq8+gXfNMSYBHEDf6+T4rvg3n
KMHYXtswc9mp5BA6LPIu62E6kMCbJCV5wpFFoCtfdQXR2bw0aGbGgUk1LCnBEcWNiV1mQbW0hsEg
L/Nk5wESQw40rU/2rh1yDifAU7YnsVn6QT3WECfrZVAQnATdrYTEWGvj66hF0IuBGaV1aI2QsCoI
VoPZ9/9rNxbi545KAQMwry+sqIBH1Qq9EB0DKzigw23rqLkV00dTetVd7kJb5j0T7BjTE+pWo7wA
FXopaHZWPdbWs+lKM8zOJy+PEFbLDq8sQXLH3ilpUvsG6jkHfyyP9Rgl0B1EgiGNtFi3PgYc9vCw
noD5EWH2vXN4oCGzxts6QgCMEMXaOCcj2MpdVlKJ9AzIOuBCJOBlvFOn7hfLsN/1NX384uo7rlar
zRkFdxaNM+055l36Ne3n6tQmUe2vKfKdT90I7Nr2QdoPJ0APFBvuuyDaMifLJciGun3HONBFbPOS
TAewPaUpHp7CUJPahC/LoWRm4HyeNu1Fm5KKrEkka4ARy72AYIkwVUzV9WmyfrrOq8I3QyYDuRiZ
GDxiQyWgG6ue+NuOKz/HOQVB7ydDZosRA53snNjUyHkC+4Nevdrc3k9J3ZtU4zt+eS5nq8vR6mwy
bvRd4JSw0JTqlcQDYap1H0gNxcHG9xLarNmsqZ5DyFdIuP43oBk0x8nbMnSrIb6Y7jGaMKhguiQP
KeJTlc7QXCviUGy+sKAp5RKnXy7LgIH999zLx/wshqKjN+gQF/AxK44UCFyKYEubeJnbwMksMLTO
YAGwpwnqFEi32Z05FCiKgXwifwAZx5QQxQwX+7yBt+1wCkTLczFl5sQlgw1pN/RVwnePtBPCGm+G
fT9QXvL8XuKjc5DscPLwMlnpKCz9IuQpEEiOcQHoYZku/GJaQfhQadcI8Yg+Nd+PkljrxwMqmpn1
3sEc6rtfQP4cDoBhDMXUKHOtebPnxRQzZtX7M1BjPsO6VRhB49XJFm7qLAsdPR5nii7ISGWWRbA9
cOvjgpnUN+5aELayWY26Ewu3H/8mA3mKUaQjBC8Mk+B/cpFH8f3tOQrHWV/yhb9Fk1fEtMNxeDgT
2HnPNc9VjYrEoczlcuCNuC2KPbpOjXdXr/R041llj48ZXxpKrPi+sqnMH5mgMusT/GEnZx0CNoOB
GNr7SdEOJFnFZeg+jOoSSVOtmeTSBkjGyl5sL6YFrdDzeu8vYzCnpuGixYltVeZrL3o7/W+Z5IcO
WDYP7yEKw3/F7YFMYBEFjtOxrsOYf+YTDNVJhd2RIn8gWr3hFAeB+MqLeCnK9R1shJRdmdN/O5mN
Uq4KA8hpnXDs5XHHucWbkIIpghkIHWBh0L8R9WqpJAEq9Ow6qwTQWuE78pqa0uFd3w4qU0Z+B2l+
3Nc4mBDDfjbrzCsCcruPApRucmWE4YnFI3IOfJIi7zN7nUKjCh8E8Q4ls/p1UrfFwAPiGJJMvhep
ToR7O9Tu0y1JbyOi0B1Hct74voTAKe21W2WQQClvDNPkx64wEYWQo+KgyRTvYDXwFjc3RPq4sdcX
21hevBkOeUzORpV85rh3Dgqagi3XcGAWJYxgrtHY7CCZEh1ouYI/IViCywAq1JoHQfXX1R0pg8Mm
c11hvV1hgHp2bv6AefYco0nEK3w4EGntvkrHWXzAHDGD3zWe1++zhphYS+vYuC5F2XeoM3d/NpIL
hm8642il/oOBaxrfTF1Q5LCZJ1L+E5iwE2wJ4dOAdo83XzJvMOQ3qaGiHG83xPyNt4dj5ac1wJH5
Sw1pQfrD9tEg4Gz6d/gTp8FIufP1DE9EKBSx9DhKrEgLCtO8sUQ+1gYVA3ls68XL/2EZAolXBlNX
kZRyc/n0HvmGmGIgyKwSVdVb2bE6TdNJDCwpu7Bc0qYZUfEcLVwsFR94DqZhA2Ee0TYtIOGlsbBW
MkHOQt1wta4RtnGGQdH7AaYIkzhv4k3/v+36sfJ/lClcMznA3Iqo4ZKAUG1eMJJMQ5XYZwSlfQb0
NoSQn7tGKGlrNzTSPXvEqZdMY90WIuWLKU255Exw1OZ1OkyKzH+otDqjuI3TPV9Sf7H6PINffTWn
AKuCeBeeC6pJ/msjGcHXAxbs0MLULhdAYpcqxJA6eT9Z66nkcNqF7H4L9d/I8WfHH1nNZnDgwSQs
v2+iJReXRwbvl2kVuQLtIPRXtVO2fqM5+oRYeN7PKiVLAYg2MGsa/hPEkMYB6TVjRBGa5TnAWANK
QUX3kN8V9f7KOnH5xmowxboLvfblB/wlFFWBgkuQO01RPiPd4z47FS4dEGHhJrGLRvZjNSj3GQzN
xyWkEdJwQOE+5kjWHVFzU06AtKV0msfvGJVp1Wm8cVaeXGUVNoXjnY4OSfetQqi+itrfvhvpB5Sr
43u/HGbBBaJzbXzpARqU7IY1WGSa45YauttBYXrPU+LgyaP728/lEMllUy3YQeA8Fx8mOyfDLz+I
IxnKi2fvn40lbxPbtvtG5/EPrTLfTxXphImTuEysyqiQ6IPWeXNsiA8mTRqpadr09WssnAMISKnT
A+SUyZzMpevJKa0yAh3H4E6PiSQorXsjlxjoappILlcGGk8LwaSGr75yPWj45m4yywvf+s0J6/fv
Wmqq7tOK+Ec+usjTeRv7sGesBgT6dAg3TxjRfgLhlGLu7BJaW0zdoxGPIe97As8vTELdn8/VKzkJ
pJJM8eZuEmrPFOqtr5TvAI5XQ3/yU+nWsmDjLk6ptZG+EIqpkzMcBidsI5aRKwflmcPTcVwHd242
YFBAnuX/hlOSG4Vgb/zEXno7X1Be08oHk5S54N3gI5omMWy1FVDEOcZelsEh+2W9YJFCy4ozG61x
PTLxoUJnPW6WlxrxPcpDBShKoft2G6NdQIM7RAulFffTM02Rca1lKYg6suEwlBu1nk1isRdl6Fpv
/zRrJT05xA2UPQgKpsREr0zh3o2QzoyCW6x4SY7H0Q8/hLX+iZkYBmbWpR1myqEiXsAh6TE8Luwp
rM8hBSLITvhJD0qwAdDQOg7gkcn5fgkAf7bSIucL2bQNNyagyKSTcrm0xJRSFJiwuUgZ7y56+Uul
zFQ5/Bj5RpV+3ulDF/3BkImzik9aVBd+/mGacpXGrfaKpatGZrzsj9YKg7jWHo2zLbfEtpBJVQao
id/Q0VJ4ZqYzNZPq9F00qR9146sy4GdvBWRo25GgHyE7uhH9gpHqd/ZMEsnhQDfP2RJV+VHzig37
B18lwHxbNvxrNMsjBYc5RayJhCdN2VUajA/iRINxG1i7GzW+rbMbingc+3pMJ+q21dQYszv5nWR+
wlNWQIKVSYCGZs/ICFZ8eLHWVxUUuEhe7uBwX61U3Esd753YqH+pebKqu36pV5m5ehArTRVvjk1m
WwaovsXDaCeWSW09Cn/c6AMG1xR4NMiMeChXHaLN3JftpmvYd4xjf0SiWATwSs+YUgxeF7QIZWFO
+xibNtJ5ArssNXXG48aVGe99QSLFsE5MoOqOjqWXhdoHnlwqj8+BmgdvfUpoVs+hbTmnyCqkuk/1
5XCGb+NIfSNXMcIm3t7yclOCXuNJKgRAqsWP7sLdPLzOVut4EKJVprEnsusZGgn0DPpqvyP/4S6t
LYAB9TxO+7TH1YuXcZ0ZqJBjd9FlNhTCCBHykF+rwkwLUMQr9rHqoCb8O3cHfLDC6YCjJITXiXmv
8sHSJWoH6jl7U3DCIeEZ8BtpbFk81u7iaJZjIR//xng8y2zeLaLEtStaG73RSkkGHDssA9a/Pk+B
vstyydbWLTSAQELmToLzBXj4ETr01Va0s7y5O1xtKYfPYxodY5InLgSeLb3XBsJlrOu9+Eq/Znlv
ZAPQgD5hSiZWdDfZEvIaaknp265SJt8/PtiyrwcCq/9PnxaUAkPsUWVYpOA8E6HdmguKR9z4aoiK
dAyvvwoCwqssUjwGZ1mRNsiJUrqcz7SvF4vtzeD38zbmFEixxpJSazVJC3dwCObBHTq5C0EOXQAC
kC8vCUDXjeNY+dS7hDFvqP422hTesbwgIBXFYOFxQNe/h9VtfsZVdxNOkQdBeZ9ZxommGgGKqpkU
+V5hHBW3DjqK8ouMYA8wByhpGsDbUKQDid6qsmLKhuszzDi4HezZtwyxuXFhoLSBGadL21fXh4AG
hoNzgw3JaH1AG4gZcyMsF5DXZTiVDx9nEiVe5MvrKT98kUc1ZLrECHiNh9Uu0eCdtIdD144nWIcR
S9qBtrRJr83fAyEapTkbTU5LOr6z5+hHpZpBdmDW6kxtsbl73cNEnQWFFf2Ql61yyAg0JS73+i26
+R098R8/4yX8bvg7RrMbC8ANaKK1mh06rN+O2HqkTJ4ARjX95b5nI9otMzTpsJleKOY/K6TETBI+
InG19RWvgoartUSGcwMFcU+g6J+9fmm46DiBeVgcapLnxOdLSS2out3q+IDiIELoZFVHFqebpXge
YuZEMzYBMdrvlDLaXCcvqt2sL/FXk+O+PYlMD+4ZIShnXoXFXGmTbwR41euhGp6CAEIF0gAys9jz
Hks8GkPKW6zljrJMD6GgfxSjlal+i1hcnOY/Cu3R7PC3hHBFE6j/J0X5Z9/Y2N6toGavb0hwS+Tg
RRwxbZWA+qAM8aQzzlOAK+zugbbtc56rPivjX7IcsjDGV2UtYB5SkmRpDG+2gyuBK2N5DZUbLBhL
KhOClgMRSO39onnguBXNiCFTyxxrbaPCUucoOmLeNj6h9K7mJcM8mbaOosMKSJP63fb+vikLjKuy
PtiOmUzUnAdRqXgoBm/XGhu0VugYpKc9KurJ0tIWPdx7Et4ObR9eMcli0wP+gfvldvir6Yf9EM9N
1rQneeFL8K5FRXEys88EBnZT8UAIBAxh/ZZffrUm1v4HE8JsTSTkw4I6qDTTCscUHmjqJcBKhKrG
wAS3DI9Njzc4mn1+dw9t2PqtNlLfWbf8ixycxrmPgM+xATmnZjCcvPbZ7YOIkaZPgFC/0hc5QPhc
xhGPzM9T1PCrtKzUtXUI87aL8TsaM6h/v0W5Sc0Crcz/uZ7ZOsa7uKPUziDvvTquCtjmvZSOuMt7
OkTIkxkcSXL9J6yqBbUbrL/0oRshpVho0Rh2CUxB9CvYgn+9072nAHeSbcZD5fXLVlF/tN3Z3guI
8AcXUqmgHo3nBerg3oKzUbdFIl9mDEy+bzgDqY12MQwe+tZXjLr9O0lTCogteCjG8ZzJtCXlaUfq
05/XyTKDCPPLHHyi2S2T8UprM5P5e/0zNdO7VlUG5xNkbVFojOlnP2yzT8iTy9GCQqKcCWBjsFVF
3COhRc2zthKw6h3lm5Do9VV5zHcn7yLPiflioVQ2jSrtlg7IJCM2IZaItvzQKDCpIWAVkDxEoMMI
uZV4ASuqaiOo+pd6fTLfFvYNIl+07B3h1fhxsSlU974+OkLHqKaTu+9B+tcwIFYZktHQaYbqt/n0
e7DOoLO374anf3UBPzGD4f4Cu+ISwXhJr5AIMP+86kFEq80DurkEwP7gNeAYvnXzOWRRkjNC/ueu
A3zjvsw2A+dub8VSxWkanbfqLVPqEmelnVWL4/W9RDqy8RT+B+pKNuQo7n2pcHgbR8QatJIHSX7Z
mw+O+89Scv0J5k8CI1RAbtIvhF3AFNtbgmVAdh6NITnSSy4tWWg8A38LLAEkBnSDhpkAaOZ56iqS
j+ZxBydmpzzNSXt61JdTvNBplBYCkJBMS1I7GyzIrdIjC3VVxMpdVmLB/QmyDTrmsCeN6vBqwwZN
Ar+AxksMhs8leGRckhs+N+VyywsWL6xAEvODQDzUu6gcFdNTonNLUCIdEpGJTOm9cUQuJ7ahiwjU
pNm65h6+lnGVefkG1MZma91bbHYvQgOzrBnPfdcamjt1wCXSSCOebb96DAvsNcl2NzeIIEu5myZ1
7ad0CRXRNx1Hmr4HTjGAdtJS/4VCMwRHkwpR9ef9g4gf5NlkZ31Xr6an+jTh9FnJi+Nnk7yXRSiR
ITig27ldztuNmauOl8FBAyRwfCYyqnDrIS0byz9Sz9S8u4dbY9rfpToXMwV0Ypms95M20wXM4/7N
/wveLOz9gap0MP0KPZhLF8el+C2ab1/yIbpsk8OVmQydWH1PotvwCdqhzDjACocUnBDfN7x7QLqU
Ihyq7MxZk9wWhhghlhOrB9rSIcXY9UUlhpUVAYBNNZHOnLzIWqBBsoyCrlF9sZ0qkZENtuOQUiax
0Bea0XNXISDZJPi1CGO/90FVxgQeJtUt6K5HWAnhPat2XnMKFt0YMMS9D4K1s9KnLd1FQo5BqFT+
W4dOf1Xy8gPndWt0yirqRXAH38pCp93KUnAm5K2QfxYP8djm9WJ0m/5NtnSihptB2gSlrOBh6BiF
z4ZE1a3c0QK/4HpesweNxqqmsXpJRReGr6Pf3nZJTjmuBwJdfMvDcECeb3JUbYykuiX7glkOx9oJ
P/L6j+OuVnBMxLPF0WbWURYSGQhyifGRShig9RnIyrHGWtyogod51kF/FZu8j1sP9qXBExFHeTd2
oXl0dOsSRSQJcojwdxnGR/BdH5dT1ijC+Nc1NxA2oSLXll0892x/tPQ+WWlg1rCA0q5vakOp23er
pOEZgLhDmkfD0Wv6uXc2roWPotYB/JhMvu+EcL6vs2vGoFhdKg7+lbQ2vlahkS5z1K+XVRFzWrmt
/xegaZqmpm5EUmdx7jZB/dEUlbdQ5t+n4gDMvx9DalrHrCnZyqEOfrRLzA9Lg9VdDleGDv+H5Iqn
AG9j6K41PyoU4GIjwVeswZVlpgRYOw3moIzltOYR6N2uTjCDX2zSgIEc1KMvv7zh+Q6NvegY3Bfw
Hsbx5kOL9Mhxr6gI1CEid0N240KoJYwKnwmYZKg86xlPbKWxHGYxNcQ8kivNqGy3+SOP0WDnQEQ4
I2P5x/vhj65ZPuUmVm8c3vF5H3vueHGA5aR6HlKmgdgB7KkoBp02dwu4rhTfUvp4ZAIh4yNZ7e5l
IpW0gImcBXXsflx0AgGqA0VxKdUi+h6TlrsiCmcl04Vj+YD1YSuj66Ln6ZgheTpcNHr6unzyZyw5
rxu7ATjteYffDaDiGny0jKz/Gz/GCET1lCrTCAhQyz5qSi3gep53psEpOj5/PSNVWr9WjbLL1VbZ
//NQf00LHNDlP4LbjdZMaPpjYXvcGNvfHzOtrbZYmnFwAiYQlMUZO0kt4sZSNJ4VHAO4EWQM3tZz
ySkqpC3iw4k6GwHyLhmIE/NWIHGLX+nP7Z87/9IezA4+rSTiDyzKxUzzkdoc5bWfj0OkXhtwSvPa
DcZHo/RfA/FPT3ojpbYRLom0q2U9IDSD7EoT85A1R2JdP5/MZE4tEdiGOTD9Rk95iWjvFN42n7t7
cy+4nuio+JPhOZLlTkhlRtC9Tphp9HFfHwCGDqQ0tgl71xUGFl0FF0KXDRE8UO0UPmAZQ9qd0xeL
VMB61pAep2xQw/rB7S6A35j52zGTNrBv/d81OgqIi589Xv3QRZwTyOPqHwz4+PNQKKrrcTHGerPh
MfrPFSV3gztc+42ExRliYAmL/4zrea7pgwQ+dyX/zZkTfzqGpPkm7tK9RjauD9nx9ok594V4bRdC
YZhCNxlyz5lbIui99X4N2DscXeGO0lB7RFjSoLYucIhIv/k91TP5X9kTRlYmE8eOsNZ8sSrWl02m
7nTB/hGePFPB82+mr/0zqi4pxlAX5hQUzV7hA9qrZ+CXXlQywRASOk/Pcf8YgyT0elrdk9uOvX3f
EeFS2QZhteSjwEGJX6QHVMvHVlq2+h8osLm79ZGEZc2v3Av0pgQPRHNbdaDGnHzkGo1JWKBh/Cdb
SGCKC9Brpoi2GwYnfXHsuL6iMfyQFFBad8dHVRPCBszHRyBWxujmH0DMoA3/19QIyjSwhxKBCmza
MAGqzYDFpCTrsNW1RbIgLg04TOhlkAmbDzqASV9x2Y45+ZxF0OB1tPDYwDlhMnd09Ctz/UTrkOeq
HoUPLx5Qj2aWgEjMUIH/gtaCru2ALXr+aIb80y2vWVhj/g8CUywbUpG8TT3kgMyPi8J6H6H7V3bc
DBLJH5X7WYIFC9kLp/elWOibM8memQR6Y44DO4scYWPYjyp4/Iq2GDkS8ZYx4rQjqf2vIsU09mjj
c+4lV50bj0QXTeHRs1Twc5CnTDvK49X0IrLu31w3RLdPr4irnVIQUkL9hRZ45BM1h2qvMpxnAouv
4egNB5YkT79MZgH1FQmblCRRMemlQBHa8UkBMNwqudEp0wbTp/qA3Rca3MZmoFMt64y0w3HA1zi7
G2uWI4vWA7VFvR+IwdZVadKs1dF0XNoj3d9ta6NSXZJa/FDdDFUwXrJ/ltMl1rH5vrw0TSZK3Dim
taqMX3O1NL04WIx7zJGVT7gVGah3LfvJ07SsVOU9Y/FBieRo4Az4yAKxNCSNecfQIXGIOf9Qlcou
fYFKuz+Occ9ClW4Q5ggAWjgEoGhVGWrXf6Ix6l/rtUsXxjg6pqgLtT9jb/5aBaazaZDog/6ioMUb
4Z4HRezO0AP/uLeUkUnDPCNTWvePz5dR3KL9e3LLvcMv0e+iMkXVFIM8eNCZbAoSoXoWF+5Rbk/o
Y7dWALl6FVgoFvf8WWkt9pscu8k06JcvXfTNk3HRgEXdVmb+qmLR27iX7A8uhMSpNns9MxvNtw/I
GCAZlxqYoe/WteCTXRPK82awCSX0mrCUFhU/cdq018UouiXlIFmTTJOAcqTwFet8HGW27a5pNieB
P+VlkdEAA+DKHCi0TZESnYblO1gkavyD/R+QUBmk1dHkUUzrz2wZQMdzskT7qybOJXdaRqFlz4Su
1wvotnhhYtk9rvyunfgaLw+xUJWk5J9C4qOUzX7Pk1LGxfOl7nqugpaDGPzTcVW/VNpOmgO7eyQr
kWMpJXCniHF3uze4t1aJk2fZDmQ7XI1ltRAiJBHRgLXpqWkhGloYe87bCOYcWL5+d+agYJNCsDpN
tuUXeSvMrTq4bbCa2w3MJLXdWfSqSZljjcfEZsZeInCt+Wkr1o82D8lIT6tZFMkbxSghs/x4ELkW
LRiRouM/fWjKNSE69wpjYNirF1fllW57Kk60qX5yj+2VNGhdAHPT0BY0SsltGh+uCDiVr/9DC6mJ
+UECZToEHPRKc7UJuM9rOBHmaSoiN/cE7PF2O0RaCJ4MxpsvjPYd3hAWo14CHuQiUqBHhV9Bh18x
zo7M88HqlkpbpRrXJu3nWI4LNLwNRWoacZLJ/6aa6XxFxrkC9SxnuJkyD1HM9Ar9uRESTyXfdKLp
dMN5oWDJNbh0ceHISo6BsqpY/sPCUF2b1u9QYh3jxRXJqCJDGk4lCb3pXcc7zAgtsF8ByPmEf62+
2/D5Nkvme8Rn1pNirPwMeGnBfHJz6EkYXeLQ08MHolNrzq4YtXswI4vhSShsJlrXbd0g2cgjV25y
JSrWf+UX4tzmswnjq6GCnOUiAw5llvrV5lfEwdoOhvpOCkmaU9usz/eNb8p8VEzSAX2oK05J8eTf
2qDKNpz2jdWAdhiJF0cY5G5p0CFX6SM0kijZKkm2GN1Os3j+Iyet7t+yVkOAt9afQTS0IUV5UOV/
YncWYw0SMtSKitJPftGTf4baWXrKLJkarj51Wne/NkZR4TAhpDA+mXtDH/iQo+pVmDhogNljMHvN
sFR9c9p2i0g17J9FAhq6EZoS0yXtTsvrvRKxDiOCqjytNo+T/AR+5luKXUzwISPafdHjKq41dj5Z
0F3xOtg9sSrW+pe8Wxh8lhfd/laxuYXqT1AUvzX1lZDvtIdxWCz7RTtvNZrSWVG2KChk+gunZJEO
wMYbfbz0PYxCX0MEgyNRFlgpue8mjVmNnbwkzcUtnqqqs8gxRyyyog0q27FBz9fn/IUIdGISe0fF
c6sBmjVxS2l9FXOF/YiOXxlwgPi5Y1a8HoWzHg+5cxbIYBFqwHxMsHv04jvJ7qoz5prtWlHyBpdP
z/FHo0vt+V0eoRX31clDuJlci+QgleV0jtaRz8JR3HtDtpjjinD8iL4qauMEM5geDU6Sk+Z7IwOX
Ljh7y4jybCiTtYj33wEsZEZAzW6VH17Aim0BmFUQSoq4oQgEt9kP89hDEBWvJ4v+gFa8TtKhNxw2
4bIuRO/Y8PUMwCk4P4dPKPaUrbVtptFe/Z601HQxd5I4p8b7FulEd9fdGZkeBBtXjsm40/lqgWI2
fFxyU4sUgPNXNrtwU0yaqL7W7m6rKvpWzCG7JlWb+kqUDsvxsiwAsevEN5Lqw0fBZbBu8guWndVT
PzSCeMnYqoHY8J/I7JcL7KinS2ZPhv7GO4PfY0FHbfFwNwwKORXcyjbrnl4ivLGOASjeRaUMJx9N
stNGnrBrhnyt2mla4zxo7SIehjz20wqIxBa06YS5t/elhHhJp6dhGrPH3TzsH1U76Ll5EOLD8pc1
NCnK3s09Rs02DOUph2m6AxfjUqREFmpyolF/0MjkiDTu4R2lX4IOmnBdSOWxxkRlIx9eq3bkdPyS
txYNvU57RtM8lcwE8bZGrA/hwzVdzY9R1SYAsbtywhWQJxmLeZcH86YFEqcYqoxlQOfg0pbVJmi6
Uqd6Qw/utjFUuZktV4UWTXuBs8HDDk1Pd7boWYFbHdWvBXsjCpE1++LQY4QMuE+3Em/DwUx2rM7P
OJdIKUurNWYvvkxlLL/cdJFZjTgx8DJCXGrPLLxyQc/FTRpjGen83a8GDiqzyzgvBegcHcAePAQN
EHZgz9I65RQrkSfTY7aXFFSCfP2btCLEf0MkwD/nE3/fPvkxlsCvdXNaG/bIZgZ41m+tocLWoFT2
03fflKM1Ou5r5oSDAwiIZimUSuZw/8cmaDLx4cUyN0jSW0EUaVW0rd508tLESFwZ5qrENtvVFQQO
J8yUbcW7bZqE8Ibp1XLhr37hH3dlY2Jbl+bDMpDe/Yi3Grg3hbn1xX1iMz1JXzkxcU1aSvhV5F+p
PlkK+3ZMlSAl33AREPEDpcQOF0e4qccW5WdBWn590h8FaOv4c3zIgvb7PO/qOak7TS9tKo+/kwRR
+XpTUvsW9G9yDuyGVZXUtkIM6lPl0EOOFzlTctca3wEVQbOnlbhC+tZwCvpUj839Gjfq426I3YFN
NanWgBfpbde1ERFWlDhTzVpoN5GAdjIaOuq4xlHQcmSTRdf1JwbgC9Y6/NPlY32W5xoyDwgqkrm/
rOIX//kUVozp1rwCNhN+mZIALOUe4RF0dO/mzmgqYYPRqOISrdXmqyogbONm6QOTLRTfZHErUq0V
pGeJW1RzxZVUIhdAETNVtWG+EfH3lxKd8hKSTz5xWYtDC/uZrMOlAWbkZQve/gK+6jEK/MQ4Hs0y
ZoZD4e9M67CnKaAwmqu24ezXhNeMsnUEN56+qpmWBrhF97emF+A4BQh6/8z4Lw0nf+F+L7kg2DEr
RDrSKvstuohvG4vXzkzdqNF5dj7Fg6XBr6dyImRmv4DNBBA5Ld2NYpw8KxPR4chhM+rPBe60Nzio
lr3LqWZhtusdZCctNrrNwpV8xO6X2D287eCcpRPNFECnYTg0NzBYbFMgGjsWHZK7cH0fYadGCBvX
mimwY7A4P34Ef1gSvlPf/m7GZ6Rb1IEr1V8kq7udX9kBiuegVxdneMhZgt1qFwZ1bOMkHGejh+cK
Md2YOXDtZIrI4Rly+5lBd5TB+OG8qfMw16XLEZ/mHlXuBGUsDu61w5AyFsGTMtgc021pJRuyKRCm
r3ZcUE1S15/FuFXAFK7ziE8vBo607K4chV1cSpyhU+k9dFFZPBpK5KCj3Sy4lSnwKk2DFIcvYoIw
uLkJYlCs0D14LGmdrhWOHXJCisaQyCHVcGJjgRvQDvaQu2A5+JcYqrGfts2V4y8MCEi8RU77uIEO
EWKldkToWykXkScUuSD4fBBiOHpWyz6roC0VHLDDHW70BXOHqNkzy4gQHPWQwQE4goj0oz1l71Hf
N0a97eCatZjxZcCB5kWdX47cno8vO0UYyeArZek3zrmphHtAIttTOFqrFHGu/V9M+IFBLcIhW9op
jeETH7YpRUwauWzsyhHy2eY9nWGlGrrsIJG/6MDnCk5nNQl4w8deqchJ2dv8jhDo1PrJXkR0m0m3
T3OXZuIEOI5mxeiJLHRibZz7Jt1sdXDUqox6DgQQERjTsPihyG6ikxp9bAZYNkMyP864+bCypaIU
LYpECIAR2P1KI1tYV8jRdGGXpXCYFJ2LZ4RqlZe9RTGy4PmG2bPcnghfasxgYQCHb37TdjePTGyN
cdkspXCfK19M1Q1Bs7dgez4WNPWj+vgU+QOK39kvo21qDHy6nC9XsvGjWppE9/HI/No5TzM6sR51
7q11JayzvtOHExx0FWdee0WzeMOsPt+qnuHeAnCdPIx8oSl2Bk9ozwL7oFETFRVsBV+djOrz2157
upf5zz9kBbBcEGAULl2YJgIWHfMEf8psdinoXzjwZBnOi8HYFzVLtZ94PSaP8TKLHIVxdrUHOSLa
Te70MLUqrbkdCKXl8iCX2mvMNg+63DSvVAq5J+yLm+nzu/vtTrTvJY+CbJOY39m98qpiDK+nfcpR
AWkQ91tjt2DUe6aq3Rea7HjnmgYuive2cI9L7OxKbiSCQr2jMZZfI7sTWgnzF5Jxd7sKEgIEhof0
W1Xato6y77dNGPTxxwGTx0svw/9GRH0n2ViRb1HLd9W81xkgNM2y2wxUJ6+e0U6LyZmhgV0zbKIa
bbPFuNRL7EezrpZVgIDXzj4W40vmm2UKwnjxzz4DEtRXUgjA5gaXfroJOdtp4XnA/eMmQ+RBmbe9
V40MmNIM8FlGvyo6o8o3R8f+i4gOgwpB817XQEhxgnWXuPjJvDNkvgiA5eVJU11QJLJyI40nlgGj
AH9TTSb5Uo+UmpJVq6/7jPRYjohcaJdvOJM7EBwkRiaAQHHfJORw8QyM8Xe87qRHUBGbDc9bkisO
GS2QMmqGx56YBroF2ONA3q3VgaekxlAT6QDpy9DUBkSXavDJu2b12MTTxs9D5rP8Q3VSELlove8p
5gI09ru87Gpzfmaluh9kvecSH3bn1tWwxJ9b0OycA+0+Jnozf4whKuDzFIei9PcJS7jZp4QKfJ78
BTC4iMDQz6HPuXpDsJ8aXmZGC8sJDm6wp5xSvIGYprlBLCStnzcpItgUvjz0qayM+XfRm+LF+nDt
SFRv+qF4K/mjgXXd3ZaapihiuzJVaMvarwLQan/PDWYdf/NZ+e+vwhmFmb8u7ALVhy9jopHIKL+o
V9j9QBjF9drrlGFb8g1wuNWKhyJUHrDeK/NDGOoNns02q3pZxouR6CJ8ThUuQy99t6Jdmr1lxRSp
I4U79RWge1IywFx1iKFi7JdNEwPyhTSAM/YvpaLScuyhUBKALej17pdo/0KjZmrDFCRfAStvALXc
td93f9vWzfP08Fflp0qTgVozdxpYfpXHoc/ndf8n6XC/EhXsdzXkMTfwVdPAYStbuZwdqtZQn/2U
u019/LOAEElRDRWf/ijnS3P1GwpceqRy+L96YyZM+EddZ9FMWdXHN5GZogJFMUyoC6LwclwQpDH2
YHvQYhuXBWhX1aaVAZ3HW0VedvDwN5hEj26htRVpvl+BRt5xONZ7UKFYGgTmy+Reel54NcnigS1M
gTRqD4swXpkMCRfEbcvnloJQ8tbpjQOvJh0oiNr3G0Rh7P/agnNsg500S4YbRkfzYtN12R+0rC7r
cSK6SJ2T+Cmw1dXE69PMZg0J2poexXtaMnPtu9lnrqy5BYox41eFaiAPYEtq1HfS543AkgQxN7jY
q6MQP7l3yoFX164ROIuSqrX1vWccQ+Zs6/WYBX/bc9NfiSYuTbk/4gV5AKwGlZ6fWeCvd7zrc6UP
KW4ShgesYaYiUfmp7aNtjxKOZ5Bl37wAksVO8p6i+eibXes2Vp1cf8CiBXhUdveGvBPgO9s+9jsc
QS0qrFPO9tRfJDmA9ybhbah5DR3H5ISVpxZjeqDeOioT1vz4AcdBU3yvTbUe6uK9CXL8PeAggTtp
4SY0JIjCIZcNHSPZsClUEQS2F5oPJUXz4aPX7GcHZMUS3CgRg9ppCo8tuKxYbart8UHUOo6S04Rf
gtw6R6jDsztMQfKBSyEWiuydkjagPRW+vx6fyXkwWYW2d/b2okKdcET95GtB1RWkln4cEWZZ3+yN
BehFrULBA/RUfix/ymtMgGl8ZFrwIX6rPkXU4GBoVqXlIXnpjLhQEGC0MMYNogHKTyGD6KFtQnH/
Jk+VRtgs5E08JaM25UKbTTbHsVkH2oxAmmcxnTlFR2pmRY2wB4Bb6nC/Z53lcU5Knx54OQ2ongKv
/SA3NfPY7vYATmdRDGNyyrq4x77jBxbeFQd4QSZyaYbzPDRpZR9x5zg7/q2wkAKLua0I6ag6AcoC
kQ6jBqdHaVaUWxCGBAKL5SAgIsIU73VVDVHglaFwyA/CtmPpm0OZHyiTTsULpYd1I7Zp3mMfJwng
MP5yRRypGEmJ3+clf0RD+fwSTkBTMl9d0Q8GmehCjuEPSR0SWbWSwyXoMJ7yZsws/UPl8g34kIEk
2qwcQGySlznzuYMCEbKWs/gs4LSyy9uqsIktGre0t8RiB9FCrxACFutuzJvJpPRcT67NMzEye6Qa
Xkx8tjjzjrn2D0aRSJV54puandIsKCCelYwDkxknWqEukxPufS/n2QeNKRhP9PzShSr32vtKV6na
50M4HM/omJCwEI/uhtcWBYPWnQ6+6OjKa5pPy9vTgm132qcvhZ/E4WQXhr2kFF5a5hbeZ+xKFjrr
zboUeBWOy3+llIv8mH8OnIfiwq3WDmqOrqRO0ycQ5wUCjEpYbzgOWkZ7+riqDkFg+1vIxBSeb0jW
hHQ9dRsmkuxvSVEWx/vWLaseM0TxkX9e1aaEDrJHEacWgwhpkK07GtfaBGcP0NXPetnic4TI1WWP
rOvyiM7yJmXyun6OJH1aD/5I1L12OB/2YuN03caiHjqWRtzELHdaS+oWomCk+U9SmanSs++SUPrE
GRmyAG/OExyA3oV/Ig4d57RAyvVdEysG2e3UW9ydED57aIVNVJZM6CY6Pe7f2vHe+NsFx5g7nAm3
FrazJ1xAOKRYFamLWWrDqpBJk4nGCv3z178r5mVY2xL8a+ufgk3KLiMiESKcWE9OTB42sf7J/BL2
mVIV+/wqdWv2oKeM4uGHNm3nIwruXSG6n2JPwQv5/MM4eiJXjq2eiJF0H8JAizcgumj4MQ3++XXF
dKmxdkY3chbPngJBoiCbopF19R8vEvaJavzO9c9c7jGhxKvs66psJha/UMfC+nEKcPavKlDvbooy
I4dF3jQdFlv6As61Km+NzsSbxJDwu+DODSjeHtDEAFDWEcqpmgMggMsvoxFtgrQmJ4m9TmVO2lc0
XqU/z9ScIrfUIdWzOBPKuUYIYF0HdshCgeJQruBOBddTSeI1bm0t6fnb8auTi8EryXJrL4r5HUKP
+rMwH9+3AIVkNgLZMJspeqcizDHJycpkkPX3WZh3lxzQxzfH5qohzWKPw11ln5fewi5Nl0PuoHce
6x2jmFKMKqOyZdKKySAkcddUvuv0Nq6qUVrQLzPNTLh6E7EKSSPIEbIIgUU8O/jf7VB3tA5Pv6g8
nBrHgPx6i7srRTZP6e4u+BOM5hwHAU01e+DiRYswU6Zyj3Z+OzK5mLEh2HWlXNxPxxRwv23Y69FK
2gEU6zSra09mjQSz4qYS4H01i+uIM2WPzII+fnnitWkr0KuLxUHtjSHuVJeuZt16Wd8lRFDU4s/B
7psDB/5d+1EIWLfC5kmSKxUHQzZMf2/7BSc5utqKcALJoeUhKLXqFKyMOm/FBnWr188bFseOyWf4
0GKbu6lq1gcrfdxljgHW+C2WABfA5adeEJQ4JM+aZwozlpoDO63ysfbbh1RhWUvTGCdldYpBsghb
u1o+Ql0Spj55iBqg4dk+TUuCSq6PdyGqKewoydp7sPRg4lm8OVStsVV+FzfH2uA4UBjhq0UDiVE3
HMu5TRXeeiA55eh9MiTg5tPPXg4XjrckEiA4JFiy095j2JJ4C75gbr7dfqegyHtHG4HgkcurKTSz
+qijyuxt4/w3NizWhAdC/vxHkvffpfuNNThv1jcttvwWbX8rZ3tpE/oMnAyKuSG9Qqn7/e6unQ0k
woJqilREO6ooodSRbQFSddsu8jBaMHq5LvbsmPwv8mxGqKXMviiYY+/PZYEsIj2j9d3+Z3dU5+si
VhgSRDkUVERXzEfM+A2ypA7CEc0Z4ecDyYbO7QfpE+S0Afh5IjJ5IJVP5coG9mIG5Yt0XRWvqP4j
mub3FQPrEinCthJigmiRkpM4+VxngWtpXxV4zMoavmdnrUFmKQ/DqDPBaUqcKZKsMofRCgdLyXet
LkPA1B++l8lJWKWqod7CGyq+QnxW8F9s8uzOwdcNwvuqCy9TQZqmr+zAV+XOjwd2T+HWI/4vt6DG
ggZ5+hqAVs1uVTcHmCqvNL77lj9VIlNC8OwVmlKynoTT4a4GKd/wUnAXPU06GxwrNSVT+fAKevdB
bo3VqASDvV8UzIelT4zRh+DM23aDtvi+JlRY3PEwgiVOvb96EkW9RWY7csDvvQx8Cwar2A/5vcxp
X9+T9DyoePOR1a/v8XcDoTSdIl7E4AOoXM1AovZUbIoGtvOXmiRcjXIbNpCdor20/Czg7bd3Jv8n
u9n8vsqwjENeMH2HoE8Rg4FLEvHo1vr5LpeGbrgAeaywwOaxAPTsDR+fcsmEXMXn+HEByE/LN7QA
MPqmHuBTa4qulMc++xL+RdteHV0DAk+zc0irZZCK3ipnBbLvT+1vpKBgKRSWbvK/l3k/6KQATWxw
bWF+fzjk+m7oAwltAVafuLgmHoyH20p0NIubN3H21vmCddk4uDy4+oyt+Ick+mjZsddbrXO8uwRx
nvqPhLwE5bHc9gJmEyabr1t47gB8vEZPbh1Mywur0FJT6RnAeTe0RValqgsjKw2E7yzsy1bpiF9T
+gt6infOEzBz2KR6uw2t05Cfd1TAHt1q/WLXTIkh6WkBSgGlKdw8ehDgD9HIuwNC8t6GWgTHSxte
7Y1DjdHDQLej7j3HRdfXO74pXPyiTHn6dcMZoo0z/2jbHER1yhyakMgAmVW0KxOuLtSfH38lpbhA
Hd/jGYoBfnGg3Yjcd9H5JNebzrpubqGDrwl+APXzSmH1UElsYPes0CusXp1MOCCK14BMYaoVg8SL
uqs/R4YLsORAESmzGhKj9pl9bK4eYLlRATXoEirZ++CKQc/n+hBo2K7QiOKajAAYnpYkHfIFri1l
uOIQ2BWXcFCiQerO1MxjJ4KLqp44cYjfQ9T3uMiaUnHhTWVJFOitqXxxHeB6fl9chow6KtKcuQM7
aKt4qC8xoBo3QPPPN0RKuL8Llz67O8PeGL/pPQKMCylREIG6WrMTeUCMzz3wbRX2DfmZeWdNR4yT
MpZW1nr/7LgjqP8uecHHj+KqjA9DZwQQbIKsU7cXpRCmcY5ZPvpkOSEQtehVrbOASS/llaIycyG9
AXEHz7BUx+BVB66wVSjtcG2ZYTtb3jUKTtK1RSsWp8UJuqK+cT0hrLKEy7UUo2VQW2DLufdUjXOy
txYy24fYRHFr7XIRPZooitca1VG8G2BOGiDX/Rc+V9FswjIV0M3eP5CMGTFfrT0Lt67yQsOmrB/T
YkEk5P3cVJZIyAEMd8EVPqxrQdrrO7WCyUcV6zS2THMyFxCPoKyc8Oh0eaHU6N9/lX04Wb+xJXEB
W3C1MyIQecSXcCDge6VUfK4BlSbPIRB10m1rUMXT5rpnXbDnhivvz/GuJ0JjzLW0tKMcanTYj/Bw
/VGfsRZ4Q8YungtHynSMdddmCfr4bFx25XFg2LY/oFxUtZ7HCLGY5WeA0qa2KLyfIbqhooem/kLW
qLRuzZaTAWyGLKZqw0AzZRtHqvqgQylJyBWg97uNp89nQ1CSYxeHW4tzke1ih6tNX6UO30H+wQFd
LYdFY6aD9PcERqrUFVnHLPaGxyio/0jME/0zZkDow3/pPXW30+K6rOH3YjhUCW7Cgl+iVDvDYKV4
tAirdpm3jb4qwKXGAjtRHKS1dagsg4agvI+vaRlr3nvBWTAbZr8URU9QUVzeniBG6cKI5uQdgj6T
uBik6S/Fs7yahDI1+pOL8hB9IEv6L41u/Lrnr12GJU+RvoxSQXgBMmHAgbpipBkWTg15qIAqYRmI
k8TUoRhyiofT92TDqfBqbbyTHXcmABhRnkhXhkDxuno+H0GgZg6PJOHJFbRgEIMYHQCgec9RmD9L
1KKEvoDE8Cl6ro3A1bj+Ry7IpSIOIpg8Njsi08uR5M2bNSF9mbXpHIdosDVN5hWMaxdtpQ6dQ2VU
+fVsJPS9zAawaFjspYh+LO4845ir1g4/txaIGJKBgZxDAHLsaxIsYr1cINI1YZroqXm257Ug6y7v
sknaNPVaf+2z0WMWlHkinYXJAx3PQRclcKdNHoHqZqzS6RoMAaRnfHXu13Uxu3jJUb6/FbuBTgCO
7KEIUS8TezCcQirdL6JvT3zxXaZh7rcAROEhRxW5p+Mjt8gOiyxVLiV+KrapeYZpwuMhSwWpbL/W
uTmzhKrOfNcPqPhWen5GFhyqNSR7vF3AjoFTzQdRg5zfNn/z25bRKaWaD5S7I9gHjz3Z6+Q5cnn5
fpaDYN9+xiScyBgjAylpqmgYuQnfk/SlNeZZwYSGjRNyLCdu/EqEUD6wXKMT1JztQ7rd8+hc8QcL
Qsv6MHvWsmK3HU0AhqpZl0vvOm3Z6zT85VrEZPZzkJSX0wIaGIq2AqycUps3Uurd/RISwDQeh9QU
gqZ40b+k1aTWa5qqdabSzyjxUk3jN5uD0q7vCcvpndg6AVKYj6pM2nv1mVUCTqy+Lyo4Sxk955gY
K/ukerF9HhvO3jAxZmoJxtwAWf18ANlmuf9OgXDq0AXENmenr0g8mP1wMViE+6baI8LIS98CtlsP
dCkNHpP9DFoEPoeg4uz/omy3zHu05YPYDTTgOTpgu5lOx6RIxEhtUs3kNCciU6Fne72/iE94LFqx
sC+BZ3kvn9iJIj5t0DMEBFqwNZnOMpzcRxG+GGToxh0BZIJp+G0Z9pYJMNBlpZMX/zpDHUzEA9HK
LnJfyey8YBUzDa9SG/jjPuaH8izRIZlx5Cd7ZdHACxjfd+EHvjHqJHRKk2D7Pgpor3nPIkQg8Yrb
GFFOBNjw60MTtrSrHcefGAAGpJuLXoPdnylCXfMoZUT8wVxa05/LPE2l9KLPsZaRSz8oWc9XbmyX
p02udkAWlBmloaq42fYgOxebRiF1dOQXn2O7SUu4vSroszz5J4W6uuYNo9KYJflpHnmUhNtIHtkS
UlbN+uGvAgbvDsWnsGqXiADDmqlYelPggpIkDD9o0e3G1mtjnoJuMtyCD/3SO4OSsuncDWDdA2YV
Hspb2WABDEmq+BRZQ8ZwKmWJ/XlUBxLfhYP0oSpIDEwLqRA21eE3RcZd+lhGFDdW9awIMBlhhcz2
+zFYD78U4z4tQizRc+s/PZmGk4mCz8VToY4fHMcCmbFkgkEMGwL/70fKsx4X+lHxftCpD35tKMhG
Bf+6ilecvmIhI1Yvnjgh3xBSYDKFJkY3Bp1e+k3BRX7n6B/ZkL5GXLH8PWrWvTCKECLA1Hg3wifZ
CU0tbQDd3Xa4JKHdjO2+LvFyicUXqTutrZiFOkPqtfvqdYRiWbtBTTpBWhcOh25uqr/EgS/8034B
2mB5vVN/wseuh6jyY6Ms/egEfJ2KNv8baRa+GYzUT2CBu7RkFUfbo9/nSyIUuZlCJOx4D04n7UHR
qB1VMSs24NFz7TZbnRHoww3Mycdk7FZpUtfWAl4b0OIqCDsHxCqJX63rxTK/jrtFirR7CGi20XJa
uN2SMvRh+rDfPboKYjtW0/0Xb96FJIK6DYTVOT3TKv8VLI2hrFf8srj8++VczHRx6gZuBi2Hsp2I
DJtpCyW5/t/llwLYar6H2qQ7ZEZOS9I8/N4MIvJsm/O5yyqKP9Oqcr/O/ejFCxwaOtlirhEz5UNN
BnNYh3S32sYrsSHdxkUgPZbhPWJucD8yV0jeK+7L4li8i298rDgVtwxqamDu1fQTjjxowlRPSd25
JErUcCFTjTSIsGPcEUvhTtgGfwhVBFYV3uQbzEB6ME7kHjQzuj/uSXKrqbMz5+vdYWdjUjINSGh8
7zCDmGSXJNbV5mfJitAZO66h1OmhoGto/V9cHBOyyh5CxC9w/cdtKAwHD+N2mu/gLMRdti8zmB2b
dU5hSq0U+7vV5khAm10bsOgI4Z+Bte5mDghG7xj2SIlWBdgalJJixzKV08FAX7ZWIyxwju12ImGX
JTxUhO+eiVwqFsR2KVp/nuHIs+5aTrj8oN9j9ARrvU41289319bSVg147Uk4ySBw5Dmdng+zQ/MJ
7b9T94VyknnlQuAZggxaHPuxXw1H5Xi+n3lV2CC8fzD+D6UOFnj+4TLiNQTj3oSojYEKk/NUYakr
goD7Qqzq4vDahnUvLpE/q/6K0sUhjYm0sfSgP7T677d9+1A5I9V/l4TsCbPbHOchf6OuHeDCDDsD
OxhauP9EoUr4U8f4t2ZtpjVXnZThD+imK89D2++0KpsTX0iJWFYfjhHgk/2KXAQlYgdY7B4xQWPh
AZCahhjr1PT9nwwdGpwawpCHm4qzRCjZfQluF026YBwsX3lFeezO1c+90NZjsPcsF64ibZKWm25C
e0k0b8ZQRGHdyBh8hj8b/EsZn3o1lr+nBuTADogLJRPR80Bk5K21lEjBWRPF3gVDAHxuCzgfv9Cb
tCFAkBpN5xy0EhjWn7mG1lGE6OQ7defAnSHwT5T6ds4Zklzoy/JjlGAylStkNY526bmkrqEXJxf+
mM3UvsW2zPj+yFXEERWDYcnhkWAON/C8eCgzwub/oJmDe5wiBT8hSK4sXyGC/675nc8D/Zuv7uPA
eCFtXL72QFV29l3Bu4jrDM0O6VJYTTGeACjv0WAq1y4jtz8tyLPXSPBdi9vuT9QffRPFGqgLOkIJ
wqmlexWyieHtrcuEYm7LE175vKTLHOqVeCqpWmNVoWeujtpzP2A1VtHOG6rIzZ/Aj+UDGkmA+CSa
tkbHt2rvOVuF3Q1AG/VvtFgCOTo1eDMbd45rTtqIdbUbczghEGYcAcKy0FH/J5Y/cRefqEdd3FGW
Jow5iYE9j7H36TC+Bwm90ECGvr3ctf2JYUIhq8YTy6/9AHrgnRqORQTdI37YqWValQDBKqpocQuw
5rA4JmuXJC35fj04+3+g5DgH9NWaDOTjj4w5pvn8cJawP0rm/98TYCzI3qvOcDRPGfKvJr1hnOMi
YmlhipuDbyNPDI8hQm05OCse8PgbhiEZO0P3QrGjmwfjikZJR/NC3CTyCD5KJCneRuP30MNyFQ1P
CxTBrwr97eiQu5E03Z0csmH6f0g5gwwk6fbr2eSiTW1k+NX7/+aV4enxvPtMno+OYFXOnh+5UGi2
UxSSuPJ0zZxTBW8b0i31pYiREqbJMxLcw96PzP7MB//8sJKXUT5pE9qfgPjlQnB4PC2mRrWhuJHi
KQ88HQPoCarSR+NPHSqHxe4uNPWIvkScPu7euxdc5urRx5WZTccFWypVd3EbOt9Qajr3fkiI/eXx
OQS8KVJJ+GJ3LQpa5IsSmdkuLt4IwIsv+9O9myMANCYALsyQ9g0LF1ejEirxqAZz1+/vnExDpwf+
eF0VbgDZ3nmFE2aClKIJQHIcVBr1oPpgfu6pzHG1RK5vJ5kLnHYMBq6j9Vl3MN+gMTGuQUR8bhMP
Fx6yY2Rtinylf4DvaxVDEDzTV7RwPTgP3tMGpcUJzTpZbUGtnZooYfWWtBZmUDV+TFyIPTapsW50
nf1aXRiJ0bVaVtxPCd2gBK0uON0dG59u1rMcvzLlonM+PRxGlVSbcRgnxTVBaM9CWSHMCPjbQSa7
zr3/5G531x3rfcHdgWhj5jOs/q0yzygiTLnx4TGr5TVamkHlwYFNa+E+HdjDb75XVWaw9L9BFGnz
5iwjYwFDM97Er44JXtO2faPbznO6BB+RMbM5UknfQcbnJJb1U4EtJuT/HF0y3Z5VPqn3PNA1EBBe
hS1iY79C9VC5uQlwzxvI7TgTtD27pQQ073x50mC0mkDgyvSURkcwKEIMGwcN2w0DFTZAVXvRGZGL
7UTnKS1TRHKl/uZEFdA9syfj5wwSbQBU9ONf7iOHZAuryU4IEeWHMj+KiG1rlLAjr5suPXhQEyi6
xB4gU655TY6w73+32Trhkw41wo0cJGPYVI9sMy7ImzHw+M1vPEqv9ZZp4+xgpaH+hO/7tz42fbZa
jW4KcS2+l+9oz/m1miQ9MyFIhMSWuEVGzhdn1gZOF40H6vCZMSCXGmJnJLRuHzn0yzqiWR2KotXq
SQbw0o6ONUe/h0UAvzK3jv00M5+pCH66GiZhBWhymUFEDVIeMno8ZSZ6VdyxmcNfRye7zwH8zIE1
LSMpoDtuYQuBljJUMHcuhj0dk8TcNsOihktOj6XpKF2t2QdmLV0un75CISj/9ACr592mKyhQrWkY
1zb9EhiAfD/zQzAODt9Xgz9dq1jP+s2Tk8Yau8GVDJoeEqq9FBE2p7cY9tf2n12i0k+qPBMhMtwO
glm6bGS3N6mD+8QDoCFnh+7HIZYxBU0YNSuVq+L2IVNLv9iLLDBYtlbg0z1E9vBzh4i25hhosGfQ
tfIxSn9mnZwIROMAqLIQWFVaJAqnxd9IQ+Q/dXxyfuZlhiKwLiEeHkYAPDFozb5LHWLTsDqo8emF
JBA0HeQgt7slvbCJsgmYqmB7iw3timplDWj3Ezmt4htqXoWOStEFt3TNV/e9oU5r7nJXhjpqp2ez
FsxAn+FlaBkoAd5B3rvmRf0VSqbsIKEtQiyskeIwFbN6FSlRHV4EUGoS0QgcuOwcqqQDr9WEVieA
BJuj8AZf+PCwDez0TOdBuCr+XXkZuvnBsoOO4WZkDfu3dKh0sluGYFxTfyWeXhXaug4VOqmQlfTJ
SDC5rQqYJmlxgoq6OREoBufF0aar+U1hHkl+kkS+8nkmdLjfz3/VQTe0jyPYZHVoF5Es2UZmWgqX
PU6y17nK+qqwRFwTKDLbYDNedPogu47avFPjdIf7QntgyYPiFDp/4ni7qRysLGsF96DFtm8qyTNy
3aJNIEVpCg9RU8JDp/tsM0n8SKM5eBicyL7hLabKTDQ7x0ZLcs+9evlRlL6Lil7dS4pXhC6sVhU0
9VnRaq1zCp7A7O+SSOpovAy50SoIVX11qP9yWuTZN142182bvUzQng3S3iS84bArU0peNMeZrmsP
6Y6IOiga1S1IJl+vQZ3X0J4L00ZmsSLzoVEnqVnmMa9JAeANYbroKCM4t/ny+TTuEFzcbOJSW/ls
cbpcghak7haBK5NOUCXb6v4AaHhgD2+7uga0E1t9L4o08THjyO2Hs+tVGpvvyfhRxAcdKVsSq77P
NWl87HsjvwEIXxM2k/cf8ux41outKDDRTWG1bTXfLIOUssx8NSlUOJlIQmXcypuXYfoCetwg6WJH
a3ZsU9xER/Bffh9lXsOcw7t8XIykFxIU1dpoZkZP8shqpmHHljOaDGHNL2tWqWvf/OP7bbezrLef
k1xtLUBQJizjijHrI5nH3VmGp9EmMwTr3hDUltGUere8Mc6pEOM+AoTS3DxMpgOFgRr+pwt0DGZ/
0JDVNg3cC+qcAMtSMfwWMYoiNeesrZHEQfGhMKTmmQuXaIacjXp/xQPo82v89mgvcHYZpOqz4els
i2FFJfQNsju7//TPZqNngnRZNjQD2jPawOgH4pIeOIDkWtFvFVIg/d141QUvLYLFQdBWt6VVCypE
jsNgHNABwDadEQ7rrcy3L0r8rc0JwXDzRefPhmZD4GPDx1o7Dhtovd2+CwPjhsAShNrehjOXt47Q
mDtn1gU6sTp1s+s31Z3C0fo70Xt6Mny8i9E8O5HKDCTF0DN3gCHaIzCcW0MVE0XKMPRdVBytUZJZ
0qB87CMlJdi9G2FwsKkv22HwWalV19xMmRspgVX4CiMod5S+WzRzLN+TrXjIT7QGvIBnUbuU+VBJ
1byh3HfAK5sARqKY7dObPQjxdeYGj/x0nPczJvkcnn8hxv1QwZcH62uZA/lXseRozprFaCDGLLgi
1KkBBySl005Yjlx+gskxHbna2C1uGVxezRK5qbfOAvDGrm2jeRdb/ei2Wk9n8tqIuviOTOoS/K7J
9ZgjTF/gGnjaToWOkJBbRDdHbfjXItGWh89aGuA3s4Olvj+IRYGUAdKPoScge+e4G63KvXzf5ViR
AF+OyXwiQxEfV/bLYnpquz1YWx1uyiPOzSWwa2A4FB2zeWhIiLMXM7dUgnAZRZh1O9bqRXhhncIJ
a2vybI0vZjJcwejud5Cz1flpaZ2mCu/KMWPaIhn7lZgZ6CcxSzmB9TEJDk6bLjsKRSc4ITtUW3yb
TiISDOshhKYrEOu4ho4YCXr5OP+D69Llca63zk/Ku0JUDy2ktas/WfEDL3cPZd7on+Y6kR1LSH4N
XyaDymUoUFkjrGXb4blW7j4ZXPkGiSKL9m/PjZwdcS4v7JcP0SYcoGyw1ow6O1aKOK76/Ca+We0t
8U/nH7aWFTMTQooUFceisCkdVJYDbq1vp+Agc5yDhBGRdMaoSTpSgbio6WwKN7Z2xPxTdCh4Q9ws
GkvtRWuKoYlMkTdcJmx+ZKjj2WJuiczf1ubqS9HKNnhyTSSuGj6fwYE3ewJ/NtTNEo8rHbRe53pf
xneMAhaPKICJ5DBzyE4YXf8FtjdcANXSdCK/ufqsCvqfooI/gnah9WmhsVNNDeV2ygKqlwK+uT/9
IjoP3ruhNQeLrK/PmEJv7+yPj+JDMjxpu6CG3JrHSfCl/EIv49IuYVeiLaGPmXavLV0y7+iF4hRG
/kPbtqpY5wsk+w5XkanrNFl2tLIR3NzDTCMjhmNAJ+yTHT8LjUtmN1CobHTe66AKYsVy8M73rwHJ
Aatj8FDOOmlBt46fH5BkqId3yc4q7SQtZjlo2Vzd2DO5Go6wwfdMk3H1epeQkwPSWrgLr5CK1H2X
RP8jz4fiSBFq6YcU6sF2Tz3z1txOcZFtwS0TygWTghqFeWFlT+CWxrggKr4jmjMFeVECXHkptA2g
o1nmXeuOSo7OfvUKKX+Rd71ZsYG+M83f2JExamH45goEQts2vTAzGlnx8IFz9YWakAWqKrdiHEsc
ryrQzBev1kBxYuHxMWJ7x/ssNkCZLOhzwAlM8YLUXGO7STSStMDe3qLiML6nQ/MYt7QhMpDVyR+W
WfXu32dP27j4YSy7B2x2wRGTytO2mgngVB/14c8CtkjbIAzJE5AOHgpGR/yaGUIkutr1uEmcwrg7
vnU3HkStjA1PExZv764paj3VyeSPzdzosGkx5UIIVEbTnOHKDk+dc1I1NmnrscUROv5vXzjwVQ1y
qOaic+EggNsCsij7aufKWzhdPd7mmoY8ms03vFKZOsdlHP4xAfjcSCbVyrsd1STVLBgmfb4b9usl
UWp+DzvdDN2Dr71gqD74vs3wu3xyiTpBYh5gw6pikq9v4df0mgLBuact6H73f8FL+DU4+DdYY4tZ
qAybuOssBBUSUzUP7sA2TDYgUK+Z/hxTZ72njhfk19LhAXpi7mN8nD1kqlnBC2nQYy9ESgSpMvqM
dEZCEKIaB92YkfrzCNgx9mQey/mu4mWralvmMBQCMdMYOj4XQZT17sZr6agn65hdCmNPaM+dg3C2
2jSVhyeRQfGXGqAD2mCOvJAqvajcVPKgCPEkUELowLy4gfL5nJVJ+jcTf0wJ4exm1n5giMvn0NLg
/gwcBBKHMUwGTTPJS8qaTE36AXSnWYI3EptZJNFKW9T8aubSF2dbLhzmqLOPc3isRxLbyUggtKZL
3/+PKfCX7ssc4GGbMQ9MdxmIb39YcngcvB22gNBIMxPS0EStGnE7BnI3TPvh7mFK3hpCi6VvI+S0
q6oSLrEnruQ0ZCMP3oty1HN38FtOfFT9kFTqOKkuUqmaiAtmqQciSJfCJF3OXMed1rpbFDdpyulC
BSOvYFi4H7nec28r6KCyaLKCqpxgVLeWxHz4KvnNEfOH5vGMFB7Io5l4qFViIiI9A+HP2iKNIqRr
f9tr4BGQpl04RmMqd3yWNDP1lu0zFd5/sgWOskFv494Cq5PLbOkG7+R0Hy2Vy47IZt1V2bn3Aqgj
uauh7IurtIqNfHq2N1NEpnBmkehKIAfyIEddHujD3MTIimHRZRwu9jwaCdx88lMF5mwHycg6O/0n
XzYC/u2tcuSzUCY9cKod+GVmJ8q9akm3qo8Id8Q8SlpoH1whUNlj/Bu/hYVDigW5EykbsACjEoff
6aVwKMz6wQW3Xf3YS454h8Lmh6eWnRmeIMqNmAoPBRWcrR3ZqynBVV9dNPARq9Rbz05lo2wRNuEB
xMJx11YdAtxDBCT3SHnvzBM+ZfuVi7VUsjMZtohoIq/jIdv/F1GZ9f/hL2UqvosYniWPvzjP9kAW
ElRdX48peY5mqwptr6igk6RyKO1+MTcaWLFMkZbkd0TtmDUhd4GnYMa6FUso47zQeT5+DEFts8Tk
h7lyX0L1wsjK9qqyNuHyNdId9afddhfUwI7CM6UO0IV+SSj8kGCk2EL/OdRwZr1w7XYLvU83dAh0
lsAIuPgSkvfc1rEU+rMTZsRIxnsS9vUiv6S2OgQu9cbeTFwqZHlzC+35cjB/7iD4oZHLKaYhnlj4
rFhSB3WW6/+c0TUpGNT2vkpny98Q3buhM7DnX6O5t7Ee7EQpSmIZOxanSwS+wxlf2xTvWYG4hQ+5
EnmmbKI83RL0yNfSMktalnCrChL6VDlvx0N7B88Jj3rarxTYbrNDqLWJRy8bdzD1VgUa7dqCvMmO
wstNBe7aElG8Nbg12+CFCn3GJ9YPTUxOL4s3PulP3kXwF4y0XqOyV7caLinrKUIXGAsK10ABkPbO
mpGsYPVkqNBqtWLU5FzKBXn2DO10bMMLQcp57H7+4+jl28aVeAewmBTWOd99nCXSlbjIJkdDH3uu
y9Ef5aWBpyElS8sKkc+ZRRg2MLWeX8PnyyPD8ARpd+SQG+TMixmRxc6vLyG6zC5rEw0vXrE0RiLe
e//SlwUwQ2v+Q8ZsaBQ8jxPXtwFXZ9vZeP1jNVTU0fmKqtZt0ZC+GU49LMM2kR4UspAabu/FjXbI
tXD5e9/xfyJah8HluLp2C4JVXE+69/SwiGmuehIRVtqfuc4CQtnnhWu7pLOMAB2GpsyZRNTEaDH7
x8yG+wHUu6XVIdETjlTzffE7l4qfz7LaC2rR8vuWErGa/K3WlHESK/+gf+48pjS8bCUFFYkz56YG
5BukElFshAEhvIy2lPhtUV38OIaletEcX6OFJodM704BQFnDjHhteE6+sfOlvLF4H7YRRRO0rRti
IDurl6Ak9E0LKz8WGV71NkqxATiO/jFVCnWdvXAP3RJSLtnjpe33Jc7hBt8e91tITLywJBBa6Blc
6Cn/3k4CNuRODBSvMAgbEcvGQHaVIUOpICpe4izmudZWhff3mZUSStG2bG8KFqxa0V6rID5FTYx1
Ek/fmDdpWbibqaMIMRez2aVuXb+TuwvTSiIFKz5o7LyUPUgV8aBoXvQSq6JYIP6EHfDZCZ9//b8Q
6b7Tdt9vwaQ+7R2a9WzXN8GTm/sUIPNE0EZCdg1SJO+Pe5BHwFKDBAG4LqQiAXuwruWVXyuJX6Zw
Qnw4RAKhawKWWxRzGQWTWk7F5ze9yolLtDVY95s4/2zBV0CHmp8Ch9L4IDofL9yfwOt8CIqbJZVF
psiW+gGgcv0yW3qE8av+lXkRlFtFFw7qdkv1NqhUw4RsyzyMpztA7ellXsalid6iIJaHHaYZ1XDk
4FgKtRB8PuuNjgphAP29fZ5EzL3nGC+l1NGNCdUH6uDSMudvNYKKW0yuWvpN6DMymMQYf6Stu7kO
420PHI1Pu9b/U8oFb4W9ceDF87ONaNR41RCItUYJj9GlKbZwV4097SDv3OKD2gJIfTAeCRGpzTVA
5p/ED98Ctie6OvRjOeJ0/AfDhTdjeP7amIHo+1YbxoxXINR7hY7nW95ZvFEv83yKvRXLrMQbcIEu
KR9kJ6Bz/SN5Rrh9rjDNr+Oa49vwMy2dCfizp7eSijjHAd8iBj6kSWgwiHTfHloEck2Tc6SjEaI8
2fib1FaigbXofBxy+2ESiI+WXPF3Wk+q6GIQhxpRZmEHgXzXaER4Hiy2laWHrOawtuP0X1PDGOC9
65DbjJWiLDd9T3GP2TfSIlTcVvwUovKuYLbDFzB8vtvYkuhZO7XiynuvIk+4E/e7PG9GiEkjJzlH
gndlqciqZFlE7MjiGwteM1qyDbO0mrhgp0zsndxBEIzvuKw65TVxVMFs5oT6jXX/Pi0/jsNHREiS
JGS0hh8x7WnFo8AOv94qWjOUY+WvKMER27QLWTZZp/KWSMb5ZCzV8ltBnU3WhIyg2/WwdncLkB8G
DJwZJeqMdPz/CMJl+JrntnF6WOHLC7a0ruyrq1C8Pp2Z95mPJ88X/1Ma9Q/RN1EqjlhFGXyeRaiu
H73IO7tW44OtmqR0lvoI456tJYbJAryEprM06q41M70y/FlUEqAOS4//ElbHP2vwM75Zxjs+S/Q0
At0sCg/xDXPZ4vszffwxnLzb9kYMCp3MoKVDJNuLe4cA5AwYVnFRxqZJj/MsfH0KTBPdXweYaR9p
Oj6RNJKz68KaLuJ3kREmX418oxmoA/WwpTsJz1JYL32ogltdC8KKYh1T6b7poBIRHQ+rqKuBnprx
+BJPVNWl+XKxCCVjUlB7WxyMKUS4Gy/qNBKO0F464h/lDx4EVEflptBWYUWFLZ0ADLvz/Ccvb+SH
wok5S16HSWAgL73+Wpul2n7yDSi6qOEoVKblJKpvXfUJ2PljTbPkOakO+bbOxWfhnYzaXNFC0Meo
exDYpqizZPyP4wHFNqvv/bk7v5P3q4Pj8/pj+sihYGj0FoX7RNvFIW9ahjkcC7nOKVXG9o51JZes
t4Ruhg5sVGQ20l0o4g3vh4VebYenH6DVSQhyygiBRVACWgBcm8zs8H9qZWdZX4i6nPmB2JqSDkXF
u4kP80RQK3Lzc4JR8I5bprRalOAn3kPh+CtX2J2ME3whvg1BaiSIb7Six/OtDPO7IJsHIdyJmouy
l2i/k1T60A1WNXpp+u1bPG6pKafZa3bp16K4O6YxT8RpoK51UvZhTPwu6i5xxOJwhB/SqA7LHm3R
fqP6Xllo8zbYNIYOgYrhpnY+GohqVjXS8jM6qset19f7QcgaiKxo8CnjkpSksdK62Atcx7+jeEtY
1tSy0aN8ZYCICuYFLfiVDAyAILJvvjAa9OLls2X+QhbgD9bUeW65t/vpNTzw0gsVfXDydH3B8Kdk
D51FmSo99npNFg/4dGQ+DV4soyGXVyoFd+1UNgWifE1JV8W+ANZ/6NeVeEMdgFuiPXj85ru0Mlzd
oWnfuL74or0t4UaZbgX0ufeYQ+vpdJ3C9MIW9sHRT0maCsZ59hjH+REZt740sXQeqXi29QM0SI2M
+rTRQxa7qG6OF0dqjpgSXYmJjNUTN4IiWf1dvzD90LShDIKHH9Rmd2VHrMZpno/KnEFuiX6Mtc+j
64x7ceGR39SrPrzwLU9kvcmue9+/bnlLRieBYpPzgJydJ/m/5l46E5nhuIYtGj1RZg1IeUcz0ZTW
jrNGxN4iXaR9RDAiLSCVsAiRsyM+dA5/lFq/Ye7mNWPA5a2k+wBLQKTUk3gnRyfYTuMQAFgQSRYu
4Pd4TM0S6XUP8ck29yicof+BR+eErkryjekyiYn0mquMTfw+CpO7mf3iyzau5weWPbxkPIxOaH1b
4+73XA5F5ZmRLBLwvoTrTSl7YUIUFGl39ejzIL0p4DFamnU8f35Db3M88LPVw8il2ZTAOZ2iV366
4Sd0pyrfSyP96AxyEZPy+ZTBg9BoK+oAtI+/fjLCAtCZeDkD/qzctFcWPczLAEAtpufbJ+H9vS/H
9diPoby0Q5pw+3jEpCvyquLRmsNzC0nxzmm9BSESLZ9lldpjy6zY3tZzKmDN50bZfJBRsLoZ5pZc
CT7UTPWwlj2PfouHrirdRQ+57P/y7uU/HTmEuczH19rvB2yAH6YD/RMQ7cxnOoQWfZkOGHvMoQRM
ddC0fARrWxaGxC1iyi20DTnlFlzbW+P6njlRcfJwm1Ll/E5GyMuGU45n83Dk4lPpqPdPs8SRS4+8
X2p7yLVtZ3WTzwgpr81Swto89/362RsYwg3nunb1LdPMGgH4NGDrfHWzhgEvwlp2fMeCBptqt/q6
lmzvrRshcJ/m5CGaajgfjeNESfzP1lptHQbac7UGJ1bY14j3eD+PeqhCZA9VnT7YM8CZbvZtG0Ch
ZBg/rruImcznYlhEepeX6zUn+znlmiHCrpp8sltQfa2vBSGTnVK9JmXlh62YwmlVnqxjCvFFJs6j
UeKMhGet+jOKcjkRkpuQmoIsEFoLF8lyhTn8lyVoXsw+hIrI56cdg+FGY045q2TzOWPA45e5Z0uH
iKM6J0eOTfFbR05haRzIxG1dPNveQREUBxXjhtVWeCeW+Q5w2TKdlxOadIIjOLFmugTVg6QKSBl5
j3mvyXK+pJA6aQqM/jVquCBH+dXT3fjlaeDYYecOrQ8Bwfm+OXtXOvS6Sgj41hy3if7XmoOS/Mqj
NB6vLCIQskb/2C45RBqcGLIOGT5Fxh1RdCmLxHuLEz7KSHOBf88pf3nnVgP92QVHp2Vd8r8WXnBS
nYVevJl/Fbfb0EOYYyhYs8+5cHqFzLV/2f0eY9Q1SC1xc1jmudLTz96QOhzrFyTJSOjIpyxbfSa3
k1CbNZtf5IaBS+IPOwx8FIFF9x3z2JwzJN2ZaAn6yqI+00UUQu6R8xZdkR3/X48zQHUNh0GKJ6cg
2yQX9tb2NlRKnYbAOLUIZbNFADSoIHs886bGkrfmLahUU8260gz6T272CDjSw0btvTtgufIUaQpn
qYzLJJSLE/XQIUuXdzbeo8Det+33v/XX2KBimN0peTJJXZGag9SYY19z4Tyshb7e0wz+H9qLlh0T
AdbTC7Xcl+EDC5GKagp3/zC4dmsion50xOEKUi3KDGsJVhT7bN1I+KI4/rAfh/b6ozcf5zg2S27r
UYBkhDN4oK/plO6roVj8+12VIsik851WgT+TWSkY49N+pnVG312JCDVig9Hhf9SoP3qo6l9N0U0s
SrHO+X+Nk/cwK3ok48NmBUT7O4KS7+8OtQzBgZdG2zIGHP3mcpqPNnnu7eckuSpB1aQ4gPd8lYp7
ZV+nNBh52hCcnvlqgMtAj7i0ltex3HMD2657MJHUkgh6l8KP7VhgLxr3ybW9BV3q5zI/TNmVlHZh
0LwoWIRs8dThNYCFcRfi7j2nt6UBUhJ+fKz7iYTZntJywLt3JH6z8I+vvsZDoDSur1xi1Lzoexc/
C8RiRwQwUEm8TTbolDtl0ZQMGIxnLc+1BUnC6hvcZ8S+ESPJTqxhEri/9IQ/kMgHCesjov5KEtvl
GJjC9TflJQEh8lKbRHyfEp8tlp0rVmFArSJ5nYGos2j/ZY8/S8njcM8yyhTo71qQ7kVlBuWx9wdJ
a0aauH6achFCnUaWSt/ojh8y4nybzW8/FKLBriKwZT24YtYabEkYxOegwIPOU1E26s9/hVs+obMt
kcBfjpfmRIapQ6UIHdH09JNBXa4QWBRXyTbBFSrWau7VruRji+eouG1oim2QXGquEzRLbOm+mXlX
L7g7TdRQYCi9x8Kwp9+s3qzBS4QnpqvNVh9ZIzUGZsmkXGBOmMJ92tE2/IBSjq2PM3u0Y5ueg756
gzIyNllKX20fi3wOdslAcMl4fZZ1D+tf4ION0hswBkG17jyTjFut9W263cKV/NxeFbVh22DrhwNk
rkGNONgyxGPs3cJV5RYDCToAJEaxXT/0rljoXsJmFQ+IQQWpISBDTgVIAymvcptHtqlO8kkDAoyn
AFNkR8ftUgWz5Ae0Z76I9Nl22jFZSBbdnSezJ4zcOTEuGbw1OpYI5FExK69/JuxVH6AF5DOotbHX
RB49jaMR6rAWJwfxrBhC+ba/VgNLsangNE9gqLP0tSmCLQ20MuOEhfud+u5I3+q3A7IASP+2VIlo
ea3sJrecLXXkGSrsWhvQrgNPeZGwQOezM32G53WjCtzMzL05MQ+f+Itcw3Lhew/5kmnQ1rUTTSIj
c1EGto/KWtlfZ2TqKqKM2ULrmyQblD3nJFZeWKBRx/HBP1H4XyTNjG5i59xFQI78lF2ltqVogBe2
Qdrmkm0jA3VVgjiBQeWz66wDwpNg5dMqr3Hl2SWzHiLihFViXh8i7v4TGWzsWAKHH8C99D951Wi9
lE4RvQsyHdzb1UE74xjdRlkH6Q/MbD0PjoPx/7xBjFrf2jGUd8vyIYOdPf/B+m6q6N7MQ7hOvsnn
FCSTr5dLiC/kijUd+IZpSW/wQ5EAl5awJIDgev3g8lbuOWqH/mrGgVzG92HgLVKECvcS8JsIx0qj
ItfbzLeI3HmNdFuijZFZwweeYkBHV+ia1pB7U1q74ZJBgrtGEszqlftYklBuiXnFwl1PLB4S2LJ3
W3S940ZnDEb4x03itVUs+9107vyAwmO7XgRwkYzfKW4B/t1I2F8AT6EwMRXKkoQOEXSCDvmVnIRA
hXkRKCESv6aj/nKCuNVQKJr+VwArbmJSeQro7Yahdbwuq7ZISbyaAUr4V5Nf+JTkHt1tbFJwBTzU
mLc1itsg7yxFwlOdQyNl55pW6mBerAgcP0RPW5vq0bddAQr3yFcpfbstjCmjt+6FSvzfVyltsgtw
WSZ4BJ59ulqQf/E4ivqPNtJmyvUbVOSkIK2SUffBJht/dAjVr4jClJoeJiRKzisurS0fvP1DTDL8
pbASI2UJNmx/h2r/9uF7Eku6gyTUQZonYMFaVe8X3yPonI/lE100F05Ko78u1htUqyzkOCV/kGEQ
N+VbBuPMTOicl87ktMUv9N3uZs2vU4dVhRLHPKZsh/Oolp8fSsa1pG0NQY2dCVfO43Ydi/ZtV069
LEOhsoGlYBLRzqkKxE9s+yJS1FeNfqKcWYTeYFOfsPYR9XJht6EZCwyTuGMjm79V2K4eMk1O7xuz
lfrrn+Ouj6NmmZ8kTPUpeP/R3Ki1tQR9lvBjCFwrglVXa6pcb7dzg2qJgPp6NPqYUYfDzkxyRNQF
dQdz9fOr5tqAewcxoVNGon0ALcCf+XVLGobINFEnN2uoobpN1b8IgPhJ2KCClUTTo9mgjqZpbjCD
vD4GhqaGwLdbpBSJkw8SIRV6SQcNKSULVctu0LmU0ZZuFgt63fFP28FneV441z2HYoSAobyhZsjt
z7u57cdaprismcrB7oboCISxLsRyMAxlfzZt6KZcqUPZv7DxAk6EI3e3JjxPTzsplTZD0komYnBZ
ffy37TqxXC7IEihuNAv3H1ZpCDF8YvQzHNMEEZO3ZsqerxEZcJrRCzXR+pwAkLYrEtJ42RmAe7Dz
08YwfnmVQkOEaQMn5EMqhLAns7EepgMiCi9mIsakGa/yRXA+1MsSO+3eJ6mdFvz6UJ3oEKEAO9w/
i6vTQyt68mFbKzo1Ij9oALF44I8oIbtpDogvprROo5imz9XlS1jPUevWZuO7yEwxfdgYu+6FTVKd
ToNNfQTu6az4oOwQppvh+RNOUKuGiOovalywrNhLGOguHtz1V8fUuYD/V1ccq5CCbEGupLNhoNRr
NkVVtRiIZ2nRcmp0YYwR/k+m+Qwxy41T4TFBpoSqFsIwfjkqNimAuu/7mwYUtbtgrZsmI0y4EHHS
DWmkYB4Z8ei32F5dVm3l/B/VzOSBGyUJvDk8HBK4zGai1RqSSUXXoux7LHyUuKmRPrjHPvkh2zbP
0KTkgmXxNb84d9KK47BfInJB33BSdo/WPRVx8OQTBUmwTo5ULsoVT+lieZZP1SRB8TmbbFdhWJy/
4QxWFm+n8Z5mRDx9yg/CTK198DQM2vfXzX+Wv5fDWu7UczjoR/XVY/PoCHzKr3DER/lQK62u3Atj
cgfTC42jd7a8SR7jwrrgMDc6D/1BiEehIgh1r26ilSKnVn7I9KSuIbDtScsbsbW2Duk72Uywmsxy
ur/pDHDVfPlTpwMdiUzKD1Q4LYPiJr4mQFMW5Wl30QMBSEOxfypL08G/pYn/DFg75KcmpQDCxBmd
AHIOyiY+pTN2z4rTTps2YoP3wLHPbfAA3q0WFUEZnkzqP2s1aHe+87tBA0gkfmN1pgGOCXiRj3Jx
q3bzPI/U/6owmxHUuJIzIRXn0Wj1hAByXrokIyKPFb37oPLcCLM8FeRVphac32Wu5SClYMknhe50
LKtddT0p9GT4A+PeHt3sUJVcAp2idmHx3rNKX1BTBr2XtJI9cmeKRGeSQsBzIsyrp5Fi0J9hvThG
Lw/FvVpAkkN7vx8d/5Dx7yz7RXPjjhW+ym17Xg8/WsXPhUPND58RldCpf4QePSfMEFAeTTed+tCx
aOdC6lnyka8Y+Up/78mC3yD9krNf5qP4R74TiCGqdTo4uBEGvMbvu89d/+mtXR/MsYhXoB1Nou3M
s9o5khzCe03BUbjbg4rUgTr8g8qtrWiS1ncrcIgHT8LNthSjMhOCJvCXK3VxuVAbsYe5tbqS1ZpU
kwFPjuEzAprrE6opPSZAr7orEXbkUpAZ/dLTg2MsI0VJh5LNgxO0LqHY0e89my5Kw8Njbxr+97t9
Hesh51hpOL/jahhOHuZRjr7ojc9uOMq6VjPgZN+7IVPHw74drN35qQD28n+JHhAVssyFzRnEHwbQ
NHK8wsbfazoaNxQEVgfBw6pQBltcsxL7oQ1dTu5ZpEpF3F1m3mnMkpH33kmf4LboEkSeRo0HOLQg
4IITiN3UFolTY5JpUif0v3LA+ruyKix1ldzczNwdtqMwAeKOkx9GzIDEu50jo01iq+wDIKKkRoZv
j1Egs+0nvrRtCQI3e3mVMK+7AWLXLjvJRyW+BSXfpSzmQc9knH4ACZ/2Huz5p+Q79T0UWrLVD7Aq
cxKfLaPlzOiivFnJ7TV3aJeuYwGpf26WprrGqOVA1x5CTqZktWQ9omKT/XuOxCDFuzVr3Bfet4+R
i2HKa52xsI7sOHOHq3f/KfTj6kry94wFWsb9cYvI4ZXVyl3Q1UXHvjUaNGE5kGgmiUaO3thl57ax
O7p3eBSsgPFqUsncn23GDXptDpE9Y4yUrtqM/LIqCXxMiWLm7Syb9fPYhcWgWb1aM4BWekYc3Cgs
bU1uREBlQxU2RKwxARxqd0na0rSx3v5KsRUWhPG7XdM/ZocqZnuW85kCU9gSla336h06Y852wqcD
dIhUfnPUpdYJqA6iwmKuOQUA+WiB4OB460yl4vPhlXXTcbVasQYX3t6ffjNOLnzALn93WLWNOiDG
RsdLjJeyXyT+x0Qpb6lVijP9JySZwKL7mn6z6jLqZRbMRV+pe46oKvmjTObcMx43Yfjp1w5Vmt8n
Yo07ad5mCgcnFDcqmPglo/QQ7A3VskjiYh/vj0mhy4xGdp8qpIkzaUhXZ5JMNk/IEQNLvBGXVPHa
1Y6IM0xRM+yd7K+uw5iefCS0TlrKHTS7euh42cHJ+JwTKa2A8jdyl79LWsgTH3Z/c0mrrKBqTxn1
06AxUuXoH+3RwGJUkXXaU73tdmTJgc0i5OF1oR86U1IuUi53B5UN/erWVX2K6911jr0q8F6W17BB
BYwDsbwRUSm3ddyOUCE1chh3LRevYXCCNhhb8Yk4rU4GZFli1IH7mG9x7StEXhFJy/ze3/2Q628F
bopiXvn+rDqzT0X1Z6RgMawg4v8FD6DoUDuXyBTyBYZMOi8yY1nHPE5mMOYpSqGxYSLp3SEFNaPb
vEz6mnnnxXp1dqtqF8U5wdbSiOK6AVPbGpKuHRMnJvXV/bGoJzxvQ5ZRvRUNxs7BEfrhpcqqvZd1
HYJxUlckQ4Jcf0Kqpoyfb/HZO/DEc8McokVOpDLaaMWNhHnVZSaxnJstM3JQlT8PflsnkCPApxP3
ESSxXXsawZoqWUi1yKbASxUdIHTkCDnU6fj8AxVcWnQAe22iZCImDHBMzGQvbqpTtdMjAr+Di8h6
sOzRkNgE6a3B2RuVqaR3ItRFOecWF/vUpoTLNfnjvg3yAS3B8iVzuMSVhd8gxtvBTE5EbkvbXwGs
fPWEnE9h5T6XWj1FckvlqR++5gQXwLCxzd8PRI0bV6M03rYOHyuK99RZE7a4KGmi+cR6Fssi2E64
9oKXzr5FSNevnkwRr/DrrXUWnqixBuShQWke2/TNa5Rq3MZUESuIGACKKwWE6v8ZXfNr+NEJojLn
SPAwn61hxoYzE+lIOMsxqmDfcbwHk1ryhGJeIfxSgylXUG2yswtuIsRDLBFyXlNPPCxsxo1NsyAp
07rsghkokNuUmVp7VlhKZ77+2b20opSFx4rj7Mh6hn9Ea3C7jzR8qA58+yGM/mLem6n8IbioL8D8
BIluyLfuBgtPkAG9+/Hh6dWbOT2hXfng3xbNB/UKnK6jBsarXB9iWw5TLmptlR2gHWYqdqEpfoEo
UB4YWUi63DGJ54OkdaxJgiQtOULH5LvfBK+E6vItM7ptRuc5sXdZrHYt4JlLHekXAh4YuXV/+5z1
rUKDWPLhZq4Mv6gRapLm1xRYDYfNL9he4/FncJKeX24wbiuJVpOkRRoey8XnpPtlCozF8efoKQEl
aXDMWaGjoZf5yrGmGweYEr0/azCiwoGVF6/7g3gcpkzkowcclWEmVuPaHxl+Ker5IYmd8dKAAk97
gomYHkV6ur0/jQpvfiDXPoT3kVDg2AYlqAd1LGV65C6TzJ0DzY+lHYmKLB19JMlIh4kv391a5AgN
Ze2yZbO/y/WqdAuv8/tcEd1sJmKOIgZDfd+LwYS07LH3OCTW19Ivjt+dlwzfyb9MZv4l5Hy/1Tu0
cjuX7E1GSk4aGGltkCGekrkGRVrkwnOc5cRL06RrG0hNEmCna4KwR1lNfRJ4sqnLV9U4mxTIWWE1
ZoCKQeWVx6QJHL2ihHRfvSUvxQT4NrPz9zMusclh8xk45z8GNSCcFie3fCOwHVm+dfxR7GAaen1T
QLlxoX8pbqu7z1Vm8CxIRvAkJAj1EguamMDZDMNoxWnwzlq2Yz0yKYl6Gh44a3moOELeVW0HY4S3
0Q/vDSkG3AQ67DhSbaB5ec0eZfVOW+hvYccfsptEFkkWOnKnhtFS+UesfCtfI0QhOq+1E2d2jOxx
Jo0yBwC2hdrz96tIiA78QqiMdktrlAZ0PcBT8a87bfYAjWuXKsQogCkX2h9/gfv3Gyg0Vq6r4BFH
D3vBM/odNVEyJtMp+6QTnRFZ2HNpwHtnks3z4DmzrgBkGNxZ0V9Q2FPSHbf4YH3eeJkBmo/VeWvw
Jh7q4l822Odh0O0++/aDwUPX2Bx9v7F6BxilhLjTg7nUSxrKrm759OgAf8LlR6yeyUHtAXj9//m1
/G1nk60QSDDqFU/204rljSthU+msUPoVG44N0LcQr/M7OUqtjX/+d6mSRR2Gb1MKH8T/qXFLzS5e
fVESFHHtRh1Cf3bHMga+m4Rx5hlSabKxblyM8175/oYZFYQpAKK6Fh9tsX9b527sBHpHlRh/h0ca
Qo6zK4gitC0xd8LmA34h/CXEEk7LTBT0Fr1orCE4lxLbPoImJR20yjJPJ8JHKfj2ukVbcAEgg5Ls
Hl+vqsg2nYZZWsJE0QLoLycVGon96dml6wAzeXZH0oY5NNsEGRqg7lfsKo/ZtXNs/jPumpOJb/Ko
aLlHyScVbqDDR74By5DgFW77YuoFynzeS3HXwvFJ7s4U0rg3FvXQhXLRktNCqza+fLI1AVlmZHia
tLdo55gWR8mJp3fvT3f6Y895+zHJ0yUqNV5abQeJ4FEhXmk0IrWwn3biJ0K/vfv6gIgt3qTvMHRu
HYGK6bpK4tOdzYhTKv/drKI8O3i2oD/mbxZUrNCZt/w6JUc1v/u5m4kz4w4BaBb4Z+FrauGhGiu2
qlC0ySB2WoaNqLE2Gf5mrGurPbpbJspk8B6OnDVwp7SM96IxtdH5Vge3nQxd8ZJAQqalj0a5UKPW
/Wdzr2062Qb4oOQYDzTx8pOh5p9J1CgoU6HhvpbQ3h/w+lVpanavm/xA4717kzqXG+aeQp25ewZd
EyuLEs5QEdeACvjbcdqxqXdTEiV70yoKcgv09eIHqsvgeEiwJS5LXF1Dtfx7EJQYgjKHnIiC5Z45
W837DDQ9TL/1ilBzlZ7WqNhmqp/PLxgFILJ5d+J/pjJkMZz1qVsTEeAAZx5x1wiqvSD/doec3VAu
VM2Exak7hOBWuBkWSRYgWU44w5HEkYOShbWpnl3U0z0ah5csmWDriwnTqCHAg5z9O9QKT0xkZ09x
bHkIh0WoVnJAZ78QymUXEU1cQIV6n+ZpqnbA+13zgEibmkayRDdHFPE8nsXB8IXDMLJxih/wiDdq
e9c4Bf5LL5iLj/Ck/EhF2N4djItsvATSgFpMD/bzynKdeqjpnX7sRWIiLbl/TnB4pdO/S8ls8HJa
CIlJN6ptfgtHWAYsMildWRrZtbVGaJ+6wHV+yrNHdTiXVL4aVnYHYyEd6l5p+kUPIxLuo+QI7X+Y
aE6O04+Ofrgysr0JV9wZ6Xi2ZtcHi9ZdB1RjlUc2zHeMh0hjUig+tRcVtVIY6RprPZainU6uns2S
xPpWzFNdpQEyWUHOhDdD/BVbuYyKScEqVwNRnKmJbd8daepHW0hXF7Oar1GgC52zYfliwbB0Nn0Q
o9/iZnL3FgchgEbJgnguvMFOZyROS8Gc6bjFmFsD7Cytb2V4SjoArFIrfRaKFnpvpo+2RYtIyA8s
k+Yyft5WdZgcUuYd+6aDMxRORwKiplBigNCavMvYodhpr85pBUQWmQc7XSODsJvP76Ozjq3w9Eee
vI3IAxAdkmtdn4rYeR9AYkc3uaqsAyBU3cLBE40XzMUhctIZsQLgUCJtCseyITpTO5JXBJnXeTEn
Kzzz2S+FHOPtSl5YaSU8Pn1lcOt1LzFy+/wyuq9m1d+N+RqsxA8fl/fWxhRb1udBndUG/ZAyXd1z
oz1F77OAr0EsmfIhN6dyPX2YaFpl0bhW7XsvL9CO1d1uoZt518HZMlTI6todHYwLQCGdCLBaWRf5
H3//WoC5RaDtPRrQCikgEjVT87IIfT2lza51g+AfjCTFhmSN0dgAoVFe1fybUs1jHlNrhYkNZqXz
b6x7QwyhVjQ0Saq+q5UGzqfYj1Wyhvx+PJGDpDP2mLzrsJYF+lx1WotFh19mtf3o19SaeC4EGGG0
A6SGxTNpS8hPQbKu+bWT2MMIBeDcHlcujNP85RULz0GoJoJ4KfDoBQ+6Wii5qWlV5sVm36735W/4
FOhW5V8F3H/WWpymV2vsYcJClxLqkaPGmZWQe3qsmc3kwDnfa8DxrxKLqVtZ2ky+NB1KXPuxPeJi
XVCa2eBAVmU8QOfZDjAgJLwfxQuyY9BTod4hthJ96Ck477Pa1NzhyhGJLqwDrGw9SBexKRfkyXTh
O7GODLdR/xTtzsZQ+YXGc/5pdKjq7/frnT718uv/LuSb+qlNR3rj/cwZFi4LP80MZrxkgh8pE1dz
4MNdf8tLzm1KMgT/3EmwGNjSmHYxr85rlepMbaZsM7WPlZ8Lm93SIw3BVGq7YvsvVcNqUTha8nm/
bW5ccHXc8YyynmsmIAm6pLs6kBgFsaOeX41MfpzviSqy67FNqb7UJxyHeJCW+9BzfxBX1Iw3Ykwt
a7hHPVCHsqKP47QwfN+R4yXf5+fiPys/w5UDATaJthRgktPFlLHx/ycH78ru3CEKUHh2Hbz/ZwEP
Tq3aQ3Z+rTKMG7pNnZEFPY9RQ6M3fzElYL1deExJF1PDEyP60ru4tWpKrSa9AJXCxOcfukZpjgIu
PwiON6qm3+Gc5zg4yxzyp5/RW1sBX0/G4Ibi+e/UuD/KkJeMKUxy1JSXoDfBrOin+ZIjb7z3xnDD
OX/ebK3XhSpbBIZdo/cvoNUGxLRnrkh9teF80nFFEnDazU+beQe4WarZiPfOLXa/7OxLYjv8foVP
omDZblMNBKbG1wguRAot3Uf4MuSfB38GPiQWZlF+j8vXING45ehnZD142HKWUAnPAX8YkSERNTlM
jKaktolwAv6uZ1p14LdHnPGA8DzkZJ88IoSlc4k3AINXBLZSaplh4HDDuj2kTxhdLoihQaSuTWN7
0Uc+oT7SqRAfBhmQKVfMA+1/ma5JuyTP4HeRAMV5ByyWIr1yiMDGWGPPaWlZsCRa71RiXgXz5Zwb
TKqI/lYTB8WSFufA8aloLQS+3ZArCsLYtQgyqCzgtX/ofQVg+yYKOunEkQTsZgTlY8cNdm2SXx6h
6Dzksfaxui1IsA6Cpqgct5Npz2SbVcbQHscbYkTD0Gg4CB4fun+3wfigdTvfM48f7pFt2KsKsMtR
0fw56+dREsU7JPqcuAGaBCqDrHajqai0OOpziMptE5HqmqLHvc+t96MltKRoZO7c6MGGew+sCcb7
x+KQ0psp7l729sOAKGcRgMeSjpBcTR5uIQz+1eeSeizN1KxYWlZm1J5BxynSEk8k6XfAstQzFLmn
efha9HVA7ZzT6khw6cWSdklU5MhHJWFA+QPyDLrSTD2wk7a/ZzLoagex9zi5qIS/Po3FoS3Qqhhu
9mxdnzoaA4r4/vfr/2DAGnCQz90iG/D0rHFjdnpjDmsYXJFsAto+sI0PxfbgXL+cLNMXFGNMR80S
qaMoipNW/+0yYAEUlJ0sdM/g1QYXDYBlmCKuykiEHpAPzpU0p/YyUzDkhvtWGCBLQ0MjVgOaHlC5
bcZPKJdF29y7RVFtQGm3Jj3DfeES9a9wMwqRSjxrar2kGZNBAjTGMle/qIlD3PhX256OOiNGM340
c0BigeFI8JdvRKzcUw+B4KZuYs44x0atNvtWnR/O3c2096y0fpybCNWhZvmGNE+FCNmQDKmDBSwI
NiZmegBViYR++hifvrkpKQn7PKtDwhSmb2dp3vsEzJ5xVbLWFKX56fdclJlRg2ghTCMqrH5jqEHI
A7YKP+aXSxklS94HhH/nBqhbAVOskYgnfpgwZzSNg9E3JQpi1/6tU9df6x1Wwl2bYiFavJRSi+w+
gs/V6VLxinCzYQ00fpgIqrM4I2oO6YrkZTO+HM5twD5K+V/SW2lbBhMagU2CG1K9KMG955wLlzSw
b+hFMYthz7RX8oMpvRCPkwLyR9VWJOgQBXCmkjiOURWeVVMHjnvdPaEkQQTlDJ0ds9K3h8IAzkje
mDOF3J2qA3NFTokhKTzexFf3KrpkBZkQRZd8qQ8xDovKr3qmmcSiRmKVo4dJjdI9dJfE+d9v7Y0g
xqyW7Q0IhUCRfDduOfWBnf05ir5nZdpl2Hi/lTwNw+JegNiuMw7/o+IaobXRyD8IgE1OvFRC+vjO
QYt85kg+8Dmc8Ud2G0Tn5qjduqRPmfDWOs5IYLgOYQfQZjbuNG4MWz859glkhqokauM2ggox3qXy
tlpJZVB7zIHY4F8ffHbKQkGlVxsIZLw8lgsuumzOszzCPEslVWtXaK1zGiM2zz/BkSM7Wolk/x8N
Qwm5yLhZkYv8Q+EuBoZdfNnDdvrxJAuW2RD0IcATcbo7ZICvnHOZaQk3b2+eDEFo9U6pq9CWWxa4
kW87i243bS8wUiwDId09YDLy7w8dfmJd9bad3Y+TauCX/HhnniTeH3ReG0RQKBb+BsLWKlixJSpv
2I+Ui9jsjl6SmHy6LUVv974gcU4zQPYTN9mEKV04RYOZbZhfmv9DDVU2U2WXOdY1ROSP1b3Uheg9
/pUbN2lKjKqBcSLjL/bsBSraHUCL0j69v5SttrEBwmr9qmEzxdaqZJd3BoNpQO9F0iLKqTNWg2cd
J6vegvPx+YLJIDY+59LwOOua8SY8qqfXpfIeu+bv0/7SyBqhfmQzdjdzg8GKxr+QXkVRqHDfnDLf
5p7skVG0+ltQ9gcUQfUFqt12BxiakAhh2fRlDvIfH/mPZ1u2eb23TdqAvs2MZU0kOOVlOiZfsQ9G
W9KaOglvnEdJiL0+JGX6k4W/rPYuK+PNmZ0QRBiJCwOlS/g2n8CPt9zzAe9NlBKowR3hVblK81Gn
Li5O+ESJRWRq4hwfXP3iKVvAXdRJfFjS7y1Cc9fOH4m/GgGttSty0AhbvY/e5ERTypzT9e/z2cyZ
F5NQmpyajWYtmV3CqLMJuy1tu4q4aCXDQ6pPCGKOk2QCx4EhSfmhbAB+fOD5XTCMBJB74q4SrIXJ
XGLjasJ2+Kp6zDsFXWDkae2/WhlpFyHNOdVf/+JPft2c7RPX5CaaUyIMzwuycvzfDF6F5Ro+o+aZ
ol66joYn9U9TX/XWLM5Fef1HtDgAdK5er9gqk2YoP7IlaZfXolncZbnRplbdKT03TrCe+pRpeLDJ
Lo2A2QYuLJGSBTVrcdF+gr3FMiQzIV0ZFHGoV9hx14h5Pb1+MfJtx/7veqP83Hg5N/IOVtU0xKrz
hyT9hOFfeypOAplQUeDOB++kFysJ/x4jWVSN2P2RZ18yF26W6gBI0IpDpCA+Uhkt4lE4Rm9qeaXG
LMRnJOB2OROyQtiQqvcmCrAgdO48GfFfP1ejMqRYhXlWYHMTxO6voMcpP96a1ZTLSWJwXec96OD0
nscf+Pi6UwjGO9Fp6hxoUzV3hy6QrtEa21lUmS8wiHtkj82Q2AqcYy/WKAxDp2j8Fu4Lk8Td16Js
9qPzEsvEj+4pDmLhKrkuP8WxCvjUPXIp86hj8rloE2HTmvdy0EyQ4SArhpqoxIIHr2ENLXsKk3jt
kLiUiY8QVQXvtLThno5u4vxaxw4eDIdTWsx+J6NtamwaJX5ByPzc64BVgQl2ghbm9XdKZaP04PDB
26ZsQSRL0CzWwxowkGB59G+N5ReMQRFVX0XnHO6CK7oGyJHZ14G7zx0sxt17niOZ61C5pVyHRMby
UsdhajhV6XgptpY4LHPZhxoh2lj+QrBLFzqhSLccakFeO2H/y4AlQIS8G5/e/hdU0UsHlT/SaCsa
iJxygJbwuh8SMdO7IRhaKCOAf6XCyyAYMuA64Ubzno055IHKGAAnzy1PMfjAjisGJesbA8O2d6hg
nfVXGjCo+CmtPsSeCTUkDgr6jHhYHRRPtg+hC4x1w26jL/tXo1fVEH1sTakOgA4BXHSML6Bt2AAj
IDth3pQISPRmBQ8d9a2rbowwRFnaCx9bQ800Ud1+K1U3mK6iwA0QYhJxwhEqHeyS6s3WfNptXh0c
rsS7KArKuAtzEw0uIEMpO2Hrcayfjk7AxNke0f6Jm8xD+975DPyYU7zQ8CdaLl+NijmEJgi8MES1
d5ym4KUD+3pedcqanwXBwU3ec4kxU37mNIQx8uVXaCt4Y2rT4Kx/e0VmnwmSeEitLqpez1a+EFZ/
PT4e7Hp6Toa/W1W590U5RXLGWh4+hMsFzDItDr1wJ8R8DlFtXAGuqTSZb9zcbwbgcDsjMDP6cxTJ
olFhBQ9TLtvEjjHvrbbXVM/Vn+9KQxuLzpdGPeOZNQt9zsZen7M0HnGrwa5WxEux30EswLycUspw
shZE24jlQOPZTl+7gMv6knuTSqMq2STMJmBscQfSwbcWyIsLM0SIN9V5UsxG+N7R/bjY+PeT5xB5
ooV93/EvK7jjPuGlNQFLci4buWtB1CSl/g+dpcAfeKEK306WkR6u1L3BKoFFHqDFLMTGuITNX/n8
ti8thg4JiUIx9HWys/QU85UBDkiuIYuTKnRFJzzjpgVZEnMyPXsAt1TQIBukSChbnuTjXLB88stE
2gD17oPlamyffNpXRevIWN9G6cW0ohWixJq1o8IluWbQxsY2b8SthXHZjSldoNU9d4M7iAxaJ4gJ
iqrpgnHnSzpkRwP/Pa64d0bOOR0ELEwP4MYB+r379dpkXvu3hY84CYaTJP3Py/tvtWRNlWO63SKZ
iW274QlVcjoMWyiTUhcHNUIqQaJ6l/6eVQWrTCIbQhExJYwpjdCCeBMqqV07gzaY4qvmIHRmp0LK
UayWUWVXl7kzrnVEPFJSTTt+TFYeRudM3j8QEMDc8LyzTNl3N5O+nq3mJQyM6ZPjU3JSZf55ksNN
rBm19pe0yfWdv0wRNsR6d58GZ1JFXvaUOT2CDaitLOQbOrhHLHLCs/6TMH8IwKt+eaZrGBIfG5JR
caojiUdhrIShMXBrMIjGOhi++EwW9TrY0Q5eFFAyu3BxvjYyV3N7CCPjlxiUMvGHzIGNPWklOHTH
5F5RGE7MhMiUqF8M3AQi/EEGis7SZl5+uoXlIs/E6PWRwZvfy1h2e4kvE6mJzIJ52se10Ll4lf8E
wnz+vvfxcZm+u+60ktT6XvH3qHOCVu5oxSXA3czfE9Td81NOuBvYmjHuqiW2BqxQreq51HGVFoqb
X819yDl9YHV2Bms0M7AZpSz7AT+2p/cbeLnvpAJEf7loLoi2QtGq1E/0rjVlD+LT86cHBG/YDtun
3LURa/MOSiWp9PfwiwIknFfRl2ubc88jrvNuEkKZFwjbWQNUCbKYUl5rpvpnyOnbYEZYEG0McdlX
0TKUdnUOIdXHByywqGPC/lYAFb7Ggz/bUh/ezrEbE+GgtzMUfdKECBwsd+rb0iyQj+t5bSyQlJVe
7QCd+MmwfNVQMzzauMB+3FYgNA3a5rBFhgh2DQpPmZB5vRuNHk14pp98N5wFOkNdkU+pST1RHXlF
UAT6f6LhM3h767ZRIfC6CcUcr6FLbVJc5GX4SYepAtWfS8wd9KX6FZ0D0Ds5Pgjvp1IjUb0PzTQb
whe9dDW3dWvdXarv4b9ooEBPnTTeMpdVK4hS5hFj3EdpzotYfGbjmZ9Ese1dC/HitiJ9aIEyyvzp
4PIhjNRadywSDDEdFo2VS+nl7RYS2moWPQezSbvPnA/fXSwf01bBLsj1efJMmwQWKJpXZ5487Db0
qUu01VIWOAYprHBG2qn3PpBRLNBYtmz4DqIfLqa4fqWbDWHzSD1mkIYHV66CAyVdMtN1ZLpoROMn
PhkUJx3P+NoW8ItPZIRaPdPC4pE0iPlFq8HDzMRrgwF4qenTu/Qmv/siFL6ABXFk//dzkloKj72z
QFCLwwuNLEIos2s/LiQAYQMAlOWKgcfu4QRCCH59O9hqFXGHJscT2gcr5uK1knKu4CbvP0gYwJxz
dCo7lItsSF72obGjDH+sGQPvS3f0NZpeSqxf4OTadmGW1mzCDVTpdZG87HKyXuTZN77QkNwi2gVp
tUI+5mG1rMSUtASA9IaLMLmNj5BvmsLT2LNLrSFkcGsP+muANr6sk8+xjf525Bd2DqSraOz8VA/k
QXPjwLB9MBTraX7ugHgnQ2i+wqzQFGpe5459FD0xatGguxq/XC19kwMRIhCS2l54xPENq0vZlPnh
hDcZbXUGOZvRxUMN/jBBKwymuhpxjzte/ja/9o9ZZnGQAQtLL1QIiwJ2y3AN0p4bGcJOIKZj1JzG
DDpIa2LVwkn/6yz+JXl6bxm2Vumox5czMbeqqLKJHeFKk8QDUoaI+ObcOWFSSbUEKHrSPA/x62+p
PxqsfLkvazTvq4nNGSvLJ1Zn2arUhNvxRn2Rx+zkdj6jVM7VVe0BNfsVIvGR8uRMdud8XE7UpTb0
EXkQFttN3IrBlL6YQNy9ys/5DiyrONTQdyMo/U4y58EwZXguUNcYdxl6lRvEhX9NC8ykQqByhGUD
yzFrbbXu+Mu8d9lVxscOmwL7uhOXNRu8VXA2ZHShjxCa+FqyM4LcwUkhlHu4abOzFsnVxtb5WgPa
gHNKBSsIFCeMNWO1Rcm8f0HVUceB+s33wkxCmO13MIyaKwPqTIrX/VqkdSq0zkPJxFgzZP+X6SUa
Z2hnxpPAU8PPAQ6nAfAmaOWQOL15ZGIOyjizCTV+t6zRmXOKqnfBZchvvzrq/nUBbfxLgeIddddV
H+YcQbLkVzjBd5kNqJK3iuBOex20qcYdufETKcNNYAW6Yl8iwXHZKL1X+BK6UHO1OZfDGKzBv4gR
ZSjLJG3dzsMkZIbpLMyROHpL19PPI5TEyzzvHZNSGsDBG7svnV8mS61ZGRpDz29rhKy1MNFspx9m
Sccy+WbcoDXnaAL6OdfnIgr203wf4Vjpz0c3riFBp1Gx2oxFpk/gObIgvd6vTPxecZWcCpQqpG33
nAjdy2tzvhRQ0MX0flhW1l2pJ2QewZrALtxfpnk24z6EvPbfl7QctOziivndgcuRNyMJOt4A2VRk
7Bppqv9OVN0Vvrq/6VCxeLGgHHwsB0ffJEBQo2rswqh42imszaeA3ivQOIl7sWbVX0AFlKtn2c47
MMurJA5i+0qpNpeLXthpPahfCHDoGVknRzOd0WBPmu/q5RWNt6Y7YisohcD8YTX6qXgn+tD0T5iB
2Q8JquPC8vQu+axhyOGoTBPMZt2FNlz89/om7a9qA5LvqCKS3ME8D0VZxm8XXDWoznuekkbjw0Si
FKSjE4nqgLOpAJpYxBOP7dE1FNK7Yl11d/2su/8LqCIj99NVkHldhOGCCS3wOefdLyo6hHowzkks
IJ4ow9CSATmFqJScEERh0/334syXAsp6xvfVMqDwi3IUaqxbouTRvilxbDDoRge1KzgWMyPjdW/v
B5+35S9z7R75INtMblt7qd3Cv5Rh5TtLYyAQp/z8MQqhovtxve2qOixZnDfjixY5wUXnPDI88af4
Two/5rN/9vztNRQtHvaYJBdDgM9E2nF5tATZKZ0/SN6Fw8/vASzEkJtudZRzSKSXxNZoAlvOuDkL
+R0tqmmQmzV/nsV0rfnVRJpNgZjZiwEwwsr6q0iOjkDeyObK+Oe7eB+69Nq0vTC35he7hC82wKw8
uB1D97ydmIia2G0YWCo/mOM7+3+lhgUhsnhB2NEBw/BRianK3Ny3SODILDv4oGYlAy5+PTCXXFVb
5KLEfHPPiIgTOh3TT2CHpLgHtTljHekZJu+Uq3I7dc0ECFaaiH4QlzEfP54XEvmO3vtm9JXxs9wj
efuBzVTbSA+jFH9B+0WyOw/oiadeEkzv6PJN+0JNl/Jy2xIXsAH47gcKsSYfO0o/J27g2hnQz6eC
vCARDdI6qslQD8ukAVPCnKQZ6wIY/lZIVEdYX9MsTUGy4O0RvewfDqRQ5Na3BtGrXiyAJeeK3pm+
Ln/EKCTofTI3hLulH4O4T4QbDN7E2vRwy91xkf1xqtpBXzRpABJgzNuyBqJtCvFg/XSYAPASCtpx
/eqqf30RtItJ+xdgzcuxPYnyM+GcHQID++74RmRO2UvA48ubS3caVNqF6LqexM1wNpv3JMKZtWL5
gV5AHBR2i21ZdVe09QAd4amMZqZ4WjL62YAEv68SCZhDFxc7f01rVIm9RyklriGc4k3ncgUrQOZv
c5G9Wo0/y6JHGvi8d7V2NQ/L3ZrISA2QtK6HB2Mk8mSK+I2SkALtN2DjwfxYg5jEzBf3w0NHIO0k
dE3dIAJwSExm0HiRddz/wCuENE19r2CPxBEK/D7gmrBoBVPPnHlyn/rIOkcYFY1JWoqxV1ivTI+w
rgMTPs/3m/QV4GKg0OtM7y5GWDDoKrZQLX9xvuEPwGErT66xNY+ywIPtC5TaTs0tP15bjDpltFD4
KHFyt4cg/QKszUSMvwqqUcFnovpAbLzcekYAXYy/cPnWVaGh88XXBYnJc1CZG6iCSMyI196sFcdH
eIuOJYKhPHhTFye+VpQaR1QTQh0NuEK0yY6j1e4WRv4x0ebQGDsi1to4bKDQLJYx6hrM0Xqu+062
2GFWpufBlODiFnO4a/qdF0/vj6ER+jbxMLDOvl2bAgW/1e4ycSph40nXFiuR7GMnnkjQdhjqYvDd
XLNIIbv0tVDPRsX9SSUgkrGzXDqg61ZpsdnBXzGeFTosmwQGy31Ji9ZoCZHQTVPRx1VkAr9vFMq+
fE5eFZCGSjvJR8ZtBpuhXk7W/o/1npEXSOkyU3c3dq3G8T85wWNGV/bKCl0BcGBgQq8jGVtx/Sl3
yFbPMxHNU32rpSxoRF4+F895DWvDGPrmtpZW6pn6dBrS4orTR5EtjNFNYwIIulQwWIUPEOI7NNqN
E0PMb8yyqyERE2+iSYfSyjVwOVBKGoYO7shsEbkKzhzo9AvEC6ZZ6DZ9sRkYPWyurC6iMde08ppl
Uw8BeGtULCz1LQqGYW/CcKC/9dMiiOeg9YlPJG+AokNW4U6wYFCwItV3XO7sFClexVGOGxJeoKEg
WdESNsdkgbr1r+0e/rbYpgSgFL+kqPuP9FkUe6eTYslvyH345A9eqDZM/SbOZagK7gN5aSanbMhX
1AINOC2lm3YionX1PucO8XDxj+mnB6OKbXb2AmU6BNZz0acPmoVMGkF6KCOhy/t/1Z+JzZHuOqQ/
+Iuyb14XzjS8H11KnG6Ruvzvi0OwnwfTWldFvSAAYCfVoNlY9/bCJQ1D/cZGY/8Rnu1xA5ldSPSL
RKz6YJMrshwAXpgQZHlNMb1VS3gFBfTsxYFp4iF6btBLrhi/BDZ5KOL2reylFhwkjGM0Hin/2lAg
PynQ7QP75Mco+p7u7NiWWgr7SYLO3PMGBgCO4acavbd1jCAnxwnzbzzSPyFVEPDgRr/nuwpNiGUD
/46MKdnVs1NiNjGdKqJCBZm6k251VVDagC3MmtK3BneCCEs7E0bSN+b9CiR1/QBnGZeFV/SiYMf8
r89nWUPU/UUgqU4Zj0PDg/y6sPC9cjYILsFzoQW9KhZLzq4i06DGoDBtcGEjv3PMzojCxqELU8PI
RQrpl7ryVF8+Ti+h/goH0Xf2QbN0t2zedm09RjD2AjLQRZwBAENu6sMpJOn1tgN9W0fOtyiHt4/p
jk2qCg31S7LOR5WvYt7leQyv13fYH9iJ7goIm5eB2wtptklGaDcERL1IFJcZX5KIBZJuhnftBqCr
ZHIkHxR0yRmw12LiBwZb0/44Nt5fLwtcu/Ikr1CUUORBGN7cxkISpbHgorBUqnTnDTWl/FileKml
mbtzd4JZiOP7/GWYXLbJVnH3VY9BPvxEdTC7qInMlZzCeOP2Ejm/aKTgdKitOwKdp1cGPdRDHqiF
XFpHdNhUMmp4MpXGW9hZgXyMLlD535WKzAZi7A/mTQPgd5b4if9Z55fjkkNMs3IuIgQnfn+hS69S
S97WFs4KQdR8Vrjse69f5tvfAC17FkKQ8qeVqRy7CGTv2+M539B1UQ124sCtdJ0ViTATfKbiSDPt
9ambOkY4N9rYNH8Oja07T1IS69HCmXvswAOqJRG/9LLWk2b45asg8A1CvBUY1uD61+2p/sGgtVQy
a/XnRu2Sez8VNMJPdB1fIdroMjrlIQf8dOQ7iLwVEsUFDPmYYdf1d3gKKlS25SWrl2/1Qs3/+Dtr
EHJLXVNWxj5mc1sewbdt63yecfrC/tQmoanZaVo51TAdH5bL1Da3SWcRiDe57QBNJ1h/uqyfYxtB
rDyux7X0Ob9I5m1Wj0ZZt6vfXiLF8WQ0v83lZipOWCunYTkPTECT8G73qQ6rmjT2caXkgwJkWZ8T
wMqlFmGB0Rz0+52HzHr2k7VyZF7R/fWa7MrKfznNCmH/dIinsDBACKJ4IK1t518oh15lhumRiMyI
kWrjMdwOBGbli/rxy6IHHBN6Vj9krdLrJM9KW0wTwAhLDZJAFqDDmCvQnPrplOdW+AGYtFjQJe5M
5gpwHrdxXcbrtoytw3oDLyaAGsTx65ya8mK1eMaFsm5vJ3wQ7KPR/SxhHLQqOOmCIHl+qqj/N+4O
q9036XG1EWipgWHZnAVbnupy4fOfhnb5BT9t6xAYzXdwS0GYmat/jxbBP0mQ2hKj8FyT3iZzgv59
bkezr+O+HQG7BG86JZki32mLpCTaDrbNRSwJpYzaZYFd4zt8kccu8kp0Ty+Qyug0oYBfVpskhPVO
Nffd882QHNdWXOb/BveOlrVjLDv0O/vJTDyP8Ms45dIj1HOLwzUrFtbgbQyyhn4LJ9m1/rUCcU+V
U2fJoD/uwKCIU8ezpBwxD+tQpVY/2HCMbq9myFcZV3xXNcHT5ZC2j8q+gGhqIDXvlolsnWgNuadm
IbQ4IkD3PDWVqOkVdz1s4Ka0HJrdFeVNew5EvAIusVOivlTdHBIBBIoD0pL4sys7Z4WbbBFUtfvE
RPfViZaoPltP574UbLMoJqjVLOGzlXmdXSHL5vbzjZpr2s2hwnRdE2veGBVJsmnJ3TNex+gPTaH5
+AR0Ibc0y/ORF6rUkSuLNdM+V5qHGbVnyhdVelNIRFH7Qv2BnaK4YxVxa39IulOIxD81nh+8HCti
efyvma6To2DlyI6bXg4d1xyPfUJPwguJ/ij6TxGVavQ2k/h+TtVGFmvCfgD/nUwO1x18ydOM1fL1
ucinOQYEFuCYE2miygvhWe1LydzSCm2R3pVALGOxOGuqS0dXTDFTcwYZhslmCPMzC9qdj27yQ34E
Tdp6Cp/DXO0LqqCV25yNP49KqqtHHEL8wW6zrFyX7D1utOvB9n5V7XvasyCkKg9SFhR8qzkfUMWm
gdgS/ypfy23apXLii8TdissxwY0sck3HzSnrM+Nd80HqQroYofngN2jtogSAxJEEilgfKq8Ly5q5
FFNi/6b9kVdn5Bl3vvNy1joQyDKuPWsUjEKWUd+JEXbNUMaOg1Z1+JepskQIz4yoMrhLHg8CU31L
LIxFCppA1yYFkmBhBVKbpGEhlf7dvCH9M8SF4PeWxgM2tb8LVVn5lU9Ccn9GAGwQ3Ly6xHpTJdF6
HDxtJblbMQxwlYnn3k0g290xr4+TPpEzAuqVpbtXz1FNxc5rNJ+aM1OD3OnIlFGQQOIkVRCPp9HQ
L8fTgFfINbEEpExpukWK9bKDBRDbyEpjZvNb2aBuA5Eb3d5BPTlDMOCnTPNVyBhM+xvZZ4wUfwRo
sfjl3lqqUGUs+G8yBYfCFtFd6X5fk/wSCEnwV++PIbSDpRuO1sMdz73+G9YyFRGZwTtxzijtrSwv
jXh/aLWwCuJBr8HOCtnlL1V5Tl+uof5F5Aq63estKFUOhCEhSlB2Oyla8grH/b0eYN/gqmkWISmK
ILxmidOkDvvhn/OoVZlKxzZf7Kb+Af5rF/dgaGYQXO7i4UTOun+57ssPzmjnkcYtIdnQeNoQw6O8
kvN7RKpg8o6jcbVzenXUhyjuEE8GRdZju4HWIlRLANOavJKGYUPVS3qJi1zjODXxK3002cmR7G4K
wTY3MmaqSo4NWQfpKKSGcrcfaspx+Bo6aRYk98Wgbs+pF0WPzL9MDwy8bCKA5LQPikCASdvoruWS
+rRs1lAlsOK1yKVlfCCAfV0NeKpZZgVHWZ9GZUhk3ovxCYpP/8JeN8Yi5lqrVK2Bkpkrcb4v5kjw
eXG8RMbdzRT3COGmjkUNcPXUANJj/v+wxINL01lMZmWc3YNk0vkLoPLMrWARwLTeIgOTV87lJJuM
PVFhZaQg+fHVa9Ih0vsxmSQXtxFsI8mKSNh6Zu06mLpJLr9/AQkvBiYdILjiBhvi9siomh+l0RvI
Ra2YQwLmf7IvGgmAvBkuAbxwU1V61SE3q8je9HtnlApVKfuoo3FEMEiyYfEq81DgDqGwb5kSa0yE
FAd93XoZP0h9V+UgHnc51wNijm5TRvzXi1TOAUX7PCmag4YCTnBjP+8t//ovi5Q3ZUuHkjhYGTSq
xcBUyn0xpdfKYAgBsBlSGGolfDPD3fI6DRH4vTaW8CGraXqV1yLIY+/4aUawDIcn35HBteqwROQL
HdHKM+vFtq6i9d4heEBpi9NH1lrT+c5BZXY2JBWwfaVzuaze7xG8O2QOV8dDKrk3fAPWKWoX65kE
edjUtUh9Gft6QPT3AWxyqUZXXr60I8ja4MUgbbHF/XXgEA4eEU1ButZ8y7/pZQACCZYckgpXH//s
ePJr7imO44HBH9itJua9c8VW1kxnVV1GsitN9yMMpEyJzYV2UFjaORAzRWQTQ3SkeJCfQmy2p8fq
3jyk/P3czh60sROtnQ9QH4fed2rD6vNYjuPDMhUog+XMyoJy/gLfjVzFM1lh/pYUnYwtAl0/Hy2I
hjhiYWA0LSCASu4t5Vl3F/xSqDKIZxHHagl9g49hF36lB86UXzgRwUVBQv6zZzN6xV/Mc8hfpyv8
qkzSX22wA13lu2C+brFYSlggfnKEjNET5Sv+dRDh/DzyBpS0my1RHj7u93tOo+8jHimP1pNITp3L
DWOuxOZIy6DgqbP5QpWHGRjhANdnJmNNe6eZXE4sDBaE92luBF4Ty8zfAgDiTy3azbOniAUAWq2N
l/8605aloh35z2LA9C2DlXhTnQwAG3vtTur6DjAoWIYn2sgOEnl97QKRR0MlYDzNzpbP0VnhqBMN
8Oe3zBkylV6WTSJMshK0Hku5Ka7PeS9TU63W08bVgPAPMyMAnRGSaUScZVdLCk+3/fql8Y/ntjmw
y5y8dIkJGwoAjrawN3LZoGYrdzJXSMiJ3B8ABDxUHTq3LCXhkE/zAx+Si5Yk6zl0Ine6bYEFx+5v
/lKWU7gpwg4wfgdEw6yr5jG2pHKGqW/i9ESqs2g9UHFq8we0Gbr9QfO+TxnuiRgWJAVZLLdvpV5n
mqIg2Ey1r4XtaXugRST+QEablFx7qQn2pZ9HJCt7661GoCv7EOL1JdCVMcuKXcZfCqwdZb8f40VF
/HjPDa36XA0ZLuvo4It5vpJqDWS2EV7J3snhxLOmRj95Y2yhma/lXyrdcgskBVQaWaoekeBYSkGM
eWoFk5mfQ4U1bESbh9ibTss+EWYgACeXPPJGSmi3bgzqzEtdNxxW2VY9bqisQkzDOFUEWyyAelTr
qJzJA/2PTQ3lEKHAHT0Da/Lea3+gUgdry/OQbFWj3r5ByGkyRWVWjCasXZ+ZjMaS63Ub8aKfDKj7
ynXH8oCUgvin24avKeDSf5IUF5dspdbjoUBfszXx63EjkSjKnaElIC4vo0dB75vAKvS2YMUKpXzO
R+LtJDe98m3TxVOXzESNm9eikNRJyznwysg1QznmE93ydaZ7x65Vt40SZf9HbCOeh85NnC2YJk++
dVuwP4ZEAKvavmJbkdwrkCgfzjX/hRSzr/TBA10EYB1V3UKnkx6M1BL+vDtpI1WN1YI5SIGIDTeI
ZaEnwJEmLhFGyV7EJuCTGwrELtKsO2Xo3BAdSQBL8hrdrWlD4ZoGhRyEMjAPTTIyqvzspzeVYVLv
0qccep8pExbW0K6kXwaFktyNhDDzeRV5qGJOyZLZI3RGpY30IQ0cKIMFAneFDdyU7JB8FPaEEXHV
OYGBxJErJRgqRlpTackIWXarfrqcg73YfXNQoISTtSAqXkQg0wemPeuVa8QjCum9H1MAmxi/NeoK
rvQots9BUsS5JDTb1tNY7y2IjdgNblrUokj/gpiJXS5gCZX+WuGh4VjJ6lnZ7kPFE3Wd+Tf3COAW
cqFCInI79+L1v6N6f+s/wLVUpl1GhWlpLWpSXmGQJiiQKdqiWp/OJGVYDCR0//iYFqJ+DFYgNRhY
AyRW4IEnb1Pbb7LSVeICKhj/Wcc1PizQzcMaPOPKR+Jo7lHug0qktfCo4RJqSascC8FDvvbTI9oY
1mGy6qn0B3MR8gZ2/OilBd913FA1dDjAW6EowQMmUZdBcd5Jt+Wy2HhU2AJqaaxnZr3NKhp5gZ4P
iVMOmGoNzUPY/Yr/ABBuupvYwOYW/qORh6FOEH3iq64IINYGH0YGSdgksvUSiFd7mClSbL+ttm42
T6EYD+XNKGp6XvxDtynbbEvZiAEHWZiooLJBRfSxMbry7Z9D6t8g1vs6HV2XKVnU16rOVjPhpSRI
B8PMZCnE78FpAo7z/EVaRSpry5p2Qt5V6o7Sx1IofjkHRdFW61amP/ThflrZ9lRfawgg8K3fgeZx
iX+OZM6646r79nM23Z6lWlB7eKJLecsQi5PT9esaIsaiBver/GmXds7EVMlta2+V2mPjSMGxIgig
SqgtNWAIgqTohay9T8gPQaxvUY9vwAI0WK8rySr1C/SCvdUL5aIuLB5i1yp/G09JW9NGktRemOkS
nmnL6pL4tFTyqvKovIjYv9ijPcjtzZV+T7yI1CCZm5/SOiR23wggf5bRDcMboSW590rbLV4oois7
6Y3QoaO8wv+bJVy7eYmldZitgNcdQuHmsB0wx1gFlDAPrm4VatiKCi+O0UUOxNbucWr7d+pL7e3v
p37EweEWNKOtmno9McOccFAML0HDp6Vssl3g0Pg/Vg4EGuPMAOEH37XJDoWpd/LeCYB2yjTnf2X2
RiSO3ylYmWhyRwIao4MROeGs7wVwf7m0EtUDCLeLyTv0C1BVq0K4MYlYQ+MtrAoqZpS7g8V1l+8C
+gxKRcv7U4fq6rRewEJ9nK74qEbCkXB80knlKdhN4nNkdoNopmB6f3++6u9TLyPr8NHJAuS8ciN1
WjmlwZUDH97/rIhJwDukLIRK022eLFCue/gUwbEL1zd+by/PxKVvVw1m9XlXywO2+2+AohvKjbjX
/jZKW2zRRd+snM1NqjbIrbT/f9p5Y6gDcel5h/cAXF5MrgR+UIkaLHNIAR6JHi/ME/HSVql9zafe
aAqs0LU6uSCifHtzKqlCZWLC8iriZtKaqCISDh1+P5bXSWcaPkJjGsidynT3053owbs3ZsiGOT1f
33KIPPk5QygCqCTj9nI8MSl5gBrrxiWO2WqWceNj3kO7EkgUUrfADDAgrMw0bBSi0hQESzdSSD2e
2v4QXXyU/ppSymMC8fsmP2rcrrRVlCMYg4L6DCu3iHrZfskq4Z7bvAMnNYsVdpXSw8zjWwh6m+aq
KCCvFgGZ+FuxntxsKGlMHV/tGq2KK7WiG0BPFwgR6h3S9Nn5Yty4GshRPjN+H/MK+QM5E2v8KGSR
GLY4WIAd3SN4Mu+BIQWUnm/XVFQUF2k9ZoxLhNCuVUVaRkDDwwZpX7CqW2fHyiZYdSU5eMGecgWB
RYSy/+4anls0ZMWrkE7QDcwkgX9cfCHuNvNUHRfcxfXIQ+btFXMjK3syeXVITOfrW9KOM5Ry0P4a
a2+/Bc/hOhiB3QvtnKSh3/z6RIg4yV0JLY8ecex6E6ExwuxySF9oKk0ZtemgBpwHM9WBWfv74hE/
JTLjf7pZjHHeqMmtb7I+U3LGa6M6JfACcZurUtoYEPQFHX5WRPKOq16r5B2PBlkVOyhkXBM7VVxV
ByoBvcYLVkpH59wE5A0aP/GYD9OLnByTgFt9Lvwzvi3i5WvU6+ePOQHcmU5WJQrCidgLnA/PffMe
Xz7ov9YLQCwX8wv9Ww2aKEDcK7ir4wu6NOHAPatsPnDgiah3s9pb750sfcAhO9YXBaQPv6BWUW6R
DA+KH2/N+9YEgrp0Je9h/dYjePusGUBxFz90r6Y7C+Jou1O3hpnp4pbNaN+WTjr3iEAY9/uqxfaT
XBhWiI56yBpsIqCcjzOUCxlF1YMZ7R6Aj1p3cNCjJTSQezBRAefCjIp+3od7ivTXu2IjYfC3MhsG
aZRsdXNfYhCUTpgcMPyRZachxw4kfWX8biB3yO4547JCLBcX/GOBgBQdP9i1eka1xy75xBKKatrM
kIGuR2SA8mVmlAW3iQNzU8pZ4eZZxu2K6POyKY7w6NVAPEFvFUiXzp3uPkGbbKBf+9DoW1mPcfGa
7ofKZesbKY8ilMWpFmPva5LgJgFEoeqAGfFACoY96pXQ0s8RlQfEGECp8+tnAxBsfbLCU3EJ/8hP
9H1WSE7BfOLhxdTOvRbsaSnA0rqJHXU5WKjtGBX415Or7GZiySxC5PbQRInz5MyMGANKUUPcMlSY
VkravySI/4kEC3WQWAPUt9LYg1RtaMJRbONdL7YovzvZBSGNn1ysanv3ZZJpesmujq72YsBVHW8z
YkMlox2igBSDl0cltfzf48qKGFZphzvfu0XbFYDovLqi834z7aXKQbu8VHvt+7tiFUuwLMhCD3Mb
Mh37s2kpMIN7TjxasXo3pzrVhuLMpjEYcLKTN54AU6edrnVNhF6Aj4fLlp+rgQ1WiviFs7+Sr8Pf
WYFQDB2TbfPmTJ0MjmHhO/gh+UbjfSI93u1py/rOk1zybvDsnW5C3/lCgMg6FsitSLDRbHkhhPRq
hFbmU/KtBVQ/DyZawOgWWcJz5qDN/ZSMWVw+3y2ZYWpVi01ZYBW7nwlgYgrftAtrrNZ5r0SMEUu4
UN5qluKv4gk3/dZC4/gZnxF3eAajK9ugDPcndkRJt9waNxkubMWTtUqli6TDZ67XmKRxA4W/5bhL
kFD4OyJqo0zK1gP7ayGm2s0BG+PDIkX2NZB3Mbn0kANQ4mguAgGUOzrREaGIXyaxnErsc/49NqMQ
cFzcrhg8qYlx192JL0KIeGK87I1xhDJpaCdsDBlzP1Xpxv44+64AvUtcZa97usfG0jxUGlOC3zMG
hlgpBfg9Qi24n0lyVAFysoNkCfJIiZ7xvel9xG9HHe7otwv8GaZXEWSZV90fVIgfHyvy9zc2iDBB
8eCU571ZGspM8F41F0md7pwCJxZ8nWHiPjpw/ordILiwz7TN+S7/fEm0Ipt4ZNNJZcXxfkEb6C/2
vowAT82vJvMSpEQ0sQv/cMfCqcoffxmUvpvHr/gwe56DSt98tDDdbN55+xZ2r8LqDOMJm1CGch1j
N2YeF+4yEtQbu4g6WkN/EXHALev9bw0nR5m3SIw84DHel1RRlXLFQGa5+Xd+TUQL2y5mm8+cZYuV
tsuT6QSYIDyOnnCEtiAwhVvMb9H29eCrJDNKYEVToHm7m+G5/WuLeQTNAW8DBP62+1ipvGd6BwLZ
xNu4yjGj8kB9d76YaCZwLR08l3h6XqsHj2rKjzg1rErKtz/CcMlnvsASEe8XjFvsKAq9IsOLZ7AC
gfuP6SendzSEk7hzfNyGupbjOiD66HtlZx5Ts8NLRyfklEP7M0ORu+R4Z/VO7D1I7tQmkQYKH9s2
AmSwXsbe9zX9m7C5aYZIUJFnF0bdv3kJgEo2MAYbea2ovAWC50259LmkqdmXekTcyYVI9d1UQULg
0FHVxbnobxPEwENPQxxHW3rCQzQb2nGDWF3o7n5pIOV7mwYEYx05/ZNFXA43tV/lM0RlMLJqhvDT
HA9lzeQT3UZ33aV2I3cA4VToMNotZyD1KT4HSuoXVqjebkzez9eNNcLRvjzjtEhuseAt20xywQTI
fYbtwvkAJ/h72pW5z3ak8VRvPKoTwDXjlOe0WTj4hakySL3HkcwJmPQAwdbL9bwX9aoEU/AP4AKL
GXziuZnpaU1o8dpsDxlULiLj3A3YYbXwHq5LXJael+oN35Tn/Wuujv/vYsRhE5ddgle9PgmVaZVm
xqQCgkb43X83ho5piZcewYJD084I2/3gTa9PJaZWKc7BuFXzSf8F4nzk1b0iJHt44jWdNPAPdMN4
1uIsMjnXT+wTya83WqAt8YcUyVjQKCXnkDRF/439aBr9/QACG2yRPFaiUzxwxteRM/xAiLUf2PBv
3i6uCHyaRoovFMbWLaAfaLbY58HjBt89cTCP70XuODXWWnuqmO04PHvnC6fzauqUEPbb2qDM/6CI
X9DE5hfv9E46ECtr+g/3YTor3xzK5lPCWdWSy6NIcUD+HUNTc0S9Gf3T1jiZHspad8EnyyQqiyUq
Z/BzBl8BvqV4o+pmEMdC5aXbB6bNCGk/ubyfHOC4kUnllmydP+JWQwz51v571rf0uhe5J7FB+1X/
dXlo+EfkJ/JVTWaRAkgemfTR8d7Mirlrwn2332V/WC9YNJh1p1BuAcJKUjw/z5qC4m68DZWdlN18
EPf+AvjnJS0nr/kt0TiymxCfzlIG8bDVasHCPRAPBxjLYJVqGe+NfesmMzWlOu/uFXe6ZOR8Pz22
Ci7u/4CvrBwC+/A+odzLYd0wI0G/wOeK94G55nEr0JP/Kvm5P1NHw28iHLUKVhuWNmtVx8B89Yv2
AiI3U1oyvdvtxoeNxTOeLSvJlK1/AbXwt1KP2px6PmS+wG5QvONN+PqfNvgDceH47AMPPbeQ1VfE
dvtRA5b+xTAeQ+UuG/CfvZabjH38IG1UbRCWkXr1zQfAwBhjl/ShmLTgvN9oOvgBEdBWlkNbGJQJ
gtdkgNozNoyUFYplc5CcHyL85ipzJodVLKA9BYWeTYWcM3LcXDCQFJNhsHfrhNBWPDFzVLV1wO02
b6mEJuXlJJAxbPOreaxbVxq/sPPG82KrOcXCb0gq/xMEwQ2GBS+WoCW55UwHbqMplwOVoolXDt93
HkNHHQfUWXF/rnLpVl8UhA5a+MM+uORABvuQcT8kL9RUN5OWzamij8iA4L4bUKDCirre8ISd6fh8
aXEsWSTusWU2vFT/kNtVMiZeZBlpBXLzwHAlON8Oj0J2xniqqy45bxd18KFlzYqoQN/SnwlNSjrG
IRp00okYDHaXrD+BBm4dEzSJpejI5LrX+OgqGw7xH0j3wCn5ouiPwTcqB7I6MPV7EtLGt7xFXfHf
Lwl2msH6l7iNzeHxyxFVutCmotkNpMqKBint7Ce5aCEd9/AeJX+5DwtmfWJF7a3zOgPOe446tgpT
GbAL7xz+X/kD6yV1znsF17d1f87oNJfacYgzEet2B7cunLoPH9/m7ynovB41Lr1V/k8ZvNL08GQC
lspberSiElVVnwOYqHRkzxbeYauVMA7SmTvrRdAX8J1CWVL8FumSPe/nA5AeNpJtGdwjMk1ec6Ro
4qZPhIOC7As95MGzwOLVMkE9Cb8v1NsDqN1tx3uEaTTY8tfDoEYNkSRjqZulrnzSnF+vVq+lRsOT
0R/1gQp6aNc4180e6MLNcC03RT1s1xOxgVdDVkhzO3l3BexAiKHH4CBlAUPVKoF8I9cRBKbpwDwB
tNT3Vbsfaeg142zV0FJZ1rVahvcbyM4Nwx99hrRgrdkltOx/fYIa9HcWkuYv+eN1hIZHyETAglSu
y3p0sDyy55Uh0x8JTKIBe1KBTQbQIMdyC2qH7dpAq5fLCpW+mf8kpQrgyxuZu4inp7hAwyX5QZu6
5iUNcAbJBFYP7PROOys1oUJFdL4pdXAZbiLOvXPukc0vAOTgrpIeZTeSoQ2qh/HK6cI4yOFc//9L
ijzg9QTZbmbysoLx7FipHPALIjLJNy7h+1IEC1vNqfS65VXOta4DEOSVS5vN7ZZJRmRKg1VxwtLT
wWKf1sCihnUZfvf1qzbUrfAFgAI6lPpxxVzJ8HLc3KMr6mtu+If2RnmPLYafcd8cFt7ixhsnzXrZ
DrJbBjy5YymJLzaTsiTsMwA0MsxTfnSCbcbPWxLxEtMeUty00qukZ+F8EhU6aT1/2JRME0YXxzLA
xWGWZLZB6Moni6z2E0wn8g8HQMfjSpAAre25TIAwIWYb2/cdrZSjOTec2zG5eTtwAWrPp3+qq9Y1
kmZJtxpfbMey5NsY9iA4oCqijN4eJxFWgblngyWET8YwI1u2yllF2CRtXR4d1YQRYt8hX7aaFIx3
otZY8FGKDfvNMOdsHdL7RjW7x6KxMNE8wmBVEBf3jg3xCvIQc6r6SxvoEzTXlI7SmIwYY90ViYQs
3e5CsSUa/tM+Go5MW6Y0GoxEuY7gelqlSFSwwgEdH406r26GfngN5bU1fqJ7xx/NVyuA3gVXKAvX
pXd+53v8cjtnmDY3UKsHSNIjZBXCJJ2bdEYBTgqIBuqiF+yTHxcX6Tvr6HoakEBJZTcmL2G7vI22
IeeNquFfSVSMAPmO8Sh/R97CuhWm+1ObJVlU2Jkt8YxF0W6lRG9wX0WpzdS/nu3aVPxCaK9NCTlX
KwlE04+Gl38zJAnRfAt/WbcG8eytJZWPUTaCldsqKZK+9CPoDrv3+N7xIxrvgUD758hrRRdsrncq
9NfrhWXXYVMbxEN1AxaGrWMb2pT8yQZp1k26OQhE0jr35uqQckTFeFKulVrSPARIsAcaL9DPBiGb
UMENXbQHg8Ljy5dV8DS2oZl9D+tszKTiRcQkwotheQl7xwBivsruODvlLBwxlobgVKPAxqjAbpue
r/bGR/IeP1AEVZtCZeS5ycVsHmPSGoNbH89V+itCY+1kOAPDSBktMHH5/VhLCFYUB83YRbtug9F7
7HOF/LxIQ6zHXfsSWKZIwzTR1H/EW39lnVRYMzKEPzT9IW7h8JNCE8/2n34OWgQmaK3ygxEUwpaf
azYV/jyhEiq567spUHAd53T8qwUV8PDn0Gs2IereizM1pn8iYsWTrEN8BUQJeiYba7dQLwuBbM6U
f5buK3xozrF8p3yTu3QBqjEpTvyiFM3SuBl1lvPPzevgFpdmeOJKNV2jPtFR0tIvnOq6TD6Uiurp
MPBvjQbrRGiQqK3DPJ1/liaqtXesOMG1q+PyC4xXB212i6LQqNheyIC/LQSfg5mi5sp+M+WJh/05
Kxn+GDc+fjeDQ7PINDYh91GAJ+Whj50NCY3qUvnHEpS+g0/6EC36EOIqbrG/1VYp2biCf5IBYqyi
hP8reOIhyRYSa+XVPm2Ij8Fc4moKzhhNNaX0wG/QTQuMZlV5d4pgXGBG6fXOgYP6VdooNchilPwA
kqlcD279MzJUuSXmresjsF2k5jxQVkhACRLGCv3qw9vgfO6bMNVMghNBO7aYsIkELBV6ycbvLGmg
omHyLLG/GazNcPLQxFkOBzDBtYkkNpQW0NUaK8MdFfKPHIjrbzs/lN7eNmufhes66JL+1MGr2gY2
V3VebooQK7pnFdlGGqbNoyKyNr+0jo400wWYbRGK0Ukma8wUs/xwHCGlBnaRNovhysGj/yTRa4uj
4q/863gyyRHWfIue8RSnLKy6AAZbYmokOk15+U75xRtlC4ENsgPjYKM6H+6R4YGUXzSNlpJ4MBFE
6ri1bvxZwWT4FAdUgWPl2J7ARHAq7XJLUIDHDRv6pjbLgBk0+lUkFQEOmGWSXt0ACzoFD1TBq3SW
+2B8ykwADq7OCyhMyjKj3XFMLyO3QANXgyh0OpmN+psVZlqY7Zm4w2+gt+Xm/gHTJdRmnURZhBXl
B9n0kVfNZfAmE95ET0Hdf15qhVzBFp1vMnAC90fjG+ilwed+m6M/uJ5bQfiBICUrJkxg7NRQ93Xo
T4xQXmuW+Gnh4Z1PU0M0yxWcw8ZR9/6W44LagzDV4eLMceKmDQT1n9haolNr/7zNWtwTdmX7rKgg
w7IhKjcvVwYcaFXuS7CFTmLDjhUMtnjYAynisvTXw45IbauJXSugkoWSDXMEvH1dqhBUb5BI5OSI
0V6VLSYfB4965i3b4ThGeIAj57qtBNicof77ustybYVm3MVgsP7RFke3Ya9j/kkyZf/edIXVygvT
W/1JLDv7bwvJhFBTQMo3KIf1zThB9z5du/cRW3qAVd9hF/dNNd60APSXLK4ZTsYai5tDZVD0UNVh
QqRsjB30CfpBrBQCh3kmA8EHVGh6lYgLm8HUqZCxG7K/rjVtz8ZMJBacasKUf73+kYYHUapY/r08
ihS0M2EoCD5UrGHI0ho8gQF82SZsKc09R7bM2xYvVOVshMHPGBuRujvIZ+LpyzLIu2ikGW6xsG44
hK4SAqic0QY5J0yhYYXwgPjsXmknaBbvI5phtt6hdyX8qE0dy/ZzdLM6oS+gb7rQACKgPw4hsKVI
eWePufZVRt3GR6mgcqg/WajaDzGhOguiQIO7N7VCW/iv2cFxvyn6Jv8e7ptzLO3LC9O3r/u7FPTE
AvNSbMIeRDGSM+L1iUCUCdZlSXua0NNsyD2JFFzopTKVR4H8Vv5yuUMKOIabZ90MejW5RsU1cv6i
sUSKCpAtpIcYmo74qVJSMekDhZhoFw9mUNhLuWb+ysHXVrtXJNeUga9YS0ie6GIsoyI7vKXodD4o
X+Wck7SsTrVrvud5XaXXXro4n8E2hqD+PsnFquOPvKCQX13Id1D2ZJpe0vmPREw3M5v+ZishjaYV
qxWReg+Nt6lEG5YGFk2xt4sNEIAhhmZ6eS6QDohbtj6ZMD4zUK1wFS8upoVHAVR/A9IiqoxWBGTZ
miH2VG5qC0lx3en3YS9C4Js8Nh4JPm2aimOb/43Tcxc7OZMQUvaAMWF+Uh8d23IDa58tY/6cSjWl
Du9gXx5Ue2XjbRniNB7ZVy94m3e/ZVtLWO4qV2/tCU4KBOc3gsGNtZQuU/dgkP8VaG3D9HvY3/t7
HJurNYRuk8PdE+f3FT8FpxUFvFovjytprh6zmF80aFeX2AIVrLxzjbuGGeBX1FJ7TG+uU+jFYvWC
WoA9e+w+2UjlJeSU5yuAW4H8KFewQl85D84it+EwHx1hbgHPUaITbxRZc/eaALoOVsNRSpHBVFKd
lv9jSzHwfdOe0ILDvsMevJ9WxaNg/b9d3EZwu7mLFOQfoM2zhtQ8Ec5Dy/BJjAWBhSWYp/l7K4LH
KNsK8VgM0aRomNZy7CmXyonHyb+5xSMVFDhR1LHTcM47qkV59qHJR13L8QAIhK3JVluhqeomCtSl
4C6j/1sjU4Hcn5BZxYNCbnFpcwa/EOj7gq0PdfF/16zinl4vvpev31HRet1N/ee41tEvUgp9Jj0i
RjriRKum4iuuCNPphRa7z85V9hgflEjZhVFPT/NXob9GlB3WK72yrf9/jwePmWcAeC6NKRTX99Ni
t6EuBIm0PCN4Az4AZEaJ0LX4cBfGl/QBm13yeEr1y/9KLp+ZIKdrcUSWNp6pkOQyQppu2vg1MFkB
8MNmYE3Dbjx6PRKmn3wP5u2EXLXvfeSl7n9NzQD+R8M5wgLwFa/ARwSaphP4JiAfT8Dlci9JNU1S
aD8gJ178BXo8oHRUyun4RumS4eMcM6ZfS7H5RyR37FLi9IUMr3fgjgAUk8DGM6CznOym7KFyA22L
lIXW09oZJP9FoTDhguOlp7MNiy1LE3nYn5CAvNy23UbfxGB2bGa6eDw36OhaIJcMcJj/SKVz/OCU
o8igoegWNtGxYc1Yld40Lj9xYpTgpUKapaVjK8I1cX4a7aCTUWSJfvppHlBy/mBHhSgHsd0nSEu6
6CV/oTYnIL1Isvr0u81p39lXewlTXd/mmHZ2R5z3kC/pk5P+EPqQWgs8qVKSooOzGF7Pdy/Eue0m
w50gcUXTJbDb6k4HL70aCcw2eyUoaqRJMVpaMwkHaHY1QfnpgXj4Ge0LJ7XR1akO1gFZ7QS8KP1T
faBO1oZ9d0N2HXdflcD1LSuAaMvT748+UvqDXKKDSME3dfSxx8Hmq/QYxRX+fo814WgLffRslJwT
q/Kxhy5gwIJw9a7U9zYHB6an2ixuS7raO12+FxY0uE8G/WzVxESAOP+bTpVSH2Di4awI/8576QSO
H0xX4O0oXTcRhw2daQTbt2JFBcIaFirlFlNOxncGvxz353Dx7pel6DbvrGceCse9vE3zajhbx1Kl
Ew9Mv/63nVFWRO3P2WoMvMWi6MaYyzebITR/NOVi9xxJN3+V40k3Q9X0SOjm+8qQz32bvimA5rzo
pvlzYPBs48NNIae5Ux/ZRPCce3l+RleCIEpHu5NKO2lXTdX8JNEkehplSyBVTVvg88AqAhVp27t1
tSJ8c0Pdu7+tyJcMaxXUB842F/KO5rEzob22fnFaFqGWXYx/c2dATOmjD2cNgHJ1arbtsW/lRDsr
G9NRyL2z74XRorhafa8Et3EsRGG9FB2Q81MfXN4Q4U3QuuiBb3cFt3yiNqjwSRzrAyBo1EPBo6fD
T2jdPgOWwYLm2nL3BLNnEC5rI57PukJFq3Ou1Gdf8RVUqLteO6VmlIImeybj1K7CLTQBzqyRKcoc
gQe7WuCmdIUwNowGoeWdYqRB45/YWLz3ggoLKgm1svxEzNhoFO7C923iPB9lPlWH31ZYQGnvLWaI
6e5R7LVHlR/NdTIDrWErVBG+MQbWgzAYGoeFi3V7iTff4lMqtDrzgco4OXyug/RS1RLiQMzom+8f
yYLlzJWQvUBhZQMX/YCsGOQ/GUZQgCZxahNIOCRsSK/ETxKQhD1+jx91/2OhSJ570LO1eV537R0I
7ULj6ovOCrfXptDHaXyHs2M7eDcWCNH/6PnDrFK2FQFP5KOK0qgULl3H5BYpvMdyHbWoub3noEbt
X9DXL38GrpV0aDKnV6CIZirwdF/UzRwt7tH7rHTwrOpISuFyKKkhoSWzIBKJfbV+kobmz/0xIT53
6SOso3BwGfyhWGR/fAfz6n2ft4KzqvXRCZZTsr+Rg6ERRqRmv+UftMyBTxMyDHd0N7N8OJOpHx7x
BQfBeVZi0u2CuQGw7nX0yVjPJlBZrO3kQU4sxnP5RG2PDN7GBPPcPzx/xrjrlIca8tBXS54OEaAR
IKkqUdHcEVBdVoxldzb4hc4OFBUOKy8ShCpAhgPWrmInwkJ7KJtjY1M979V8xpGbfRxIb/mQfw+9
v5Sv1Sktt0AH//eowSqQk8IQzse+ZYZCqqIWrq6HH/5rCamViw/f2dKJHzob1XdKRP6HM6MuY7qm
vMvV24eXVMc4Ou5NYt9EzjWSeSh84hw2he7ULWnQj+5rcNYItCYjcWL6wrPGkOUKFyvaPcNrDN5r
KeTABhCxSetqH1I9uigWyTm8db/Zaw5yM5BBZvPU/C9mmd0K4Tn4iIgIw4SgFxAArNjGt4ee6e8S
x7t3VbdahPmIlKyNuekex3RmR0n2YTrsMC6EFOxm6eWAfNHNHhgEuJquOTVdQ+57pH3QAvLykDUH
5x/KeifcmDY1p+FxBrzig5GHaKQQ1SqTB7pOdP7H1MpLklrs5ju5CfDZLaFGt3OekoEuE/ftyDjP
ea3f4bqUwwbhULKm+qiX7qYmYrfV/6Cp89X/EM7Nr8EmxFBPSE8KG1hAFMHJAwdkDqqFHo/K0V3m
jPq7rReLmXdve9Ygg1wYcLwTRpcS7npcB6yBOeFdDIoyultFAigl6VsGtETCpmqiq58BUinAToSC
1sAjrm6hzJ7dPFEmvgK6oyNO3TAamz8gl1xTnAza495erYM4vsoKKAPo0LkD9CsaAjZ4uDPquLf7
qY4M6+mjDq/1DPN7HHhlH80OEmKv7h4AFalQtlpMG8O3ivtZw7v42meinY5boctyEHxikgtNxupK
1hNuLw8/sn3L03kTR9JsCPeHFZ1pBa51djzq8YgEN6e81OVXbJmjnTJK4IiUDoWg43r2TFBXoytj
7tJwGXWeHcK990W21u2s6Qb2eeh867xT0ieayI7iDYPjxPQOVjWCAfvo1zGghksJiC2+p5GrgfbI
r/gZOkwG6oLbtUA1tHoiPQ9p3GRf3YecxExF8rSmvlwi4fwmuhYNlet43/hIuWJBYDCVr59zoind
vegHPEFEJ5ILCCQ3HcfSj8/9I5xjqqm9PYMoX8WqzUKnOPmf7/JTWMBa873tQuNvTLaJRTSFgNKW
3Xe9/jOUEwPMe3jnA291zQ9386Y6K4pV9QM/BbSeiOTwAlbxqAfKuty+OpGgYiZ8hmuevtZXtloW
ixlkjicsrlBknFR+LYb1xRqUPc371BlF6VlIK/XShl2gcg8Av3D3gRMK5nDz9PGiZyTmGe6XZSv4
TsJ5RaQq+V38XtZK05Ds1396AnWqNpH6bdqCnX3QPtrfS5sz/MLykPzjJVNrzhPQGaVQ956qZfzv
71QLkYScL2LjL0te5UUgbkbaZdPkD9aRIOC7R27ULoaNV9Pwqr3GSyAm3PSwl2PUtvSAnj7FvbJP
vQ9TVUyOn97ijP263Y/zByhoii+fzIZ4eqtjZL5fbzo3lUcU3iae1jPT7AK5aDiyR23JuOYWgMTg
ijviEk1rMwcVDYv3EFgoB3fuQGK12L4/9Gs8K1mOqdXc7tCgJj/XSrbkiqCMwYOHgezt4IpJDhdg
J6Z+WXT6MmMaBjGPV4UhAqbdt0BcbN0G1t9nWS2j4W8sn9QjUAY2Z0vqBxBmqhLL5LgHayeVl7rU
hj8tE8khOnLZ6bV4Dp86sfVI0/UOrMNmjS7HVP35182J8pfPuWNL4jDm9XdAPtZeIS9ja8jOFa2e
YbPqko3DStNdbatflmRFP4WPBUB9ChaIXYczXNqCCyFalr33dpnnCUgjwD/zgwyUda6CAuaKAgE6
pebTP4fMqDcaDZeMSK8XLg45yFIH7ZEiUe2HpO+TqzwkYsqb11wRb6g4qpQqDjXm3OA0cQtMnRTz
cPRRdFLGVDW4z5//7NGT1wgr6/7KD9XrvSlILTzZq5cceKel0L4+8UPPiI+em6SH8782PHLh2hE0
yCnlIWoXa3EGdgNiItuZDzKpkSjagAtRynTRcdGbdFUwU4xpczVutsngF71J5dOsHGz79V0iBBa0
kDI7GhM+b0mnHTbBmjPSRFN0eKQRyvJopwz2g3/9K5rNVifyC02vwWEJXBlfhXUG0zE3PTAJZC8V
uHOfVY94K//YJRhM46TjUmbDokPBVNfoeStjuUunEocqVyxxYfwuHdr5xr02PX1f4p9K//ORtkLe
jp6uTz4LvR0xwZhwt7fbzwWZ9TAaqRrsIjqmRPi/EJ0K5H0mcu4BqDGApGiwanFBVqwn2zhjABQE
H6hOnB/s/dwTRKKsh5oKRZW4klCwpulzro9O1FPvVHjIWUwCOeao4SCGn/mHwe0qZlOR9ixIp7JU
uBPiqByyTX9dFdZOQHJ3pQr3br3DPWj5OVZh5CQXskf8MrbjOgFS1UNscn0rcVfdeD3zXYRAU/oZ
8D8AjKxzZ6+PFfXlnj6ZIu9ASDCGzPlNb52StbiFxHrvMaommsl6D+iRtObmArRpmlAmz6znOb1n
JtpTwjom/y6GiOPQRt4BtslP5abK8Us1l926pcAOuTOqKdbRivi2/xJuiJUOaMOZ2ILi+KDJfGYS
AE23w7YrIsIwk71gye+H4sc0f7gRh+yhBB0s3BiJ5ORJhniHJPHlxQihR0W6c3RsZyT3jFFfkMap
dnxg2nZPWzya8ZHLyd8wI2x5efHoeFeSbuTOUYypgUgzERWfmxX1pp4sHHU7v/CbjcCRu33MLlR8
0S08u3pvjfwRrUjLcKGHwl2KB1BUc7O8cN0gO+qqE7aRbE9zSFgRUm67Ws720buBwIojC6SV+OOR
NEwr55YOU8D5RfKW5S/y5WW9a4lJmxkAzvhL7CcShY5Eu06mLIjYFTCxuBIxyAjL/e1Oc1r2COms
1M0HN+/KgZreFr/xZF68FfIFKMO+6Xv2JT2n+6jsTyb15PXGk7s4S9wWL0wuVFbrGa1gc+QXmmFa
pLQ31Fo5EDwsBSAOzAzLmogl3m8blfQb8Z2xkdl2wosFdfyEVhPiST33iucJJ0YxoffDocPHTNsa
NmEkYeeOypDgTdjnhEoHo4uKKir3wzH1POrNqS7cqAXiuEs8Zpi0MmOad+a+Xa2xoHphdNGimR4B
v90SVIca+jqAxG5xZJ+epn2UvR26pX0xfEtG0NvsQ01VZ3zsMS012/+AniSXS8Q7GrQPoJAag2w5
5ffqUkq5NG0v15Wt9Q8aWKOJgR4RXVe4g2NZnLAVgU2Ml7I1DXYlA726yRlIPJUZvS1S04Gtbnlh
bBw/IVTGtBl18XGXDULl+vmcrCz6cGGNIwK8AhF84IM8Gj5CDksQlIoyEj7fR5dkIoknhN5t4FSg
Z+Xnxui1U5PIVOwXqbQo3Vv2DcrFo2dIwS3legozXi2FTDO3UeTj3wlz/wJ5zcuXKVCfRhQBEOVO
CYZfaIOdmiDTJdh2/BDKW5R/enwk01upq5AtViG0R2G66esE9MLsaoptzVZpRg0iOdTFmiznE3Xv
J1E9PJSADWYwb1h0oDjjmKZ3zNm0qiwtVGU3PkJk7x76yvmb4PO50sR/3mIu8OfsqzG0jfnj/yop
EHnCAjsy7jXqwKHcPuj5aNjs+EDX08+bxet7vCZiGEQxyPoDkKg2TxG94BemqTacHxp82wYMIZoh
uMagak8fix2em8E1aZLlt88fSZi7d4U2FtlOCDb91rpMFdw1jH8e59aSnK9mTnNZvJCVhClGC/e3
wQFJD/SBfo3HcFaJiLJfHC52vFPjUi2GMLfhKBzBHKTxQxWbqnx1Uw+aUDKf+v2Q5sH1abCtgOY6
aLo/ccajKaOybAljHrMmXrrtYKurFRCUKZZ4uOoJUD7WIy2rLqRNGUp+lv4NEPrYlDvmJC1roRW0
9z/5sgQr9pzGKnju6YWDuKKg8QwTez5hp1UmazTlJNzU6MU9KUqhwR3Q05f5W9PNAXDpfFwrHytu
7Gb57bxXZLr9Vb5iIBQAcyGc5X7P1Yb2eq/HtPVVnD6YkkcoQNHDVMsrckN8vLoMEz466as45QHn
z0FJGx2/Un0uFo1BTQUyp1zQlkhFNPHq4Elod+hhOI5HFn3LE1r1wOFlqdAua6RXKH4dleD3zjm9
Wmsrtfn185wAj79KefhFbp4bljcsXDEAga9Oz9QV81mUEdaIz5tMCkcKmbDgkIGEWsrR9pZPTE7E
KNvuT4/h+hXdV4tkVPnXwyLLuTF22YbTcLybmS6kQoDasw9n9BL1d4ki0Nc2Ti/qzlSHRKCrPZUD
+lBvJOnSWiItUXlduD1U0+6DpA4kmrUEbot2KSKcs4P3islRYKqHJxIg+lYjaBtYO+9iJUKEe9ox
9Kqd7TXGXVbYX8IaJiWI+ITFUnvmqUfhDS8RDQg12xqm+EMO0ihLcHeI1DitK/T4LAF/0VEkaMpj
8C2a3C/Epmje29HopszNJOJh8H/lvwb8LBzJDYHyjh+WqQbR8MtT56wyNh4VvjwsLdcoHBC9yS/2
XZPMoZL6WsX8pDRk54kbyeTRU7F4PvEPKoOEwcPrnOcausJQ/BdnpPTzdit/N9tkjR6LOdSm333Q
UztZ6m9hAWeQiy7dbF//bOHqIysXu4BYaIrz4UoEUiuusawA0gdZDkIKezw1q8h2xSY3iIhQLdAQ
hq6TIYqIGNZviBvkhd9o3oyzGumNJXbc+pcRYdIarYUD8o8sGJ56Es4V1QGNVDXiii0W38c7xU8t
00tamZ6zRxpFmcPhy2qJTs+Yrw+koC8yrRK+DXaSHcWiDnfSJg8yERCqtO/tSqKRfw64mulZIFJD
yiCP1kqQiAPtXtfMIZkRdyJSEfRbou5Ij6RjCbIyetAUb6ZDFX7JQa0l5LfTXBhHle66QJqMPPNh
QvPObR3FYQcM2ydHHksptb2C1ADm/vBPUfGCObF7SfWDKUP4mgiLHHxQqDth7RTDcp9HRBauZt11
bMmptyfqQWsY23y6E5j3vuPxSJPjRRo7oEDIYcjonIDGNaBQtcwf+cSYPO8ziTD8LseuIcBVHzNq
oQ5KgkWIokfm1GRTWFN8ODJzIxz5yVdwYXyNNfhxsl05De+aFllRqWh4Qje7QfU+sX8rBZpZ9+LF
soHr1NcSOZdjpBMmCg5kJWxDIMO8aRmfSipzrpzc9ZrFdMLFlLWuLQFvCK8juwxEULdwPjqdzzAG
fO6Vn7oRf5ChkrSOwuO+KexZWu4LZU2xEXxxvUbodEgs8llsvw8gjqBYtiW5i91eTw22tTJ7MTfU
Setq0Z1f+UIzapmFQYFjKIEt+WPn9gOvulPuRD6T5vBOJMO7yHNjRUscqdkuQc9Y0pNMhTaw1c/c
LiCkKgTKIPgFtyl8nRIMOWp3r+EWd6eLrxjOlKlxCCLHieARzmtp43cWQbiuhdbyODeTTkjJpav9
rAwg+tHxZC7A0PCYb3ySJcn6+9EOA4ySmMGh/3sonf6U9VeqgOi2jrwCKmt6pGrp9i2Fx/Cc9UN+
ie5Sn8fpgYgnrfOaVGFMEktMvqyTXmR8Wb6Hdg8lAk3y3KDJ63ue8PAh79i+zBkfPD6BM4bJx/A8
94CB2c6BamM6u00HOHpuEP1XY3uOiaq8iySt/bACGCXIE1WPzbe4P6PQ2dbirwbHfrXxuYmNJbub
s2gyB5jouwA9YoAzBv9zuQdGRVlzRVWgAQyvB9sK7ydJDAQPPK6LeEmAaGTX8LKWLoUKTGbYdd7d
rlu8gDToEpqewFqXS9ICdLl4bp7pg1ieSDoITlp/9GcwbjslotTqqkVLDmQMgxLEkKtFR1WV6Inb
hd4HORPeY+9boeVjpXRKjsHPYLfjSmeaexTsJgViE0Py6wzb32g1x/X192fYEr4ueaNfPOMqwLc2
mXDwT/+X33PIxz3AcgpLjRIaGjYadleByWPJF6Uu9GSJk+bR1tO1p1BDuqNAUu5oGmpxS/qmRUBY
bFK9mI8f1mLUwc2K5L/bdFAG1MOM2kdPdFItT1hdVIekchJaJMhp1XHYURWubyh8b1QrzATptddl
sIvZieheAnVji5ODyYvGlW5eBxyOtMi1qnbujtVLo38iXVG6QO+kJzcIZwQnjpQd9Zb5d7xK2AQG
hHtsfXUk17YQK/Q06tMbDbZxEtI5Z4iH9aZ3YPLCOAzOMJYBM3Bk2+qxnXjlNmdBi+rYtDTs20HE
3TVtZtt0X7cpt4f1mUXo/L3YqS8STPQ/H4BZJ+mhjTPsIzmCGGW9aWscZR9YcTTszxaNqkvSfT/w
wwSWVWcH8zWeMUYg1XNNSUn1fC/OD89f2EgRicSG+9pMULOi9z+5okzimtI0vla8Jbiq2VwAp8zu
hxxTNLjexx6noLf0xBj31T7t/IcsdpueOtIctBSA3xARLjHYNniF5lEsdIS+TCS5sjfIq+dqz81d
jxlPo2JHt3pI8JOvL1KSYv3EB5pSyI0cbcrWz27X9kvVdKxECbh9PFL9TSH4/N381NSM/xIVW0jD
KAQh5+l3yNzgXjwIzY2qZFtG9Exwnys4xJHA7QA6/XestO/NFvOWIqsX49JRnSKIzPdbWzO1P84f
afiVVfTAoo96m4dXa3g56aQyNeuN8sarktgURMHggx+EK3qY6rtSrky+bXYHdWz2qzFC820letu1
TmAL+1DcPBR0Pmeanu3Kw3USqMxZP+Ek3/wPVcQwYR35yZmyO1fcBNip2eObxOTV3ZcK5WH9KcWo
j/28MnQEMhsVP6zsWPiuAr9JICYH+2vqJsHJZxBsDOpqhPquNVSnG0gJINF2FOWWvIwfUdNXtTu9
XZbRy7aiixHsj+Mkg115P0n2Lv2TuVXoMqZDxbh9hdJzgY+3iFmRdRcR1kY/Y2hiPKcWN54zlM7S
4/wyzdUthQnb+BSVIOzHcDSxw97W6M/HIALW8yhKagtLz74UaVWi5pFBLkqSN7RfsYl+IDcFFq8Y
8XryE5oqRcaMjEtpch1hg175Wf3KQhVdwLlT3VbuGCJolKFH4dDrV0HrFLnE9i52mue4kwQhqPt0
7C5QrP7xxxzQvy3hV+Ak28oj+2BajQD2LQV3dUVUauIfd1dhelJ/1vwk2/mGoGGy93x4dqQYrcNN
BaFanMMYjhxsAZQaYPkBtJK21j2O+AGOUT7jqcvIWYPIItuNAMRzTONTLBicTBD0IQLs18omwfKN
WWwOrYiC+xoyYEfZlkqJZ4u/fr0ZhTlVc9ypG35EnIznIY4iFSxAXsDwWE3Gnkzx96mc3ywSgzrL
5iSUpj6OufWRcby5Mq7hSBOCHkYooxOhfQtDgcKLYOzZTpVv8hX8N6bnX7wArlp452MzQ3JlnU38
u98aZVeXEZV1bcRvmt0jYibaKlYJBIlaDFejRLycHVx3Xg6k0ro1WjRGiLrid7xJNcoYlRFSb1+S
IGMo6REylknzAFPRk6uty2qOPA/j2CwkCpv292on3hJeTHEW4htMTO4z6RWZCasI9X7BMQ+51zu6
DRvGfJXDQm0Zs/KK0lGmdBynD7qh8ZRT0LYoy2wYj0UNN7VKO6NhS7MltkRxoqFm51NDHxjDnJOj
2YdgRH0bPZIZ1QCZaCByoPYStOkCM4pdtIceqY96URnkJafjy9j0jtaE0iqsEm/NVQJF4+cSQ7U0
hIrMN178UWKSDxjmPXfVDXR/ljfZazJPoBui0N5xuBcQJuKDgyoHeYeZXKcjHftez8aj+RdSXQ/y
yAupJpjXz/M8SvY9vz4Ur75nqntL6KCW0mQbpvzyyOq47Ofc/nyNz886Q0HoAZV+CjYqmHRcW2Qq
1F7B0luHizRIkKFjN2j/BwKX/IbN7tUOJNa/WFX9WwZ6R3al1nAY5adylPS5JHZl2w0Bqsccs2nK
PYzZn7lUWXAVoqKVOdv1kCwi1spbc4fyWVdT+JjOkfnn7T2TRf1hLouXqhUu6yPaWkQOeS5nMD9i
XbNYN2T/iluN+m+N/y4ODEoQcXYk+rFVBZWsBJDE1fDIywYZnWps6gaWT/kqLlXRtI8UIQopr769
eW5ticQowoLeqLFMjSdfqpbPn3dRXaQiZE8/PT8n8vgUN9QECRnB/GNvzO3paZoeQkpPCkCxVMsk
T03+6FoWM1jtbytPwYLrROWEsVDKlF7BI3j3TLvHrcH6gRbgLy5xvi5wkEQbH62UIjYlkVXfAYvB
zZHcdwLZ3BwTmCYbyR7bJ7hs1buEPYQ4MZpD5CP6MnTBefKvq0ByVQA3N8SFDyUK2j9HXt6SEyLB
RQ7tTOucpzEM1kCdYm+iKHezf5dTT0YTMYEA3JJukPxrGaIGdhJLWxh5vWwxyYBIy8Il06Pu661I
+FgVPRsy2D4hmD0OU4OAAs0UU46x64dzob68fNoKRTdbY7ch2Qxr7/2onWhh5l4n4R7dU2wLx2dr
3BzLXVwoocrz/WXfC2CroeHtlfbP3N6v2Dgq2dzPJ23THTCkvh1LCTf3WfS+VMq5A2A2ZvjMHJSv
uPzduimICr8k8zhoYVk7oCkyVWF9w0RpPcTcjjLKuoIvlEsOpsgF/KfOjsCuTdTRHUu4pEHoqdmB
js4I/hqlnJ48HpdC0LoBgszXJpFTwb4oYdZQHqkFTsS3UVatK09Mx9qO2mI9349iUfqL8M2gkJ4S
B2rztbb6GLIq/bTGU2Z2U9phAim2UUaZ3TcNGEmfwL4Z6p3GBbeenlX6LkmBhQbt5ZU2IVQPGwA2
NDhR5YH7OVz7iwKfXsCtatkJtICkDM8YRr/On/y2N4ylnuhLffaG7H08clmdmxxvohwM5rfF2lMq
c4Z64S+yIvHyFReGN9+PxUEZk34gaJzzGsUF1lFPnl6ayEo/+h9awVt/T2dHj6Lu0o6OvRw67w8D
2AFcqp4C6cOZGbgMRaiyE9/sdEf3LpC4VouMSmREpt9HG2TRCQfRQYkWvFsWG3Znwqv/sBM8R7I9
1qKx/zA8qU+ZNrm+PefO36UdVnkSSdxmWcS1uBZ5QHTRy76o0ZLP0j1wQoW5q8ym144DXgFm0T+8
IP9HvRy43qQFWdC4iVxpPoYAv8n5YEBjfzSPLLwGk8lpGxpsYdTeJBopUD/BSp2l30Fp3eCYBM6+
rsz0CGYXebAtonxP2b96WJixd4yYLFnE39gB40PFtPvO4t+xe0JFnJhaC5/kbLGm9MQ3twHuvv0t
XOTUHp4VMqq0V5cZtSGHLccQvcpQR81ohNSSZANxpud48ZDpL5ALAH2il5I7/Q0POCWdnAq+BqRA
fncgk2bTIWsNjTr2ModD3lWrHg7PzrpDSopGSBg6YQx+SlVFkLR97qEnqeQWz8zp8yeifvf6waJV
65yRHHwRvLuCH6YN1RuoGVK/JTtzGOCYzxcIQ+wUY09h+2DcbWRfva7nQKrJ3fps80GZQJ32tbpo
k9/JIF+yn7g4x8zHHxnMKsp8RSzqSpM9k+LVKRuEd8tD0P/24St8ZJ8F9jxP6gIX8XnTYTx+MXxM
UQXW26uQufMcI5LYw0uQIbd9J98+IbrdCJnPhJ936jvWqlv0Jcqa3c20AW/xZIWgLQ/xFiQKGLut
JJRvg9PTVr/pAsQx0c8L98+zbGxcJIBBWXVKL1iHf8RyZSISiyJ+Ab/GgAkDAQASKA/aIsmNdsgZ
HDnIfsg6v4MKsrC8UwT2m3N8SEyKkjE+3g+yAm6F2xDMgZ2urQjo09m1qIFypsU+/JlQfOdf9qJM
kqx1fKZHhepm785pERYH0UGjzpXV7bASFZkRelzyVPmZPGWOA/fe6SdqQhyL1vce4g4YcU2p4gvT
+C93idmH1eVZD4PJQlsc6byGx89kYFH7cdpd1aWYJm3XXzfXt70ouupdCmYl5iivswPRB0MawigD
yHTK6JzeuZ9k+XlOtotwlHdMMLbjiUXssP21UNnQPRnjIUSbspxmhhfr/eJFqSaF5RDfPEuDe8BF
7wekzCPYLYCbSkvZlDGZ8qAG/GPaqhe4Fa0C7+lTMHakRwXgiyl5hOPNx6ou+vxSivMdmPCXEyON
cVhm+nxb9ov/jwit0StoNt8MhrlI2GO4cpivKDToEafoBH9uLea2kD5sJB5Ck/uOmXbZsXqrTr2c
sYyy24dtl/YMPG9r4SYXd4/ZCMI0+SfZWrr5BPOE3h/gFA2Zvec8fW2YL1lAwTLdS5PwbDSt9tao
ZLN+61IgKB4wp3EckxC81fHir0goI9unLnPEgc9wRUbvJ7IMuoaYPdAR8lkAQ0vUTc3I8Tp+VD+1
XkjGuM6B2BZVEOlYNtI7P6EvtXGdxNYu3YWedw6aIcV15RPLIivo6piL4G1aVapI7CfPnNJcqxOR
USxYkPZSHzUcpfnTBn6s71+jXSHtsF9yoKPsIFZfekfSV95p1HEgxoVoKFCCRRJCB+HbWSuhm4sj
MKEliuQT9lNuFGEgdkw9QicHCtvHFA2sM0fF7UGuMS05LGQ/dT77gJkWMXKRQeXMh6RT8cJCqt5K
dn03HDHWj3DQ044NThf5uHVe7fExba3XfFR/QcXuNYJCE/DVxpPVIMGghCqhSKHJSIUdokCp0zH+
NRcsJ7QBrp3gkByc3BFN9DlS/zvgehn2Hbf/5zEK2CuY4BhHl5jAT3S4Zo44s5dmjePsx1atwwEO
ZXpVron8NCwSL3EhNhbuJeKOZXvfXEULTa8vv9AOQHGb+UfOr5xVe4G+OVrzHHljpNIoZfBzEH1v
hU+ZwsFM+kRZ1tJ/Mh2T4Bft/o4+7PicoVUhrxiBngwc1CtBmnxbKLDb7EXYpTj5Qzv/+JtSqWYF
h8oZWDQlYGIj97kh8WJ1zLo/U2o1tr6OWzySrPem7TeuzySV0xauqUZiz3B6mfp6ynp8M9FoKdRw
KvO13fvD6CBpTbrwWwkjGPyBYBja7RhRqzy6XqzYtdozNCQCX93n2thsYuWTrzSnxD2TwqIFC9xU
OyK20nhoc5lJ9uzbeoDIvG8A45axLxCgR+2NAGQ+eEGSJlL82DMLOtKcGUnDUjmG9QBv1XItPZDV
G92j3LcVjkN3CuofhLyFNfTfVqug8URgSH8c3N0a7A7kB684//IzdDODBuNCshs8LO/VOLp0VtR9
hQtQycPsWWiztYaMdAYVPoPEQ3ZlLHS/qdgQsMKvs4pgEUtcqvUewgga1qtmtvYI6Shd5d+sEufB
Bw918VHNnWS38ySl+CXlUwQGB6O3CHN764cgozYT0KSprmm4ZsSkM2BNA8rzKAW1HjqoWsyap1Ki
WLU7HSW2J32db9ElNbTqAGMr5/mx8C9bD8W4I5Rf81CnSoxw/z8/rklC47NNNE3zXdWpmWMLIhvE
uhs5bkydtF3gW0XPuY9dmTxBneTkmmQzyzVknZU+/rye73dFofhq4io5jgoAAmqmbPq2moTxT6Or
8HY+nLS6j1sOzA1sNh+bbK2s4T/gaqHa0WE6YrhxYdOc4mKa5YSUnW9tFsRpiJPr8HuXFkwy4P66
6ggH9f6OLsT6jluf5ylb6uf6BDGMTanEEcvNO/0+81Rv2TwD3t+vLpH4plnq9LrNSs57clNy8gIA
oWvdic6S7GYlaNEDDTJ5PiQGoJuzinTwV8Mi8p40LpJFiqAvkYxMNuQWGNHutzZ006XrRkQoRdU6
+SyOmaPFfwVrvOfwfESiH1lWBPg3fCvZm4LFI0Uvno/krPECqFJmiLJKDNcNyjrKmYdwQhQ0hdAQ
hMrI5cepMlV+m9bv/lmfKJ+V1xia5RQjAXCAkWEhBWkOjAg0b5JpB/jaJY371yRHe8hOkQ10BIsI
DXPc53uxoqDIhha5ypq75hlMrus9vAySWcwYzjf2T3lWy6BOT9NE4XiTmBPNttiNri7llQn9AimB
5TcSrSUVSxSlmwf/Yj5yF6JLEDYMb9xkskH+u+41wF9pVl18whDGMFr2LJsegIbu/BJomZmNCp6L
a3nhBwb4QFuQ0mbyVX62PRJJJdCI5L3AJAdiYGcFm8f9YnA0ZAx4ukL0lcY7kds1w5gaqpPNonDz
Ub742uKgl2AVhvZIRJMtUmg7601+LRbocysktKxe26geEAq11hIfWPAuG7Djpv0i9WjKHzNkpeJC
D5ynmpftSGa89nwLzuFPBIputek6NT4Lliq+C1pLVbJ1LJHW9KtzNXtqNED26L2mFYGEmeoyJxvb
J5gg+FLnslKPNwTnVlQoxpCuePlKN1hpccL7EZJblaDeLt5E4Fck2cb4VWu+yTRoSGX+QBU4Sng3
YcDz2xQNXyjgtsUd5YnKgA9XY0/eTBwXqu9I0pGeKZPhTy3vH342NPz9jRnfwGdjj7Iyq5/Gu71c
oI0fCSCK4jirGzxyLlk7qCICh8txB+cRDXyDTJZlFxVsbNzyBdl4hWrv9IxaYk5eg93adKXEwqPl
tmPO8z7O5rYZQslfVs0/hEWMwRXh5NVvD6QW7mikxceNwWxAyDosRncjnL4PTuM7Z2r8wSWTEhxp
aDQQetIYlxYUmrS2Xz+5QuMbQiBfK5Mlrv4DfFwGZCA2SSZTYBRbO5qszkZdC+iZPzpWJyorrlYn
KlbrhXaAICRpHw5WCk871omAcUtsf+Net0Wt2GKFGv3iXPJSHbCrJNty15MLBu4p0YiYYh8wsFUS
NUPEyEhEqxFwf9DQWVuxMlJM5ic2LgvtIdZI2rMQElAEEUIBCMRFdpoPbpNvl6NGZs9zA4Hbce6I
ulm/YRLT8sCiBrAQ287C1l6AtpsLZpmIMrE6kNd4CDdxVB8LXLzjIhONsidrbnuaTftY3TH1V3cU
Jq71bNs172UVoFJcpJLx21hos0a6SwkT0dx4vLgfdqI4zaoWu0HPPkWFUY2QDk5JqV73aS/WwEum
DlZ5DOrBvi3JBD+ZgjnfkrlD3Ey9xVJf9Q04uclc4N2d/tdRr12RFcn9qxGgxg9MZV4jB0NB+Bdk
7yFJfskwF4KifV4/BEgyxDEldRa57TMktT+EKUJjatCQo/0C4q/zJbzJNLPAcWA8LC46/NMl6wZA
trvFcLroeIHPkBX1BXw49GPVvfjaTEk+ei+rev0gBaHRjqFwBtHD4aULesyA4xMLNhCls5VosnOB
5g8JnqQV/k5LtyKyAkwzyc4Sp5MB7EBZ1SzZD9rKnHpjk/oCpzDdfvsxr4a8Rx1qxhsJq+L7J2Nb
cxWFTCpO83VqB9VaQVNBt5dk20iV44R+Sl8fDjhs4a/3nLRvtRoGxf1x06wAlRxRq7tIJiBr4kc4
2RWlmoj/xIQNBEbqFeq4aHTUADhAzKnveka+izDo2/CNrKQs1whFPOmRNqey4OW7qw51d+R5p/BR
Jgfm+PGox5UsGk0YCshaWB7Shu7a7DexoW+9PCiluLXsEkyDW2xGUvWpTV/wnIEKHryo75RruwpN
VsPapMtGz7OL1NbXiztjfqfRwOXdEEEB4ppVXoMgAPLTPVzWLIvXwXdNAmiWE4luuuUUvVrcGJJr
NZkB53rmGQs6B7GCMCqha07n7I1jRuWnIYjxhdWE8MYvtRmXcgXmTDPzTCHNI7XkvIJjG1fQapBI
PzBfwZCHzDnIqYj1GB1pLTznUqK589RUxtJDU5piscir97dB3gzvrcB62HcYYxFll6xOvozIstdw
Duo+yEbh8FAgij7uC2iXPKamy4XUCZYzYmMXr++s0CxAqB0DIFIBKshsCgI4rGQ+k7opMP8DQWem
6uHglJZhRtrwQt8cvqmE6m9qSem4f62iXahTXJ0+CCXWRQWCGqnQpRtP0UTzK+CQJFommo7Fk5PY
qBv8gSCH8IOhvf4MdkuAbIArUJ/2EjbuhEVuzeyPzZ1z6iPFE6AOL5yxQ2roaw9DH+9wkQGT/K/z
Vvb4gQDufKWeBrIFl4FU69Q4Z0ILmIx+OKAEChQkzmNVOgQgoPjPHo17P+OBsn0o7FZ75sSAQrQS
vNRp+HK3mxWLSfekAtpd4ZWYmOXM/gg/VC9ViFtiZD97oC1rcVBF5/fm4aDInpF7hjNs4nYWGrKs
QRX2KaoqoddVS8A3zR+JZnqh/nJCRVLzcXlqW87OVoqkd+Cd1klomaVTYLm12Zqu29ePtMIiekBg
mrOWjMNNo5lSyrArv78xkHcgIkZeWxIvMbOj5Ra4w/XPx3xiNKmbknBYCkwbTeKuhHgxorieIuxm
6PLwWtWISWhzzpP/pxcOkxBtOKQUVUvYO9ya3qWiR+qtKItcy92aHDNRlzLyLXGsR4O46gDMGWp2
mQM7F8ryoZsboLpGXlPUjIQPDq3azLSYC/EMUWTZYwZfA27AXqHZn4MsMf2FbUFcfRaDkWij6oir
w0uwXqBT4RRnnyduxJqmqByfAzLxkAq8SljFrmI7yKIpBtgZVjzfyrWXr61D/t0zboVhXke+RBL8
sJ7QQPPPJFgXC4+V+CwGoW+mKt3U2LjJ2XTjIpjGdOZSzT9/o46Td7dEhDfHoDy8HJ9mqQvtSlk6
BsIp7C3+TPUBGCYxLl611mbwfefS8t4S1rZfA3sFHUjvJTdhDKo4FiXeDIxR5BnNV9s4/xjwQ5iv
PMX5R1IQloKdrlYlOCM5haBLAoqlMdYGet04oTqXVY4azGXaeND0DUhbSEKdt+P7bzX+GvjAAgOT
LqSFDxmvJTqHXFQd+ZrQ9Wp/+Xws36VYQfjiM7h4IKyO7dtySZMAVPOB8UpuzAzlVVbT+9agDRUx
u5qBD4Lpi9JWuq/r6K3gJ2Lg4VVMOinKMPtmkErQzOLVBJgBiXluYI9rIBjmZ0dvan6q93lCFQKv
ff4eC0PiJmaSo0bHIIXIJ1DIiz91Cq/hZbsv7qwnwx2MlObppDP4jyttv9j++mY3Tm4x3Lekx1Q1
HlwDJE4p0DtLH7Z+esXT1jniyTR5myUjvdQUi7MMwg9mgILmQuUsT7HmYuu4NPfHcvoKtBIZPwDm
o1B0D3o12vWNCgIvC4UXQ3/sda2BYbHBnVeGdGYsG6hTIDmzQAuURQutUuYxdipQKTHa+lGllbUw
5j4kzTT3+dBlHfPzf4Kd0/N2spAwHkA/XQnaHDicUxOgnekWvY+ZEGQhifxwe7H1yAuEqtLZLLmW
qMfGOcoXCNoj2MtI1XtfT+Bcs3Op5c6Hf6VSo7iQ7lEbqMVc0rr8+cTM4GNuA+DwEVrKXLEAQUwY
+Rb4RCcaxTFxfDxsFoEG7oHNg+pTKpC0L1VCwyAFuuo2LJtLUUX35Sk4IPcBS7MKlDyEg5FP2KqA
gB6tkCugqkZDTmRKirX1J9Zsuf8nIVh22vYhzR1iFn5GMEqCD2jl8WZ0nhUaSYvK6EHQ32nrdZyf
oh3ZtUfDo6FYAhX5y7QY+qFHLtaMoSfzfCMF0ZLFwrXNVBGrkxPLC5Q/tBvbiBuvq3dX7IQW5LeW
6JFvrLNAWKzcqaPnxA+qYozWTzj3Ygsg+iBInXDu9gLTWGaTx25e+2QGcHWjTkIfFmMx+kz3sP71
TtWNMC0NLuCrRMoJZNmDp1FJJsIxWcVTvhgROZxmG2xDnRKgsVCWtUplnuvZ8/fnrH33Ect2eQ2x
iwNjcth4Lo4Vgm+pqYB7mY1LUK7Qig8ifa8062sGTt7fZvu4nAyGHbS30/nmVqYqnST6L7ZT6h+u
M+B0C+tfOlpnyRwxJHc9P6uWNm5qkeYNtTWYRv2GsXmt91L6XBPybvEThlHgHz0qNp57lFT825Kk
z043pYvZRQoMF7NfG6YqT+oj8fwv1VcFPExLUHaOn9sFQadj2l9Mnulby9jCXOg3kord6bN/Vl+f
s2iqbhRXJ7c7ubz1JhkjvUpSAioGNytz+8kGj6iQsy5sfnc7x0Rx7WFSyUjGt38+vsga9MujVmob
qwv1YUsnI5kC3xOGm5KEbsaSSrVOEatA1sxahBcFOT1x3q48qT9KLI6Paw8VZUgWOLVfgK8bBfKS
GFwm7qy2w7XAN94Qvka9G3EtPh0AT5dqict7SUnNU/iY3Ii8p3jvrWvumxjY04dNppsV0TAl8UnJ
qq/64WIFBLezDKjdaQXfQmt+qehw+xniMy5gz3Lpq+yONlvy0hxfwgFL4IuIRlq6Ha206CK0Huzx
HqweaU2a4LCLhk43GAfDzgOMYcUtGuB2jqT6R9TKfeuCXbjB1lhHi7qnE5eUgnhL2dEGSlYDrege
r6x93airWoLkiXZTAEPp2Bd8xbkatVvHwnxmXXC4mvveo97pS+mRyX/kGTbtaNU4udeK7Ks1bTUW
N4mNyHi7Q4Nkour1ihEAaKEJiHDTkEs5a4THInJmJk4eR+QrceXTfgtCjyOl/mC9df+oEOSCJsll
UEmToZw457kh+KcutJG0UC/eng0ePqPJqv7TY9YngjIVuIO2yYaYbhARnb3HCSL9xel6x+ci7pEy
l74g7Kid1YT9n+HPZxWrVo0HiaVF/vlQbJWdjLa68i/aEqLuQQTa6+iEh1NvimNdvE7uUstOaAvM
5oT6oRO+YSB0YrcfcFKRjZdu+bRaCSfDaCge506Hf5ZCyQls1AaCaDR4+S0jGtzgpfTVhEhswrD2
U+hHV9xdSUCyiYClWEmCPCTVTeUXVX1c5ZWkVEV//yJC6iZ/BXDQ7KYnAMMRHfquJsLtrthpVwLu
FUU9uAwPvToJLPIxgcsYEmFZ3lJpZOfbcMFBLYCGyNmofbTa6Lr2yHZbc6vkF+qFFxUwnnYgbpV2
uYgLeDHFhhFToSAgQ7G2iDMfu+jooLW4DVvwqjTZJvwHarq+teedRZoHau6uJAkaKNsD7fH/Q6vn
xX3qVcP1r0ZCpKbNBTNSjAsDbMZdzCMW+bDWk/0YGfNrFCp6wfW3cevRdzxWVTuhOy3qTRJSUlZG
xgD9x7TCNQsoB+ahvklUdFjc+6x+8Z44ReevO6yeKu/caYh3NoxwLWUQun88lL8aV0KOuY93q/Ot
FNyI4M4S56kI9mbK+jURVU60zJ3e8tMBsBXcocT3KHZaCqdfRrbYSl7kdF8voUbc6xse6G+5tgOB
ptSceD8Hee3wgb7HuUzmBWnG7PCoH5jVJFGe21rrPmXE7hiQWRQBUumV+7FD5gWFsr4bBSigj1bL
gIVY5X9V0zHiVoSUd3CLoTPCthPYCLI3hbQ8NBRsdtq7SRN+HBiueW1fFZWmcyU/YjXDb+sQtEad
ukE9tOCA6gC0K8Qz2BtOAoqdObALcl1mLK+2vv/P0gyhcHoCWiK1JGnm9Ax2xEkut0LP67rr8PBv
0LHT8rfZfrPBQE2Ys1sjxoRdlLWqFmkxEhnllyQpmFvut/MWeaYevD9KHBG4Yu0noidd665Pk2MX
OgBUkoyz6mOxXd2oeeFD+1JZNgOYx2GuR24ZXB81Lr81Q+GCmc+zk/VXJiJ13cIveFLZ8xHE0A0X
EaI3FpyZCNR8UeHXNk5Z0qjdOzD/ZTTbq1IRRs/xqxxEB+do0oqpnsu7dGnn36nhg/AJWcy/872v
HHPq8T1X7EZGL59I6f0ErgXkTavomlYQ9q7NgKN+0DInz25j5dhkTB/5vyryvlETG5VTbYPMKSHE
TkogOvcjYyYXpAdTJkp6niSR+BJr919xuJSVkFpgrTOunuQ62MhRohz6d2sI1elSLw3rRdYbPmpA
35EWYuB2oo9p0Qwa6sgQJcszOHm6xKN8u5ZNdhIljAfg25Y8u4993Xp+SWhGA72DpiG8RLX9PWHK
Tmv6zKhL7w8pZTq0kza+bmq0W3ivWsYgFaLAidbM7NoLE1zkrIdyy5O4jZa6D2ks9xls//nBdNCk
j1Nant5B02ba0miJidmDfxcOEXFRQd5yT3ahpOqFb+beBtIVki8EoMERLu/KddQbJ4MRHD4kAAbf
MBjeIXHE+VQYZBaWxAjm0fN20tUdlmpA7Ol0kfmue1WcXXzvMQOyDANzJhmBkclQKwTdNfEzHlME
70x14ORzPzrrt4Spnaj1ugIWyUD0NUN4NToTGOBgQr9TEwDT1aP+4SsM/EGLwCVvFpuWpUQBb8nQ
APOxLmZW0XgBzb150ZsncoNad5eI3Y0Tz4zJvK50xwPXnEQPPGeyVi4WtTYgbANlJqrVFaUDGUWY
dXLhe5yQKnf/V80WLETG6kOICBvjy6953qLGee3mblsvko0RNSMJReIZ8y8cFx0diCkPAiHfVy//
SJKm8RJlZc2mruSCfM3kFGQgb4SIYeD9wa413zDxTuqVu2X75zOTOmYZ3CyaTwI+0xrcB8MnuvuZ
jWUJ0ivAYfoSOZWnU9f3/J5GXpQ9czPGi9F367lLo8fy3/hOCTIkaEATUgXJlzSjyZ6YjGsX4HYh
DhFSHBEVxfk4wEYMLdklHFz/BKc+UVcNTGh8BCSoDw7qXsklWQnS4GF4SYXCmZO5eaO2yeKzuJkT
CLgcpx520Yy64Ofk2hIwDBSPt6lwCbi8wFYb4fGHFBeGwZx7VsJVYbc7WyvNOZaO2nbOeVgc7bsx
/z3S4F3b9BEyvyEW3oEaDatu4LwFxRTaH2AhyWKO6iPBBUyUWx0vYnf9nd/UFbqsZTNXd2s6RND/
1YQYUiPadFoM1Dvdo+PyPA4WPgHcxlyWHLL1+Ab/NBzsnB/ZIDE/UFJZo8hd0aOZdZjRjByZC76q
xXRFhujfGwVDaC3CLXp64/AcZiUQdIlOQWzxs/yV3Gk4XQCL53lYkTK3PsKqL+A+q5oKVpHpZk6l
PxJqPQvN4X7IL9LCwKCs78EtChAgiEdsoVhZK1vYcEiCBUR9fm01C+Gs2U6raHVNZ/rd7Sfhfd0N
Xf4hPEuoWBUrVOWMZSTONCtJkCtmFLLdCT3BNfvgrqxw0rG33ojT6aSlGVq2+1lfHMIiTGnqy3lD
xDyMN6Tct2+HlRDx2NSb5h54psqv3JChiIOhPg88CARnghRm6gb+zMGCNocjc9QbPrLTeZ8XXZ5x
Ix65Nlm7p+tknAtM6A2Zz8MK3bJ5oHrkmbTt8SO+/JzTDnmVuSqaZJLw9plIj3UDRYKibPlmaa4S
6QdFSwJVYIwWl7zD7TXZ+UmTPYIjPnV1zBHU8DNhNoPX57fi77ATLCLq8917Z9JStcxPUYqjSksR
dbkUKpx88NPZLlTjsFSXm8g0861XiQkv3fVdWQJmJR6wds3DyStwEALajQei5YDplZ59eyaxgAmp
cOvTsyVfT0Mz3Lbcn245+3i/DCrEVcXcqT95G0YrloLz0Jb2tPBORcODuqjV/cuXyWhTwVJqg4wZ
RcdKsil5Bam+vKmJFzjQpuvjsoqDAv7Aq1Z7fBy5utaeMvtoNFw1S2TLlDW/Ur5ilixmvXkTgTn8
6YLB27B0fYZzEes/uUSnYE4dZMOtJVssAdYL0evNc4hQqiDlXL10iFrK8ex5Il6xNl9ERXGb41bf
SBYf5HsFguIq6XIw9rZ2RUB++XexwvKrYrFLGIrFa7WLK/NjpWguN3RIqWcxfBdEj36ZeOzFGfTf
Yy8EZr/wAyoKqCYgr50S3+p0ERFITNI77Xf2ymW9fHHr3oVorWRxkJWJBHrMXgAHwBrYFT76/gBd
5EHzFPIwax7fdm4BXh1oNHp+MkCyWQ6AkpA+X3YXy7ICUaWgNv1LYpwgnImzkWLvqFCuCrq0h0gu
YRWd31dFb9mx9aeO3R4Nn/ae7Yd/9sruXmfDgzf+9K1xImJdh4WPIvlt+0SkRFrmYals+ygb6jEa
SaGqwL7HvmdjfoqtoZdjX6v1Yco9YLC+PZczeAG8xFkrv52dAKQdCvXK1GJzKE3Ua6gOoZ02wy4J
DITuNqBEPTEL6GfPL/VI96ebnfbQg9IANE8tpmDfT1vOv+O0qct1VUdCTW5R3YaAj70r77BgP99t
cEJCRbRXI08Yj47n99sVpdNZJmauvAKHu3kKuV6JYroq7tf7hpwZp5xpVZewlTzzdHalttf0AfD3
C4K+SAEl5NT8CUjvOVK9Y1zmsTWnrlNDb94DNC2ZaQf4vfBAcM5lZBIrn7ORV/SaXYBZoYsCNpRr
n5WhtrUu5N3QmfvhfjJUMle7PnV6b09Mg4534n9BhevP6jXLf9s6vJrDLUV2YvUrWrNkGYU4svuu
2NbWKgMRwoxbeCShJWs8+d2i3/DiZy9EMAk9NM1lPSmIWBWY0R7Uo333PIbPqy7kVn/xwRa1CkDt
HReJyXwJHO4qXGoTGICaVWULKLgtgwda7EPKho5XrrctQJzdwDl5O7W1RpyyyZFBK72xXy0wQ+Qc
rRbmyy7pue5QKY7OLv1vGyChPJRWOZQPOGl/l0r4IsZfhI1Dd5XMrkniLZ3DQTGZuQFgKGMsEa4O
zUAM3nkIk406i/T4nn8zBxOrYxlcheze6uIxKlOKpVFMgR4bppJqxZrdw8yEVLB9TZZ1ON9JdwRx
jTspRamw76Rxq7lvAto/+M9O3NF7nEEzpINKiparIpguOp3d5OgzVC8nFOgUCp4Qvn2wI4Mqup+s
UI3vF2SUE/DaLtv6k31dGsaOnf0yVGaEgOSSSk3X44oz5E+x3be9Gvy2XXbfUwAmrAXHPrm+2yNd
WhyCEEMnR2UnuwOLMF1+yI9ACJ7/5qXjUEuUsvybZi+KSZQqcKU+JtRgISGLIYDyVfsPH+jekgGh
OhqNAV2KE+M0TiDnx6wNeAWzEdqamLKaSrCTC5q0VT3vKVWSQ8EzNE740Nnz+SLzXBSmiTjtC5F/
nNJ1fzwfX5uidyLctRksu//B2OX9XS7SdqffcuRqp2gebaLXYU7isvgctJvq7HjRAZ5HLSpK9jj/
XF9BGPXY3qVjBvviWlyq+wXxlHUqB6Nb6gAGAN+cmSFWqDx3b3tK/uI5ndkfksSnra6nAfb8fhWx
KeL4PktoyBzaP/+FZlQ+rJutI3ipoc6/rx5Ug/IwvJM+CVgjgcX4aXgBrVJeHPFGJufGaZ9dVT2B
aacVA4WPiwCgVB4bsNWq01edBNWfp5R4B4VaXaPOUv7Q3GbpI1pVNQVx+Lhulg4htjpQqa4mbEl7
pjRjsDMiTI5EpBeJNanlE7wj0p0FKhRHiSVBrGLWCAMD+kSpGwOiMiBfK+6t3Q8BV0Fo9oFgYwsI
GCLu+pJKekk5s1GGY48U29fy52cjIZSsurLOpHCMtJWrIMDfYJ5N2Q9I0+TBIzzZqSL+JanAkHv4
e/aJ2Dzr+Dt8xfm+L8mu5is5bhSENAlppb/Fy2e6/BZaHAJhafCnC8bZk8kVqkGufbkT0CLLGAkr
5JNfn57mcTYqFjtsuvtwh+LnYQQc0/7bRc4/shbUZ6hLXhB/WzXVCmD0KRBvSXL5kwOevPbyoWhv
LJomw/fBz5A3TycuUsfbwkibRFfKa4ch38gWsg5j6P2drC0y5/i2NchiBLgCxekdSfa+pghXizNc
JvafwStBybKxj0h6ySKrbRF9aeAH5hL+V2AJlkV4VSsGepwLlyYKY0VO5Ew59/U1bBs3my66YgXW
H2HTFPZbOtPO+Ccdepj880VmveTrqz744Fw+RI+CTzkiiL5OubCdyxc5Ezg6ZwSMZ0tMGscNYLH9
ieIGQU1qQXeTvGoWAf2GwKETQXioiaJJfHdxyeesEpp7CLQPHD6mgi94vFQZ1fNTNWDvGfjOx3kS
VnnT42OQdQUtLijFIqje3oJ0vFQOUr4X7UeTtIc9SE5gxXQVdlE+KLX31kU3P6lbLgi5kWx/xXHb
EL9w5uuazWNBTH7Vv+BSd0dLQi5boEM9aPKMrGXTuA9nPJN00CUm7vG3rgj/GKwBsXbs2yc00Er4
BEa6HBHa+4QM3Ja+HGc13no2cLDpaiLD4ZPZOUZQmrm2+V3scK251bY/G7J4DleeFnYCb015DXZy
ec1HSE8YrSrRORbKzNSCb6gfxe1fTpogkVCA87tcKGU2zTRcDtjbjAm9dDQ5rtKBTR+m5AvgTLdS
trTS7yqgSkxCsWQoE7As/mZY0f+oPhDVhMOI3jGzro1Rfch/1YAXmrbbm9NcUyU6ZOX5g4am+XW5
s1b5lfplTDZwNaHwCqmdr4WEBKRW5Z4b445PBfIeuGVp1QA6vHZWaFoMaGWJxwWLLuYK4B0w/hzV
uszgB2zEUYvH0+C4RoyJUYJhWwxTlqUmqs3PryluD6apr0XQpLthLm0+SjGsQt1dmv7j8KNUWJQX
EjYOVKFPVZsGnsgJfU7eQqhVyAKE68XY0D5kT/fcad2HhovjJFoUmDLCGHqlatLj8FkqDpNOYdwZ
lDw/nkPghF9Ww0deFqPKiVDClLCFfYgouJpXiaPDGRg2/Tg6WaAjfR0rOg8g3HOTJYcwHYGJEpTH
qQy+upWN9kv14p3QTeSo/nOcI6E2twXklxqtT5qs2CApnX1MTSNBHsb9TdMkwp10NovPeEtEloBj
A7apT5jI//InpTa/2U4ItByd62ImeBaHENS/w+Oi8jIRLOY/7bp/5lhnju8DdEjQbuKtE2/vPaFs
gTLgtObDuZvROrKNTR7x5oXYrH0ad13iunUMQ3ntig+29QX5ZKGSzCpSGk1TrgL/0NLZcWG2hc7g
71jv6vZhGcTD1MQaHiEd/o5xHsvrZ88v743I6GySEEbuy5gtwgyyUHd0P+hEvW5wKkAWnw8J/Q6R
I0o0fwhr40wbDGfD16DnVQcESvyaasDBBjlLKH2g18EYcUZF2LOBDo+RZL24QnGsaiVuw6Iy7+uR
sC2vkfyddHbXXTZKqVTboZyyhIVH3HSaZVHLPPp3dMJwr8tPz+jAOsQ4bt8paOR/C50nawp+6EBg
xZz6dMtS52h7TrUjt7IfBSKJ2aCeilRtoAdwMcKXHqFkiMyBJLAAaJq4mSnA5fj5NVqcTEblyisp
a2swE5df7cCHFmC+092Ne9UopzdJSlREmBdGG+zTsp9zikzYLfpCNiIdTU1VQdmmEHNYsfDakWpo
m4DXHCRfQ7ZcnrVjOxTPSCsX3fP+FMrTQD1eNlCPZy7Q0e2Z8p1F/scwAkSNBbzXgPgg0u/epjfY
+F4KyvpnP9v26teBRzcFQQVN7mUSWzx/kXR2SNAdzWzbhV++2atWRuNpRZ+SjK510tEw4WVsgvP9
jLt/PFgkqNpZAHlAPHGNK4jLfSEGNwaGu4yLWD8iMUus6GBn9xxADox1mblpgu2M0bSxH4vkp+0+
SDX0bs+cd4xcCOg2R/OxsZaQsLXCoHWAbjUpL02D0DMpwO3IvyVqOhuQZcmtLOozPFRqbfvFUcRg
ZySq3BzB/17XuGTnMwiG4yPrm/ZDvjf58vLmpaGhghXkiDOW6scuQVSLK+u7bVOxSwDawkAQUSky
CVsRMSUACOFU0mnHXcx+TbYQC991QQ5NJZ6b3rQOphW4rQIunJDs1zudGkyTGDaAWC/Bceo0bU88
B/W5UVfs2v3H4+/S+RxfpZ0reWb3lKG+TnXltw3AmwbcjYlSGteBssahnGoAooyqsy350gnoAnf4
bynJCdqdYvVaBmC8dSQV2f1PEE0UfoM8XmZGXo9cmvWJQRebb3uFeU76GRDGzRWLZANV22hMnMkg
4GsdtoRSWv04k7nccb85QBfb/vBrLPV1TDBrUub2LnKMeAg7tO/FMPqwxcIo1E+aauPWa9QzI2Ff
cKbZGqZFUXtInkqNuZcJwqSF/wWxILlaxgw4oDTCbAFAMZ7uU5clMtVJIeZf1DgVdd7dajaQO9xZ
fHZTFAJ5FWG4wZRPZAmJgxgu8OvFsOazctp+IfYFWq7Oa5LWyoDCO26rN0sUCsHumA2/Qm826as3
HkADcoUdEm78G6tcmUceMqoJ9D39pTlLCJ9JdE+v0N8j36yuV9tUEJsxYMtP0Jz5Sm0bbxdjCUzk
ajK9XE/knSoa529Q5Da0W1Nr09/LRTYWXhadzI8hJpKAKl70dAPqOzOxGXBC66yucvEpMtxfC6Cm
N+/OjPQWMIOvmgwd4azCfK+ItFOC+UxlJ/Qz7wIJ9id+mopZkA8aOS+Yjc0PkYKedoc39ZFKnO8I
1EPnYIW64rABNKmqOgPFrKY91NKJ09zDVYTP589RKhqAvX3qyBOAju1mAuNKe+XrE8XtO7vOYaLt
fwqaHBPEcjF/6t6APNcgnwrSLGMppNqUEVP6N20TWyrc40LnBuRBiMGcALKIqSxIbH4eXyj3vgrs
HGk56sojumfw+sBfKxPHK4TMxjjuJAcpzEJA/ze/rfVA3gRmAvkX+ZUiqu/ht2u/f45R4Kfezsi3
T1xkbGaDZCRvj5R+gMWYAjHTQvpeV63/Y4xdZQupoJ2N2f0zVbTtvd9ajHnvgzn0D6wb46OElOSY
msjdQJM/yaud+93bQuedsVLYQzOlVXzjrHmv5zY76zGo3J82ZCCYDD03wZXJchXhIliWYKB22lDu
CTVPAwIoBD9rxuuCBR7lpBmvKyE2YP49i3BgtUgV2EDCf+UCFrU/w2Ewqq1o5KXW/7sUYKyDiX7d
5M4My8me6sb+BM80KsQ4iedp1GaigxZv74A3uftL3jEym/rg4hUH9NXVsE4OkwNTe6eQ54DIIsl3
C/uFt/Ql7dz+20vYXoexjkiqcIEU5anJrFcWBp760tWnng5NVBsO99KvqgVmf3Bc3EcqXwZtKyKM
d942z77/rFdDDyWP1haVFPYUwtLM+x+V/DSC4pZV/4XJsyGupVcw6vPw7GAnmtfK3v6+aaPmPeqU
uWoi7iPttbyix+7bJDgpX6d4iK68AlPlRp8KThAt85vFe/aov3ykQjf7HFtrz7U9x2DVjIgTITBv
Fp/DDHF+n2bVsiu7yT9e3mRhzTVwEgFJ++BjFl2dibrQpxMR8+50sFh0fFsUWwUmPW5/HdO9bO7y
SPY0OKrl4TJqveoTiynVdhgfeQpdY9xWdcEMnvkpQsQVEnq0fhu9Hg+Jfiw/mpaxljoIvw1KQuGX
RZO3H+erbWUDKGyiQJv8NbkVm3X348UxXPX2iVj3AZfYHpdLmdoH4jV0nvc4My7H95IoFisLSOiC
UMSi9eFLNFnvo7q749KQQtwBXny1x36vEb4l3Ro+pVwBMeuv0fRZ22Qk3Qli7WmPw++1SRkWTrUr
JH28q2MzUKQkYYVYmfQ7eA5CyVoFpdoSJulwLnCkUILaHD4m+H/NN1Dos+uhVTEN0UTtLn7ytEoy
tbSx0/6WcJ/Rc1JVzhpg+iWMgVAFeuNZ1NGtsc3lpcBKg4RkHjGNsqM8rUVnpKNsWPNBLfCf9oBU
jRRtwpx1zYfgTn/MtiRsiPyhW4vLallk4Z+9c8NCPDmdn207r9hM3/sdkwY2RfjHi62dDF5in94m
9qTtzRo83NfQRCP5E/RwyoMVAge68cegOWv35xSexAOv7HBTNA1d7BNBZQc+b0vJtMeG8NEY6zBP
lcTg6na8hgpd32WKEjLOez3ocwOixGTlpBaiei44S+Y4KiBgJa2heIFfDzZ8sNawveiReZKBkzPc
1ffZzXJXHcgGHNvay8bDW/Jdvch4nuWplueqFsVmOTBUcipScTQzFTeYBBaoKV1zHpAbyBZmen9z
anuqpq6NEScuDbe+79kTFmLCGO+VZjELYQ3deC68R8nKEvvQSvBDYj06KYths9oz7CKyr0EyeUaN
ZU/KgXjAPGeLFlSa4cuF/lICI5EVS+HgaW5/wWvhfCc3j1zxIJiccZSP5u9jUKBNCESTZ6G4PGdA
WdGRaxJRa/uyloA1BfnPW6GtLjYGJsy6tl5Ts+KjuYZkrgzHrhyEcsDVLaAgnvamWhXburjZAmub
lq4VThIJ/XocyKPVQdZ+6uWJ+kaDbrmX7SatxFvQpoJZN+nO2+XdNyyBxesl7n7M5mYAdyDVY8np
+cMKUyEE40vAlbznzH3BFRvDzKSb/hz6z1xuXY1NCdiFiw/wOeDoD6bM3Brodv4Z5Novr9r+RVgg
LnvNmPWSnPYTbRbzE/U245TS9QNp6lN5VDOg+LVw1Nf3nWUYf3UAkOKpEoy8R42ohAG+wrG2qZTe
3vgBLYQseWNxux2RqSK/EQ8e+Ux+872Gho0JXdnyPA/dXUHDXTizgu2QtRQAT6G1q9hqBxmXA/W5
UTo0YiMdDja9P1k3ijuqieZq4Dj5eqDEeSfHiZOGpnLyVpna+7rGIyak/cFhyzxSC7ziTKZKP0F5
c1bmSSzEySbiS0mbLy8OcwWO8AT6RlHwbYrEfMVE8FDz3NuLItcGZNR6gEfBnDgzLHRJpjvJggBz
HfK9HprbJkUlgSGDxXXjiGUjTitsXcBEIvGkEetLETjxcW3tbSOq+ol0oGqimalwI9hu0faIVnws
lJP8kDWP9A634t+3kF6dKg76buWEbY6t9b9qnFoj+7VpEx+bmywqqQ1Dit7nrHqHd4iTpBLnn4Fn
dhkxI2XfZbPykOnfh+JaoUiOLFmn53d1kNmQoaKmJe4oRMWkaGMdCrEMolf6R/jVTIVkmbwyGicf
UzJX4nE029zvKWW0OMvsjJjiVSan/J+xC+vMP+Ozfez1bS5X1mJKaD/2Vb2G0B0hUhy4SEJVD3tX
aeyZjFPWAwcyA9biWbetGAPd08d15xEPdI2ls/6ppQmniQBIg5YyYhSTzuVPsKMIRERcRHeCgwKm
0m36OWpeJJUk+JAcdpIEuFRv9yWU6ZND7J8ndeLapKFAQlI9RjCj25YOGEdp9wiqDZM3ZaBEnstE
pJvooLtbE9/5bqBToHlEx41LzRg6al4QOGEeAV7DN1RP3+5V3Ay/dpB/2C4fEI2L9WsmPxxItA/n
gu19SwU32kx0dSQBlDGGBVtboXakm2nfdQdDLhhPcb/ChR78bnyIMXJbabRE6hoIDrQWqG1GSPMZ
5CSnWIWH8Cq+mIPeb67wiw4UxYrtpXGYLjiDctSxQut4OlJ74imLFPmXYKhFmcRbOTKVdUSfMHIR
YQ8IQRjDbWItG+qofkKuLK67UgTGByJNyeF/xfK9gA88JRysYuZlWEjY3At+e2w7iZZzGTI7Mycw
hIpgqSbE5noNu/aauYx4ILc13EI1I+s9ic+Xt7nmtOVuoWVtdmT9WW2ncP3RCq+vVjWekR8lAGRS
9wTcsmCACsh7LLowdxDd7/3x8C9gX2eAdFrmt66j6/K+Y1u1wsxGTzmhy0uoL7EfoIoDm5hkdXqv
FBN3oR2kZRxNH7DFQoiB2kn3kUIOYmMmyF7ong9tBhsjYIcPjJc1vdPK4fgHszVIt6Efw2mM2NrY
Pk/WvE9l4K9cG6vkVWe1qRxui2S7RyJguueoZ8mqVVTWTjJyhM4ad2cIXcaDvqR6DGcWgg+SYbqw
clN/vBr5vHyt5x0HEqJhfno0lArVrbf6ApMuyjEzj7M0NKdmJoeIHlkYg+psjKvoCpQRgKm3QFLu
uMNdcdsLGi3LH9EWIm5WYU7e5ybBKIg71ouPom+NTXaovj8ScJoq0OTYNH9Dwqx5e/txqC+/F/1m
xIJ8qT1o6ZMvZ276LP55Fge3l1/cjtwv40rVzuLmZkkTrV/aLCGIyhPMQthbp0NyeEQ5nAZ8RlLJ
Ko6Dq66vXtVPS5Us3ujOFfcVrRTI94KEZhP07T3RjFeX5q1F644gL8Zb9W0WrVLIfQTnbTU/WGjh
DVsNT5Gef6cIVqL375zJJfs43EgdV+1z3CHBuqKUXvGMLwzOsjd01tqybuQ9h3DKfcDuvvhDN8QR
R9cPk73C0MIQeIZJVTaFYI4Ctm6hgVTX8I/0wQ8rfgu880JGocshQEirKoube3s3gR1PC9UIz+1r
Vfqb9ICp37XiVnLqlUuy06F57/nysROD7vdexgAIFBsiWLJ2XqOHmdnYy/ObfUjyfOtWEMvU7fUm
/BUp9g2Hj4B8Hx9PMBJJje76HA5JeBAeA2K858Lv/OigzqGZPR3wwqMK1zA7LkKVbNRX2IgWYuQa
dGvzZ8tddnlMSvxWGRDrJu11/BnFDMu2rOFOQZZEj5PocIdUJ9wn2SgbI1SRZ79ZfPmYCXl5cG81
fUdjy94Lp9RJcSzWvdirQWt8581TVYwDw4ZDmR9i79W1ip1p3RD61aWR5nj4kcd4kztAWx0xfuy/
V9MlEYi4vyfcroZVyta+ssupFMHseTDUrVQzqM9dwvRSEcwh65w2nsRmWHckp8k/fOwwZj46GKF9
99l70DLl2rGMbgs6rA2FdAOjizvq2AsYdJshVmYSczmemWx/xwyYYv8CjOHis7hF/WhoJWEv71LO
jc9mZkkFLG2WNWxcupbO7UxBL0K8n/qYSqmpW3a5WOLUmOBNFMf91bMkU4nP88hBkxNh3J+UZ481
F5TNlPdW6l0NKeo4kDpjc2cgeHcHxYDg1hOdFgXcgZC+u6kzdEQi+ZgV6ca5P6JFhkpN9cnyEpOl
GmjsKrc0pu2ZCPZpj/CWsba8SVXkEf7SkQEaXOVcAPbrVtsgDkiGttSj5D5MpN7hZvZ0p1ms0fND
4mUC7NtWjtBKWSal74ytIQ9nPbmrhPvGfrhqAyKe5DdJn2KmA0TgpMF2IBwFpRbe0UD8zjj0/zEH
bM/TdhMs01nkRvuqTFKhRNfCZzbL5WIp1Xum7tV/LuHf4Sjja7nSTfkcuq4slYRm/wyb3kwgqc7q
PC9KuA5t1N5yPzZ7fGMUqjRrV+IWApikTdBxn4bURnG416JHChhtHu+4uWkYJrghERdmFk+CheGr
aCVOXazbsZ3oZTbZjN357JaXYnTXJEqJDi5Xuwt0xcCix2mK6rQIEkZOjDqAJFN6kACEnCnqqtwz
Ts5EXT1jEDhXecal5YJ+sMyjn+W9fw1G1yUcYk1yZZ00uzd5O+CO1TMMjFVnfiLoY6fztX6t23Pt
8XsAse7F7JeU/GHTZ52ZZT+RmS1SsqyqhJHIOMp2umgeuKlwy//5uO7UtPUyOnAa8LJWxCUP7/Ml
yY6ojfMNsMKCWNvELLzaL9J7iFjS82u+JpDSP3GQbqJK+lcU6xgNfjX2vm8P60jzn083xS6q8jdM
iXhhTQYdZSqtfmqe6rJ53t3Kor8yyhV1ji7rTGZOkLzt9waJfWqGe1zg66g4mYpJqEDxV237229n
3jz2hg+vdjakdP4MKUWWTd0zuJHl7AinlQskecDFILQZc3HE9HzyHfXiYv6fh63ZqQ2dYf2GIoKo
lEytHyP7YtIYwUddUYOQtHv2Q356adKRtY93wEC2L6nGm4HxHuzL/P5QAdEOsFKZUb7ZZEVb1t62
54qZYGNOQ/ChIVTORMyofa4VhIZ1eQVDlp8HG7vCvSDNFwQK2q0jGMBomg0j7sjgiRIEistyGNqP
lK8uYneW0KXrezQaaR9PlIqr8QBtczdtC2zhKdNpv1kftMQ1ixrYTX5xJc2IaJIluMEu5DtLpTvz
kgyp3GXGnVkL7mNpegbkdQCOXDAoOxG35e5MBZ5XnafO0Ga0tNbq/BVLCkzkNG2Id8KHz0CUWKLD
aHJjGX46W2GQsHoHzzfJOBViUgxqsvfuPhdgzo25WPplfnWdrhXRerqjOm2WD9AdQheNfw6VYU1U
oZrCFj4OlPe6Be3R75ZyevftZluk9Ouvi0EXhOL221/5MJ8qJ9xDv0K6qbnmUACWBHl4jylpNsRV
R/mR4YhS7lnLZYaCSxLBShHmiGrPj3S7aS0QOH6dWpym4qlLJPxr+gQHMF5sFxiALYmOeyqz44ed
quON6ZdnLR4NO48UPpTP0neArmgu1pu5ynZFHroNYDEGYVs2Fah0p1A6QMA1Oz0FTR1cV5SQAVk6
SFyBX1UtGuUVGQRnOloxnZUzwUuUpAxaB8k0oh7YW6QH+jDWburb5IG3fDG1yz/gmpNVspN10+ZJ
mophwQ7LGcjP6e+sc8mUCVSpZvWoPecrXTZk8cQqU8lcDIOq1Ek8T7SvVmkmf0eHYO0M6W77Noqx
8QxfS94rA67sxilK72ijs/pb0314+k4cfON1RruDMxoOc+wIK59SS23Q1luBgMGGG7RlbkVysjRG
IpOudfi25KvQ0cOBUrJjnzZwez3h1HygYKsPy4SOGqNUve1skkPNcZEm6MdK8TsXjmNrRjXObPkV
IHkopmBnZbCc8vqmFd9PXVOK8yzmezwnR2E4XSOPZeyeH+RHWWRvKndPRyFU1KqKAbjm3ynlnzyN
lMnhhruzgq9Xl9ZGGlD9mlkTgg2QYRY1CnLyKHcPN89iRnCD6wjAKo+cQ70FKHik1wG0NJv3eve0
EyUDkqqklfn6z/+aaJNK2Kf8g+EotuDvGJVJEPlbz8ybjDjjrqepUSHyWutVx+HYdZnvaUiGwdE2
g6rUUg132WR1MXp/AWL9L33xnkR0Sv/+jTa426zmt4XZyF0d4B+XhuSH4xWAYtNU2oqtafMPIRF4
nB2Pyw7trsypYfsjl89pe5FOdqP0GUt7hh2acKin0ZlmxhlmG7dHj9Gsy2HnnLeJLgYp1jnyl2ZV
LxalhZVNf/9s++u+WEEavWLAlyA9nySY9z/buO77dL+25pjxjbAP+kDRlgjJlCcFiRlhhRiPoyt8
ns/Sh6mqWzG9X7gZTkGCz4wlbatIdGOf/vAdFtPQYtLLDfvpEQWkt9vT4KXJZRxGgTJaUs/mKaVa
sye5BMkqYVBSvHPdBD5K8Ls8AD4PFQyXElizKUtOGm77yskMdkqKKj8jEah6MFne+3xKf1+jRpkZ
cEmDb/LLA6qBz9B9nX0eDtCC7LEkgZtuI2wMjs9pSANne3TjWsUFR4LE7xFagk3C5gYoVuUtRJS6
WvWwyYObpQ8SCiSJzDAJ56aMUEq0jL3LMSmZvFnV5ZQxPPLHu4UXs4REs3VW8Gm/pAQGTK3+vDnZ
A57hz3GmMlHf662vw1F1lieKa1TWB3z6X+NZtFg/AN3qU/MY82FEjd+yp1jSm1lWjmwSmAHRCVlk
QyWPsIjtV2AdEnkJVBC6pciOQ4G74JDyYzGCjsE1kx6n1GPMr4vO1uv6LtMKBfg0locRBlfdjHKp
E7vaIm7FKqjqn0nwwF9EEjTj6KwoyaubL8Oj1MsEDtFTxH7KaZNSjyA/8HqI6ns0wE1uoSFZaClI
GJQyJ5DwBDm9HLzyBETQThlBOy6fAQTmgBnyC3nGj8q/kcTBd2lA3A/7jmuKVgp6Oyj0rU7WbKbe
FdvclTYupCewXwKeiXDVPsLWM/lrIWYBpp57sL4MorMhkibmJ5pPBe3SKd+1EMIeB51+fGB58H5W
OJVJYyB2Z8jMgV25bJQiy/vUr8u40pAL6Po8UT3/DZjlspwJpZTuOEyyOhKu9PURmZTILiG29pbP
S3vXQtjzrhVOH640YHUZbTxg2G0mTZQJRdnLzn/B511em2QDV3NHq8ubL66UyIOwL+KljotvcZVx
ViQ+NV/LygABcJz0U9lvAGEfuMQUF1Oja7fyUeInrXGB1LflRz4SvgOBiwH43RZBFoP9JUwWcwnW
xEX5FmZr8mPLq7J/fOMWni9rTJR4jMDiuwtiWsqKRmLkO2n+S+dBVC3PR7+kWeNHPPa5EdMM9C5H
khVW/xIZPI2JJ6Qk8HNVMoTNDF43RRwUjx5I0qHlDpqPsCZ/ByCJ2pUcxIhT686DM9D3CubP6ozg
2KVLOTJpdsjtE2+igwedbb/V92Dcl6FjY6hXqj7+neJ7FApX9krJPaWFDqNXoZQBQwjuP5l9NWgJ
3npimfANIGpWgxmOZeaHRjJ/pWQZk6WbtdMG5l91CKXj5XNRdEw7Ah7oyNUbrb22rz26f239PQ5J
f25fvcivKdd1a94xoK9k3E5fmz15nFkPPvh9cbDracmeSm6mksMlaBV9c8vjf1wgNFQMkbRCAlHa
t8tPqE2hyHquTV7HGKLneu7tzYOW1r5LenylEaMlIadfbTSP5yuLbSVY3uD5ULvigKVofudBicBY
cM6dRNnBKKluLueiHxItw5iNqb7JTaMJUmb9GD1JLB/Yriybex+FkXRMMScxTx59x2U3qWQ+DnPj
zQom+WTOUpTidYUKjwbltR637RpmBhLfTy8JvQPXCLgoXdjpMGfhwzm4pDd7LddpbIVb57wuZWB1
t8VKSjF9hSpSDZl9a0sn5cSpjhAYWt13lMAWNYoEf3gam4DPU3xfF/TKzmNH9bYBnl6M6fiuM9j+
GM5rRIjkyYh19Bf3n4MDvFiZchWmu4pCO4mQpnSR0DjQq+qmPJDAEZIxNV2LjLLGTj88QH+ZsVwp
HENPlEbOkHm9Zc8KLHjXpXgrnbhK+PWwySyUgGL/U3f9cOyQuOtj90swHA1uwxT8xFJhmln+g4hO
hieBpE9UduSfsNH/UmbJVSRJj/EXFAnb/6dovxNYIel/WDO3+dwc3mkBlVdiFF65T+Rsm71LsOl2
EpRMVHocfKgT6X7SzrpIE9+4iCrbd7DrChhzaWuPFYYKSjt8nJWxR/MSsp5WL8pb6uRMxn3fkNzl
YH00NPo4ac/wTfpzkorSODnBaKI+ijH/Zvx9VP7TxaF3eu90VmWDYwEpqJtonLmarr6VjwxiFW/t
iVwJ41BDf3tQArJ5/5Hm44ynfXNqfE9RBZM5fxWPrGCZocL6xse7PYd7vkvzCKx+bjA9dZFDk7I/
+7M9rFQuS51f3IvZOBHD3LUKi8rVvaFov+QlqA7wpDG6skrH30hZh5GisAdV7qU/07Q9SCFC/rBh
nU/kAJqJT2bfnQsIOAw+REJocd0+mVMisYc6i94A9ow0SknS7BPHM74bOy/o/zSFftNtERpb8WK8
idh8EdsMKSiMXYrRxfhC+fGDuBPrpM1PoCmj4Vn7JtjgLap3ZeZ71dC8qHqNGhul7vOWhjZJ/Jxr
hFa5EBBwB5GRQnd7SYiV8Bfl/03OpMcsvy/5fcGpgxRLGEmRZ4xF7CPl0RSTjShXLiqhezgW2KzQ
Zkuis/F22qvm+feXs/PNzSd9Hl7ZyGO1yP/ffitt7+GCUDuRN1ow6Ywy6y77TZhYwcjF2tiEgTMn
l3eybYuSHe/T3Rq/leST/ofhe3J1mNWqLrUrDauPQ9KWZjoNujYslcR6TOcPy/mNsecP68V41kzW
zbLDpNggZMsyS+RM4uIY6X73INhOqr4WHBYL0pJ47q/iuG4o2lm0oEtMmOyUqIASaorkye1inVdB
M2NMzyqFaLcxSHmi2XVzDVvngOjNZY9bcDjcd5xTDes8grQjA5qaQHxKNbCX6idfBmjc4TyFU7au
MVcifyUt80nndlXTC0DaryxwSseIIY0v46Som7/FfjMGW835Hzw5Ri39kS1vSRk1m9QuSvBe1D4y
Wl5mtaCJNZj/tBwWAO/HMSW1ozHlaGsLvAnTbD2aJ8cEPWx+y1b/bi31Ex7hPKq6qBTBlmB0BPHR
FO4J7/H7/ExiIU5QkizibQ1ZWcAw8KeRwobjs4Zz81XJbBxTkBkznGE6rzzEFOfoUfpZg8Yvk9ZP
SYjRBEZlj8ac91fhr4s1/IPKAnVKEpDC+9ba7ecd9j6PZpC4PIXk9Qq2q1d3uZ75wcui6b4YZyzR
e4NjFaAC1w8Fxd9PswOxsD94CnWCKX3EvF1nGM7adcAgJdMFpP74oMux92gYsq2O8PaCbToHi7aZ
gw7NJXxvdJzhfR/QBoMVpT4W07EaIdXoMk4Avb3yy1sHcCSyWEtYZBWEp+S9mS2yR4XFAl3E5FXz
KuWyoL15kc7w3+JdWx9QE93KodRgaCmyr7Ju2t/mgLUXTXxjcd1jN7/4GdL9i9AH6TIVCBYN1nfe
aF6Q6h7L1ig8ftRiGlvLXeviQ2Mlbv5IZitSBhlJFPghFsfasaX9R84Lp0xCm9XtaBJwHHX7IXm/
KWZCS9jKUzu77wM6yshzmltNlfdfWqRVOKiXgWW0B2+YR5xX+W5vE4Fituj0Z33DgT+L3jqsNnHm
VUktKuUoCNnjwD1w/oMK/fJCE2tv60LUKvlX+x1Ik06UXBuTBJDp7cG1kDirKKLsDGUo24QTN6k6
ql1S4zOKH25gOwuvD6We8TiKS+M5/OgtawMziKQ7uYDpiwLAclYr5YPz1/tJwrXvq7SggGdHNdoj
Xkj6wlWcplBtAAeizAMVJQhcY31LXTqdRJhY8B6W/JxGGSAPcekQ1f6J31Q5O52xL/kbuQ0jc7UR
q6CXmfPPHXUenSD2qBS4lIKvCxwz4o7UIJzvvn1gpwoY5qO1Aoxg+ZbSt882G1MZMqNCvRr7zsUL
sJk/Ng8IYiBCxhVtitRnIWjf+LdjeyovVTWKbM1uzPdW+nrQ/0mGbiRXB/kuXWmuxj0fypDs8Z95
6Uyf0ZpW0CQkWvHYmCXK0/DT//NGxuWTJv1DWAg4KC3vVNtl66U2k6KG0SJsQzS1hbceF4Xdb0El
tZ3cmsjpy/qaUPdPJYktWRF1G5DhZKuxMvsZb4mkc+wFP48SleBGSZ0wh7Ipqmi7i1znu0RbanK/
jqydNGEKopplm9FmY83/416EewWBlfud8JrTP9abxzs2lmWnzR5Qfxa0v2noruZ4xV+JnSbbhwov
nJ0ecvxLPnF1zwSb+yMMWgYmBrT0yef277hkcmNHVlVeT35TJc6ZOpZib4idEa1ALmyqbJ84tDOI
9tsNkpqGaPm8kgV4pcD5WLJTZrv6RgA0wAywna8GC1MwqoDSAUUunQcow6BsdBmKgXob6T4Uzn7z
z5YDeE4WGYaO5hYnOr3rOgdGxd0wFRJDHuw7BUubcRjpQs6VTp6FwZLzFMNBmhg/LQfm67q/Km7w
Gy/uGxfAPpE+1m4cNHtAHLVxm3LaSdJJyYQ/BxWaLnMvd9BaI0IHqVj4Io6mYKnrH5X+kCqnmSv1
AolJANiLC5SC+dSKsGRgpOXnpXQp8prZa5rPkZMK24xwk4gIkBLUGTXFBLXCzKQCygZyu1ARKIWL
1/0eBngbIj5KYqZABEpPfkf0rRfAravMY70ypLItv/Mx+0AcYt/lIc9gGBBdcEqQBg6dbj2fIGIP
xETrHJz52yAxpxTcp0kM5uL/fH+T9ZI114iHRKIqvPpd/NFvdk1Ke/uOriY226YdjcYtfwZDMcZc
MsB2xj0bC91RT25C853VLXdIi+h+AlKtavs6FsjnUyNM+iUC41Q/MsLz+JOTyuksLCQNj0Vu+58f
cZoUa/OTa0k4ZRFfL+fstOtVQWfch4jrreiKtuNhiX5V4OIHpqxGDkyQagOJX6/htn6qRBh/HMd2
SZ0duzkHwi3XfAk7xxXz/OnY4vNP/zHj1JvnObfFHAdng1Kt5FgHBVwl7u+WqHS5L3bJmgBivmnf
eY66NB73lMs9IeOg/Vd0ew8gMmq70M88YC8OtXTRWYP1XTjC1q3sZZiRfAdRaJ3/mFhNQXYfbPtw
c17fb7aqUzY71Sf004Hu8Bm/xQMwCRtA6J/1wRA+O1prLdl4PYvNXQzMwFHIat49T4FnZTFCroJH
yBz0nHmHy2h4anzaZBHX+XzZiy1n/VNc24wWpIrZWQDzp0A8uBG7PJ1hnmia9Jmh2U/tOeR1fwdE
YNmBO3CrZIHRyhIFUwUDI1EmNXaLWGTHhWwKi8u3aIVvnmbapYxNPmGs/+RVNKTlZ5ubo0a0wDp0
NkQZZGG6eA7IyPPBdvES+G19bW2qTeg6TG4ImY8f3cSk+NbHpZP5WZFlAaP5d4CWDJzPMJDCfayz
TpKIQeEtCQKNvejGSeGsXKmzJ0Zjt/upfW1auVarLHdrJ9lcG2523dc0LGoo7xbXlCDXxz/3XBmB
WYSNfkL9TXATQeYuw944gEhksM8WGdmUsWe9IWI+9i1cUz60M2yEVlH30aduXk7NT08phQ4fP8Uq
WBrjK0yO/R+rBqaS1UNUW9aBGdQyJt/9Q4xRFXs2V+dUAdaa0BMH6laPlnJpwV4XCD4OgjUYtXoH
PVtaZw8Q7n71hHrMvqDLVjcCU8WH64b6PtJ6pDUtkpqGFtK/gV1vDscQ4PLa9qPzuMvn1A39xsYB
+SWnqZkzhVsOtInaDiTskMUij4DhUNRHP88A4J96E2rmI/sKXBotrP0b37A/O76zl4S817DdznuZ
cfEJbsWfiGzPl7gK8H8D4+elylV5h0+CMy3Ckb24FX5y2AKklOimNQkLhFUukKj3yT8G8JNJqLrZ
CKoRG8wzZCsriofohXww1ORPXRtWOzC5PweUaObo7NJoouZR8KDw4LY9I3BAHF+rL95Hi8zadVIg
ZHq+yB4v7yRPkN5iX23mBkhjBvjSXRcdG08/4b72WiTls46ZlihNYR1zKap8Mmq5S6XRtGMhfRfe
JLt3XzTpKyfzS+krUAig7c1Jj8ARmjIfcLWDn8zx4JA4V0QbAHZ+n/9D1wHfi+VHDJcDXmUVFGcW
kV4zEjYPaZ7bbjQVBm8gC3fjELLA4vwMjaKgXM8jPW5R0DERv4gsgG8p46IT2fu9S8pJw3gawBDo
EIM3NKaWeeYa67413K2vsueo8Av5bAAkrPjNhOkwWW7bGGOPU5qY4F/HdjlWdysJhwBg3ktz1Gw/
HqixfD15Mr7n2nuenMiIpvVn5sPiA62UUl1b7CTf5Y3s6p0XCPGqZt8SDDzIeqLkYlGx/lLv7gP5
WamhGDgmvQBjOyIIWmmeFzuLedijNov1mwjlz9crVYzvFx69tZdSxniZIrlJXe/JBUktznS/QHZH
mQTsu0FgTgM0jUdRvrWSvT7vrduj7U8v3mz5x70hIq+ZroXIyoJXf41f+QFJ7HhtElkhG2eF+g/e
jIqAQtjoHz6D3+x7HZHkVsA1C0tmjndkAJksCSRn0bgggzfET05rj+FL/fuISGA+YzgX4K7MpPic
UdtVZXt8snxKOpzqaIyZPORsniyNSuoW3ypBHsNymtK/HvhFtFUOiKTZBuFwQ/SCIv3FNjJG53qU
MmH6XRk8AlZZjk+aGxm9s+ygI5DhDDOwPSvzRkzhYHfvPWfQna/nvnIU7wuHtnAp6Dgl3o8Dajh9
BY8/rwNUzYTo2P187nT89Ar51NVF8pAVg7wSsqiLrR0uRd5yfKQM4qweDdhFXgzHkVh1dupnQZB+
DlLrBPFfnHLfML6nTYNCTV1jjESKYOjxIeV/3U0JZvHrND1wbCo9ty1dQhf3ODBO4ido0Q9L/WkH
tmOgc0ZDGX4G083mLKuLZReYvfFHX4aW+lCAYiQsmVhCPzBPzL+Al/M3aZko+U1DUx2j4fwOqoF7
Ie5hr5c6yt3Lk7MFFhAGUbCMJ4oJcjCgkUOTv2UNJm8N+ZPHb+n8IObPmQY29L+pSBYI+xIuzBOr
2qFXi/Er0VaHCVnpsv9YJLJb5+TYG9Jm7nq3HpWCuzkyTtjyX2zU5yCiimWT5PSbgB9vgxh1AS6m
CRMQS2rZiO0fhIvFaCqZ/O+kytYIlFd/HWm6LT/pImfVN/6se9MynIObR5F/92zyAUTBahVS2yr/
+52Noy1fzR1xH3193Is25xgvJoNjZG9KtHcQOSWRKy9UBKncPic/nmoSQP2xeloK1H3dASeJxQfe
gKOpak2EjszoZjaLzwoepJ7Fj9jw+yxxApQdaN3UrTRrVWkrPvllDiBLC1VWhnCdey56cBgZdGZr
IonR25NA2zDqB3Q2Ge4KaMOnO1KZMJAQVFZbjP4c4rm4lRA1AlGY78z0V3/x5T6R3vEGGI/T1Ryg
9tAtYVYvM3cKm9DO9l+cLbdI6GtgeEgvhpXi/W3ETKV8LWGIKLq7SYy1Dr8rtpcL+MAR00gpM/w1
izEF4ZbRmXMcKX/kh1eNDBcj52Hwlei+f4maNhsu//ZQsqzbNaKMDiwFj/3JQiZEuBJVYPbd5YR+
ebHjrI3oFNgZlJeLfIWMKoGE8q3NlGeHgO65E1pTyMgW02gffdrrJFacpTK6QImUZ4B2TpddVrAW
MtXlIv4jU9HHMne2V4sdG7LfSFrJ3eZutg9R+WAxNivwIxJfoKXM5XNziepbWC12vK4c3pbs6KDS
ZwKftWuljX6lpz+rlpQnWBZsmB/lp+nk3e69l6YwSosduRferS0zi0K0vsELnro6GBNp9TAZMdtN
C2vJnjZiusPXTVG+qmJB42YeZQLtQWQNSGmnxcZltKxixSxmtZI1DadhBxQ1F7ya1gn8Qea/KICz
Ox4uVv1IwLynfBGngtr3Di86mAhX4GtxrAfMdXgwSv5ca9kocKmm68MEJY4uEkcK9M7rZ228hrJ2
jZgBIs2eJURn/n6ssRosnpZRH8x+dyfofYTN7OgFTXeoas6vgTBR2aoCGYV1kxINvG935ofG0zog
lRUpYKLnLCH40T7WjAFNS0jIem4UJj8Y/N7jteAmbGqGRYQ5RstmIJcUjQpuXRn5MHSFk1aiyA5G
Q+MaMbBBu3N/HE66TLg06/DWqWJX7zMKPnHwy1L7osyvoFfpSfnGa/ibt2tS9muHJWsKqMrRsOTt
d1Aa/4BN12pdrdSkPEyXb5MeBaHqyYBxNRFCY0iJutpNul3PQCRNMwtCqg3Q3UkIYNoFq/6ECgdv
Q63+szrOfpSt0rZFqXhRPUOGnxIr2Kp/o86f+u5sq7POU+q0Oou2wn0vZqnKSo/hRmLGc43dkMeH
hncKB+n8TENkquLlZ/KXcW+Wt8IvpLwZPI8iS/XZT6GQkX2kx4S95F2GggTTai8kyFNJl9aK94Ac
nnRLIUk2hyx5UW1zOkt/iCxW7LaW1fdOMGlNtLgB7NvZk1zODGr34tyW0pmbdMz0DVAm/l/E/n3y
rBXrVrY6c9JJsM4PIwsYClUIJ+gg1Yhhn4Z4BB7yvaFYudgYAeUZ367aKaxbJv7OAUm7gOudwOxM
3gOYkFF+fqFqZrGCZxxV6ttMO+OMHUrxVbiKnesKYLMZ1V6ne2X0sYlR0xp+Xu9aUcrekxLJRWy/
UZavzB3DTlLy/0Jvts0fM2d23LB7CRtlkLzjyjrTeZWj6Vd6zn3LKRYwh2wZ/eXs4TIZLPZDHn6R
roH2BlQNLUsaW4OqdbDViPSGfSUbirri/3A/ocG0FuZRuOcLivBKlaY6SbleFvb96LKxBW89EaHy
UMWOG9sFiN+rjetgxiD5Lwy/EuywOYraab84tlK1cRDK5YJQ3sEHbts0B8rtKMH0Qb26GJV6LU7t
jFZ8X2X+juyKVCXKZNBFeQytUo7LmEbK5UIeWTk+LonMbgIuB5lt49W4ZfrJWFNvD3FWuTDEe8G9
YM4Qx7RL2RbEb7pSBMW8BkWFWyYT1mjauDCqDAHMCTziuxPPt0LEHgwow4FvnpkpqAo8A1Mtg31N
M9BAlKX+Qf5hbbRsjAamRMLFYZA2gsw/Oe7tdyATMhPo+wD9Y+wDxda1+l0Ii0w/UqnWjAsifA63
e6xJrUf+3HIh8ndyjz+GqmFFPl0MW8Y495/tk2mDkReme/wRKFRIRlQRyTB5f0rGAn5HpOwxyNAZ
4WmXYr7wg6brdof373n4jwqyJWqWQNSUTD/OvK8+xY3yzmR1/4fxETIUrJ7GfyVVhFx0pFhTK0+S
auvu+ObE8okLTWUHfQIBztHOttkfAdLqYrvnboE6HDjbMGM6cc5BhZPqhT2NlbYYA0+LZq2Yytan
cWZWoUHNnFjnXf52AMN/1Wbq7hykDDP17ZeP7t1v5YWx5b3sHE9JoKCGetdxQ7U5IFX30CsbASB2
geJMXX/0C2PG2CudigHO+TaX0yaLhlOiMWfBsD9kF9Am4Wt9hyLRI+4Gx3WIfnu7OaBQfpcBF+2I
ZHNiAr9nSbfDQDt9GNDxD0wkCZdcKGm7MFtUD1RfWdj/GHJJRMZt+VgEBiiGjbOTd3kMNh1yHRfY
lHQYgqZupvcTtLuqvQUlSAYVfLOVev8gEI6ARQtoNQuKIc9xF71YjBS2EaqGDMVnOikqlSfcJHNf
Jnfgu1e9PUT/Agdl19AAgr5ltxSIYTZyLtT20gwEgWF0Mh4wSmuo+d93VMOd1oQwme9meDrQ/M9C
yQ/WpW9zDadPIqvFgywUFB8Lo6inAgkbo1BTu/se6jbuzKOn0/0j+s+W/NPhmUWTtyxHbfOrCKa7
MolQ+yWAL/soY5xhlkvY0K3edpGG5nqPbRTD7JF2btY0JneLPHfYWy1sSm/9u3GaGGbutp4q6G2f
LJZ4vIevvb1H1+E7Pd1ggEOMlrefCX66ZmvWSJT54g6wSZO8EV0/ImF785rWJhZXoGZy+G8QuYzR
wgcCIwooTXfME69BFPocSYXk+9pMJjKheFWmPPP9Bx9XWFJFqj3+gDlK9Lbj2GbPP5FCmnf1EfOc
CnN/gpKqaZdeNSY2nDx/qC3z7l0473Zp0EYR8vtAY95ZtegsrEH1MXPbQKHoglKP1SIK8nkpYtIo
QxAU4IsEO4PDdug2eDtveC0Dd6wHnKNLbtCLxq0z3ZnkzL2VIl4uz2rmXRJvTqvCiJkZHCDgI1WC
GjeGHVWVDY5fIWwjB6zBpjQWsMk52s2gODeeVsBn/C3AGRj3LmORy3y/fnPyva1ehLhtOfrwcrxj
wbKk0JL+Xdd4ekhXqRPiyOBL2GXEcqLXvDDvV1GgIrS7dh5CFSGM98oPbuYvrWdCZVO8VzCA9Bqs
Eg4VlvIV1+BGkVBQbfji4XV7biJtWmgUm8um3dUhohxVlLODaUdzQQGp6Eob2Nu8R9B1fdEFozyP
MX1lwZKhAuRDSW1gD9Y3m7HNL5vrzoTEQAKI+aSIvAadcLxZfV5EF4JLIgx4WhQou4yjZpSEnrT1
l2/sMivxVgeEX44HZfv8AUmZYbyFr83p2lfsYlsz//uhYPhLdCou2VPsRz+Tn0DT3k5XoZ2b+ktF
rHTJQO3XzDoihtG/3m1wT+RTJKl2IKn6R1lz0bGiR7yieYIKY7LB/mH/XDlzkgqXrZ1I8vdn+J7A
GhB5lpsRXCoeRU7qj4x211HoSiTRRRHGFf9vDeAYB8mX93CEGo4RSimWxNqbqS4f1ZPTeYMHt7fB
5+VkWjd8MJHALSMCzda57FQjOak5YWEAC+0vq5J5mCL+nvS1xdajbLYTh7Vwk6bRibz7G57R8o/X
SM6NhOzNzTDrmXNyLnzlPZ+FVNG+NDyiW24QS9EQodOzQEbINbGnreVBlPYow/tXhRB+wuYlWnsZ
kQajXw5hUjiIpcwWNG3zq+mBHAo3HoutNioEWrPAm3s4p/d/ACnXtniXAWlnzCPnDr8tNr/3HtxL
F5dzegBAKTmGMCyzp528p3V3f8hDYJq2LXM6OCZanc+XstJyKUfL8h9cT0VM+0pKAiO1gvZ8PSWy
wtmSvLnmgXouSC/UJsf4AM5wxCFY5KNZ+FcrEqNxtJJhSlvAucaEQDB71vIv81XVE6zESi8vDKDy
dNaFzuq2XUS3WLFxnrZ15W/RD2NH5k2jOK7NxgF64BTjQmSNjQJEcen5Sdg/McKqsCIjIX9zWUQ4
zoPGRV4TG86SCv3tdOlLcf3tbVfaz47zQSliiI1gaWZ8e5kH5CEjf1RYv5YNRIh0W9IQhQwudm4R
TtC8PLAWVP7SRngs+iRbBmWp/CoCqM6JFBp2Mj4vuUe3hG3P8dOys1T2JAflUo5TMsxLxjvfR2rB
GBuvMrdrQ9Pz6MdTOxceV/5tgQYZXlNNcgMlwgvwn6eRP3la7lO0NIF98xqXxoRba7s8vg8TRHwi
uhdUbtJcB5iT5hIPKfVh35QaqdqDmZ7JEz3tYumPnGGJXMe1lZ7DDZMv9xVgI1f19DHVAcbAjT1p
kGqSBILiodMxAeScL39Hkm5Wwpq+xbmWI5oHwGq9chzJPSAdfBm1GYvj50eHzSXAsuPUohYroqC7
mpNAck84Mz6RqGJLYQnIWkYtawmQ47R1owHXpwV9k0QkJluwOze9vmiPZrq78i4oHLt+OnSOGIc+
FXNYOUraQ/ruNE1+3j8S6KNvexfQcHMPntZis3Spn5RBupv2XbkZLvXol+qT1JIS1wwXICZznCFT
HZH1VWYC5iijjCeDoQLKhiZP9OzmLqku221WAHddGhSolqZZPzf9wQVIyqWil7IRSm2A0VEnWmrb
tRvovRCUbwtF17ZN/FCL7o5KPgrWr8HuKV8NoDjKONOI+xH5cQ6s3MZVB1JaOGr5sIY72k9gMB7j
ZPQQkKhL7RnXweVQxw7UQK2cjRoT8dlM53qb9U2D2X2JLwChF7uHZwlyUu76917qtV6+zcdH+tMB
7WkbgQFlt4M3S6/lzdw8pi0GPZjsXfSvoOPYspW2tA5e2cJ4DPN01LyT5rmnHvgJOJNRU6z8qB31
+tonrvr0N6r1uJKw6zMepjxKwP/H/USfWyX9dLTCmnMEqiQVrqRb7I90iXcyJALS96sNmXxd2qB0
XXf6ax//3bKZ0hSuC56pgezFJMHlVn2c4BHqwpA5yVkEt2pZsn9zZYythnMetHpY+MsQc5DVnPM8
Ub3KJBXq2zpxMXW1AcplA/NpoHCT5qe7VcGQkFPdLAwT09y+q2VCvFuA0qn2dNEZOvpTAZoL8kQ5
olZH+RvauciDCx8lqGwCu/eKAi0bWzt87YTSKG8rd49BnS5Te8Vbz7MxREerZwfM4wymAmv11DlN
c8ngKatv5SzXR3238Q6FpwZY66jxAGbRA0zw26klW0Z7R9KAl0AFKWOePVqu0VG45nRT+BwcM4z7
OR1hnNu7bS9AfEVWV4wqsJ0EhSAEgei5uvJMcIo67oRr0TF6wm96AXktxLN809Mln/F+IKEGDyNJ
KDseNZUi0p24/LSyR0RhZWv6Koy0SDVBoehKsYbhuSMDEx38idneS/1c+mDOR1P1EUiTJcabtrg0
lKkoBof+8t7q74Q4PKLlMH2ffy2AQ5bLv2IV/ZzM0QeYEesaE/+vDZ0+Ysz5XdUYLGU0p8AH1MZY
+roiZHPlj0PzyMmc13uu/4et/DYyx5XlPv2I9FXpSEhl4VR2CWpkj1CcRg3uNUnaj+z2xo3gkM7X
NHIm8AUsDTb2wp1pSzMFuR7uqFnoDxMZ2r3JE3fymLjc8IDTApIpzmgY9VUN6YY8cGNg1bdJszdH
gpVmJA1tjVOnERyujIImdtOWCFRmjYxNWQfXipH9zDa0zbQgo0iqkPrCtNSeGWeVzGBKzqzHQ4hL
UxQb1QXdjqf7e1O3LYzDqL+S7B+v8powZmsj3sPcxi4htzBO4dJSEsrX2BCYFc8erqzH7D3N+bdo
cBpa8E8fsFrExVTjAWgOUXchuk838UZ86odPA4SJFPT1h2WV9Dga0wMxClNJ5Hotr1w4bIjesJIa
yZ9Vk/X8bP9E2vUm//HvtZmUFXhE3LjrQ8zAPfCl3OCCHQofK6b7a1TffTRllc6DKaKX/Kkc6mTy
djog+uPpzxuNFYwua4opGJZd/pFeQ7/7KaghhqGVdOH1y8F5cmpM92pMuDxsUG36LKPRMUsAfaI7
DcDwnhuffDGgZY7WdIcKBlb+VGoFPTLPuG6TkUtDzSvCgxRt8vz6QU3hUrVEQq1u+lupT5sjZyIu
TwrqQa3E06rcGI2nGfyxUO6ZA7JNe0fRBOWxTY7lJ94Hekj1Hq9ri5k56QddrPeM3j8H8jNeclU0
uw9oyexgUevlvnm5D2XJET85vTL7+WbXdt1311PvkRjFU5Qg/v+juWbArYgJnwyykVLHYwwNGWDJ
WsefkS8rT1i2a53x7qJBn8TQDcRvE0DBFSXqIEg45uaZ26omkUA/w3Id/RZJy4zn5Gt2Sg9ZeO7p
62U8B9Jei8q+6Br6Z3mAG8xIBqR7tbvp0aipUd7oWUWBblP7VogvYP2SGQ6AAzjPMPnMwP7Z5s92
E9ES9KE5wOGlfJptjQCIa++IYwFCit3/A9GMDdhzDrwHElFLeBslFj19KeqVrPspAzDDnV5rDbm6
co/bkX5ZeKoEAEq3t0cpPVkP7Du4ZZz5m8zJEnuu+ojwM9Ibqg3NMei9RxTtlbMeDxB4Uz72xf6i
Gx7+ZRu1EQjfXYgTQoxuHk7SZNfntMoeOcxzj1xNoL42es1/MgzrlK0LpPTVA40I1H2sQOpHK2rP
1n4JR5BDTF+9E5UaKekxi9KQJ8Zc8TYmEVDvB2O0B860zmWbnY2kkCIYzNn2XSSAZhvXz7rDB915
vTKQ+9cYbPxaFDnSMWgGurChqwJkbRyYEybpnsejYH6ofbYpH0jyr9k7pgJWOD/f4KmVNYey1UKq
pOmM5tlxnDlY3UvYrKFFD4fFFps3QzKCP8ybqhIEcPWGm3WNlXAASOv7y33xLlqKDD8+6tzCqdaZ
kubiACFdthOAf4SF74XLiBeH8wX5dd5tVF3o+Krp0wnsmfyzYch0qXWo6ujw52+EizZQ/kQ04B8E
TI6OaU9TctOHEhtuTsUS9dYNxNWsX+pGhQag6kq/nAZn2DqTKHqzgNgkh1qjph820TkUM2Do7Ozf
QWU8DAWHHO6JVtotZCPaSVuRSXVF/WKPawrVdiKYHVb11B4499EeDZmd2ZZ4UwQmH+CzgEwpL9ZL
F7obbIX2hjR9U0TkANJne8kg2iLq/NSmg7kh1cOM9zVfNZVPZnHruaQdYw2xkmlDAJ/8qll3thrU
aTN+VdAEihefqstsqEAnF04fRdvrOoibXti7Pk2jXkeeUl/v0SVlLeZRHucXyXpDEdo1Ib1syMiV
YcirYPqsHspsRE12Rdvb7nR03/4eYKroQ1dws7x9sIZf+Na2r8fm7MvF/sVfeWGIcuczQ7H27rKu
3XPAi0I1vrmjW1u/hGrVNpmpR8EgFrsiHosw/eWTB4NMNqFLSzdFg9VW2hRGEJYHMk/GU0K4fnve
d+Y40ZpswI6a8ikEro0y2+mIB4CRytZa+iDG1Wp3c3vIGUF2uDpEQHjHkNsMqzRY8jt38TMfZiKf
FggKRgOh1yMjdtDYY12S63kk26eWTZTwbaE6tTH+1Uoy+xSX8Z4mgSsdv59OtZ9zrmC3DhBskiLk
3n0y3MNnjsV7X3cVQGn6HGUvj1+HwpkiDOEEVVOynTWFpldq7vESCqaQe0amm0tP3ZMdOjwJ/AYx
NNSAcb6cYHuUyNj+Atd0x4iF5bkomLEGsXM0f2dXyEOAGLvUeLp1mW6dhxSP297EqJdzObtnamJw
wHR5S/o3Oxu00G5sAVfFKXmQuKxFnD5qZxgrQAiJco/QwJupf1X1P/xHck3Xcn9lYtE7uOyIA0zN
753UN4wbFxIvrac6I54DYMPwVxdcpkkA3TD1zWTHKAy0/8j3wSabVl2AIKDjWuBYi5ZIihU+h8G6
P637pV/PQfVhftM1lKDy3cWbKhQiYV7bGK3fAtVhAvCOoVZ221mA6R5tsmaMLfRgfX6Qr6Tq1t4I
4/yiaICzvS0DpJG0FPzW5w6h5ZdWHgrVeMsrJ9Bdgy2CwtlFs58WsdRuqbfh3NSKXA9lnLYIwnnb
5Vzdo1QC/yrGAmxcb/gEboFbkAOSDtUVC7FAdkRmrYwgeT1YIKvJ4MHnyi5j89HMgvwg3JcmZ/ch
pfZlVdmfC8mGmzbQGvMnAd6ljTGn/xFjuBPKikQhU6aNNQmM3bDpX/IbpINKjVd7d5ZiPq2+ow6U
NoqivOnMJ2S6GKFPZqh30QQEBlqSb5ES0kWsQnAE1V5yQ5fe8nbXxa7wVY3gnC2mqnNSM+nXLIAP
Mcbag11uK2EOdq0a789N57uCtiu57nQDQbpNyx2ObW+wAd4L9uBBPMXN3EYvL2OyEtrwejausYaQ
8Lj99A3hHvlBZQcsGX8LvwfPjFAh6IP2Et3DtheAsfsqQ9U/r6R/UB/45BLnRy/tcumFCzTC+m3f
gRm/M76PUrM0suM4hJnh0Ab6icWr6FosnOZf/qsqPvft0FKxubSk013sJkJj6z/mXs7aGeWD5UuG
1XMMTWCgOTlLvqIhcBsB+wzYfHxbvB9mDXUEqeZBqOKGWB8ypL7eWg7tcF0XhKD+7lYAfh5G58EQ
B3lcaxNoGj6Gz2+x6V12MeQV+vn90GiyfVPVqPnSw93QHhd1oMmHrpaO1ErQCvVAjArhQpoAQTjX
mK/wmykOrbB4qepFmHL/yAq18rW7P1tV9d5RcMgOVUjESjiJhrnXHeCZLuMT7uM5DjA62MovCOSX
/LQ2lwxcGd9x5DjnrN76PGuAhrQDyvUCcgHCiOBfVzaONHiVWPd5/FwPbTOiyFWEnu+XHbvst9qJ
wgOLzHl7q+maXYDBk9poqyWIKyD9WAo0I147EY2pXEtgo2xqg4qCYNb+UytffufXGQ5jA4PiD9AC
TpPw1aY4W7sd6jQYE+q7MOdoE7aFDhaXduZdWIwvnKxMj6xPf7LcVmMoY42bPJD3KtZ0jOXE4/Ay
G5NuPLRLqCtxx2kDIisNsn8NkaQKVlOqe6glmi7505Ifgv9YCbkjAX8aywG3R15q+1c8br8Y6UBE
+aH/+T+kex6h+QkG7yKziGZuReVvckDZoLbbn3tp7nhMRaYLiZHICAaUiJI5LTNW95a2FvvY+hNy
CRBdFzSgPOANaiu8J5CjQpSzuwqj6BE/xcM6SaJr0foT8U1OyyeM61Cu3pYysQ+HMxZE2AVqZ93n
Kc33j4VnyDtiOvdl72Es3SzITdtOylDXj+gx/RX95xpEs7xm2rcualWVv9WHNCBOnbnS5hmTafPb
V8SA1uN0JY4h8Oh0A0rJA/6qaDtrzLZSba/o0b9YZTEr3Vfs8DyofNjJbNC8mC97htD1cjOTO6H5
ua6Pe1oh5oIbs4X21KcO8HWuJXAQeXktx/8kC15UtAfj1ZzUzMPtU+FHiux2SFIzMGzJAvmmTEyp
RcYlftXwqVsFjr8CtgDbj+/dAgMd94y4Prsb2kTMra/2QsJm2ltNqYoEYKbEEh0QvCWP6Mq4AcYP
YzPEolbUgWe/mTnHTopk9Lj4NP0jCBx0c7YRRtzHuTo0rtGhF2fgFWWj03BOqFv6vuhJnwdhf/oM
1PYJ1gXVrcxNiZWU7O36NhoybwYASMK2eKgtEncGBqefoRRyK/WLcLFhN66SRQKlhyImjQUbu0iZ
sTAn0EhYm9PLx0W+j67eK49iHh5ITp0f6fDn3lMpgtBD5+qVNPRO6K8djw97B0l2As7kmC1Ipx0f
WPXwNKm+zZat5fuBjZa7onNPmihfa0YQvAIPrMGlJrxp4cmmZP7iPC9s2+Pk8gucHJTzQudnh49d
QUXyRFndJPZquCKY7mwjq6OHu7IpYn/BCg0R3Fh/c7E/kPb1Cv1kYN6LVGCj8CvTARgpxzp1bHqk
qCAiJKB0mxxyiOgr4MM4v8K8sTuRh5ZZy9uaPfrtDTBUofwJBbeUjxfr6EABbbRBrWtUfnNcuhOU
miVY4LJVH23195ZbQ4dIMYvPHWWLh5gVzni/CC8LDdwLJVKPWQFKaB8/gfMNIP3S2UEsAJ3laDYP
6qPtibd5cTcCIS7rzZNDCzUO8MShYsPY+Hk648E3V5pSh+j5CV5xWt4OSfghqhk81zfmlbpdKko4
6GktX+8rvroyJeecTIo/PKmXVMho1haw0TDzBvoJtbe7Jgb9GRkgi0qwCPm7kzSqU7yB3lC9gi7b
iYOXCmOY3v0fn9gTmHz+tUG9iC9Je89uniI+QMHVIDaXeccAQkF7wNUFmOmXncmEb8Z8jedBYcI8
bhytY+njS7JifPzIIyzfNNk4YswGsj+Id7CXCtaoccxQUzNo8iBkOrYLzfZShd1sAacSNjDbop8B
jP3gALigFhF2Gzsos4HdwrcKGYaP8LPbm3klBqg9BKx8wMh3wfiBk9wpvr8+rf69GelsCRVPuXZP
diCWUzJVG31x5pmczjIH1iKQFh+qs5xJN54EjFl0yRm5UlsUmP4a1LnwS+fIlsbySF5JZeQTkgh8
AVmKBmD7w37SQJZYo7AI2SD4WWnhLbSx3cUmX2uRAvbfxZu2bHOc4Ng6I6sg86bb8CSra8zQtVYv
umhJSAwToqIybnjdZs8veVm8zuL8S6p/1W+FZS0qXsTfgFujMRZhL6aLVQ9qiOWLtrF9hyf2wnDd
TSErnYbVSBx0W/2Kg6erXDfQrxDYIEvCn0nTW7ePWxNvqo3qnQK7XLTsn5WVxkEiKkgWfkneSiCk
D/24hngl4IWzBhRgaAdZK3dSnHGhtwB9of48Xr/tVz/f5m5ktWywarKIZeUmGT1vjU1gsfc6n6Ss
AzZM61cWwfFIE1QFZqRWuVV9BseA40sK86xbVLCkMvAB2CnQYDLnfhblY/TIESsafbNbQ2o1gVsX
mEvTJ80OuXBBqZKZz3AcEAkbLhrqg4ptxdhtdkq18Py3BX9jHEIbbhig8AV6erbNEzkfs0Thhrlc
AwkXgd+vlqtRrAHCOCakdiFCQybVAR/gvT+MqtAEVOtd3XDIyz0tJtI6a2z8WG4TFqjlU7RrEPW1
bOyFDw1We1coauoLUEazBLeU30KIRkpNWzfD2la+V3FGKoqWFcBKb24eT5YtwZBJraQzlTJLykA9
bg8gmm4buDL77caz3OnT8wvi1cYUq9zZTwN2pYrBpKkq4FgkEh64RSqQl8X23kpwvXBAy1b6NuCC
z/I2sZD0nCDRbDjPN0X4ItCYXzLNYvY5VNCRGGiAoOe2AW8uMl3ehq/KUF9JhTixVzOpWS2veBBB
OCcm/XNjo1EPWkwHy5esrOq1BYzB2WFbWrJEIh4K9+9X4Ty7si+YXM/vtoowAl1w5VdWg9OOV2e8
YDhRaqFDeOru/BFWRv9RpdFEhRhQQLjW8FVDDphTTK4+cSR0YWndbpmmlwSpbuCjUq9Sm9lI/0gd
YE3RGpc4TDAdI3aZQqii6EBq+eYssFnPdBSrMB80VP5CtXtjEQTDuCQOG0GzRaj0fpi8OfyrdN4d
Jtpd3xJ4EWAlPz8m2sRfYjMmLnzHzaraRiSgatGyGWHEuORb4DfuN/t503Rpu9goMIRfEpBO9hjq
5T4THqtRN3u4wgp8NG71amc94yHxWo356+2M5JkE3b54Gys/Bc9PFIKu8//yqdjj0UlKxhRVwR98
CTfLSurJeXEvDWG2gQoaqavraHsDN3FmBTMkosHscw3Cky4H91FZ9oxB5yJbHsA99Kjkwfe65zao
w66kZCWpmVKIVkyssMwnFNSrjVEW1DDBWmoO1xaHpQwAmofAYUFiMStP+sechnEBCe9f/SgJg85v
p7p630S21rzOd54OPS5ddEFWv38ecefQ7LTlGPV+pKg8MmXBJrGUso2Y9EbLIHX5ig3C0dwnjyDP
tsYF4LEMhA3RLk2GngRRIL88snFSdRAGto7nOWZDFLSztAI4qEOpnDuTvLiEdv4FukZystxI/SUT
xVjIWuQnn6Q5VjscPVRW/yfM7U46ch6EbYj5HmWmtMvg8tDUomdEJ0kFFXOT5UBpaJrDBYhqfZwX
6PfMAlMb9PLgo9BE+EFEeWuxmzpdRg4SBrXPnTrbMawA9JCNsWunX0ywr5rFqUmXkoHvEF+Q+MQ1
T+pKxP1xkivziIPbyPg01BYnoTr3zT1Du+PrCd9pgu05W+F7OsDueDXhXa4cVHJaZyPkpY3ErZHS
wZUpfRABR/qI8n/+64TLfhpC7Y72c4ajrSuNNRgNKYt1W1H05+dNO8TOnqV7rZc1cvLy67Jl6peo
R78yvi4kP/4BRXou4s9C8fcXQrOQnv+Bi2I3nCcZe7ZcES/gZSl0RfptRqpA3dXTZXJEHWKyGcLv
MX8/lGvhE9WJFQ7kqkVHWrz5ilnlAirYL76rfy6h+gFtNbSuqYBtmCcQa82feSCQVUE5wA3hfR7P
XFEhbyYSuWdcreYnWCP2VhTrfp55IqMKtjT2j0hDigyNcvVB/NmYjY0MB85afVbJJRQwZfW7OS5a
q0SLMm64iOiH7O6IVQksW9xWxuo4zC/nrj11CubPlTNELyoQRKZ4zwHroz5hfm+0ybItAFoSimk4
zKnCKfKlb+zZmHvZYw0pSNGSCuPYj93Ct12bzCA4ViezI+29TYhro6dIuclR5dvvkDxNY9nr3k5H
lrc9ujdn35llakbAeMVhP/TsdvgbbYdh9W71JnJeC8mRh4l3UX4qRVlycIKoEp+W/u7hzit0soNk
RBFkW862uGub9BD9yoh6ie+gD6JDRgMZR/r3k/TG6hzIvg8NWuTCpEMq6xncMLjum1ienG96ri6Z
KHyGxUZrXAWtSlIaUctSJ6ktZh9VFv4AdAQuXXFS033JHOoeUp22RmS4fEUSAUFq6Ld2eCv45sup
/6OZPiFjnJxeiHocRUJakeRDHB20Lvko29RwQ2I1XG7pXoMtW/uexdjRlygIvRq/R0Wyg1v98LUk
I0JWLSSjKjkGC70ZiQooFLplY2qurCN7OuWA+F22VN9IzZnzF6Q8wBDmobq9iCAXkfzcnGF8qvK2
aElpNBeZoegG7ouVj902CZjc2b8QoqmGox8ojJGg64OfnjSR8076sz9P+AzHteddfm8In5uLqDew
1Eu1eMPiq6f4gpXEKznC3fp99CPr2pvN9Q7ZlwEZVSmGm6VS/bLn7IMY5dDibf0907oAy1dzG7Ki
r/b/qCXaFwSZ3NAQDypaW4iKyXfT7NPXRYIThQcMtmaw9sU5KC5OGP4TgUVMvb2D7Oc7Hv3t0O0Z
6V8q8n1BqiRNlP1kCJzvmm/k3iuniJku6/dX7yrHH3NtsIeJQckSdhBsYLnPephcIn6aZxhXP4Nw
8aOjwDzfQ9EoFgIznLl8W3dCXt9CGN9e/dGxgyGI5/9wS58FzlBLN0UDgsP1NiA2jH9qGfZ8H+1g
XFK9i4oWDifjh5OOmJjmV1c4byJOQ7VTJa0D74jOHVmmxUa4DA/od+uRDZvV4VqumSjiLOVu48PT
eA1NUnhP5BCdQwWgWvyuQb0w/hT3Ns8wyx3Eb9S5lt2esrL3WG7TJhEBpEVq8AlFqe7gvIXpF/KI
ZPxnzS4OfpgTO6U8PxXxPjSLQ6Vcz814TWlGeWYD7Oh7ylSun8PFu/+l0bLZz4VgaHKF6g9Ux2iq
VrARWvafdUrtvd+oo3G4qjXif5FMAIHHDSniRwNH9gTmvd2y5SZq+O4fgOFeenhmoI/qwXkCxy00
Xd89qJHSCOxqmoJ7G6KXmCr5sP1k7vvpYYxrAzCAIXa32dKWyLwOiKfOtaqzmErEXDzdaSVDX8az
oa11Y0d6zNiecq0F0Zop3ka+ZoCforoC4CLNju7TeT166r+Ga5AIqxzMc+h+yD2Ab1vMPi6us9Wz
TlbGJT64D0PE2flo/hkSR96ecsoVR3UJaQpDNkRfwjCibVaIpEEsuXKrKlTdqK3NkQ3gxJv06P4+
qO/BDyV25D4AlcxHjnGzY8fZv7P0T5Gl181/KhrLCw8FAz8jlPSeC+fqWWTxIHHfIKaodZ1y11cQ
Oe7tB8OGjWhYjNRgSWfrCnH7iM2zYeZIqTfpJtuRXNJzqCFfrSgfawap1aYMacx7D6KWW+1Tpu6q
lr/ZYYAKb2rBBFJjOiLLhmnR75iwdrVGWurMYg/KatNYLBGgAtAEDVrOYEkjyB8SvbK1c6NYbRLK
NV3E3T//AVCV0nSjijAmyHoD4pnXgtSFN/HkeWjW2yrbrHegPIogPR+D7vEtlXHgOCgb7eQE/R73
N0a160nafH/oeqHonE4LXL4rFJP/90BpeiKP93dkZQGLBm8UqJNqZ088tlrNM19bJ/d02OKr4IzD
8abampnTUoqtitJhihksxn+dmkjTlb6Zr13PbvLPFFbBrqQFI55O1Fzm6E6fXpIvpYnt0UysSQrV
ev6pEFwk3HqAJskjwYTbt8gvZ8YiLwBesrDAAVs9RNjbrli31i2DWkRjSM+RGXlDDuADu3Z0Lpd3
xdXeOtBZCQ0d2H2cPClIQgmu7/iP3DV8PReg8bAss9Ckf9HSmW/GJW0cM/axldLIrLjWEFGj5gbj
3rCHQDvZKbbsfTvkf3dQ+zfWR4o6JanYtFpxZkDvhMsnYRuBcrvHJTpBfvLfKO47FWFebF9Ia2Lv
swzERtIR4dRJx5SM+r5IKPRoR4f4XkU8ZzAca1x2znWJX+D0uhxcBl7Asv3MVI6YYkQnzOgKKgYh
CDLpZK5JWtOcyEFQmwwBZ8HAIQKYH3dwfTk756ns+VVuiIoltwTtXzz/eloXgmAQKGvILmCaHjqq
yUIawhU1KscnLtiyEcL0cFYlEt10mZ/ce5JtLVnj2IaxMkCsHBf0sbJiDCXby0k6pBJXKsefjtKD
VjiU8D73uW7bFvG+jpvE4ppehO4WzlfA8mRpl9a9+7b7grOwYQBQ8mU9fJI4z2uzll/C2aIcsG1M
jj9U7w13kuok7BoeRZWyv1jz3I/7ZrJ81UqpwHnLqkM1hGM1Iz9n6I2L8MiUOOu3RH3XXjeK8Tkg
TjPxzpkDmbK0UAy0M6wU+6Jpgbr1X3ADu8dLKE4HHk+yQFaoLRM+mp+6WjxDHE6rZji4EQ2x7OBb
Ye5GJIAj5aejjcpUrYXyPJd6pQwfBuEAFzX9jneNgu+nrXj6kw88gxPhVqn+L5Ne54uyL4ycBpBJ
M//nbRyk/4I35fOtupxJSeUA7a9e/7VaVFSnPkhkZ81XPjGVplUsIrqnoas1wnJd5ILzEaXlhoX/
29LpsMZkxphiwQ81vOyKEtXdKIgk8lKtHHMbaOQ4QonmPgzMx0ErcT/Rcr6/I2M7s7h2P4DxuyZa
UG27aJH3m6smGKQrJgReJkck/WL75pZLBvpnCbwAyGYmixaBr+mFFljfA+/+vp/EPpQhKSnGxg+H
I3SOF8FsmXog/lKM4P4v4w82r6+UKsTPtx5IWCmE//fdYdPCPrgLSzCd0EhMG1cV2Jc+39ZJlSg2
g2aRAczAebjNstvgEaS5WegLqGw88haYDEDmI8vCXFjBLF5pX2OHN/afopwyI9P//E8btePs8MD5
md0kS59lNbWtRhCmbQygGh+ILi+FO4vI4M8My+SYGb3gUUijkAaw6mNe+gufYr27+Dht2lfgFnxU
4woN4IniR80S66i+YmXTckUNV0yJJ/CEdb9I9FRbeAjmWdzk3oizT6iXFMOfrwM5qpe0Ef3jdhOG
3Dwl03g7xT31fHI1XgwynmQKj1TiA/ypgKYdxnWWrB7AroDf8iInw9d741Fk6Wmma8R7EcICB/jV
LyqtoaP931Dc8dAy0oJ7x/95WYuBzl74ERoN2H2Lzp6hI+dekSVq2KTTPIdeAKspwFcPKwNhSarb
C+n9uJO8X58ihX1k/vbcbZvzkjdua1IMI0WWZOTiezrEMKO/MxuyiURtPgj9qnG0U6jfBQXGjSD0
yyMxCfleJ8OdPYcXUkb5wxWnZLVPFjqIvSM0T9AA7SE5UDWB478XHC+zN3aAoEjCOghY0sCWq4Ro
GVb3u9ZNI5dA0GTnmpXveNeDm8LRJGZw+OtNHq6FS5s1IClDb2MnfibNrhd3jwZjZ4J/yMMGRUF+
rGUgjIabm6DelYQvf0rYF063neSj8zCvfBs/gwftC62JCEKiNuug9uIR5clenZQ43j3T9vaarykr
wvAT3pu0Chhjlm2NikiCc2SPGF6oGVM3lz7suttskXoFqTIlOlNv4gXBsCLYSDiyTtH3VZmGQBQQ
+xrs3bGFwzk4LUud/PeQRuSZni8HEUEb/s/1/l9A5//2dmiXRGHaR/zNIcK1XZKAcGHxm/l+dpCX
NpLdlFi70lWFTgtLABO47Fr6DodCvm7vV6/sGcAh7eRyXTIlvXMTnWUN0P+SG5+ZXl3HM2vqHWTg
m2ePuTxphxMs76dFn54NhJT9YPsKTlZdY6jhcK/HOdDK1quCUkdkQmdtuuvDGhcIEDlnofAt5aXK
AfqeB2utFSHSVirvdptQ9hCEeTKbuFUIl9wEKDLeJrqwIDqrcIQ/Vba34PHubPjiXWCoBBNYeD2o
hJIFKU+uGntktwKyeB3DNOE7XQigXzWlf3zK4HgytnJGWtzkXRqU8I6iRug549tqhpMUJxY0KC6S
D4jrQfYbxxdMeC4YF0/blX7LZT9c/ivd2+TbacmbaBNri3xSjUYUkNs4ickEU4g+NgacF/zq0oWj
lFkw+iXQpKe5KFOklAUqHFcdZ6eHRvoc+Xa/vYPnQUQImmHVjvHtR74BLaALBB/lCGqsPy1+Z9VH
L2R48ygqhFO8JxpwWmL1sAdhwycwKzhmvw5+vXUcuY4rtKYI8NG642uCwU7DV0ydpUHxnQHCdvpa
WFlHFCs/ZhgB2jtYyiPrDzLRgGCLEd+MMNv0tKleBfxlBycjsPe56GieMZGkOM7WB542KtadaV9w
DPjHcunumQXGtOr4Nuptqokbkv34O9GHnrE80bUuxBhy7IZF1IexTkIWuuST26lPQr0e/7jjKu3n
crKYQWWxCTDPRSrM2ioHH9ETQfNzsINPME9H0lPxAfhWZo7u+cdrXDBVpDs2Cj2X5Af5nMHsUNjw
9Qk37pUXRig5vGFa2v13xhl+uxFkKnQUFcUJBy+rBXAtp86wNj9Sva+/WiBKR6jun2hJG5wVPsHA
V+tcuJZ0YZynaFWN54O9fbnAWk0p8VvOqpSUmW8Js8tecV7h0+WyPal+CegP51AYl71kVm6wvFzA
knxnczK/37vqQjIrZSxT84bw1QcChCxoONSOMsAFywSwsytabqn4+ENIwiO5LfIx8sHiav078daH
oQt0HHsuC2IkjXCuLMYVXFzxfiLNtlPVlPaydI4RFteI/MqvUnHwf+v/8n4DoiAoQakRD+JHpN4F
/kHyN3l1Xv1R6fmk08efXqg9+IqDRKcPrJRZS4lglRs4GXbRzOV9qCpgqGIKFCNf4qK0ueyDhjBp
oM3vmIsBRIgfYd2tZAIup1X/mdsdOPSyeuJZ94dOrHbMwBRqc4GSt9tPAGyuhCyKNI36MfdITObF
nrLFvED0yIuNlccOdL83X7Cmh3UDTgS7GRR+jFzALeLner3+NE2z8uqXcL1Gj1UywJFUIgvU44r/
wcyi5UB5h20lsA56R2V4wfKeqaDgiQbVW+HFel1yTCEzB0lhnJSAs00M6tNCz1kAj2Ji/5H7NPoo
ZQTdjbz1dKJRPnQNCE2CsMgGzYbTdvSeYAV9doIOULaduo5sQ4G5qMKUxUleX0i+08jxKj/Pzq6O
82mn2XEufj6B84VOqH+UpAdmYSSrf3HMrsMNKNxs+/b21ip1qWIc+za0pGaOnAnJeLGiEHUxp/V5
Ty/XKfrbfy3cB2L6wEPoDL8rjhUEPFd6D3FJAkayxf48DctNLd7XRLfp3fZmA3WaSxqLzs3Khr+S
7kuUciytJVObNgzjQygYqT5XaVNYsr+snuyQ+sSr5Y4Gc2hd2JLDekUaYQ89UtG2BJsS/o2HmsgY
aiwCzVGEWOqsJKw07NTXQk2leREcCtr2GKlE19p6atsSL0RJZZIKpQoJq9Z1FFQ9bu9ZdsIw6C1q
dl+ykuY+ZqK2OIb8b87z1i5kKPB4CznAFw7KeRsRC1KObH+nENUdju/ke8QMJbhnoMh+gtvh82Hz
vITbzOtXJxjaFCS8JZ3N19V1nY+6rpOz7Z7KbdQSBmh7ue87OMSzuCrMgt/n+MlAoZISyc4djTzp
lwIADYdG5DSRpYFNtAwouVgh6pH0JqG3Pzr3lK1upoIPvHfHDRNFkuLWIifFp35Yf7LZsGOvjUDj
Pp8zn1GTPa0yh1GjRv/QVaLYXHS3MtFjzzwJhxUjp3SRapt25cnQg3yY4+EbOodYCF5hKUL03ENn
2uGy/qHy6X5nuOPfvD+jO+t/4zeBAHnKKU9dvcqasW1/VA/IwVIlNeDzy9PgYOu+/9qsEKY5BYqU
DVaCD4rH/C15wC0bt0nd9ahvTE1nl7lnqRkf43qU3nXDGDn+WqlhJZXDeSJiyLG8g48pG8WbrGW2
P25+15fiIhGckMTfMIY9uqRnfJCpca6hJQKME5Lu1ON0+kIgl7DHuzslT/vTgX/L7gYOO/boVZpP
s5GOB3N5X750TDR/sksMNAT+b4NJTuRl6HhEQ+dTv32GRsCtCBkounGmqvhN2HdbwrfIIfA+JxNI
XT1RsVObPZbSZKsP/3XysbRL9yrADYu3E7LnY80uzvZzuQw+Y5CNY1O7EzFNBth79iL2lTlTVMOu
SZ7U/zyECDOMwv0IimU85tXcQ4mtQzcOf4yHOuFxyZnFyvF7nBnzmthvHyCGeuV3rynrxiZhHKtT
mwmWN1jN1K0cJcosFiOf3BLk/HPLNmmCf+b/Ti6I9ajDbO1ggVV/oYnbCcE37TbumSi32f45eT6M
ztY/f+qjVtZ33Kry4EOemiqvt+38bseFnA/Q3A/lsBjMQxfr9CJh6OKn/YBslfaO9AVh2p9bPJAu
pJCqypewVnVPELkowb8YUBlZK2jlTVei3EsmB/kJHNkaKl1dQgUf9fUli7SyRxpNlEyQvaVUQn9D
bt3CvU6PdCThP6/JjzxoqxMi8v2qHsDNX1SbY7um7kAWaDbOwXzYFNhLMre/luB6inH6/DL/qDOw
LLDeY75UUdYm6l+ao7hCGHq54tElQt37Hrb9Fud9kEQmIIO+s+nVOG1Hcsvm8pdDpOspvAQpiL78
mhI3rK8LCQ5nqErrX1JKAbMkWANEGGclox7EhcTVssQkg+xw4AUmG0vYgS6QiX7pYB2MbrN+5Tju
7kI/dlYepRsDnpJamziWfQleuP+U0orwfuYeHwey+okmhGWuyX+UA+IzMpOSiMGukXUnK42l4rWI
38GneCFLlptBD0qj+EIubTVmT+bDS5ieTUqUdB0UA4HHjr47ZL0ozBYJvnEGWhfjgz9eLJd5Cf9c
QzbO5zjjAu51wypXtpds86uP3hKoelfzqbgbokZ00z0psSBObVsXJ6M48tLYC5W646wwcI0FuZLZ
jc4xAoWz0WGHc85Mn3MHJTZQN40XKgTjQFoL+61+NPU9IjJW7lcRByQrc/jFVAMXzbflPWEqO44P
/uis+lisIbg1ZrZD12lfnRt5tsyEKnT4gdc9VZ2ilb50M3ZmXPNAupCN+E4G7TxnEs5LhWfmQcHP
r+lXQWR9WlvNQlWDpadlr3bTAwzLdplh+BkAh8FRFJ5cIU32jfCOEdo3IESZK7vDutkr/9Klm1kA
GN5YC/Lv5LD8p7px74zPhdiI6c1cb6ffWuapN5kC47IawlUhUu59HInYqmxAdf6yhul7TZ5C8rPK
uqo4rp1xytVIdYZretW/6IiAIhdbDPXQWZ5OBWsWCQEjcxCzuA2oTd+E2ZOcnPc2BXJeynl5GFPF
qShT6N+X3Z7t0WQMQY/9rDTDVC0JZDJLe07q6eoAeDaEH/iQelqE+E+t1Saa76SEpGAl1fbbVLQe
LGdBMofI4mDy9x8ux+1jgoG2JRhLhJ5CTnvEsz9vDa+7ang0fTWfgwe3SQkIh5VN8mleIBAPkSH/
Chjo89Lzx8kqksoX1Hb0wJkJ/2qexxuUZ94ujZ+ztL0Bd+7cafxsWTSfDJ2il4VT2uNpiWx8rhed
jbFT0Vnqdif64PRCB2ESBbowINtSgSrlzaPAo5huB2Dc30Z2L3D8ZvYqvK5pyhkTWJ5Apnl+peyg
9X2H++nUrCubA4AbCqkJnSzSVJ2fkzTo3/gHWiPVkU6CS73OoQuj9g89W7+xvFCr2ESPYtFAQyPx
jtxG63MZQvEBHkf7OqiV42HCi9bZLLOpUJvOQ8r+V+qR67i4SUlci8In632eiKasSOExOlxBzOWz
3qICDjzjI8M67rYlTtYVywv679ahYHN6yIhx8n+n+eAxKl1zYumrVnyHwhw9CiASZVeJcWPYgCas
J6rvggupTwaJI7GQChZVqac7b5jgBCWp7Sa+YlnrKPXcJ1P8bOL1gFiUT7ZN9oyZbaMju4L/xLmk
9bU0YpoCu1sQNspRSDjr8RLk8edsiJCjAP+XuSSrvaoxbySdaVxqLqd2roLoOJRQWk2G1G/EjU3M
hvCRABvgxRjDFlZ8sK8NnI8kGANV/1Weie5bxW7hMY4WX9Wkd6zLl4xpgODyZuRY1w6r/dZefB/3
IllMSzbR75PD/vt0vwYl17YYzkHwqVVmkXaaR84/02J8z7Ip39GX860BgdgeNMAMCSxdKTnPKr0m
RWXDoUKGUe+Fpxhlx3ZrauEIA4amPDbetjW5xz56298EWJyZB6j0ho3gJWPkoHR4dory/MyFGnxB
Hn6TuNZRjtQ6wTCrQhXN5Y4QsAwSVtkfV0kFwzZ1f7VtZagFuyOy+ztwrDGAVv6En1aFIwxxHfsd
M5dtFSjGW2ObfnTJSZh7f7RlwpIgYwny3v47vTM1GebGY8glcYWmOKz8HeQ96XYTRQx7T6mJSeDY
1ldizK8TnHTdoV1pdXp6wtOiFTDh4e6JD+o7LKnjcF9tKY6Gm+Cwcb5VOZnD2vkix1mRFgME+Nc4
6cs3FyWKCaAgPxEEi3PUWBF+yZ5lKa3wjt8UfvXKjEoJqWCz6wb6tZkFI+6KjLfLmE3YvSDisECU
vc5DbfnWIVhZLb5j42iMOZ3YDCIcCTpNkSatq/NmUFKX5Kr5qa/UmbzLnldsyFrYWK5ePTelHK+e
qK8c2g+5SaA/57ZDo00b3eqaGo5guKKWS3mBLh9oQcAOcYmzETPXJDZKUhgyiu35/mdQ1wYOxLai
uHOMOsKKHmUN7Ue2BRoweBB9LRNIoaQc+Y3ySJYD8Lgslaj9TUuyLcFWCkVb2uh6BkKLjH1OgTfe
j5QQyV13wewq/CB0gYuxtNmynTMOeJ55hH2o3qwQYGZ0ux3KeQFxwmu92oscO7dKLaXFvUQDszhe
9zKFAk23JstEtYd9GfaTktNOohrd1AHSeqved69P7Z4mwN9M1R05S60jaC1VUvKEy3SwwSXRxRs3
K4vZSLqHOLkf9cEBG00hfWaiuThxmMuJ+86hMJSOn2TOM+aluZYl6XlLIiZj3C4593wIOTz9y6gD
8Pwp6iYabl5yEfSn+XWMOvPCDLWsBYBIqwm/4EI5eLNwkooszvuW+iVUHrMDtMFi/eoKDQalqFav
xx3L/lJqKuU5xGDiD4OTMJFHQyZn3yUNjF2EANpqHDI3tbcygAMYXRK0t1IWiSOKwodRgYgKWj9L
EUOuIErpwC0yViM+Y0VN+Mj789fKpIFn4p0Zy+BKz+r9OtYc/b4jTWwcnBQpvSCtOyMMb8z5vdUl
NoKnmLCm6PGSgIk0rXDDFyLKjWlxfDTt8Cg/0pagpuuGKo8hW4yd50f92IlWY0kml2oQvj042m/X
pI7F+TXzEUYgnsH4Yilk1jXKXNuHQguoIaXi/qMjvOhyAvKH2W3Iu9OCUNizzLmsXNNCErRjDgoE
OLFjlNi6LlLADvNSoNnMnFWDd4Kt1Y+yJATDDZVl8PMXiq0l0NwSt8RTGiEZuser7e6l5UmHRDXv
AiKW42/NLNkIqTeDvEbvTIkyy+hbQuHFR0ePE/tucpMfeZLEtJdo0Csnoq0pc/9acuWqEGGqbyA/
jYJF9vzRXEuyj8CqJO/IX5K3u9/sxsCPOW+rItwk8iIbXzTCnu8PTMEu9W70JZUBgMvYtsxzJzR5
7cxW9F3hLo3ENNmM8/jxJpDoMoVlYdDioqjaGcmDWRq+Nv+ascqJ04lvg3YJ1z2Q3yqNLG4e1CRj
WXtXYON6nPUiJDYQIR+CMyn2CYcSa3nnaXCPw2Yh+wRKptBC4hjZO5S2QKUaZIzGOTXstVFdPstq
vamM5qt9GPXaYX2/Z7Sb4UiiKGo1tOhGqa3/RQRwJ+aiyYED7MhBdM62jv11h/WsLeUEs0daM2bj
P6wgPFaE9MhtPeUB2CmXjOgmtjLYvVl4kfPWJHCcPdkyh1NrGbqEP+MRSt+1lCDFC6FKn7ytha8W
C+7oc3WPxnhnQ6fYeEgFZTZm700h7C7RUU1HQQaE3gmC8X1NBrOmu1SRsNF94ZHJuBqayVK96L/F
UQ5zJE2NVENH6GPeNetvVCHfc3dysZe71zXjGz25WqINq/rQ3hghsrUecSjJpN601IZkm0+zJMxV
YNMfRG5XUEkeSAuLIeUbdwGrTEOVXkOdLnpTkSdABFs51oEnTA86Wt8a9hXw4qg5vig/pe1WQN0n
JznyXxC5GHCGSwoP8LJEwrS5C2n1KnrBTyczSz0PQQdBzlRELikBt6mrlNqIwnRadsB4fG+l/QTl
ejO6J4NmD65UTXnP2h/O0wNQKmvj7fYYiiAcyMq/j5x4qEWDu0RUbKC0/Zkl3X1sdZ60ZM0B150R
qFRGRTb/dFkw5aO6hdSL6bClfJqrg/akrmMjs/qEXNh1NnqiiomsVN5hB/NyaWrNQsZ7owirEIDZ
7XX0rnHJONrrf2NpXUuAd6jQXNXCLK37oLRWHDEgh1NxUXy1Zww5dHwQDVakhx458UrWLurqrTY3
jQl42SbKUhGHG2wx5X9qyJQTeXFnIt66KtvG/haYyuh6wBNck6X9K13Dcj9ZOZtKMOSUb9vnUH9t
ucFtZX7FJSD3msb3hak/rD6uXpOL/NkjuaG81JT0wdVzBcTdtTitkUXDA2tixc6gxp7EKD3R+5NN
LLYj/pWygN1/ZPQfwyewvfxnDy41/wA7BQbSkOQULQ/9IcKJihX9QbllxxE3s4hLX9v9lbw3MLJg
NRSLBspcUJ52A3MsUKFcWO/noxLEqq8LcdMDcHaP/FVzeRTVxUkQl1ogYsN4mXz18jc6Kkevyauw
1VJNGCONlfBC5y8E2+2TXFEAbM3nq2idPsr/DU0Q6nhNLBTElFfpFx4QUY/C52FObP7oyCLyA2kC
nyqO6crZQXgj9QdZ6SkxDvBu2UCoQalHkLajVvkkiVrSQNY4o8jbzhtWX1c017rGpH3NqTfcTgM7
2xDKX9f4b84grlojd8NG5e1gRvTia90otAd7JQH7PPcavybkGKabnLpcPq4RbH4rX5yLwuMYPTvJ
qJ06EwW3i09p6WbKTFT30gNpmM6QN+hzjiG6v9bUtvN7rTcrpF371zsFEych6b0kb3mu0bGF1vlg
ieyk5XsknFHDq9p8HYZchLepnJw2tCRwgHl8TEhIAADMq1kfRhcoK7LeXoovtoGR7pZE+eMtfy3v
pKs0zc62z9pAHbhkzX9x43nULR/69r2xITMzltVby/0skWgl79oF6TPsTUdOZqnaz0Sxl/vLCY7x
+deGN0LRrFOtpEmO/EgjJOwzT99HnfJ8+qiWOzWq0vHGjNJE/eAioq0vKQF4e2MR5PwujrARpA1Y
ZjWbwmz3AHW4SID92YzIsYab8UNLuA66mPuuYmf1JwrFADt+7mVrAcae1OfUdd/Fs5MAvNwcqrYK
W0yxKs6plDGACqtiVQh4bX97arHPwJebEhpvz2fqJ8638dlYFr+JjabnmEgVfOaDBmwnCUuimb4V
OZpHI5sE6GwTMn/kDfGPyB+0ibmk1aR8l3W8I9h4Nwwqn8lNkN4ojGgYUT38Ml6t7Z6J9tXL0dqh
AfJXVamEUJv1em+Rbphyqf9Sc/GqZUfwrwQz8vAC0qxdc/tS3735UONtBg+1EUwPrh/EXIoGze4a
BIZeMt9PF39trWziCB/jlY63QjIb3cJLCYfAYBTaOY8hCxhxZ4JaqSM3Cp6kb2lp9boYhr72EgZI
vTRGMF2pSiznEC2K+9tmZzW1BQ5fhMTYdsDJ5umYLXdtsJFUqFHMeIidZfZQtqTD9cTNEzPd6Js2
EcHpt10Zc3nzLm/uVO1B3Ao1oUDxUlwMmPNvRSMx1A9MWVhetKNXlN655EA6hfwxc31Qicq0PtMO
ciBHZj4qdgDfRCTPLT5YV6d0NgDT4vs7NShHS6p6/zyJlMAQ9m+t+GeZRBXr0J7huWostSktzRov
eTF61NiS5oCpKCZNJ1+roA/opQzt4MmHQfBdCaXqDwfFUngjvpSb8CW+ujwWaB/s+Jj5hKc+zazL
gk2X1tJv+pdZVtFlaJKATDnVTOB3biyXQhD7sJUSrl3PPQyCTIPfwqyqCXq1NsByx8qmgE5bZjr3
xH9GCPvTzo5cq8X6woNsDN94rWJDpaqxzbIFmf5tKra1JNcdRAXwSp0XrprRn/ZwiGVBDdy1zG1C
Qp3BUnqVqk4k7poOQmJzmTSZAQdatYUQYx1qwxzejXGx/OtJsE81S0rT7Ymh1ao4nP+siL+cbFao
D84Il7WTqOW3GdWngUu4EzUPSvefKVa7xWFkdexvspqyFWO/Dk7WJkMbfD3w23RqvpE9BO8gsdH8
jrzMghMI/bl2EbWMrBtsOj1q9LbincZNBQ9ayaAf1EP8nSdy+m6zp0qBHNRLV6FE2BdJ0rtMB+Iu
qcwP0+54FIRJjP/Iwv76CKKrMCWN5c//JJpBkHkt55C9pwHpnfqmxirQRsFZlKxiznZiae/JxqGx
XACledAjnMw4K1scWPlOd9npX0tjHdwIYj7BTZBrJguVY1LyFiG2HmGsn0ew1g107rT8Mk4xKfC4
tn+RKqCzcBYnxB/OjKORo/kVWzG+kh4HAeNqZZgyrRujSdJDoG1+lO5hRj0rmONClR8dzALhiDZH
v5lS1uXl7C1f9l9kk9iENLURJ1M0zIlJI6NDyjhLHm2RB+FOmXp+hYxWh1MxKKh59+z+tETgKSVV
ygEvzMqtK6MUXHUBGsGMX3nI3Mofr3gCVdFn6xRtCxmJmw/hBAuhivQVt+XT3YBzazmYxMYAMoxm
bBGbJUGyF5vLT4ymE7O3LhQDDuhjJdItMTStaniv/zjLlSO4MDDZgUGvR5weIpCTGSheYjlY57vr
Ljl+nBBJGgI4Cf21XpLICLcJCciX6rPM4B73tFrdvVLm8d5kL0Hjd8z6JHWOlW1D00G4DvupLKCv
3QxBLf4rZXSc7HH32Zr6GesN8m5rAUsG8zzGlR1mIHpCELlkFbJ6Jj3tneU3vDfV+rVi4p/BceRE
qe1dTtUjruiXhB+EOYOlNCA8N7NOeBoAHeubLc9r7iox70j77p+/p/ixpcgq4k5XcAnYlFtpPN6v
sAl44DAbSYrYi96aWoQmECEouNmx28Tf8nsU5KSn2RHkeRlxKQQkVickJdZ6MGFmGVbPsoJE3wQN
kwD0JT0g0b8NRZR5bHd57AkyYCJp/1P2QLS+QfOG5nU+09scIgypmv0sJB3MZ+LG4PqssXsmi8sW
PG/yRmaU4L+ijx/0GH6RpD7jNkEdg8eg6etEUvJx63G9uAClajGQ8zrxNIyfnamFvQfVZ/naX2lA
3QlMM/dUXrey5JEcbGcl3VBLlVHiqWjQOG47eTYj07km+ED98W1R/L9PHgcRfdzz/7We3fifO8Db
NhWu1qEi6X6Gk/FD8dJKyw4euKHVH2onPhOaWTguAKAa2QbjVzBAh+MWd5EswOpZ+//1LhrEgjNs
YBz6RcNYBWA//OwjSxNc2F4mvhpHX3bskFgqVpixf0jgHP1b6QTdCtpLkYkjpSCny8xeNE4DS0iz
Toyit3NWA9mgXk7EhudsQeKpKqsnsB3xVKRBqmJmXaC4yrUrPMSCDMoPlIgOWvP4GAezhNgo4B7y
CL/8X2K020BAyldU3Ul8M+cq/08TuVfAUoULAnTY7h+aLxTpbvZIloWoeWlo9hinUo1sbqLgr3z7
5XLCJwEPEJPqkA896/8rV0ZjnXussvgkT9po/O/TeUnlsp4hqsaDtenNeEiYLoHPdLzPJObIeVYx
CcXOIt4EDQZWnMxAQQtEEUWzz5kVlgB860gR/eG0Rcg9Iq+YRpFilPzQQgdL/r5CzEsmUPb9z67H
NbTrBt9CcshvB1JTvScl08X5HelFDcckmgJhqOwR3NCyhgH1B+6jJe41vaqwPmNZNhKm4MYz3CEi
8medYCptTq8f3Y9Hlof7y8tQmLTKre+3S4pR0+BKz2OMipnGoOIxGWKJ3mXtJ6iwRj4e8ROp3WQC
1/uEPV39JjB2Qd4M7HfqFkFYcg4Tv2Yvp4lmzVFABt8odtItvA+kUUOU/pItLqvndomqYB6RJLE/
TUS/n4FfNY37LtALUgXGmFHrvtybrSx4/I+cwzd9RDeL8L7Wo+SlKI713CWRyUoLd7fwb+C7AEbY
jhZ43IV9uLVMPC4WD/HFCJrobMnjTRyjMN7BzjquowS6USyUqufRsBPO0x5Py7dVLrgRVFdAmRYc
EGdxo5r4yU359zxb7sVW5nR27yhCUcerDx4ZwR79/kiFf+qa4JMtn+z+X9BaGV+ir3/gxYcBCT4L
gMt5GH6zQyHpBye8EsNK3+zVEt4/C33V+HmzK/1IUteLS0KXgiD/iYAVaeBdZpUmYV8Bctw3kTw0
uyGtyFrcBaj1Vazdj3TFV93rQqcykOtbya+WNGBz+d/MxZZEnWVovNbj2WCqYbeztlabvNa1ofUJ
fH3Om0rdDGk+/soBPId0MFMqYygs8Yoi0KXGFq7H6T3wb8SZIFRxniGRRI+4kEV5b7CY3f4AB2LY
XVhkli47sDoKpqyWZ9uxHN4LvvJVyMiB7SuFXM6Uo7jPMVxXnMpF9hiqxUM2espvsPqdoD/Z5US/
AMShP0ELHI4jb1+zDBs9oPSVcAFYztFktq4gt4uyHyvj6MnLFOcevfKmbYm+ainb/pA7rjU4Q6Gh
0FHCVpjH2T+d5Q8T4rLbGw25XRJ2BQm7djlSYDOBiwm3HhMB+jDTa9W9GT3Fi0VQUOxKxC/baMXP
2YY3qYSNT/XEDsUtb5qjk4ln0BedUjccikqUEOzjO4qKL6X4HRD8M8cAffCGGWlxNEpQEgHkMHW8
iLXM/PEp10HKeEbEp9CyRh0UfH0uhLryvFMe10QFfVpOZdcudYPhjcR1tOtEKiGoE+UylYzst/0U
PKWG23m32Y4UXUYNbJ6WM0GTGF6MvbaHTAiafBUuboidenvW0MRDFNhG5FNG4ZyyUbR/q1cw1nY4
WCaTWbMb3+uSrZG58+IJDhObhG8tKsq+BLaZ3Y1KVFlxpSZqT15Zl2yJB8OAGsBQkf7sXiGhMKJH
OVexMQ8/8JTvzIjywRSqXBIe9Ffj6T0SJ2LP5aLTMQV8NVhk6mzKW5kB1UjOGCEx+AXrrpMJXj4Y
MYyayaqG1ZRzDgNVn9gBNIv+hhh0y/B+ncVXeFNc2v0qG5mVGQmBezBnYd9kk5P7fFrokmmaTTBu
yuOiAgJwSfZNao8er+DjOm+t/1+pxm8ZeKX+BtxkvEXweziV4MGi3XeY4X7PoSUUk2ujfB9jiGaf
OnCCWQ9n4qceS9T1CxfjjohrEMtF+RksQNDC2wqvrD40QCySo1AQfBzquP2gJmN16frUrKyZfmU+
hivHC/OYY8D+FCNvznIDUSt4jBtfWycv/G7g+8webTZdfrd6UZ9rC/LF3pcjg7of8jCH2PI0jXjT
AfyyoKmrbT5g1sb5gEPfKtRnRjyS4Eufbpg+9/DEMdk4EQ4yZBVpYTurjZHx49QqJF85r2fNeWjA
j30VShLrBIuWR9rpQrUiSUAIZyD3Sl1WB/ltSk8nAC6Za/dHJcGR4fPb2BX54+wTBddPtYO7kzZo
USb0wZ+G/KEe6L89fu3656ko8J9FYPp4lFNAMBsa1/ex5EEnHJeDIAYDdXaYjnDP4r67Weo85R3b
gzy9AJuU0yeOjXHMzgT9f0v6dSB6a6hN5rQ3Y74s548ARJh1lbnFI8SXoBdz119ZTUxl6m9HKVZO
Lrox9mAaCi8Fne6djTElhUA8vRoM5oVRqmEHfLIiPwn2ebV9nLMRja5f9gyOXU/QIolXZQa1p4wX
iXvVhmXSIsHp2VhHX7+VIGr5PewAcBXpEoyV6mW6aIls4A6CvJHs2ULGmCQwglACM6mVh0CkrTh8
VB+b1wnrWfIEE8KnajcenY4Q6NRqrebFFUZaK23xkobnRLz/NGdXdGjkV3/CLijGm9rD7L7Gtl6I
JcoOy7iLFskIullvrdV7pUB+zdO+aA+VvEAwIid+Pho/32F5x6A6FyTo+3cdxsr+SwpPXkXv2MCH
BWAtThE9UD3F5gJJ7AWpVP7Y9u9sJPnPxVIg123vixrgLwxm9+Uu3GmoLhjYInlhjkQ8iEtvN/zf
wn2xVx0o3HZsfnr7bm6I/hDJOd9/aJtDyuFWUftxlYYE8l7SKlB3V7FLvElpvBoEh8AnWHph7Sgd
jmoJP5JI9RozkPLFEZ9QGnw87yUBbRzrCiHNA1Enkol1B5m99icrtZNtf84nLLQNWyLP9moc9a6u
ux1UBt2aNzmgnH7yyYBlOnOUrW/T2G5NVHiUnCADpIuWPYqL/C8CEpn+nvk4PzTmT3ZvNbojQej4
VxDAOzF3h9Jy/OJA+/7U2VsE++ameGTFQvK1/7oJozgAqnv7ICNZgJKb6AugDv+xBbCsDJwC8Ujg
hxDyCeZ6RJGc4HWmdX+pZFz7ePlzg8kYkOXjqdX8MaN2pRJXk6kmP3dhX6Ei2lEPexAa8YdRtYuf
/9bqn1Ns0Z+Xbn5Ll8eMn2IYLHIL660lBDu0dMOuP+pIk9PGu8dsNQPq0rtpZ5YvL9VSGW6zVfba
t/XYT311RIODBuVLLCgylO8WVp8LIpgb23Zrbl+HeVRvWD87cNFF3OfM+Cy9Bzv8rruBub2/wgyE
iNlk1CehGml2qHrtTFs9utbTsiguxpk8+gVuKW5jdQXJ3vB+l/Uw9msrkxsFoyN9lDhh2R26UP2A
5bD1qSaXRKCHbxLGKdUFJCuwtQBZOMXhZwKvt4z0HyatR/rDID6VXdrAwFPlkCRLjx254PPNBzy6
kGyY0KJTVotwSzeSWoqjTSbfdyUbP+l1F2SVDCeJeA7H1zos6zfGXZYvQj4y2IeXIQFl0aaNZk2v
ZnYlT8+LzokkT6CVkaCqMY+0rfgB5PWpHKUBQs0RSjrqPnA4jPdY4OZmGqD8wrrVTBAoKlGaNZbp
ojDLL4fj/2hsH314JPItYI1q9kRp+Ram8GXPoe9MLU5NxDWbSmgIs4MsTRmljXm45meH5ZAePTy6
I5wImt3O84ooGeUmb4HeTEiLhfltH/0CFpom8QHk4FJ21msGWaLT5NRuqY/wR8FQr9bfZCCqeut8
aL6um2tXsnyKSuA7jq420V+tXncoTXz+ACYNGngdUp4cbFB2fwxpYFyGO3H6/QLx3Psr1IAMgdDE
4cx23GxDBs1sXV4tiFuh3NQWfRv+1cyTEaPSNWELrOn7KuAedWlj/oSMtE5lMja37F3miGRHdrps
gOQz49IPqivSQGgJ4XwYVd0ibU6aB4u4MdbkUrjE3zt29hKKddwL/SMOCmy2xHOOSkqmPIZJLPRu
QuwlZY5bhKFPuCn7oT4zoB5A23GTvE4Wc+sdHZnCz2Y1c3q6b7jYW353Yeiz+gXKOtN5g8jM2SlE
l6hWm9vYzeKPhrc2TODVGEG/ndRy8TTizl2eqyrNM6c8gMn/r3Fmh236kdnX1m5vux8/UV26iZYg
BEIs82FFIYkIrNVsnjSacLECV8pKLMZZ8+JctsZ9pYlrq2pgZLD6oYmcKP287HZdT/6oo+uo7qLm
3MEN3HhrwjQu2qR0MdijVDOU2zFwSY0C1/S/9mdTmxP/MOtY4dMziL/jOYMLjZBCQTh2QlrpM0EH
Zb23UlbLA7v/xdi6TgdsEl70K1qdZQv0NYwE5rbbLT84QGR4seveiJW9/9B4Y3LGHExBu6K3AYWW
CfCAOD+2RfHbeYf71YwHvKBLWhDhN5vg7XfoIv9fmWDwglglt7Oq5K8bchqLtgerlQYkUfYZpjRg
KV/SB+v04F/Y30fL3kKrYUL290mx7tG8LueTAmF7F1hiLCoEIbPzaRoMj9i66nnz3/RLqWIgfenc
8+LVXda6aQ5Cz7kcp1js4qSw2JHgB3uddSST9sph3LU3EnvXo7xcOrsHgfRAnJBNcb7ogBpbbA/8
wwxM7BuieP9YuSLpErzQ94v14yNQMETdIWkUQ9r7DeZSYVOYVztg/di1SEmAN1YVZ7srfEGOC1Tn
tZ1gDH9+M5dd5CmbdSQgiPc6L85G3BR9jV8B715X3NDXlv2+GxmKVgnO8jQvD/Q/j3j0ypSk4y1M
dueoTbncufDgl9hkxXw19CwVQ6LR0LTcvYNfiTBNELLdKy6ZBYQ0DjN298lkpxhOQL77Lsm3wVsX
37MHTplqsWuuRbHvRGddOHOHMVw8uzmD2pWX1mk/egUhqEP5/llqQRMfTfEPTzhklZ+M57mduoEs
+nfV64aatUkogb2d9B97o4B/rxpQkLthbIghfupzqjAFkS8glOwHdfLDwa8j1SjeW19vzm7ikmNP
N+504p/fsbYAUvFFJsKj2oQhfoI5BbPPnuY0DI2gr8z33A630Weklqq9UlgQMDk0A8E8EhbD6AzT
+3Lypb265p1VdU+UGAsaqgexFEShPGLbYq43W+nKlR/udDKjkafnGitlViWkQWcheMmYd3cz4xJG
ZctZZnOR3r3p5UxuEIchySdzZqdn9iGXztUKM+VJDceNU2+9Z7gU2ujuoBOUcLxADItFf7PzYQWg
M/85+FT2VLQpe25jSQoVetdCG9+8nvcOTF6w6oVp3ubkTn8YHtIJGnM07Al2Mxk6qvPAnnSgA4uQ
+m8m9o5YcOsOq7pNz9tsHlboVfhvhYBSeNO62aGwUljc5AC5N+qrR1vSa81Wh8mRyLUJw8JCjZSb
RH3e0uMG/teAThGNqCLBP3Zg5u9PFLXONWVHD7aaQxY3cKO+6LNt6Ek59k8pAGkaU95x9dzyG2D7
RPD+KdvmU7DnF1pZ8B3K59l3zJFOHy916rGEPKPRjGygjQhC+zVEoNNstcmwN6ualQeGlIIGAdEG
wqpnMIq6x8ItovVhML3SflDIlXZNIZ1dbusUogjN3F8ziR3K5bAuewgQCGTV/QrvQUedJlUBnU5M
vnQQZ9MSg9onpsd7rNX2AdqHawEv4TtSiM1Kj+RPQFdXQ9HBaa/W7zpAUd5Y1++CxT8Z5Lbjjhjp
/WpQ/8Ee5F3AwIGrGo6oVBGl2LZr2Uete9rg+oF+G8WPIStZiA7qd9UAYdaJkiDU+0Z3go3Wcmw2
UcypbrVH7OugT5aZ+hyI6xUJ6QXne9C7Ap5whER1tY1IFLsiH2hmff7I7NgJD0GHUh6ZodnHVsgH
Bu/snl04SUG883tApS+3LikyyMeDOwNy3b/8/1D30b3Tlww8sE6ya0WIoSNbb2gb9JMiyENlyLRN
t33TLF20wYGgKg461ZvPIQHSslsjXSSXuOP9aIXcZ5WCYvBmwLcbca3cwGb+ancdeeYDvUbbBIiJ
E5wKMj29BdXlFCc7djsoSkhYfTIKeI65pO8as8F3VGoM2Qbu5bDkKL35x254k8Gq69L/r8x3nbJc
c+siPdZGNO4Ac8qKdm+gAf6u+hicYvAqjwstcEeLbUXEom7mH2iCA+Y8rUelk7MCqIj2nZSTjduc
uhPF2Llyt4JFAZvnz8+rYHG9No9Bd6nKuQoX87wEjzhENvgEGBEsLpQFGgCWxqsVZqW+8fly38tZ
wMDcPLjus011lsBeO702iweOgOr0Wh87Zs+IGUoE8Po2CDeVbTHqt02ZPQBkF+rycTeOYU0Xv6Qu
SNMvOFyMwhCh3wJgNmyo7QHLS3krWNFNYMs3BQMcw1cw6JGGDiNREuWo0si2MCsw5LOilUELamhX
9fUvR1LZis37WbGCrTVMfo9Kq+856vTU9U/Rcgwa3/fGNs/wAZBAN3rHOcEwlMGuK/TSqtU/PP/R
GMWxIYVVcr5NAqCB8xrGvFaINu+m2juRd6NFELEzdv9eBviqQ2yOl/Z+J7rCxXHLboy26gZByvN1
aRqtKS0yyvJBbbe+LXrDaRylWm3vvHJaVsAtQ3R+Qre5u2HXqxAXEdM491AD7/Hpx4+70uoKx7fa
Td7yvxjHyiSOQwkUZqECUo+s7cOrukGmBi5bu3sgXSWZxnlM/xzi83igazKvMFIRdQESrDNfPGVp
J0wZS2ZUMUEu84q7G/12fbq2mdUWALlE+h7N0uW8iG81ckl81fhXwIaXei1GhlnTmzAHsf+z2hG4
q79ogSzLVpT6M0o+eXOe2la65mQ17EAhw6ZhO1nb9vCJ+AowQa4EVUvLgs6eVmyudb677N15IKWS
xDsR3kpH8vhCw8qxpZyDL7KNu5ida8yR8rllUsOyCdyjOPu2igsTbDg9OWp/QRDZWSc0Hl9gfLCL
NkdW0WomUft5krRoLw0xeoAj5qGcaZ4eACgs+KIOLCErQ7J846Px5flV6mm0RJXldGhz+4YF1r4y
/hmzafUWOC4jn4ozy2uhWXJ44ZsMhSMQaKJBOVf6uCIyx551SBh8I0PvESyr4jonN0l/YFR+Wmc2
UbM5Ye5Gkh/pOKTTB8iNBTiGno1JTaJC5gpOgvBZb0Mlp2N7GC/Cd9yQFKWRRIjJkJdNJe581wTt
0Cgc2iO9co9HePzsgWA1MboNcGD7bBgK0hszqncc3OESTS84GIeXaJytHjFaddGvk01a/N71BRkb
0hoV4d4Lz/aMlszLXpQWj4kyDBrrWd4GQYUQ7GlpP7VCSqz2ZeGM+mkJJ0D5X+rUntW6kooR+tMm
WLzL5XMIGBQSrXStWhVwHvk0ks8xzGTqYR7s63NDz+h/8H5Wegmm65wCTO4eeWcBM1apwatZNlyB
5M6oN/gWKL9hgk5FMKP30KtlxXtniuFqIUz/7Lqr8hvSz8lqW7YD1nQDCpAvuxd5pEXrgUFCMiIy
hgbYbUW+M4M0LHMJFr++1B+YISdgjosv7wyV8cGTVKY5sJOQKRHbc6TSUwmckhmk7NAfrsgFfS77
gb1+V/DB8L8J4x3pHPqdHV5M+iCTDYW5KA77V/jnwapiN3ozYzT27hhqUuwhi3RcN2pQZcaO4NLs
mf1C8z6xgs7N0v8lEpfniQ6Lm97rnMemcT3WeEBJxhuY+lk336bO9lod0Jzq3c5XW7aGYBktUYVJ
Vm9YRp1PqqsEnz/EoG2ZCeNjoWo86Kb0YnLPVI2QyUdoa1ixjDynihXHRP1zBGgTrJiZ4m56vqqs
BHKdxTLFqlUeVs3tjQbTpHY5ZCXe6bGDCKaxaXMYx29Ej/j9HEr75pD9pkgmUfBdEOsOy0Y4CFx4
DoRZ5VsSWushpE38OVfUDu2qnOniFG+KsmGhUYpa+ZL5P0NpgI7oZcD5NgOgLWEb4jPDiEvcZxts
xaL47OYBo+d/o5zLS92MGrAJo0RCLBDIqppzG3F9wmHQHkAQpshPzJEL6JLmuAPOGdU1uJXWHRn4
04AOYqQ2XY85e/E18YtAfDL8Olx+sJPEPOaL91XWtUyQhG+6e7XWzToYtdqUYBbqi0Vbi1yBc7KO
ztLqp2lxYPZRfmJeiF0Lwn6WWGyUxlM+aDph88lxocQk0soFStuhnnz/23kaCWhgsN1CwlY+o9Um
ddCsmaEuLC4dwf8zJJu5ZWOmDiSP4vvZWhDg/DmsICj0NAE2XNkanmmkUAmuUz8V3CQVpdlkIkSB
E4kUM9tNiOYW7e6pyuiRYoH9vC+sMx+03yujs3j4opK/nlWVujkjbXYTuIoacCm1RACQqsfRTBX9
cn47dYmN7CaJ7zfkciaMHXOWEMMHuzYoz6/MKXsMC12TLzcEKHP15rE4MSNeulAOnI52i6TnG3g1
rnOo9ooS/tNgZq8LQjSLCFLC6ay3Dcz3PSMs39x3UBcHZznE2vRw6kO3JLc11UEdOIBqykXlenYF
k3l4QV9ZZPXPbG/BpDeLDE3YxrNFMvIvcKjO/M04gZ0lKt2d4wq/HPnnkQv3aSPmNOUDCZI8X4IL
xSNp6fGQFrFrsbZeY84zD2CSCOI0kU1navkXwZq100gImSSfH8HEKzY2+/1tHi4oVjrIK27Xgej1
fod2J/eSWEaiDmKpfYEnaNxVVQ8fh8M96d1JHDxYcBo8+kB1SiWp1Tpw45rfhBWncgqIjPYaKfoQ
eg4Tnv/K9BO+TO4ndhs1wI9ma43+CvuhUWBz089vbSoo7N3kWP+b2er9ptY6/erhUahgEqQuQ6Vn
28/r1KlNk4WPnoay7ZTZjEmMXJWT7L0xhM2M6IiRgW+LUGufXx7DkbE9e3astK8yaGteI3/yAEv1
JY9aqJp2DVRMnvMKHtVzOCkNP933sjCfE5fNlQ0sYR6AFPTyltEHaMh3iMJ+UirG4X0TOF/gTgn3
nv0WFcSvnXufPn4TnlS4MOem2kGH9IntZUNHCUldccUr4jnnCjBQVZD+DEAAedxCosqNpdmqCTNa
g9APIAvPYUInFNXY67zVkspq9PhOBiJ0kmTYnkNu0/cpcDU5e4aIpB2om5uQvrjNpzKK5/wk03mp
oBY89TiHrdxB6sr2qx9U9Z8Ecl5qjlFZn3MQLAVJYwh6utwcz0uhByCjqwdYGYI0FUlnAJ+kOmk/
NQfHI0vkoe7BrAOpbZEu+jfNrirLW27zhnOJ369xspVYiK2g209EP2En7UDTY7/+OF7fIVjjx89s
74VPZwu8PKBAiR62acakZnQu65RJaYyqfsrMgB/eYKv0qoP8QglYFM6lrKDr+EJb6Dta/oihArpK
SjXGWmhUrBh7sOPMoelgh6rGtpVf5zhqe+GQWMNdyjnsky9VpUZu0NrIKM8y5f1jZ8JYd2BqWuUR
4npCISnPdvU3YMVPfMoCPMb8J7il6d0dq6GO3pep4tlGGds0JA46P7h8FgPhe6B+LGvwTG+K74qZ
sOVEsSKAW5hm5BpZAvxGsb358U+E7UU0NUoKbPdTjyaphGhndb+7v848NLYMy/alrXQlx4INTI7x
TJJT++23+6iGuApBp8HLV8kP5J/F6GFGOtLcPKnIxbphhZyEOQ40ExIPAAM3wGw3uZL0J1kd34AZ
cc3Si5IlHXDG5fqxT4F3qJLyeUQmb1yROyEJ56AMj59d4Lj+keMIf1kOMnYAIU+oRtpa0efbLxhN
kh3fWJulkUBZ9wjPueDocRJR2Kho0MdDBWXXXTpIIgi85X1wYL97S4u8GHOp4qJUWlab+nB3Cqoo
8r9vyyw3TzdPIytDK40SIAR49eUyRMoeh1OSZtm44uCXdKhSuHLDvnw+3lQmy9L4mdkx8RFETJGe
VJVpbW4zWV1HOZN4dYPGm4YqZv1eyDaXnf1HfKWQUl6yBRjcB1ZA1cJyHc11np86qjRrEeWQAdHi
SxNkAyCV5OSzRZGxvp0lDPPpEBm4aQxalM1yXNHLqGEG8aSeBl3AGytPVwKyedGc6r4i79rI67rF
HgafaXj02vP2VdzP+5s0p8NqeV1AvkxgIkbdVoqmzvlc2wx4hisL+IJOiMPwljgJMQnUUdNKIV1r
lRErXGv9jxN0OyFKiLiRB3iIDNckIw8CXA5WIQSLf+cHMQBbQk0AwFLwrb0SX4L5vwhcm9Z6SgFY
/YDC+vWUcW1nkIHzUx+70sf4LpLxquoF9IKI9AUI2B3WqbhZwMCsHzOgHKKhgMdbQ7paZh+NYoND
uJdicSNXInjYbPLoUt+uST09w/itz/JlCCh9lNPy0lFmNiUw/NdnoTxPAfPnDS+Ne/SDdyzziiXY
ZLnfZDyogPPJ+RTKFHfQBQKUG6RpXYSUVQd7O6ff3Biu+7zWOX85UdOI/1MexBculGfkgULLPuSB
tFzZu5yy1E5a84DJO2bp5oYxZAg8iHlTm9GAOnUHrGGTMZvfx8qwo6SgvvtkSWif7EV36mY3aQWJ
fP/m5FJ7djD3k/db/YU/ISP0lLUuU5NcPN56bbCgk6Y5jVKzI+1KS21yAGpA11PUJ0ldRnBef+9s
lwdWJtTK3FAH9r5o9J0FUB2VJh0kXxBKShrU0IfmqZD/hbohOZd8rDCmT7e4iyil9zpx7d6Rzmaq
+CQVB3xTicmV+BJmXDlQSklQ9u5DajNZvWRjnJ8XCi3Sxnkl8YPfr70Z4DccF1igLFVT/XF6m8yl
mW92XAaVduDL+cXVm0nXojTEKKuWmmZlgH57H1sjhhv5is1+Y2giHsbUrQbQrj3PlraT5Z4WM65z
+T8lkpzi6vgtXmyGB/BXaAn0Aob7Ll75cdmhI/v2x6CPt1g8W0ATOuJKEfa130Y5isa1GZaVCo6A
PeiCEeda+49OpQYYQ2e/GOVG9ZaLxRNL6L2ElloXcRqfPQkcM0gfUpYyBQ3ODCI+Jfp74/74sM63
FrxV2sYKNFjKJ0/XahFW3Ctd2p8C9WBRsF+wVHpBUb+XdYqXlCBY8mpV5rpOHOyFRSHtvWzCbewB
tyUMPCRqfK2z/niYT69lWm7e5Hp5xRchma7Xu2aS5WZISZb5c/44Yn4vOSXqTGtBHdKpAXojXOoW
PjK1cWObSS1R2jutaYLnrF4F15/EWBX/y8ME5yo65nZGG+jzDCD6znJntU45BXn3e2+hBtBPwABd
dl5r1YrXiY0GuKz4r7//zWdZAY+AFY7poYjJx6CsyRvj02r8DS3en6iCVz/YfevYGKwkhqzUEvB/
58no8um7XQdEFf5BpOSWM5cFmxtDW0i5ZTOeNIyDe1/5ulLak17xCHuBTM/k6VrSYK7mt+J+o0JE
3MG85mdc64sdjN8geQEMN7NfrWK7PaF/cbUgZrqWYVEIXR75buiz7ISrAUrYLlU4dS25l+BoOf9Q
qsZyWDSlUoQp7HrMo4XNGEDOuhJgvNZstwZLR7FXJSXtSowXTlXMwDJZUEz1JRDoG8RpFjRYfsAF
V+tRGbHQy4L4gIEa2tGRU0SNZNPsY06Tvyj87ijQLMucini9W+1BdQFHvboJN/d8yTxQR+h2ehlu
WGZuMNiar0sFUoDiqqlN4xBAWg6TqVEDcDHt5nJCtLXWIDS8ppep8L0/N37uNRhxvTpUucYwqmF8
LkUBgOJgva2cxVBYOeK3t7QMG4xRliyPTPe1/sAjDiDgmRRiUpqK45fOO6fLUd7mWtm1SkfDfy7D
r5lGabdaQ53715efRgb8ALcVZ/O+2vyTC1OEI+JsbF8wXkpHq7hHqI/yWRgpztqVK1nnJsKFZALK
o5H6MtGEaOwkhzYrEfvnspF7zlGtPY4ABxp5G5YjPI5m3bS+4/+YnJihgIQkOFvLPxlJL7c4Wzmy
2VaY2nOFMH1rjaOEZf4Nf/TNlxAnLBCxvEYdIFgo+/bFn3u5pr5MGhSbft2Dfo+eONlaQGWS6Wtj
fj4wxejggYoIOFRTLmlJcnLSuot41HmEX18cxhZPuXC9YojAEFiEphis/TC7VFgVBiBFFHBp4SZj
37lSMcs3eXOzYk3xSXqeiAF4zBd60Q5+e7zdlPlack/MkvPUCBVi/GBD/YRw5BoTLoweG87+W4Gh
hmd/AnglsZ7DdkwftFof7XnZxFxfVdh8xqpjTBYjK5URWXxuGpXHJK6xjlQqIK554Fr54jCf3S9D
AYVXqRCRN0Os9BtTXh4+rgcEm5SUDLccbW6qVj4rN8vCoBMcXqqU0gMwx9IFiF1ZcAJWdzKPjmJd
FNpH88lbLlFG6RjKVHbQRaUQKbuHRT6K1d2p8mGHLKo3HiOoCqLqKjt0j9D7cAAFoKJvJSaXJXdt
Zra/bAikDuFUV731ubY4WCaxIrYcWjUgNsxnz2o9cld5pRJYyXGm5Uj5c6oQfcbTO5/ZL6bns6w6
biahMGiFBG6wsFXjKPquICgYf04BwI24frU3dkFKSxmgvLjt/N8gQs0hc+9eAM0D0goWsakUGL08
6u30VmpVVGpdZmsSf4xMdZBEsINfCRYeu38JzqnN/wqhQ/sP1+ptVZzpOGjoJNGgAhDdEn9JDjbM
lXRgIQsD+xnCByGnow+rkVLulXBE2OydyTHFmuSoeQaMDJSAy6tAUSuCpcU7RWot0f68WzY3BWHE
kA7J5GLn5Gcw3RtbwZOWv00u8FtvVhVc/RPv9roONwgRcuWyQqZl3kuRQH8gFSg3wBrbB3NIrI/N
XFCB45krq7jWoJj++aeagFdvK/oQFqrgyPAhAxvpGGzVU0u/AV5DZIQtUt8R6guQBFquxnEp8p1w
+kc9pASya7FT+1tkLvdtlfNzxi5YKIzhFjcp+5FD/UlA9Q0j1sVPfdOsyz5VMWNrDP+eL56H6Zki
n+LRoW9BLxJanCwRdr9ljrckPYhq3DrlrldeWm2NgiEQ9gIhSr3lt9Dvro9qRk2DSLiy+peM4iRB
hwdx0vd4kEPndCQ/pvxOVt0VDiw9a51d0V6LI8cBS3elp8AUkTJRrr1rEiD7OlqMzoGq9MQsn5fP
bBvnB9TteNHa14l7Mhg5/Py2rbaV8fO8D/8GwmPckxEmoYfzRdUdYv5IUcby18k4SU31fBi8zD89
VGZ+YNslTgi9n5X0r51z5gUA68okNpJ5d+KsBfI6tz4ORIYFh1Ot9mD5r6IQqkw4s8TbczaucB0V
ag9HEHWPy5VuIed5hX0V4IgSy4RSp/WLlf82EaFWJKPUP9Fncw26YJ0cPz2BrugyJYxRAbCMHmg8
PYv4z9dvoqxDDcha8V78lulz+Q8cFeO2BMPoM49042KShTNWLNbhvy5nWJl5RGXaha9gWSa+Y4G5
Zt108txmShZgfvgQSTNAUqEqL0aIA60o6P6TvYZVhDHIknzsrzeuEDHmwKgeRpgSZHbR5bkAwni1
BBI69bee5UefadlCPMCpxn5+S7s7K14jvvRsvmmcCc2UcCvb+mjRqKUN9BvISidpD/N8anshmQxE
VruhJXwgeNWtKT0GdzUmVArtRYbPTHEeLkzMu4V7PKC6TChb6cmm2JxH5U4T0p2ycT+i5F3svy/6
o08aWbqmTRSuWa8EqxPjeX9O1qeBVTFu0zZIA1NOSNHwtgFJHtkefQfOaet02oLEas2mRO62vDMe
LtNnJ8lSHjm9kx6Ax92Fbghz2XbP3tonb8Cpn9UrgLZrLN/s6G59AYQB0hIf5uerDYVpizNLLFrz
zzCopZgUej95wj9GtoiN+ZTsOL78AAm62r+mlXyeDmAuFMp0A5zKWxzuxtF3ODvvkDhlyGbuNvmK
RXnqa1pGtrZxBGXKBvtN6iF+SOJY6+reUEf1Xz0JD5GxM2qAiPe4S89PgRAwVDS8YrEag37hbEl0
1P0ke7tAO2bqxuBAOnTJ955IQD9M82tIreP5TCFZ/GA/kGbjweR7LBo5aivKdonqFqFX+cZUSWUS
+Xlgl4yrvFGPq40/HiqAU581f90RJLOju4Aj7+hcKMQVZ6aGPDt0M8Itgiqxy0WSUKph0LOIsoXd
Q9XskVE5zw9FcbrUqFbDPDnCa3VsoWPIkDaXcicYQgm8XRGgzr56cFncB587NEF9tMGqtyoXOke6
v/u2ZteR57sZUD8iOiTM/Jne+Gk2tRNOQHqK6THnDdH7OnvuOq6C+06rFK/upEYXGI+4jsml9BMH
aUCR9drEqNPx0GjkG0F9EksCnilIR6B3WQ4lDqjMhTAwzTCaN5ERL/1TN4BJ1/cN5e2jNXyr0KSU
LL+nGs3Dm5EHJZk+i52CkXMMBtm34Yc/8rrmIoh4XcWEoMTmAKyrnKttuqn7zkWjGFD48hHNw/u5
UsXINPzp9RS0YmCU5Ki6FGpa9AZEGGvKHMCsWVZ70pfLHeT2uUSm6kOhOoypzCLkeBBMuz5cHGef
qC+gTCyifKlWQUaJrgLxqJhcyJG02goet+Z+F5COz61oSFmYcynU48h9pReyupdWRl1afgKDDokX
LikA0p41lFOOTDyqh2mZ7WOs/I3NAl5kKnf6alHLNyRhMESU7UqgVLemcbxRBEb0cxxFyfdKs2fV
kmQ2OFbguvqOm/XBh8VKoUt9a9syjYkN6PsFw5JXYo4sOs+0RbKugbld6tpeVthz5TyhPLp4/ZSv
uFImt4ExS6dRrwjq4gFauPzSc7cblemVIKJlFBLVBxsY+vMNZN9uya3+MZh59ufPJj1PU8eQfnNL
9Rrpnrsm+zkVy4/YBIQAOhvVPg6qItsCoq2C+jr22kV4fy2SFAQqJGkh6PzEcQ5keKZTdVS9lVXf
J5pxj4I9BESXv3MmK92XUwTwxRULKJer/ehkLPd2h8JtFvrl+u5BiU0KUSFU56R8DF+pF/bGF2ot
/UYAgg62GVdcGDwreO0O9KB42QceWftVX5r/DoO/MkOZBBjyOL7iqaLdiYgKFBOdoWYJN7UNExbf
86VrAoTy6HqHSQeJsFfuX233ZLd6n70FsUxXZBfBMkVPhpCjBFWBo9UmYKAWKWt74daG35O1cSIr
39lCRlOCkw9tQ0YievMyZoQjY0ynt3gj3WlpcNYnt8SGPmd+Q3gxGWqwFi3YC09TOOyl5vPHTm2J
purgBdnS4AB+0kj3dbkR+L+hF6N7o6tzQFwhJnQ96eCM2D3RTG9n5J1P6LVxl9EmYASw3pjmevAt
jeSecaHcoaSMYYv01HOkHJs4gkWceyuV0WilT6cjI6uKdv17DEuuSkgD3gr8tdLPpUdkLzufYsgh
+Xr/QHCMcHbkL0g9zjLy1DFmL3ixAasoTAlbL+ls2co2HnqG6TcrxZKOjjvxK8yW+S3wAcZ9NyW9
nV8yACIww/LVK5WIl51N+Y9RFW0Pm7HHBqR7CF904YtC8ETY71lDA184LjY2ypI9ERZELZkT339C
HuxM6BKkNxiePrpjj6Yt/P2gRIbIXWaFRttwpaZ+rgR3AgSAKYbi6p+UKIST3gChk/cDzDYn8qmK
qf+V8U8xBwgJJ0DMuEK+LFunj70TV/C1OpgGxFI4vF+nBUCYb1KtquXtOqIi5LZgqB9JAtbdeIlI
zzDOTGCjYvAQNtTNYJ4J+4mf490LmkQfHmWnGYpqXIOltFnd032ogckg5Mn6pC3th+qczImCktGj
kBKcuH4waohRKRyA3lE8CdTPO8AbhzqWH12KE2WS6LR2M60h69UA57YL63A/ui1xh8c2Hm0KDH4A
jIxDzPh/DaRytA/BD0I8/HQjnHT/pqAuTqy7LNjqfValvqYneJnq0z3rGlyPmMX/I9QlH+Wz4WYb
C9qOaj9lCDM4kmRWw8Wf/GQ0rfMPl/LQXrNYuZJu6p5cJWf6g5kNvw+NZg5zp2R0f9Mg2jzrOWa5
fykKUXzui5F08fhtkRswXdyudMDDunXH0KHKZVZY2hBaF9elBCakBwnhjDHRCzkZdnTn4KhivQGp
TiqCxCXb99GDEVDfO0PreygRASIOMdqtYDaPPDlCGkCorSh3CV2LsMm4DJl275JlY4fBbV72y7SV
/WnOBhh8gaFXc5iwuFUbJHnizAP8BQruF0RWrKsYg/5dzMflDzJQ4L3f1l6dNzcsjTM245ZwKS5Y
xoYGDDNtJvJFW4vbirN8DU5dKmSaEV02fvIFczZXq3UfK42CXwvoxCE4N4oJvzWwmHdNgfaAQaRo
+VnsU61YBcrKX9Et8HQFADdXzLzgqTo5+ZlbsnSq1cg3KWmNRiycWyOfIkqH0PbkyLrWIlW+Xn+H
z8ttPcEDqWOyI5w+fQBCkk060cE0e5veocr/peoKSZyw6RAug+HjlAvJUZ1KJnikSG3CJSHNJzxY
0XDkGhgOvQnEdco2O3xrArJeLXWATWXj5J26gm2m3/MQcw5xBBfTtl21Rbmp7RmQOht4jCL7mFZp
mNpsYwgVUk1w+4kY6zSj1vHi9mpBRQ8wzITHiE1P4vg/YJOZkRJF7a1kPv/8CJcWSrnP4IbaVwJl
Y6pbJ0Z5BHpVUmfyLyywalyaxkWLOQXauwVUPPcxkwiohRJA/Fk46mg6qBfqeG9fv2UtJGip2Ywr
vhhSKECDkI9iYzY64ExI0hCjpjrNjiq3KcNN9uxh3jcRREJqOgk5PLREysG++3yBy59SrGwyXY+f
2eKEDmMQPKieXWrBCENZirCIYJJ6sfwAwEOGbuaXDtSecHuTsFIjEDTTv7sko3brwN1X0nrpffTI
OSaDTCKXSFv3UAKx84MZMyU1KJTcj00kP43810VuvJBL0M7Ya4zhS9UUp3UgIGpQmAymfRXVeQ7r
OS0BnfirZ+SDa5hmE+uieTVY4y9kPqsc8Zc5rcR5D47pozTuPSdSqG2DMwojExLqhBxkhlDIYMJ9
KYfLFatNNG9w0byQnm91DW2zJVm89/qBUfGQE+6tl39vdaLo1XLDFP57/WCaHxEB9CK+Wkdrx8io
vAKR358kRKvcICLcW5axHljRjZ7bsVCEk8xlE7AJNFtEhjCrz3PXoLXfcUdOE71ZV9YGexBEApXr
wVv6pjKhdyMfDVaVQ44I7yYsvKdq3GbbIhA8no6xCHwJRy4bnc/O8+AjdY9jl6xO6dkf7LsI2vjC
RMHHhGN+ArDUMJ4weZrhREKp5PhwEdPKN2SwjEdmXezgnM6PF5KxpylKonGcL+nhsiZPwcg8Djf5
YTbKXiGxMPLlF9QOme38HPV6kbGfhZNwkD5Re8kqjXOpWmSt1BMN8c+kA+LIRIBwFF2zoOTXQ3Y0
OjBKtE2+62BW+AUjHt908JbndQAgZRktgbjwfJDEOdM7xAltoXnCbDKgepy77Vd95pQOEWWkavgt
CRDXNt1Kp1jdprtFLHMavBPC1TuE9l7vYhFfUK+rgM92vGY+BYHgWYw4WIkAduSDj180nBaw1Ei4
9BQID8VC/1xiIe4OQXVBblY+/ZVitA4ogSuB2JuPJL0c0Rnb8ZQvYYkfkoXwysGiT0TrpnzC04Pg
cEVu30xrGA+HjPdm6DA47hE+6HLEc2sdp0cmnBOM97vJZgZkCJrVWtiHO4CSI6NGbiOQCjHyjF0d
T0r7cLGnkfkqAXfaVKt6J4/PEnLWcuqFSGXU9UfO+ppso6iu4v4AiFswj8YuMW/aLTd2h1rAZeV/
3G0fxN8yRik64OOnaXTRYhlF7A6ieobGleMDJgDzRCxZeTlFTi7R7t+RX3I5xcUoAuUHoH2F8Yvg
bSs9aoGCcc/bFXyp4q8eK5o4gKXiaTt9uNvpzScb9r60P+9hhgPcgFEs/FGS3PZFGIK2IuI1lJHH
yRajR2HgZg4S9C8BeL5W8LuAadwSGNHoD6ia+8NSjwwQpK1RLZwrd4M/eEZIn/ur5wQOzBEeS+82
C4cGIuL2vdFnYsRUsnuI64Mw+6vwdCk1PAv+Z/4MbVxSUQiP0q5P6O7Q+NytKUmhrvgFHpe0NkyB
X5CQhu0w56oV3MC9hywPERXMlV5wMk7fVsXeMXlBpUH8QR350sjSCSj37i0LH1ea3W9FRgMJPsXH
bhqyOewzHNpAUD9kaY607fNK+eB3sN90Or0z0qcP7BAoH2eXY0e+o6babNNXcnKUA7oi0mVouIlo
xIWHom0KQieOB6PuxDJvgUK5N4aNgZTAan1D9/hFekkOMsVdnJLbd04ugCC8veRkzO0u5WDCgrNV
Iwfe/hCzYht1qVsKqGJ7B0BNODe/5E7aSR1KsbPmM98rD7Wj8MStpWc2OPVU0a6AE+4CV14T5SMg
5a2TxhCexoHA3gNQO1mVp6ZdonXlP1ZzVms4s2sJ8PU/6gfnOycpSqnCjp6QILwkpiU+J+S2DLBT
95IkBmG4P0FJZd4i/5ZXk3OE/nnY4Wk2CQAtb4vIHZkHnahJp/atn0xrXlt0deNVzwnGh2faHiDN
gGkF7836artAACmKbzegZytacwyuO9qfDfsCsjSEo9zT9RiWmdjqIR0+OMPLC8RBYN91qg8AdMMH
H+Zmsejs81QGSHkPCIAD7hOqhpGZ/lxTtLqEQKyviooagEZrZW2YbctuMDoOkwwZwzWUzZvKFOrI
gj0fNU+i+QqUjlc8/UnSBK8jx0HWVbZunPtzDqZ0fKZzoOsHTKE5VjGxIefzt49PtZUah0JpXhaV
hSj1AL2Tv3zuDyOtjyoPFH8GAWeQPHpbovL0cIqTRBF6RBsJauQGOS/v5yZ0SnEtYFf+IXsMBVYq
iSTE1zowP0eVYoqh4l07FWmZ3JYDL4Ek4877M/BullFj11OzTQE+0aGm7qUU2YdtAhjgJeTnswnK
cHlRF23U1w8CD+cOJjm4DQXX7T7jdXiBKZMxS89JLAmsPaYqJwN8O/U0dsF9/iPJXCRCdvXVS06U
OUi935D4Q22CILYGzBSu4NrjkFA2/Pn8VgpeKbRC6iygahCOWprT/NopWA5qDAyracSe+BaUOzmw
Jy5JL91tOtdNnldRm4n92pGVP13Stoh/fNs5PAWKgrFyMHYVKHFCaSmVfT///CC+HGdLoHhhijxz
9t9zP5Wf2ULBlEQSHoENgauBH9edQPgSC7n1yi7pMXSEl7xCvTVKSupob7c0wxa0hQfctgXQfKlb
j0s4xeKVKdne6T1kMrwFgIAGvZJnQreB7jHWnzAxuVgws459zn915XKui7nWjuiOXaoyz2zS4YGe
kALZUEq8tnG8rbU3mvRJxSv1wzL163qftw7nQfxICm6PVX+DlcUaSuf7MA19rMyGgl0BWIavQRfU
t1SFNaGYBabG2IlgdTPPd78WTSlUrRGtOpTNPAOl3CUh2v8MtYXIlRvmCcvYehewt0DWxo8xs3DK
bMV1gQ58unuEOCz0qCYIEkVw6aoV/wwU17r26gnvp02J0zeNW/zYI1nVgsEtYeVx5jTFkimSdoNA
YvhwEYAXpuO9ZzuRK4vcpDANlYbEeZhGVGdUE/ggYy+Q42B9nNv7zrpvJHQVpE76TQeMHlhkACtQ
DOb+sQqBTgPln0Xlxx9lAzztG+x3vd781ZSG7sJaW2mqMr9GHWskOt08C1jC7wfn/aXnRRAVgy7d
J2cPzoORKzue6TYNHf+yZ2TB9pBZ22FswcJYSsbg6PKfQrrhTfjKhsgrS9N+WHhxCKTQ09IUv7M4
T7TvnnvsXzCb/pLAilvs138N6MDR2rA72Rph58CNj+AuJi4h+HD+RRUMQV0JfmTQjhlrEAFIMiyy
n8fJnehxBF4+IVaV/oUcTd3YUj2QgC6rCxR9psAW718jpI4QGK0wQjaDhFPt2HjWQ+uooDGqjoRD
7mBC8Wj/h3DwNlAmg5Ap/W04B3h3JjrwaaHWDNGs9ZMcYWEANLg6Mk7j46xl6MJfSU214CT8UIFA
xBXhNHIADJnLc59lu9vgi9m6hKZN4zPL3Rdeznrl8mcc3+H9mbN8pzG6/RwA+boLp3RaXQ3IibSX
r+7iZfyNWZBinXZRgLXExiiLdVyj+FjCrkjTbCek5t7eFX04D+7IJBnaBObd9X1ikUGCI3nK+IKr
DWDODK4M1ylSp+JwLCriAXoqqIzu9n0Qkh9RdI9HmYTpVyU3iLOzkTJ+CIOgK1I6RX/XNoiow4RU
YPZllVZRdqOquiqto5tIAZ/krWEqoRTo+3IcXwcY2O+FDYVPWoeVNARuTaD3TcoAPvYFKnYV1yjS
X6mJzwWZoQ3uSJqkWk5TNS7ZZ/gFvcOpYXlQJI0h1UfvQwCi4+7Dhc15x9iFAIF5b/icwYdIbhKG
b+gDsvbegYXknaqLAsMrSLCHlfbt9JxVdsS9MtEn0ZRzdE2D124h/hH28eWUcGu8bqZ7zislr/Es
9yfnW7sTClE5hEMZAq0YaHLbF2WKwO3ZvrTlT5zGVRo20o9W3UeHGLAwSZF/osHhCfaMbveItBC2
4k8RLmwrPxVTu1D5+IVW5vYNCZRD1b7ZpJZ0ea4SJNttpDJ/8evfToJvFbJWEDFidN/btpUd5SDb
QmEfsNmBHqKn1ta/RIEpGsxhJ4e6Z/VqmSbPnJ7WaXVP9TunQsZxozOpdSdl1KfiFIPCwR0OWooc
XXJfKscNsfSNdqkLMexg8BltZEAj/MDBvn7zn7490rFR/6JZ37u3QxH8Cjug0r/7jqBmH2X7yESi
Zz9tKe1NSmjsmrymuCA7i5KQYZfj8fra4dxgRHtaIqR0UKEB/I80DY8dlBm5KKq+egpwyXdEkuDH
p4LAMcW854yN0h5cXLeVzRPPYUklT0qheZKyK5wgNJmvdTAQRPUJj8ME2R0+S6xHoLwAqbvG4dPG
TaVSq6tDJt+K+pHHTeCIpbwsvJsPckhsrTnkZyk1WS2FV9Y63AvvBlTuh2WeC1s5MYF2D0urdekT
nBwiCRUyBltzL7SuYqXUILCG2Qvg5W6sQzMB+6ERdBOuOwnVZzhbUCV/2U+d1kJct9h1pqhqA4lm
hGfuVTR7iyYsQu3+E0LpkTxs3WqXYXiV4OG9OsdkagGkHM5Vuu3m1/AZHXy1fJNbJJ3ZApTdzNKS
t7SiueVfcCSVwTTSX5h9JIhusjNysh6+bmqsfnuJ6oa3Z9hWyeQEGwxmEWxYcoRdP0ltdvrb+3Wm
pzpaT6xSxRO5aySlECGxtFBXFvWfcfPDLH3oHFtn4YWiCYa4GfXMJdcKZjRgAfckeYQzh6dvPlmO
iGLvRICxKJXqEdfRpoUFTrRMRuE4iNTHU9byRhL+BYjiPt80Gy2Fo9VMAW8OYfDoEf1mWX3LVGDm
gdtEQ7ntUJUeQRBRdkaaAvL8rbsT51nTmLjvpZqLqW6Ikge0SxSi/BwSjJd1iewuYmuRa9PW41bO
46ABN7x5X1DiNSj4RB/q30mvTE+kggW0EZvBUrnqmkQkRNgxJKDKwib1ky6oRAi41ZoCee9nWxwg
V8poQ5Uf4OEKXQaDcRHi3ZptbdqnhEzyYw15nzgwhg0VXUAg5k5eYw6UJSzLxlq/rKWuIswJTdAT
JNCxFSS+qDOJGrnsZSPS479xejGtutm6tk2AWan3SkFw1Y5hc4cuStkz6uRsRw/bxR7sz+tn39N7
StDDvxDGarsDCYf6Stv0BaTyTK8EiZBsYB4XhUKh91+1XhKIrLupeY/vNofShV+4KuSwto+XMPEb
L5XnPI85Hc7aCRRPuEq1FspApy4nSoHZqrhT0Zn6hntT2u3tReNwhUMD7RU+jw+I3H1Y+vlb/2WZ
2I8cht/KaxbnM11PTsqPHmKPEqYh9+OLYdJ0oH9rXIQiwdOuccW55FJEFQ37UCcu8e92yovHS3Md
9H5syG5dPQbwsmm2Ew9Pd2KUMoRi+19JpvRprm2BhGu+qtngdozr9LYEQ9icuEvSUKkyyFHEIPS4
78RGSB0CSuXgW2J0nFE+KIV6RqhfjpiKyWn6Ho9lk56vHPbS87lkDPxLIxYd3WUhzv+7+s/vnMU+
AkFtVTzzY7qewvlAtwSmxacMuJqYNJX725pkyyiSVfmz8Br7i8GNWerQPAK+5vORGqX2yIaDKr4G
1iF3fhacnEkz9kGjeXoSvqMGXFp4HvR9JIsDk6BaZzF40uep4NX8hqm9xmcdu2Anb/fn0NBBMPS1
hnBnH6eqURjuKnjt+h4txc0HZj1CzuM1k/TZA5OOGYl8//ddRwVAo0q5Z16i42AMGIQ7lSWgCZse
zkURFlytrkJE1+CWLQrgcD+YoRBshazIxDOFe8EoxX6vFp/sTWX8Hz9y/r0t4NAdcP3ejd5wWJji
UuZQyWEx+C/GOGo7OnWw1gcPUk40BnKN3j8e4W536S3oAIzRCztkJiSnpW3Xe6gpH7kFx02e/U2u
eGbfvdk9wnJxDqEteUhI6/Af2vJOJvcAxe7GZO1QekmO165uDSfn/8W/el1NufuOaBei4b5luAcN
PV2riv5iKy6dvoMS9G3a0j6z15WLKcxLnrdleRfMFw4OyhtUxjTzVgdjXMW6VRNKEtGKKe8XBDU4
2PgAltE4//j5t0kaFw5oTHVCfpfW0gghp+XjW6c2hC7ahU+uvlu8yTW1+vKX3h4+nAHQkbBy8iWJ
aqJ8juNHLr3pl1isjaaxvDb2119KuwayWZbb+s9pCsdjaB3BjSn5+CAg1OI1g0V4ZNSnjJZ+cFL3
PW0/m+1fFHmPiFm5p1Db96ZPAKx5XYWKFQmTkVRtb5LDx7HW740fOClv5jDfCihtTUEhYNsaBJtC
3Pl2jt5E41Dqe7U8lqmxzroHfQcMnd1YMkHhHnPmpnqeRRofzVRli3pR++eW9lIOuwRj1V5VdvG5
pi8OB1IfEFh37VXoPKzo9DpTv0BZ3P1qlZtUi9RW/TD0U9OnmSzPt+9CWPRaegAQiXG4DqI0eTzd
Si8uGgcG2pLzZYDqgsrqFrQu5GRPVVV4WH31Gb8vYyBGCAalHGwy9PvkrcBRLyzkcAsVDWqN1cX2
WIG9wgJMk9TkQp3QlozemRCI1Iu4lVBqM2TVMGWrqfUsQngqSFzPux27R2A+NLGeuwPoPNSAGRjl
ON9aAKOnsd8bJh4J1cAghIvnE4BMALRFyLT0h+97i8ApbG0QB8WmpJeB6tWm9SKN3DzQEmyoANB+
MjHb6o5bWbyw0aG2tDkqyLsYYWgKw9lAJOcGj1SA7d8K8GpTBiJpYdlI2qxzsJ4iWlm288M1cGXP
I2lX3kCJDlV+YSNaWkK84FJx89W/kI/XlBc+E48+bFH/SGEEVPpFaHt8g3iekRUz1hkp5uxzVxzO
LeAsY4fmI9xMCsvoa4PFFhVQUBMQiI64KJBXygNF7GhRjry0L2LiZ2+4/4wW83stEg2M0JqNCnuX
D4rDzKIP18udP0nR21JlC97eu/m1Pufh8aMvyViKZhATpT8LdSkFD6Z+NkpM9xCjOCxilgMPEfwJ
3SrM7leVUTwpzdKbxH4lvkuUZTowcquxJ5gwO+eLtvxfPOxAb8QnhEsiWvfbGavPOq+y/FW5abTU
7UpjO3oFt2ydOCTbOMUTI6J4wbTuNoFTY1fxcr7VKN2XkLwjvCz1Zl1JUsWbVPDYSFYW5d4Z3e1t
Q1IclZfyNq+tjcJyPU81/xgM7LQAPai3B1NGF1Yzj5Pkkbr2OXeyHsuw1/5NLToMT+nNxtbuyqWk
iOs868BKyLE8CMeGkvIijlv7DhITh+w9/aIV4g6OKvs3luYSzgnozW6fu9LWqLPKPgpmYO225p+P
dgjnmmTYia/H/KPv7Lcu4fmWeVAdegqjWRvTCPI+fOxo8Go9wAX7vW7qdA9EiFptBy1vJn7Q+X4q
UBChmU1n6CQfTFKlzrXPLmG1OwWlFR/70DaOMI2xeh9QWcetOhB8T35Le7w9z7NlY7g9fdr++nfi
2DJ187+gij8fp0VBvNj6ZCcb4zo5feew7ox8NQ44CnpIJdB+hX1lBJcdcO0lTskIbFT2cy1CJ2+p
vA3vQEtOUCb+h5Vv9Nj5pBDISsHD93WEXNBq1wOqHw2zwpD4YSt/RUDTNpzIYWEr8hyUQnf5AVHu
Dpe2f3g2MM8VDxMBkqnXY7Kwf94/ILlaNalUN5/y7YdfhXyIdQmc9rH11X1qY3dsHWPtfhCV4WBt
ek7rpjGwhTZjmaZW8WCcDgG+oItlrDu+C5JvvvBzZpy8GG+6RHFBkV9Vz3OLDnapIA0YgbFWDj8W
EntyZ58NjpP5xoTZ13WjWyHrKeRik1swo8zJTHzBFLdhgWiJlfJSYRlq17x/nnyLIhnVS3FAtQGa
7Flf8NgM8yTn9K1QqiPMcfDtD3ttAXEi868Aw5knIeE5RN/uhQs0bwlmF7wFrsN5FREYgF/Uy/lP
D+jXIFc+4Tqq+I+RYTuAUwSHGgiVylvzc19KwFGU7q0FXGXNZQU4Xn1b5K7jts89nY3FyyP+mk38
3jaZntkn6EJXrnT/j+2StWGg4y+GglcB68J0XsUGKXxrINJxQiA3oU53fGW5f/Xi4mR3j7FeWoE5
8m7/zlMJWOvoywsnJgKU8pp1o7yknjDDibU+MmuxNw7MyKktWFRyI5AJQfDYqzO84zwZ6BwNdQOJ
DEyAhBUmeTfXBdIct2l/VXTwVkDcelFYAOLk0nkp5B8hdvZQSECCT8TacX1fKA4Yf2r4pCmQhldl
0sZcpgyl3r+VRpebfy0lpAbJ+almWG4WoFeCJOx/ni6j7TfcTvSJrOZI3y11peH4DcMxA2tpOsNT
zGAOA9kG9mxuIa1SlT/Q+1S5T5zKroA0bi38sIdLLryUDDzVvbKdjMujlEJpIuFSDL58K6kQpRAI
hwIbelyr8vNuz26YXXVO3xxgx0GjfDl/y7xnwYfUhbP3fpU5CPCe2LsL5E636QKsPuLKE0nyO699
DRCay0izCWp6aJ0zeWNYiP3CKmLru1w0Nz5iSJ8FzYQFVzPpbJkBfg/SPi85Bqji4PLIp5GCyhIJ
kzbqJc9FZcAWGsSHnjv7jKhfwMRTuT6UxoOVeA8w61gyvytiGU3b/UDj7RUCaedO4s7Xdy4geK1p
82AM643MebaKke4P8zSq7OAHUdyR/IwPDDoJFTB2WtTMzkI4nyZaSRe668FoqEPMqvyvfEgWjXoZ
dbs2HcPBZ+I6aAt0aUoP+fDLS8x6IzSi4OH/KxQXd6c7HorcPlDAJG3+pM7yBx497fukmR5yh3Z/
1tsBb8b++gL+WVjEsKjXTlBh2LCpEsms2J7XXbH0cZPl/5f3ygnrhA3njsNpMZC2meEeYb2BMn4R
9b0ug7tNuYlBWnuZNLMZJ+xkDuud9JxDbfPijjkt2MvAZ7ldy2xPgF/Qr52kP+knM5MMRtinQShv
Q4Fdrbo6UXagPEpbfzMBXlX7NYZL8g5IZpVM/Zd5ozWTgFo99okwPjeNWFFkURsdBdyjVpE0HPq3
YQRjCnsZBA5stFXwPxLMXyWcRP5xso4BZ2vMNo9i7iLSf806NdT5/w+hsp6igDa8DbgBVeMMQz5u
3vSZN0JHUMnEnOE9eR9Uo6/kCx8xDq1WYdsDVunx/1pxCIOTG0IXYsJLuwdWpcg1O1PWruSFQI9h
CKLU+2flaisnXIhrosmBWbi7PtkHDApa+W/CHPYiNzmzM5yC6gVIJ4VdOgZgKkdMAhHmDudJlS7J
AbCMt3mqcv/QJvevY2yjgX+HE7gpS4Yjohw9LkM7W3P/Tmt1fWYGLKUE0UZQw/lirIhA6p2bgKDe
lspucyf382Eeqr/JQIaK92zKLr913SYQ919EHAKi1A44ct3drS296uZRUjPNErbreXB+CpLvJqzu
LWzGDP4lqUQVO9KEyqUAyHs7PxWmG16hyaK8Kt/xjCTb2XZu3s8CvJI+VjQQJAb9KCYQRHu6+Tah
jCUM5BjwoZ0xwRcEXixri8csxNBjiuuYruRIclFrwt4faowABvNTyOv5TKtbf8AEUF6wIRZUY+e0
rejdUizxLVYb8itAsQdl5utIoRNqb7lVBgmAVBJsR3LaHafSw61ikuBs5M2zIiJ4wDkYHmaT3yeW
xS9cQOkmlmmBBZ+hoOGJ6M2kLuRBJCF9Edw5dkbimHTL9Jz4+SnTQW38oJb1qtMurUb0UJUD5tq7
VaFjJG2TJ6ErpAlkAPnKeHoUzUpoWAiPC/N6cm/Z7nN6Rb/1O3dGGodZceHIR2tHNWbnikbkBuJ+
Dl/bSTFursvr6lXoW5rupPqC2b5nJkmjUzfB2T4kEAfzP94fpr0c5Jt4eM5JBXgn+oJlP7I3BOpP
WWVcpbPbHEEJsCs7mYP5HA9FnkKWLGA1nqdD/lWIQe/paIh6v6ErRvfbzZvWz4YqDX64wXHyQB9U
KwCMgRqL+B29/5Q7F6eeu0N82lL9kk6sMVPvOmpR2SwHbjXdfP4NALtBuizfYy0ouU8ph9NrdGw5
B4OC1/lVu8U9x3tywC8La62DSqHNcrxzmh907a9na8pEcre7zDgh5DiHbDM4KdTwFyKarsLdqgwp
O3ubyZ3O77Xby+SrqXeoamU+z/i/9Ih4iSvsOibPQkq0XRP4YPD8r+KFalpWQCTo2TVpRG2kUJI6
Nl+thOWNAspcNQtpu/gpPDKL0zLoUbJjDXnbXh9ABWo6aoXqGE5v/ZH0jbZXUIUv28VOt7s9d53n
TJrXDWeQT+J+oEc1ulwUEJirfSmdAmZi5yONoiwbrWGQDCIk9QvR0eQiH2xp73yp9EBunKeMA+ob
8mQdQylh25YqopMwQCosK6iRnKPl7QdBCSlnEeiMWzO2/wTOBPZE7hlJtw9eMONvFOJ0J8PodPUg
jfznNmOyZJbq+82/4OYK2HgPczQkdXlLQIWvQknroW0cKqOaWCO6G2dhw5gFSmxsQlC/T+doY3Id
ZVNyVSO0vK5+8uI8zygR+NvKavhbOvyZBbnbJJlGksg/dVjZBK5IsauYUZb+dA8moWVRSORQltnn
uKSy2udjqErtberfjdE3WLJGrAFjMVISBsibk5AQ02qdfuOjK/An37tgsTQAPCzrhuyHVjUNIgar
VBJABc5vCQSqI8Lu8Bqjphnn9WLpEIeqm+LefXR5OCOZDYZwdVEkO3gzBwHEe0cWa+HwuKPfszH1
EyiGOCBnIxcs1jRgPeROeYCXzH84DuIvRc/faWRVoEysUsAEJxZe4q3RezQ5MKfmU5Ssu+6FtO+r
+qo7q6tX6rQ1UkswsoD37ixizu7IEQXpljOX5P4io5UR0sapBTnA4yM0GBAWMG2lMljnesAuX6Wr
0L1ta/QefJCzwZn4h25wQ1LD4C4RZpnsjDMfGQLisGJnf1XEaG3VtpARaqE4/0qL42UxgpU9RbnL
3wK5HQ7d4FBwEYftbhwScsVcQpPPsTnWr85gVRKNuRjJo+Fv+5o973RTyhUKbNpKSnsTDYW9GGFP
oX8SX9N8wQZaBgnDvhMMb2cBjWcVoNszW3aNL9dXGbrh+pDygRDaas7obc9O68iT24RR84Pyx/z7
CJpX1kKbyaYxXLHSWl6GBEPNAn7IWhx4t7B3tTvuGKnho0wUs7BhXE8DoCcTOBQ1PyzrGyHAXDx7
bJD1GRakABd5RIWJC/DrLhIxLGCsRlBNRIfwAtWSpwH9Koc9PN8/6+sEFYMMRV0zPN4LBUYvMv/W
EhbYVrHnP5FQS2yDlCIhtFPvZ0F8oh+k5t8kAJGsRK5eBBqECPG0NxPOfmzehF0sOtcN+yNfRpNe
j/xdhiGXoYkiv00Ai7MD45wnxriBwRndyRFSHBOSlNS4OoukFz4lSGqbrAGJ/GORGCg1NQm0ach2
1jVSp67YQeTU3TBc8ExBGUuuzBZeC9/QSBFjyEbdvWMDKyCRZcho5o4TtCAXH7RvaVIdCwagE9EV
tY02P9LXqwK7lXP/9IfIS84xy0SZkmSA1XLwFKREgVwcN9XOoyyeRtS8fjusrzv3Z4z+h/pghBwF
e6S5Ze1kqqRR3iFHOC18fOQKilUYSzGwo2I+ArJG+DCCQHXfyhgLC+eJciz4ntjb/fstVzIe8PLl
JUAVjQuG/OLVq43PRzOP9GrXWO3seBKSebjcw7No7BDiBRlpq40P5JXQiKYNte6PKlVmWZbXXMkt
mrWVfwchojf8rjZsk9nKGQ72PSB60HxPgeOXBSB61u+n+jTRL4E/x//8Q2wlKu5t7OM7cNX1ioDZ
ooVqmdT3sHfw8R6K/lH1qET91Pzs1KNDF+6fFNUTAA9YRUVhNH1vX7OGTQXgWEOmDiRjn3d1rCKp
CtL3suhzPbR4ensfJj7ncf6FC23Nk1DgeLylDckwwaszAFILIIhRzb0i8ZWRFxiNdNnMH2B/xcZN
43V0WTLMmPnIrnPojnslEc9dYaExvPMXjaiIDONhGwrVF1nFrZG0HEMI6h8+cUVju0nMdM9ZKTJa
7eqDQonFT203p0LOAnhbNOjwQK/eEM2HJj0/HOYR5wizYkSI2Gvu3YK+QhbpAgtMpXo80EHOYJOO
YZVggD63mKT0IbVp8crOLfxbt0V7dUKEZxDIHzRXQmFUl2AFoY/IxVeLC7yuIH/i62spXdCcEocG
EUvQgNVrSCIIDva2IF8bPWCWtg1iosjRTX5dJtkpHCf/IgMXjlSLRBt6qX/dNttipQB3gbnrHkT6
9Y21H2Fad/uck3kRGO362hK4Pp1vEMK5ONurw+xrVb1TPYYFewTzD5U792swRG0Q/kMWRFWZc6mv
OFGrnbDkJYbDlbAFHW5noXjn5hNhdkDbcc14GAGdR97YkHkVPzvtCrn9DqpMqdPttEamV1sffeEk
+WhVxVPzUEnNNQY+bTEqWxuwPNk7IBaeDcDaN6BeXcsGaxnuS4zkM3mlTnRzaMVFeCjR5yLHR0Cr
pQr7onMh1hXP8DBQZwhhNLhNfNhzcrUblqiyz5FKkrk+ucp4TUdJFzWFQBMlAAdEKdg29rlInylj
YTchEaEi3QzcElaUdGMXcsRJbdsc5j0in87Sa0cEEgk6EQ23lFzB/PSMl/N7ynQFr4J9LGoExixy
ZtkxPAXhcMdNHicfjoO98bGSBczZopvav0M6iAycaOgqfqos11f9kx89RN1FbMWl8e9U2DWlzLCI
N39VsgMO3cIDYkxwB4cZa1r864oXxO01lAdDzzLDv5VYRbZbmxvjw7vGFqlNr31QymtNKd2b4x6z
It9nVihZBbYbLkZcfIq9SP/qYwSEcJEXITR+NIHtq9J47fZzMhDaACWMQBVj/ds/NB2oSodRnxT1
ZFKDGNVvKe9zXGxcAf5epXRIFPkSLjr/ZiMRc7yRwJ5G5WrzFhrYrUwEyUnWOgIlvHetJaziQUTK
Bh+34xpimrXyxT+N6ui7MTTbLQUfWf5om8+lhCpr8AN2JK6O9bt84Lg1lAhLa7+ZnfpILPYfcwgV
VG0K+op2rHecBoKaPJ19tZDgf2Y+PevGOs+hhedB9RmfjOAEV/4U6flcL394ET9crOV/9Skzi1ue
zk4WEUIs+jhAJFDECf9FFMSumnm3yMBCrQZLahEYcVloUxOkvaF6T2szrFWzIPlI31FAM+5e1X+8
eYDvRCskyWzuVCColKeamrkl2BPfNDHCaWNBGFNGWQa3Uq11e6W66D6EKBdA2SP7FPxiBM3oIFb+
MXHCq0lC/t05lV1s7/O8bBzfObJLsv9IIyP/I4mWVl01mEu2oW58A0WB36zzteMDfWMzKW5wJro/
iBikM4/U4+Di8lvln8WqKPvrK5vijn3dAcX3Qy8nTZGUc3p1Gl0AJyZEJdyzHhUhKCkpTkYWPkCI
RiRSuSOHB/QVVccgcoxxk3150UV3YtQfYcJzdao8BpqpWg5132v5ydJVytTwuXLrnn85rCQg91J8
4T6Uyfy00ozcYTbmMC6zZ0TV5XGGqz2eF8ipNFGQjm2auW6ywbauCjc0K41PZjLHS+PF+n3KMpKq
t0EX1hUKWXubVC9Clv02QtJpuIv4qvhvWAeW/uzeqIKKtOKL+zijv93cvB4vQE7ZKrfP6ZZHzLcQ
QuHJJZGz/xMUWyfLSmNOcrVq9kwiDWbs6xEc8FiGn9Q6YnANY9Kt/WKddZUY6V3IldLd8nsYSSH1
61lE85bv/wIVNwmrqisMjIGqbA43ovYwzBWBVed6N3Ez3XeD4WQmMX5NB3jLIiCNxFZ8NoCAiNx6
hHbH36GRNANO/wuJ2Rb3riOz74ZKp/cgPHeMV6xD63qsCI6ETCUSlYWtPE8mot3cO2PDmndQTr8/
o7d7npDjO5ZQVDxTS2KNFABepcFdKktZ2r6ygtuMfv9rdfCmPk6GZBtkEbQW8J6mkyv63gb1ayJE
RTOq57VQ+7uG7+4/oGGCK13TKuWZB8iZT03qcLTAsrmDB1PrTeX1SgPkDq6V4qxOxFSzXXOc7wi+
6CUdZ2OUYrlT/LKIVRjpwZgObo3YwnIs65g09ToZoWQgmdv/fI4kPcfE1r7mgt1b1FkzVtLcrKKv
wFM8v5E9ExuNiW1Zm9FKcjBzaHaaPWpSAMtgRRUEpTKgaWZxjrP8U/MwPAdxu7wTn/ehMLQ6nfWm
EOrXlt6qLapU54Av55MOw61v0TA4hOiK53ECS8/HdQ4rIhF+6rZRr9tOemsPZAXHo4MdnO+OUEDB
bPiNH+wrCO4dAYa8GqkGKfJUw6EMnPwHUxa0NzsW+qNjfVdmXPjg3U+DGoeQ8kv2XUCcyFudU/Cy
kihxLYQ5Yo4aTR7NOQko5SOKhb/8CjCxPzLrDlRNumdcdIgMnIckg1tzX4k/s5vXNmPkBt72g8j2
xTTcp2nAxvCJqeDS0vYGu4jOCOPTRJksLe1jl5CSYDPAGoiODMIc9/3VNxiMwt/d6mbsA6JSvI3b
dGiXyMoNL4ogWO+Wz9la+Ks/vSVM8sdQgy6xPEJ9EdIrT3HqzbBnvHYDCnItDUda/ruojzSg0oT7
y+guTOxmQM/hHDmXmSAiB//rh1yNLchT/7tUhAsaBJl+Fikc5wltgkAYbmg1pPJkKKIMBCAmZWf/
gAyrcwA7SKWVxLSVn1QGz+nHMUdLnjFYiPmih3KyL7O8c89S9Q6iZyyvKc2piggqFRxkGRpzZcCj
SXqFNAT/Tm++DDHj37cSRTQ8onC5HfSwX2bma0c4WijfhTHTf8UNma5dg0zvqnKuN9wNlkOpbPSX
pkRyCfutaBC+fnKhPpCTIHdHsbnBJWV7bm/yY7sKc4U85zPyw2Jmbt2t8HpDTqRtv3qbfy3a/SRQ
DcshuzbqsWaYnS1iOiKqC/dpDYkHvmMp1t4GSgFLnDx+sDkqy4HjaLfY7q0XtflI59R8k8YF8pDQ
wBDPAUMjASkWJiy13TLEkjIn+nbhJeh5wkk9JFepC3JF+PnrO9bFIXXwKKMHkDCohEPtfTT137qL
RG/nRaFyTuulK/iuwNUpg9Ln/1AY8mRbtiYhCOho3g1H4X9A2i73mMBuzGYSzDVNPxIaYA6jbftY
Wjss2xpgogEogEx82/HrcPDHYlSrjEjdFzQGY0PSJmwJRP0XbOiJdZXM5ibCRFUvVEtDn860uReO
FyPCY2YZwz1evgVxCGm1AxePAVm14mHTsz/Jr4q+su3ypIkEBQckdgo8d8hVZsVIMZVjS1WCwosB
WRfhJ2SGgO+m84qhRsUOEV8dKOjY9z0geFPRUo5QSrsCvB6ivFDskD7ciBgp4BcV8sqff92sTAr4
bzfOxA3LlaDghO2c+OE1J0myxDUqQb2vuuqn3KBNFWnjopLwakI2DTByhA6UZLEhMwwQFNjuNVCI
IurHKz33l4h2sF5y2ZSb0duzWNhvV57kVNKnbXh7RZcw89VGcrOETIE8g8qkNx9aQi8laJbxA2Lq
aY7UyW3vdMydJLc0HfezVn+IVUhF3QVstgvl6oa2jdu/qnIl3W5gyJ2VaRmVefdaS609xpr74LQh
bNauO1/rlloN8RSZjxiSm8blDuK7rJEBQX/UjI/GKkQ4myKfa9qw0wpiUWpxUt1tm27ujjg6fetr
JZy+GYb/jiC+52lSNwFjfcEYoE71ZWYmEs1Xl1Saj/Kme07KjULCQk5j3FLx3tixZ6F5w6xAuTl7
QIQz1m3O1Ypy39iGxMjGWO24Gut0F7ro5HWakv3L0TizzeTf4kZQAA0NmCpQxQfiUQD5Y9T0FQNm
p9JX4fUmoDdQnPMtQsrVGAQqjFHMZglAraG1yCZf+ng04NfI0t1CV9WI/eybUsPMSFrcQNTIazuo
zeEa8Zzv553Nm2LbBXTnFf+5bmf6eLnS7JBabnIM/7SIBRnXPZhX892DZ6naKjCoDf0ggGi7aN3C
PSP9xOkTHYEWCb252GlBWI118Vka2nnCfupAnRz436jrZ/LrWIWDmBMSrUFPPz78eqetpMY3DeGG
HQfiY/AFYmGg0i4wqGrLciHrSI9NSDBea5R0UlKnxuKVCDl5B4XLh6o2YogTtA0KIuVlo9sx6pKK
BgWdVMFHC1jW+FNbUIjQkhgM5r787KQTL3J07bZFAPVepzevpyL4I3g4ISX2OXu1qAb93x8febzp
QWudNcdVUXqm2rJa50IGCnpGz68monD66edWPzc9j0VZdOh2R+wfVluZVEQyEdF6G7Z7/h/i30WU
CGyQ0hY4NkGzoKBBE4LgnQfdo0qSn2GvbUJKCovq3tJo7SdhtLYkNkUYFPHVjDiN4I6GYwelzBMp
1KOfr2erSI4sPvJqzEZDoA92BL1zNpGzb6OiTZ1uoeZMioWu7NczE/kCkmpOE/EtdK5StXRo4ImH
dTPgxVZO+7RIS7qMPIPXgyH3XLuZ/r+KtpCZehzpddNU94Y0gAY2oncTmmSnh/dX2NjIXWzb5opa
kMWw5ErShnuFO34/sJ1oi8knz31GtseYbPWa/d4kIcL7FFFBJWJZfDQMsOIL5oaYnrJeZJudd1u8
etSC+VakJAdBD9HT9mPMNwYV6hzmBGqRXRK/bKTNh1u/WHtakyOLLkC3XXY08cgoB3yapBsXmeXs
Ai9PseIVLZNgqCUStoUjiQe3/6XXwTQyJATyXDpEJyTNtFjxDuYy29y2rG/nnqu4tvMQYoEtIzLk
KD/5aIgSY4M3EuOAWhBeIrdKxrA1RZTdiNtTwvCvxQLj6d3MbJelVYPaJKAMBPxij024Yckjn46e
6zKgtYXVyPqozTnshXac8rqRjnXkcG/+tKn5f4B2MYS0q+S0LHGZ0n5Jxe4vGpqM22uJnSjkftDn
Iy34jKeVmdmAg5blxJ+YNSeNnSdPAnIuoKxH2QD3wP7QJxm+U9Q/m3126PdQgxx2OgkXqmgDEnym
tCBd35tsYxs1GxnSlHBIVLPo/FdzbXRMcxtVDn03BX4LkjrEN0vAfXyuRCU2NfS3b5b+m9JoJZey
bOSsNrJq50MmXFDJagG+GfLgu2cjWVdCDcqshsGX/JW9Dy00y5fRq7zKBJD6hGvEhtyYohvKtZgp
VHA4hLvKGBW0deHtFKtdn1XrMXHAJeEAvHOU6Dmp6lE75I3U6Kk/4gF9T3qOr/gxL6owJRQVgEk6
nC/8Rmv1SnQNDfXe9gkAF7SU2bY9WaMF1Uc9E+dP45TQJ/LLDP2pEImQUIyw6ikncBEyfn+iB3If
T2VJXQCi6e8J5ZxvVjpJF6m4ct5QBG+kN6CE8J/G+aYJBR2Y0uIWbtA9vWTcSbvUkl3EMWl3DWwn
1QARc6STdi8CXsOT2EpE1wbVeDg6XkRo12Al2C9Z7fa5j1m5Or6UiG2nxUlZLDj9xKwRp/bTd6Mq
6AzvdLPUV4TEVoe+RD9En8318/2mhom7kR0jY6CNMz0+e0vP8AboUOLpDVI8aC7jIeu6kWwOL+lg
AOANgolQELHU4NYrw8JbxTtxOvlMeQdsETyjIB6Wbf7Xh3SqNvI2Q+4MxJZ22LEfqoYimFGQDdKg
hf+TfsqOTwPHKcfxQjTht2Zj48Rl7qxoaxWWPcbQBxlZxhi+ZB/jWMoXGyCZzCP+TulXsG7zCmeI
l53ihOwbLVLZ6t0/0AXKCxA+sN827YL7jqfEiIya8PuvwN60y0OHmiFNpE1M54YWE2vHq4XK9qzu
9K/rPYzzcbuq/BSKVbvUrOXibKy4on+kRjGJdUzZZzzeLbMvkOpwMQCEmuUJbx29+r7D9NEBW1DF
IP2SvXsUv75NH8xoV2IJJZ5lNnVetmOf+GE7Fbvr1nAbgz81OMdv9InUCjEa8KmlLTUxzUh9rQZl
/jaiuBNHhtAyNNvcs9xnTn0jcGFs9PllvPG6L3E0p3tPaydtm29yWgvSuoc7lYbSbNmQ6f6rj32u
rD5nsDxPGHRulBYJHZj8b5xs5G5WGC8Vvfl9geccAPxWpKN+BaDlhjJMnAL8nTQ4j9XxR2zqW6kJ
9YUPJw4F8Dg7oFOzVyl1Y/bUTWgioOLmDjVviUNmJghwx+fpOYA4cAifT4RHT66NZ+38eGAEivXR
GolI/DkJ/a9UVyPELEnD/uOBsCMn8/I6yUgIwLvCAIQ6Ekg0Mdr3zWodpkJdP+z0UFhZb0sEfnIX
53nsWk7xWZuH4KCHaUZ10eDPCMdbItGW3jOzka7Zs6CHM8okNI5EJ77z1CW2vZ7HWNSpPYHZ1GMv
bqZLXr1sr9D7eaI8OoBFyxYygF+AkKAJMZvZRM/xLhCBwB80MkNErpC5YfHdIinialLctplzioK9
gMqZCREFo2Pz//ndnxgNNmZbEdBIfyVAJkGnUz+FaaDyPdsHq30f8RBmZXohJa4+nHmc7wnGG0hw
Xnd07Dbt/WMRNtoK5xDZznRRmUkNy6YUC8fciRoDIbYouXS2UOX+V3FjcYVMbj4n5SiaKC7alVck
Buv2YN0WSsZzmMfGlfiFpcrUllQpft+e3TIjNKVfZbqJbP9rnHo4vtpQJ8o//XlFqF2rioqGUmvr
AK6w9Jvfa/CrC6yfseCRCzPHcVFjAOzZ+OzP6tn/QlWEyv8O5eQ2xQ7vaLsmAp1TaxnRaZJO9yqM
Ol6Pq0q/K1r7RSCvI88Mhdj6UZ4V3x5lz5mqCM1NYwc+mcqALz18ckRM1l/+CoYg9hBTrYH6mk4+
homQdy5Pi4gfLmgp6B72QwIxL9dpuwFf9Om0qcwRtpBwBjPNDNaWjcNr32XLdHeTgKKQ9UVDjAab
K4+CgB/TKBXtSFXmTrn3rYO8C9loQ1qPxtz+ylHZyKIZH8kfIPedcUv+xv/+HDU9BPGBJmAWRQlq
Gre6OjrcEeFtIYDYucHq5IfKjPIMUXfJsGI/bc7UGHoj7/byinBOhBb08PZZUQCLcSXyJDnhsHOP
MIlebvW9VZHG0Pd6tMi4G1bZD1L0B7/eWV+J+TXcDQuXZM2shePtFrQewJV33qBfDYLAyljeLVFJ
0r0sV7fM95KAv4F6LSeiuP7xbJ79FNIqj8d3C4NuEQra56ovFHY6QVqPCWFnYcKGEMqOpn0Su/dl
xjSOxxmMZCAvA2NwIFP+JHBn+luTQN7Y/ykPI6IxvWSzYpLpX5GJFjoAwHH1gLhvtkJIL/UMgiC9
27gGPP+URxX66251DAGIluK51YGL9ZDoQ0qkvhCRR1mBipYdZeqodqNuwvsMjiYgVkLOiD2/paU7
ogUKGAYt9mikFcCxqo9alFGcRbe9Y5xvKrjCRqqDkPme9a+5rh+6zTJokxqskPkOloVl9Pw+vtYg
hDNa/LYYIbZ3SLCutvYfF32lOXipdcpzkGFNnH/E1vxkKt38V6kAAwS9HX4emGY9cdXg69ARhSZ7
tJ5x3GWOFMM+X0RwschuT4hEyttrl2rIpTulfB90f6C+JWgmFiEaEGZjytAurxb3WJtfqbv/oKs3
63HJVfDjC/C8HNLT/mbmIKDk+xKIY6qcVD1UGxwjrRpIhlxBeO7dpxx3WsbXaufpM4hwcnMwt1RO
ZliCesNvtZFCktK+o5WZxp2+aWVVySLbMtauDmQWhNh1zRDxtsi/SnwOpvs1bBwJIemi5/sqkdQ4
fEgnlkzzgcO76mOnaL9gF1Lral3bOhMTLAWXT+6V7VKFUvNBr8djiwDS+wngPSIrWDmKjaPKp7G4
CUv2q4N8dDrGjciF0M5Yj6hzWw9fEi3jrZ5Esao3CMKvTUkDjw9k4voCgE5HZymIQZS5G+0Ejhlc
45FHu1Rv8vMF+7OCvQ+/5i32HZIJWnq6HraWuwSEq+gztLWhnjIY/3h7nmPGNKKPINRnnD1mS9tY
88/XKNEZjR8GrryZNIzGZtbcIMjkwl2KOTxHRJAEISjMmxLxUHkzM42wGvF/6M+AA65r4VITlbgL
wJHEV2Ns477Y9i30Yrnf8v0gLOmvlHNLELmg7SV/kGgLFbKSMvaTUydbKO5YMS8OviwnmWwnllDr
7GPYPbW6oR71yBRYPjf1YcTpNmq8UFIGl9IURC2GQX7BHKptkqBbLIeVIKR0e6fhk0jtFUwHmpu4
9QaQ1gAZb+yFqioLtMR3y96UkjNLyh1nAxCzW9b+f50BTSbswhuNjGpFtk/ihoQ5KHmudnBx3r0Z
PNmkmvbh1+Il4xwE1cEGM8nselXzNZ5dRalWQiqHzRqS4PVhkGXlMTULhZXM9Ri0dxc/ynfMet2k
DIhdGgktp+vK6bSPSabwDhZ9owiVJZvIZVA1c1JIfzuX2e4yGiN7rC0wFnM6kHLq1DU1qLoCcC/p
YkeGayYVDyPXNZuAXezc7PQQGJhdDRPFQAOB0T73NAeyNPNFsOn3oHsetb8QaU7kvA43VMXUhwmD
IVNPIrGjIwyexowxHXWSMJgIOMVAzOMWZCIGss60CNYofScpCcFML9mJJ2woTRdz33Urfeb1JOI+
dZyatpnC7ZXUsWJDJ+A3hleALPM6c4fLb8tBhbgBojFy0VacdANLgFd2RTqzBR/KbvBqvCPJXF3q
7ClTzU2ynVdUHwDSQUakwGZuT44GvRIs5m9kKmTpJo+9xyVj2YrY47eolKdTb2E2V/S8lQtim1Hw
IholOTpfu44Xyw1bDdDChs0iO28X8jem/2CpRtLcVaeRf8cudHDHlmCPtKmitBuVP7gijMuOUMBF
IESanxNH/Bw8ZwBNnil963Y7uUSK4ULdEtPBqTo7mQBdO/c6q+qRkmO12rQ7AvjxlDSVQ+pgnPFY
YdBD8Yz3LfVuOMa3Q52L3fWaT8w2A4u8/5d4wcIdjVBQQ5VfbRRUStnmfyuhTrbLQuBWfMOvPbYF
7hkzW+56BGfSHlSq7y7eFK8wshquGXHvc/67ZeukghjwdgI8Ju7z8WcgT2rLgYvmpslTePdAlwUp
7C8GeQbB5nQqZWY+DTDtM84pC9spCgfnd096Cu++40e2p3Q1owpijGOYH0IH+UioIl+Z3U5oZ07E
ITx12AaqoHUjMhDl+GTLdKEpxcCTSq4ro5Uw7o81WUKHrBV/d3+FT+XHffGgh4z7pTfVk0guahRa
emu1RpVuU+ewuNJb4Nul7Du8ngCBor0v2LcI5y0Ka4YDqkGtFoTyGZOPZ0cGxPxbf1E2U6UkyIez
mQXa+Fho4i3C6eaJOsxXvaDDx25sTOVbX06AMLXbpqQKzKgT/9TdysJlc4fsamQ71xbo7LIMxLVe
RSnZjsp5bIxUQWwMqVPpBuGHm8Q8nvBVLDaE1Amnbh1v+VYg8lmF7ZlN1kDYIVtQ4XOZ58HtccEX
xlvfKQFYn7eIS3wUyT7eQGWUsyK1G/iqq1t8mib9mClAoE8j6x1jzqtKnxaNAUcdZz2BXJioWdIR
abZ7UGD1eOo82sj98Rqtr01wG1oTxmscrDllU5FC+0GX9yF+eVH9GWj7ZfcsCKN1Ehv6CqyzYazX
8VLbZbAyO2j7DL19w9PAcXAKCDYQplL5zCkt4m+k0MddnS5bhtHdsJwGWD24QpYIFPTf+zpPkaIj
ACrK+uxytKNWkvdGvlIr+1ASN3txrHsXxIPnZdgNKIalT1Soi1RxjCUp7jQbm01Zt8EwQEXm9FXH
JGnYjeAtz04Z5fSf4flPFV6FZBg4BPCyQwb/kFFZWfljvk92Ans3qK7vFLSCAMxSOo+8cRz0zWU8
WVuaupfjYoZxJFRQTlzQjHSrvgXORWAWEma6fTJ4MNQMSUNQGbAeowfW6/XclOCwFjK7Dnf7Y0xM
5RsyHhxm3mDbzSE75PyTQFHp0Qc31//LtdwymDXJXYZdlH2aloO4j/FUkBSyAswyLZk24qIUI+/x
Z4C/NUE24NT12CQmUkdXWzMvqBiI27Y/VZ0midkHUGPccsbRcSp2NfsTA2QfaaX11V9wbEbgHb2H
YqI5KTIECZDpLmumL96kcOPqKLSgGHocBbp1pnAoZpdczUEIhm84HOtxuiel5FO/rmcdi3Qj8oGA
wocVRKKfwfTlpkLtL96RBYrxJJ39VgBSmf7LPKi+FGj1Ma83vfdRhB+hLkU7AmsLZPDUwlmei2Qq
KV1Uo4f44lRAPu7eYoXKzYN8l7hB/tsLlfE5vwtWhMHLRGIKkWkt/fI/eRe9hGmpLoX2+IO8cFJ8
XML6wScopDNWsPtDBjA7HUQlBOmNM4KvtA1L/bKFX2jTYt3Y46OK9jhzDKtfpb3AqZsJSKQdQTPg
tewtizSy/1j3n6dEVNgqfmCT7sU+VDHDkCt3AuWeEGcowZ96k2j4yfCn+HSlRDhKDSPwwzIULEKu
5MwTIzyjXvtg3u5tOpliDdPOsf/jAIDJuv20D2ggnLRKAe9bqeT3XOWAyFcueK1ex1I1xGhVlhZU
e2TilXEIsAqTwTSXafeaYjBdsGfCT/1cZh7TpL91XcHRNYY1EaUk/dIcWq4VkDGUsHBr6PJt+sdw
uoqrfqOKrBrBQDdRj466Nk58t7UPjcA6wYWfm5/VyKO1twp4ydmlu4DM5aLXLAdO023HvWZbwTN8
ggGhe+ikiz5m49zpscglHq+XCIrc+URYd6oztkTRLtm2K116Tc++RarehbJ52g5WoDFt9bynLv/G
GnIIfuMp4ny3NZdDd8jUyrHZylTVOYRSiUPj+dWPVwGnqHcV0ususu57Bj1ayoCzhOxiDGN71dEA
zyvSr5G2K3RcLRQJpthdLMkpqcHqNm26mRzwUFMF9Ar6XjtFBwLExCsAotw9f2s2gCaa0nLP75s0
0tTWSVvdFsDbysoPxnS3Q701XDMFwIt5glkWwUgOX/+C3Ozj5jIo8oMOy5JC+vXdDHZllOxJ06gs
iVDjbqdcVCgPudpDs7EjkfNA+azqEInlUQ6eaqyfGOez9XkQAYfXsJeBq2RGMd5ZiaQkEgn2PMyh
ku7hsnVnIoWmY7YKzCiphj/CVKxg+ILA1JSzLGzrxNqtzq/+NmQ+G5Oo/6FXDfbIDsrZqtP8C1Em
jU83nT9kiOUb2UK23uOa5xiPqZqCxc5zMHDLNrsSQXKaMOsAbQKBxUTluaBs39mnVrgVQ6DYbODr
YufpAfBDgOGOCCUgLLjRdA8Ml8hQVTcKEl1g58zG7xxMi+C/Vanub78PHaur81QXeiytmiy29+5L
jfR7Rx6WAg9KxzNHSAYg94DbA3ZTYoFZsJlf2mxpnhKapqqBS2zpyaQx36UZN19AjgV5sCgTf1NX
wa0w2fkh4j5sfnzMJE8vZRftzg2+TzSEB3YW41mW8yNu1OzxxyC7I0cdFGw+qvUaSoVjRVqrRLxH
8Aanm8e+mx0SIUNuKZ5HWQ26V7rQ8YIsMANATLAlmwnurCZ/LdVKCStj3oOGIQmGPPUt+dIGuJGv
ZiyQRIPHIvCE/7m3Zkisxg3YzBDnsniCpOOeHtY4BMuo6Jx9+HCAMFQPOmLhFSnfIVLXSXToRqeO
tJWxIXurAfk2L9m2PrOS4AZ655pFjXJfCdtLBHS5poInfmNgGywKphCllSA2EnbS04uXFICuOH0X
gAMmvmyRI48nUUGt4ZoYjd0MXu/5ZWYEQVMd6pbOr7MFpjbN7fvIwIDErQnyHqZlziUEB1/aA3m3
Np/qHOUj1beL11jjzUWt/9CcaUgm/YLjqVMGfS0ZYFJv6jvYwaBrqzPcUAQub50UqwiubHBo37Cw
nIHFLqEVur4VBfjtVOoMo4mVmncK17mNBt95yonQOq+tjt2ClyhaaYc/EdpUNcsR7cMbq6PIY4jb
ZIG6T5v1NbS9FWYZdiQUeR5uLNKdS6TbG15wYJNrJLZo2eZy36V6rD4eS3rWkfRa+MdzFtJhG7AZ
/myuM6nQwKVXXXSi17WBelhNpmFetCnehdG7zarGYk5G0P1lTCrBCT4gvOovSOIQce4+xEuWSHJ+
sds9PAiVY2DyAv/lCLMfsuXqcPHimGb4/x2k3ANk+IEyYdEpMMYnSlfGPFzI2REEb4pR3iOwCDGo
Mqwx89gA6IbKdsMqb4f5Mls3MuZGIOJhlOVYTewqhOnGpmjpYj4/iKKai0bvPt1sfvJ4uyO94eXn
CS8e6685lngWQKXxgTV6WLrn9i/HBisY47dqmhiELCPXBXp2XXsEEXPAOQg5n+Yo6IW8ZR40SgyR
6hAmymaYUTY0ZKcQs2pe6796GdcqQH+DKkopJO7vGgEHTjc5ruaH9ViYOmXwLFJhi6UQlESVL6pL
mKP6b8g89q2IZXamLUaZ1EW4dvo9CANM9cVNE0qo8n6PCS5lqRSxcjM0cWEBdGEKZo1toxU37R1+
GnB64a77liDuMA9OZgvsN4v0+fc+HsoSiK3bIq7uhCQRl/OGLXgvDbxGz6yu5PGzj4ivoD2rqj2B
eZD38bNHL5zKL/sO7IojfnNVethuMG9AIcDRJMqR4q+o3xNz+hCuQAqIsht+OH78oJ3lsfIHDeo0
uhGOk9AvyRWKtlds1fEHV524lJrsYCqyxpkBvE95nWDCrFU9OsvcRd0fIPqijF9feavJxmWNYqtx
+Md9LrYt7Q3UD3tW9Feab4LAUvQu/gbk7dkpbHHJiqBo3MRx47jDC1SR3prkd3HY7Tcztnyxtk7e
vQR3nyIYV1T8MrPKMGwN8KgZE4QMeMngMvhxJkzrPwXro3yw476o8arLxk/TeH0e2yCI14DgpPM3
eC98VbgYEc3KhnyUT5KpWDUdDZ5m0lrRzfaqfktI/yyxojWLygg6aw+KXad/p8CX1mQusSis7dhW
lKVHSkTUhiVA96o4IpiLQcX+uKGZIV5kKoi+ti44mryHA1qLA3YvMS+hL2uvp+OnA2gs5LyCY3IK
qBEGU3YVvgZzchQwPRxtm3Da8pUSwKFiqF1ez3zFDdGpzqKIelxZ56W7UES/34NoqfZaOpzToLWx
1B6TMBksDhDrfYdgbB0rZfyPw3IybRDII9jkYxo+nMggVy7BAWljyDnO3sHpWoabgPuv8Kd5lJ3Z
/1qdzNvqi0ckv6ucJcnNKDg7qAeyeR+aCYwb/dPIr+N1h687BkFq/IhiQ2AiEpHontinLOpx/Tvc
Pfva0FFiLdtMdsHNorGdMV769VzHKQq6wCen5yanmPTBuNSGclCNs44rl4f5pXTDlMta0Nd3+ssI
15hVyGjGCE22r0kXCG+N/zuJuFKDrExENwP2yCGTeBAiqfBLUTojQpTBGH3j1P8s9Fhmh0hUtAyn
7LmtxYV6wRHy8nqlxg+1hpLuYxTaN1orULAXb2gJKV5iHXkdZhCG2ylizV6L7IEH+3j9CAE383rs
Lj74BXXeiYdih/IPlm0ZoIEJUVB4txeFvXwg+QHaVFHbaNryNmRFVmtLih9ZTSm9aQ+R9+UctXJF
LhLADtjUvPuOzdX6gCrHcdoE1lGCzQLJ6FZ68ycc2mtgyQA2jDDtxdpwCRmdT/zcIPKr0ANBZ4/E
ZjdyTv3Myn1APz1cBVeJbEXxMV4UaKWJFesK9f8MNqeXVSIGfnkxTth2AMbKhPNrSOoQ5hD5rg1H
d4TvfdeLY8Ockhl9H8qgHHY42RKJ3E+QM95dbEc6QqrunbP+aTW+ubh+zM+vR08/V9eaDe63JaXx
IaP9MzadrjVnoK+zY/NZHWBKTJVziJtVPJYP3D/shXiNr1ZOZJDh3llfjMd+IP7wPR9O4XH0JSc+
NtJPQhpgSB6veRAmfh8cpTqJdGbMFif0DuYZJiMEr5u+wXN9DCpWPGmWBql/TnwBAzD47YrvCdiV
iP/BgFR7mNtTgCI5PHsZhhv3kihNcFtzXpc8lrpmNIT5TH8+qQ73RndxokSYNwmYQBZZAUEGZCwY
81WncRwlILUxPYR9t+yMVmK5kmYFSO7eKRvV3nVJH59zUVAg1TIeft+cDTEJ+GAGKL5ZiRndS9V2
VZS7E6nlKW0k2OqouBsCKLRPJcLms0RHjsfEHVd/V59+Bicppav+HcmKbnEIWxQX7YkTImMuQi1r
hJ4wkM/6gKhF8J5pacIiVOncThSNFK27+LD7Z7fdKiwdi+pjKOhTScGakPCFRTvlN7ekbSKcu4Ox
lvowfpVHrQlJ4S32q5ZsVxDGd20+gUAiZhYgBNexTPP5cZ2DawXPkl5SdTo+Pf+tHDhaeHsJU0vc
osbOVaog5nTwYow3s6hnMp1Qsx86DVB+9Jj+iLdNlQatuGN7ZtS7xfewoQdDX8bERjZCSyEZ3wWO
q+63odh7Rz27NB/0bMurkl152B4TJCdEG7YV6lDy6G0rMC6UJBYsDIId9sghCNiY5582XY6jyn3f
1Wjf3ll1nByQB3UvK/YS5x1KHTM1goF5uOwEeeauBXaj7qoHzHuj/uEA0FeZege8yOeSWaWWGNvE
5st6xnlxiB36OnVmYj5vi9dI0v9UfDbVJVSt3TdFOyU/atm5S2GxMtlRHMlF7FJaISp2RJEMbfox
F6V+fJDVBAaJpLs/fK7rAERSw9wH4nZHO4xVR8fxdJ1xaivcHQkMR55aeacZ0LKQ2CUwpAiRvvym
UFEjWTga4BoLH3NKdudySbPVydaQqQusGMxLPSkb9zNhKjUhcoJe4igMk0bOsxb9U1lbYPtJ3QCr
VWmWd7KxW8MKj4SasEXUtTxVZQH/TZmEyCwshAuyN/ovaPPxk0cWNRBxyDluQhRVZeE48lrnBeft
udmkH4FUrm2hnERN/KbVXOXF6Xdc3lKRsElDjSA/caqSspugjpjZ7f9IVLXnJFHRHPgopYvGQtpE
TMmCAiNDs0pFii9/8zFoJxSTV3bESwd8Z6IHOPJQ8cOvMwYmiIgBwZcNKWtHwUvAMJ0u+cgV5i0K
q8eejPl7wA3DHHO+nmmZoL+Alll4XgOAsrI5t8QwFK6j740i+ZloMaKFnOMr62+phirfxNODj0Ri
35NqhmQJHkNNBEKNPkPiJUIltPbzYBZ7rEYDMwJJPRaVyGC4QR6evOf9BKxWYn8moahz/g4sL+PO
aJFBXlJjIAUft2QmbnGqEXi2pdHaryfN+Pf2EpL71CFfeFzqVzPa5/aPlV22Om25vFknLEGSFNke
Ta6C44ACzdDu+aLyawVFvGtWUq10Oa9u05e12XJ4rMNPvRJDQHvhLUOx0qZx8cCVOtDyaAwAXNn8
KdxsUf62HPHqKKau1tiNAkYte5H1s3Wc6zuo9G2peR3+4/8M6niiC6ORbneRqzmnVnYfCCwx+JqL
gLgSdAqTVEXjkQaM/3hHX0XdCdsOzK3IX+W5oK1zUxgcbDk8ji1Sgd55vw59dtIq6gZgkBKt2rwo
hpJhojR25tsLEjR/aIGFTcNvSlhzAEL5C7yjf2KFjycUudBFtom/RefCSmViaPPZzUCGDW0Jvu3y
/mGJ/RVmSCz+gV/qpL6COC+uXuUgpYJb5lFdXsvTgI8fW23JhX3jbEahtgFFytlqEwnAdN4CFQUE
Zi/b+4G5yB/R+t2QbhHligQ5GQjWTPx4FT/u6F9maS7ceR+IPzInlyQkRdCHaNiuWZ4zwSSDIXxu
rUV1n8afrofhC5RLUBX+G31iEoJrMofXAzpJOh4vTJKchB+r/pai1McZ2oAycG+tOOjnWsIGhCRR
OkxZFwYjKW8jtKdtfJHTIrzEbrZH1HUVvrBzDtwIh9491N92BEQW5WXc06AkAAK9kQWO+1QmXIJm
5wfab5YRt5qetIfWF92v4Q+RHMJxvIqkZTdZQoJ63H5rLJvAgEQPFXF6PpRmi4nFHhL0V3Fz+8J+
C3mOBYmpKfMrtXhoTJdsC2PCMuWYyoEWpsoB3DoJSe235sZgIkb+ETTWnrPq0nbgRHxSPoIGqzuw
hv2CU1989rFTQBoM4+FjvYHzhY3FFhini97Fsry0zV9a6DP6O6iFse6oHyYn+aoky9nfraRWV3uh
v4EFhZlJfHpLXpEXLjIlZshiUwZRUc7190Qu9lC+Exi18Vx1dgmUzFBleO5yAlRWoYxDY0JShg4+
oDfvr/icIBHdIIcp2Rir6SLD7yW2MSiDJplHrBdqCSUkyi2GitsCszfYa9knw49+Ly512G0x6IjR
QKausP6UYHQAJ5Ol91lM69hoy6mgeSBGN230s3DKu0jMGhkaH47/eyY90mmdmzCYb3oHRbGFAczy
ZDOBG38eYJLAuRM+LhMah1dEcge8U81UApJzrfe9CK343qiqvoQyK6eUyYEwZ9usMBMwajeKIv4q
VelZWCMW3UvjzHaHv7haYqQox8gmJw+1OqG73p70f3lwtEQq9hwyA5eq3XZfR4G/I/eKUVFFo8nd
+swmaDMJdubZPublLN8QehxbAta8/DuyXU7oXVuFGVgS04gSLBAgXeV8OE3FG00ApBYeHOano3qe
JI0JjE1/Jfuf6xS5tJiyWKaCr6tJbQoGHlSG7aU8hq6NJdkWF0DTXLlGUHQqm+sV7QAic8tXdwSG
vSVjW7VvBGrR4QRa6A8CQKCgwulrE7PRcmgvKy1y9hfBdimDsseekSCnIPtiI30HdPL6y/lasjPk
pC/CKhyEaYZmeAZJ5nzdTxJkPFQjO8HlztUSvGhH9t9a7i8q4xNtqQEIWzZBCIJ8i/50+gQCClmU
Vo/lXXpcIz2q6rICrzuv6MMJvdxT5IRcKv9yp9Rvf5Orbxpclap52OM72PuZSCGaG8wD7g93dgVM
Amciy9WVOZnTBdydEj0JqmibJGKogQaIoelmx/1kiQxYHOs3PeWUEZalWh/Xa8qVz3t0mZF0pP0q
jRHjdhaJ9uNVuNbBI5VYFxdc110cnhhZ37hxu3BOYfF4ixOtE261pkobl1BfsoZ51/CqB47LQxVx
qGy3dJ3v6JkcNRNomqzfVQpXAJ6FpYfw+VD/DDuMp62KF/m579kaySSYdZakdyNm43Bnxy4tqLE1
CHrsFQypttr4/fnb6MwwN15XZnvH2KxOitpYfSHjEMKQDbxiKHX6TvgkSFOKQMsrzcZElHuSv1Uk
EDswbmAqXjHVIHkCa1mwmx+qvBJdljSoVyqB5a2t3GDApxg7FapTXGL6OJ0/W5ppPbfwW0FM9yWI
t+Lni0IbqDp2G7D4ir+Q6wIRjZlArHAiQLjm6pebwzo+KDaospzZpDwcCDrazlkiW9KVD+i1dwiX
layvcwGHetvm24WBB0e+eZy0yhu6nc04PfYnNsHSlMya4vGAiBfAaPU0UlnJq43BafpC1m/N0yqc
5dSHkFqFxuXlMZdQzJdGL5ufJPufqWFRobp3pK+4rT7ArJqVk/OUsFTNn3LRP6ClO+cBJZrGRIGi
rwDCQj9CxNhTO2XwPCHC2veUjlUid27YVj6c1UdzC61sVqBk0+tsfh2LMUc8+lx7wrZ2lwFI/0Sg
q5wGLX6qqUNKeE4GXVAVaiY4MReGSpC11q51VDxlgDUKlz8qjgWd7mrmDboxuX2DZ9PA2mqKuHQN
KzPMSD9lp5M2vHM5jRtoXYzSEMHYd3X4i+ULJ8bwToMzIjgQkYqUlHp28LaObM/enK/5vt5IdC9g
qFxfW0rELjjuR5+KUv3glWgrnfkO3H78D2Ft8dSwgoJp/M/OflQO8+VSKJHEM3xndUUwEvw/UFqw
FnGYVEmit6I/gbCjDXBw4x6oswvgjgyqws2ic3/naRPpef56JsG46vzfH+V5VWDvz2f4TGz9venO
p1tHaQAHOpqQ/N8HECo3CwS5MIpG84xI9V8NMuAmwUSMoMdlf+0KAU+OreIbDeWwsaJkz62fnCtT
9VeJeRe5/oSGeVWKiHD4zOYJwolEbA7zSgofvuLZP7C5WdZ9D/OxwNFcFAVPg3k4aG6e06TEHMRy
HHjq2cNNdf9HSu7+L4yJ+hpGPCvUiKw0gI+tiO+Br65/iSEoGP1CaIHHuFGVnls+gAw/Ei7IPgHq
LlGxH2PF/e/tTixw85AKrF/XwSXBIksH4nkyefDzRO9dViEjqTbKQSdOv+o+zeL/XIML91PTQmuX
QlPXWQYC9gv66ky8ytu0jI1MsM23TESc3d/5fbJts8IH3gmZZUN2Ds4i7dItTY/uFyZGFCHNa08Q
CyPs9G2E+6tIYBpVUdlSyDj3OWXvXJ+VahHuc1ql9DbOqFJV0n1EQMc7lvjYlu8BppRa5TAXJNY2
3pKyDRZ48/i/NyVEr2M97893LWh/20Zg9n+S8/zSLAZerUlr7vonek6KX9IYYMkyZHFsVC2wPGFw
mzhrFdn5/O0boPV/0Y0+QExfgoS5K7czZz7JnIXqtStKDgZGcADKDEehLF1eo1MOxOMy0G/l3qsM
mp4P+VR07oWKZwUeBXRDX50L4UqMwDjTFJfeAkX0GGfXVX0JVElENhBtTM1tgtmd+RurY4yrpRaB
FxUtp4GNK4pF8InQj0O3aiBjJeswdUY27aXV9EBeuDJ6/5Y/mGK26u7mOb4QozxTeKTPFmH4vFrE
+hUBp1IwGWwdY4AngPWWHjWMgGy+u5snNcBxy9hpK79U9PfAGmTOlAv5Is+5OYr+h+0wdIBFS3+7
eUD6auO+Wy+vCZ79j+SlCR6opmMzIGNHt0sr8jAB+o4sWrOBn5KWFA9uei1mJZSzYURF6z8zSK/q
YHBERuzxExhV31nYCM2XB/oB3c7HdpkUz+Pb+ZnkzmBzYhJPacjMxbQ9lBhQZ6oXWU4iNyT6IAoJ
t1Hco854a655towkUR2ozwN2eH1CdFKSWahhQGqQnClAHMu/hpIXsrO3L5p3YFab3F+p8/Sl8937
EkAU706gtLtioq/tJ/kiF7uosAlwYf/WKTy1eVyeZ0dWct9aH4iEAFTdPuJe7+jJjNhh55v620Cj
p8f1tWR84m4dRXT867XfeXwnEVbsRW/GcGiIQSjBw1Zb6KhAULh5b6r64PQYo2A1QqEdUKXCeFqa
G8bYD7wBWBb6HZNtETGZzvjqc4MOwD0rECrT5MAOxgu1QD3GLwRhvdlyaKQVYsd/2KEGZPGMUdvS
4dmWXF5OCaqqUE7MVao54j1DMQ2YrHGFwC/tX4ikNZz94UCGPLum1g3A58EjlJ+zPQrveJQAw+3C
XzfhTtJFPW6SGd4e22i0zRocw2QqkdJ5FXl03ZbrhhEQfzAelEGoEq1q3TND51EX6JhAYzBAt08C
regY6A958HJ6zhtM6z3j+/d4qyLe0RTQv+wjrNrl+YQjImhH8iNNVz+ZrQ1BrXD2h+rvqDaEJrSK
6cmkyzHWh8tov+hfkDYR242ROcyVieBfBfqJmMQSB5qIZ5ZrfEpqnZdhQjdEOnjahTaot7EXOqxI
P3MHee6WAIEwsySsw2XJyjjN+17i/Q+n6LgIHVxiAOn5VW+7YNwGy/LiR0ApVSwC25suBh3W/ijw
VyL52Yl50xL94nxEL4v/92iMBbFVox6aBKgXhGd0fsN/WVpZcOoyi9Oxnfo6mSOVZiL5wvrLCGJu
Pw3+Kmxlrl/2T0U2D9VYaBmlZky5ejS9hFaZBCC+JRJr2jDVjDGK9GfgfATnooSuCCyXiPR28eY4
dJZ93KNdp5jfOlDCJYeovSkHVGxnMbDLhQ//BVlAdJCR3Ey3pby/NpQ1hVGlSveiEqkOHTEwUUfm
Yasqr13cFRGRKF9n7ekoz0a5hi8bwAfcPJCk36Wt5YLG3Do7yk+LvLIDK7mtqPhZaCZk77phuAwA
uCcjXSpeYSJfFa/20o1aX8Ks/zHHeveRr/2BYX61z+Emi3Wtqz56JYFam7XEV+8GrwuSNxIyV/tv
xyEm8A0ZNeBX4Qzq5ftZe2++w13H5pYsPPOHGJjXIxSs9r4qVo4WK5cNwNNdmRD25g5YADG1ZVNn
MQoWY561Kh1kO0WQiXUUSko5fs5PhDajWOJ/Ju70voVr3QZl0T2ODYEnQYa/czK80DMj6ybJFOj6
TrNM5iWhOhaqHg2IpeCGtFxq+0ad9K7m3H6Z88OYZclQjQV7ApSWby48mdCBE2AQiZnsMpKAW9SV
f4SrmSkK9QiZHfu7d/UBLJn8Z9DbN9YJTb0pCCrQdQ4P1K1NJWHSd0oIaCozDOzVknAq/WCnVZ4B
5XlZ+Nl8rchUjC8dlPcw0mgS0RZ+RkofBi/pJ2CB8Cq5OgHNb+ZV4wx9DGf2syv7O6ODYeYY8cta
zoDlQmBg6Ucrrpe6FaRwtSaJ3+8P8lVtlLLnNqi0c+qtDwjQjw7Zw9Dj6vrLUImZ2DPU9aw++3tw
0j7JmdvZAxhTHfhQcnFjVCFyN50x+7Qm54rOG6+fe0saKGuFNPdphNy0vDEvIY1OK+iCaUB944EE
D/SYUWXEgTtYdpWKFAkbpp9IQOipqdnP0lJOxIyZgSUKXR4aLEL38lJ5EyaVHnTfWE4Rpf5YvD+b
f18gKb8HjwIzTJrAa1f4b0m4Z1Xmk7Y3aGvHzalkdjpataYEOmboKsAfhZK5W5grSo3EXEwSbm6A
XenLlg2tTEfgRReES2CKnHdIWOdlij8TuVUJHQMmv8sT6QdPUixU7ug4eljf3c9PHQcrKqt0990D
koiu9zNv7z/j2LxCEgHs1FFBN9XwfZvJ9VjVhpHR1OeKgSPt8pS3vqQMQs3VB4BomMsfUIi8bUi0
UY+CdkApFnkCyG4HLWQMK0YwCkrh38qMyZNSKODjso6CvoOWoyvMmw/DChF18FsLJXv+A13JKHyD
SoSejichEIYbFiOkJxDBVefkwtqqr/WWVXZdrkaBFVgqMlXbv0c++FM9TwbEFfhBNuWkMKCJPLn4
YwjBnavi9NehnUXNY8zM5ClyjRMtciSm7XDSMSYexgK9RLb9PDqTCz8nvKWd2vgy1F1Dm+nz0tZY
B3rwwRMD/ZRv4HK91Fg7wGV0uOd9vIfI0vKcVJTTi8zQWyVbuk8i6evDCDG0wwaSu4V+okCoc0x6
1AlF0BE5S9taXQDhisxw65cEBSAzgOfml62ZeV+s/OXXtI3ZUSI1kpgRGfX4r9OPzSiFAHLGxDAG
Af/37iSR9zzDQS8MlUGR68Ba4sUgiJnPufHQk+0DqI7emhXxEfy3eMIevI9Fop4OSkeMEiC9O+nj
0U3YXV2fCWGKMkVN2xFxXLzlRcwBJA5jbD+f3d/XpzuThULSa9WuZGxoMoJUgyag8oCLW4LVQi5y
unokPWq/LR3niW1JHW4kR+2IcmwKj4UmWoAbyhxt87XDwmN34Zmx3Ylna6/BdqrV3nyGxClN7VK5
pe7wUe3p21s04Rww/6TuBw7y4eY5UNsbxKnvXabKXOlANx9OIThjkcCN8ZZEDxkk6AL0lC6Kfvo2
th3w/3izhsGsJJHtXAryBPG/I8j/MjJeMdewGPkZ3GR9pdEJ0CJft4g0IRVdPf5KQv4mKLr+qO0f
yiy5QHhWamHEr52Zgc5uoKHNh8JQBNXgDlwvIiISysVnTBjqlrfzlQGrV3Se0wQ61L7Mp107CDGP
WrAJihzAB2OJLqweYqApbsrBdm51J0vZq/gBlXawZUEe6vZCfbK78Y2QukzKQaAWrcKEYd753VS/
ovgFYPVPwMRSYA7fDnrsmpkV+YoHYleOzI3CWQqPge6DoPnDhKixW4Hb49739sISOvCHZ9amcytm
dk7qEFNdrip59DvXnpKaVA+IWHmAEar/6tjITNnOVSwGNc+1pXWp9jHd3n+ay3AgOkiXv6+t82bq
cIDFD7rJLMMtRWnXO9PI0wx6z5rOq8lIFF1SXjLgYIlHgleqfLwvS7bm5OcG8eNcu0AzHiwPJ4o1
ULwSDlLNfkejl2CEE1XLg/IJjG9gKGnInKR/a3Re4GsbEHnBqhpCUmxI2LnNY3FjvQqjfZJ5Yj8S
ZjCnEaAexpMmj+1V0bpmR5pcq39W8MWxM4W8zZiW1k+n1VQzMns0XjwDjWIERttcutVGk8UZ1k+d
OpXhGWZJxVdm4asz4mH1f85gIGHaIOOsN4/UMHO4PqZWpDZoKx3L+tni+HhRUAeT/QUBk345ethv
DAMFX6NEFdRWMPRaht7jfQgOM5Balr3MSPukw3RBVIL8KEZx7jovpfFIyWrzroWU3LniTj0QMMXN
jHcaWdCPjDqBo5//EuOD7N21iWqejt3VHSabTO3TDxyzCZKyFb8w5DpQ42aw5LkbW4cEaDKhBl3h
pNMbcnLP5sXaT6LwF8aEJNZAmH0FrdQjdvFPJFjKfcVEbBCT8P61CuYlUPWPXho9hbRMsoMi7ZlQ
CpNe/ChNs/G4kdhk9ckoLsYi2e70bwZvoBB8N8WL+1mRQf5amV+oeVVPW3nCcobxJdAuZDvgvMr0
lFoDJm81PvTI5k7RJUYom6GNZRugaORlLZYDT97lif1yWmlub/3PeFxRmmSZn2nlpTOD2b+GmLzQ
smYPsVi3Q/X1S9WQS8A8btA5kVID6LHVubAUt/dPu1+CHgPU5cdPkdDM3KlEQQrm8nHPYBC9Ca34
HIc/di7ia6bERcgEtbHB2YtvRU4JTPVXloh/YtGWLaaL3ZuvPuPBFKfLKydVC5wpdq02FD8lwa2t
awNqc4RbAzgAxyKEH9J2bZaq79eTCRBQVqytQwV4G6AnqE0T1PiQiggJ8craKlJx2u9M8SSGTx4y
8Hf9bBEXfg1Kw8qdG01HP15j9uS0Tq230IuOBsUQ1RhrkRPNo67ri+vXaUpYzlvot68sN33MsGzM
ovNhI8o8Oh8emadQkktp7VAV3hCd5zLMqaaAIzNlIYrH5kdj8+IICA3eXEtvGmTYU0DYfOC7WNBN
+k5qm1FleNdZ3kRm0mKIAdAgRuXWwLcNyyeFZJ77bdWiaiyBKaArUJ8nTUJJYbZWV4jLGTeCy87F
1MuBP46NgBV8qd1eICOMZ2mS/GtpfUU3nQhYvAu+/emXtAsRpTxGiZOi4powPfFN4mLSBtVA2fTP
s/ytrXrbVKOk32tikFxx5kNztXGMXGjGErCSRup3DyEbSBPZtpUeryUvS0DmsFH5dobPBUKelzHZ
wmtjEB9uAbV/Xt1A11+IzJYlhIebh6EyOGqzjQfe8xp6V+IpxjbiY9akW28Vw95xy6iQHL7Gm7yF
HU0pUq/noKcgGwMQaoKRHuTpEoHT81TivCkz/KUohXVHchAUbQsnc9SrwhmJDDkoLM6oIKMZtcHY
Gbcbc7ill9UXKlSWA4XWMXcm4MsyFOlVK0xdXfoieeRxIXUxZLk4RU77LlRLqt+4v+ovcMeFoRFf
FD1oBg95Sm93dO9ku155xQrL25hzY3Xl/pFUNGMXbJ7OX0fkiFuDTTDnE69FgkgEo6/vS3vCZ5yX
c96cjg1HGXeltg8Jfqpg5aupw+owpcoa4m/SGyIgF4LqGiQJul0hLP4Xs/pdw3cIcZ3e2D/qwwTH
HmVozMpCyeqXIf3UcrGyTc/zuDDwfy0urOyMelnZHGoZkJBNKifeY+COWjqtjjVjy7NbcAsmEg/9
H3o3qh7sgQyhMaxneE3SI0v9Ter4UfZLtKLTxvgVReSRzZfMQGjG1GW09BD9PdbAgdrmDuavD5Ho
X8QE8mro/UDZtckxY6FjGRb68iY8fvdpA3yR11GB0cICLGMq7XPxYsd5GzZEIz23IyadDXuaotcQ
3eTR0GweCSbD04/bVZ8lHa5iSj65If6YsDBJHtlxPXwB+csXQ4drTDJ6CQORWHby4t7Lbrdm62x7
+e25rCOkaczkd7OxBxGjI8DZrNpbuCKvULgQz9HeK0h4F8tFf9YNC4sN59i3nHEmuLkTRsADgzlV
EYMqeup+uJCI+GdLkOb9iDA5sJDoCOJyFr/uKyNWNm4jWtXLJIlOZVrEXw3yn7Z+AepAwwpFqlPO
2LVvninAuz5xutWaFkSf+IX1dv5//hQ4/G3pPYUT3lbvIAKoDXDrbescRYDtYjcdWbHyDOPVTIbc
ERBQk65XWiOsBtgsIz2S/SrNvU44ceQLY+kav8L0qY+dMv4kTAtq9L1HS8wL9Bs3S1quSualTSVa
R+FIQP6T+6SAKoPc0zmZQOcbNawj0paUAZEh+IMj1aduHYP6agLlxSO6gLlCSkuyGrPCIWjdhunJ
sYeNIAwN9lBXqSXBjq5Ogy2KcaJ3e0UvXeCJMeOBrbK4YyCdOok5mxaoRHTT2QPNSFVqfMwnt2oA
sTknqN5J+mdnJYvSGVg9aujQHQs/eyKGT/KZfjtTjdqxapBoxZWV7ZBq/nkc+emLz+DJsTwXdh4c
bArcWHOtgUo0m5JU3Kcqp4CM5vhS22WzKEYNH4wWHxBJ8iQbtLTsIuvRcOj7ov2mMI0OiCDdRJ6m
+t2LKJG8WiOa8BYEFGPZzISUBRNTfG9HkYRvAPXbguXmRQBzwFy4eEHDIm+3r9YpGMA9tJA4bmYs
uDWeXRys6D0SDRqd1nZlg6Gz4E8yr8LaOi6jckmScyVFXXknsFNvmcS9UKnTy/e7UCgmW5rtYnYz
KeTK/shBsbePU16pu3JgE/58wvy9lAq3//KT9JqfGJwUVxvU0G4ql0cXgVbThiTzGmFNWTO25Mjn
PG7a9s8iVbZpoIQ6HBGsxKft1apM8NdP7D76JK+kr4x3cerE/xJVTh6aKq79En53rFFqlTEkV83l
I5k3yHQlbWlcflsbpJOclpAiW+s/4nJSge2HZU1m/k9z54+l25z/A8LSzbyck2tW16joMq7xq83E
qorr7ueFFwTssCs8QrKOK1fIcTNnxaZK2ErLphiC7EmSrWSINUx4hsoCPoAbI0lNo5zsN4HyLE6L
yiSFXfFBbQghZqeSa7BBPAKzUrc9TyY76s5zCFQs0zh14T5KK+CXut982cb2EVzZrbUvC44eCSjb
/PcyPJ5ymCGIV/UXQ/v3dZRrsfbim0QN3DeV8uNN8qoxJFwph6kqy4vdnlIpBwaTfo0esxtkynbg
ydo7hqrGiZQMUdE1k1JRL5Fh+4FJ9JbZClY45h+UpZc6dlN4cO1gsOVifjE1NksqtU3p1Gl4EyHY
5wHX6EJSsFu3eNOeF0niHdo+eVs5DoxhHBzp8VZ8i1M2Jxd6Is+WdYq6eO/r34PLF6EitV9QFaMN
79KnwYJ+tvHB0NBUgSTM1kcLHOMwjeObXASnhrvUxDLH8RZ1gz/ECKPE78OIRg4taTSKBKWeZook
Lk64/hmG2TZTq1pgXbfvOX/AuMLUfoDKxzANfQFNJBlrc5xV9NM/RDiUJBu0Myzy4R4MPN9VfH30
hNxM8VI0Z+UNj9ZSG1om8pCUmZLjzIQhnbJPtO6oRaTxyw/hCuUtEv87pLo90gaMnsittELyKLJp
IA6LoNfpqKFdnlhw8RNDJBcQncFySoSXyR0/JGdmkm7hQ8F/EIHlcHSZWsCgSiHkZYYjewym8jQ6
9/sacpvXtFRK17uee9E0GSL6GvYiR44lBPoLjbaZdISeHxMB8JgXpk4HEFt78sjCHB4Pp/BGlh9V
RpZxeb/HXhm9lU7Is7t/1++QglLlrlD+dRHL4W8BeUmXS1tA7V6L6vNMk9f1gWa2uvREKNo85Raw
eNtGFv1owGF9m71PY3ogXvjhyXpH05sXc9U6SIcqOgIYRF+dhU4ZjCpPs4citgOElUxG9qfRwCJA
tRWJTrH2kdTi4pWAHCt3Ngk3iy3yrP6N3SIhPG2iKaa2d7rVv3LuZgJzBCxlHU6/lGNKtAI+/6XU
xE4l4Nq+XO0Ig0h9GR4eYvHRfO0gum8qDxqTG1UqBfygh09CiBvbMVqMI7XCfU/t09WjDKUjsmlr
1vDZkPt0YapV2hHqj5dMBGRZJF2OjiMjOawrjJPDoKC+djWoyhW+QEYceQ9Fa3M9zSgsPdnmSpT3
1BVStpkc7YSAVhpfn/yR9LU8JEa5GZT0LH4uv/AOsLK4xBAmEQHOm6sLG9U7jwBBhGeeb58RnVf/
omVVQUXT1k08XpdD85yS8PfQrT/s0IcUPYjbDybDtXgwYFNkX1utb7zNZVMq+dzdCYWRypDwZFbQ
nU0lMp9Sklw84DcLS/mavT00ociBTGlkpCUMIV7GM0NpR7czkPy9qc16CGoqk8dT7+0ZlWw8Ee8X
AlXRhCKZgw95a+ywPp1o80sMoQdjUyWBBxGIp5fGcYMwCyY5R2lxg0PIczqJoOscQBKIBe7JpuAN
hor37URvQHPo5mb3flZgZzSQGDsgVaKxFjj5qK8Cul9cSeQj5hbevqnITwE8bgyJwXBx6pGUQw55
ZoJBrN9mI5wd+7Ps05WfC2aPvU76shosW1wR15aw+ahNQXv9stAxb1FO1tGQsdVjVn3i108dmfye
js2PLehlXD61d0BKN0nijuKozZMJHE6Bc9U1/sdnamJdope9mpcVnN4rw1tcrw61D7Rht/ce8fAr
wwjkeEwfOmF4xHwM4DBX1532vgfPSZ4xdkD8fomiSvcBHj2CYTNfzMjG3rv2GHRshlrsifQcnt87
2IyddN1pMPKzQ6mxFzGLXmVwExq8LP0v1iJBYM1qWlLVfG1/5ZBRXZjAWqZNaHW02SKs73G6UhIR
rHs4MLUex0HtUv0jxASog8ga3RmvdSseoR13n1uM//T5+KNKgD3TeGoOpeG/4fHFoj4rlhCMNNIy
n3Wu9yTdYt945CAPWAfFQAp++L/CZFvBn0yEKobdMlgZCKKa7kO5V+JNrdcH0qTCkmOcjAW0FHSq
Hd/3274y9LhKqXM7UrNKYKRUdb36RbGK2JTEEqhiHGU1Z2KyExy3iE8ipXtZ3XepzR7SMNQo7b/N
96O0+t/dnpgg3LJNnh98i1iACjYZQchAGkTX5x9nl3qklRlm0MLEJNK0ywnYIa+9Y8oSGLugBrdx
+uDaysr6yD3p/a6YLvZbKbgULo2pEzd5gIV+8Jzy9X0DJnMMpNcrsLUyZRKo8NmRvpeONyExGct8
aaAQPGIhpnxJpuoUyxGKP/rAWQkGUe9UbO33D1uhuT4bEp3PiDetQZUCASPkvqT9GzG9s9U65mMm
XoLd+J0J/D9NUlgsogCQA5zgHBc5NIGP5m5rdyuisdvbjCiAZOkQ0trWjCprwGgM98SzS1d6h+Li
SZ+Ha3FsYrdGESgHAaqxjTw4M+w/+4y8OG9s0/E8z1Dy44FDpi98NfcueD7mF1dUS82yUVmHmnRn
Vyt+xnrZR7VhXAgSiDEJIMZ+Fw+V9Zqw89INgODY/1MQvSCmTMOBBRE7SUdGPJGlUZYy1Cvs7RAb
18rt8qhvN17KWTsoZqjFzQ4H9lurwhstUkT1eIlgGpeFpOrSJS6Cn9oiTz1ctJ1IgwNu2jz/8OkV
IDp+A41hXDcs1noNa+sgMGoVGe8NwGVHyXmuXD3u1DZXZx9EWXUZoY7q7sMTF03syF8qgdc/83lW
7I1AdHI3um/kK4RItVWGiDB8gEuYkVm29iAN+k/gx8R4/CnQjpl5TdcBLmIU8h+FWxReteKhZCk9
zz25ev42lR0pCHcx3rFunt/DO33FjIZucnaKgPs5a1Q2pu6LLFFRjurH0rkYM05s70k7WTsYCsKq
oOlyM2soJXr7G0VYcWn6R1wuLjzK9fgLNYSBzTZTLVXfKpx/YUl7uOjYnchB/Zssu3pO1UOgoGqj
v5TTPFflI7g1C9GFz2ScwHn7L3nbv3pDd0o7TVrbkjgmSM66BZ44KEemNCzeF04nTd/QxBmulODW
3ruMx/XenAo0zb5ZopVXnx4yt2dG1mONwkyeb641TiB8mAPzEW+OBZEtX7ZTFT5mx1YFnDz3kRLD
gLQSBydXKEWuJ7kfr9KCxkUih2P670Aw3D3hxmPSoh+aHhzpkHRGaCtuGWcZPyHABonXTBGtBGo8
m2wCcygPkLEmAB8WYYp5aWPZZA/kpyklToX76nFQc+n1clSE/eS65ZZlSFspn2JTuRogG8AviJ7U
xo6YqaDf5ZDkMGia9wSsew1uDnUKNqwF2oTfmLrXkKzq9icXUWZgZb5d2zU32PatopVBwbaTCKWg
C0orxJF8fUkkp7aJCz8D/DtzIGkk/FiONLDvRmrnwNC9+81KTqbQzNK13/yixjvBRpC574uGYNRx
qbNHggrlBnSPwO+QpOR8ODMbsUErWEKXNXSv6XISjYBiWkHkUcJAUfgAjiRkmMS/MZyZbL2C087S
owkA4DDWDMW/8DHU5vXH2bRUutOg0pAXGyHjFnjypP82ntkNBIZft8aBXlX/aQDk5FVoVByfvjXB
GJn0QtJDA6RI147oY9v2WyXTrZN8ym34MBzEEIfUXkJ+QqpGJdmsgF4jEzQl0GDIVQyHdDaSOKxI
jLDXgcXb0ui+l8lCqAQOTAXlch7nULMPjeFr8Uha1oz+QXxZVhtDlZQGYeMgcUbUQCsRHDmTlVTk
lW9wfNYBwNT3PyZ7grVRL/IN0RbIO1Jes3qLOp9WBaYw6jcgjKN/LvHz/VetYQekp1dc4fP+P1GT
fYFL9jjYNVeK17ouxHL61agR9rTdtU64q6alqMbjwzYOpjeg8o4dEFGlatdiVxCRM1nrtpDOczl5
cWI7NXKb8RNxhQLOSjpR7uslMO+1HOh7CywBWbGiSvN3p/pulF+LvPqL3VGd58FW8gDEKrA0Ejqw
Vp5wWQgQpLfSteEE/ZuPV5rxRwXj0FR3XL8pQCuKgQoD1LywRywSdK0tlxdnU3lkQvX1sOawPdBz
aDW3sBqQHQ+HoImxSTsR9ESnNPF2XWP7YtsbouFG+Po0Z/tXcfZYCU5hfzviO1nHnRfxB1VQthHC
r8V6vxZO/7SUszFkXrIngAe5d3u5RQi7EPOusAGnwwxlb1EqdvyvOEBps8s5r4pPjwpq5wpjCpam
3j59/80YzltXowy1qSeetImPxKdwNyOrD1T3h5jyapzGz4AE2y6PXmdX3ajEsIE+sydZWNU8di8x
nNTdkwn5WPmt6CUbaS6/H+v9yH3C2Me2DUsw9yaMt4fZxAB4hDS4Nd8keWhI8MzM4M0fe8AyLxGJ
YNbo1+qTshHJVu+5P0J+SuA96v4ckydrCruqNtQwj0kU2+NkXlMZF1tH5Iblnz3VPnBBxL7F/t+S
Ton6/dqGePfrqrCghb+ML9fWhpcBLjKZongoYc6fPbElFfDHzSGaljYoX9XiYgc9/hrBg9hX1zKT
HcypVRb/ZAzOomg72SkDMe8SgM/tcMKxanTBGJwHvrNgGOvncfHRb5mnzgdmDzhhpNEiBHJ9t4kT
iYkB1TSm4Ip+9XDPOSvldK/hGZrJ21zuphMmuD+V8eliPd4+RHFHqHYcZ13PFYYzM3eqsCqhbpfy
63UwykjEo/fOYVhMP4a6uN8ItiUj6PjpL62c32FQrDWYygjNyWJRY4o+3f7RtQ4X2ilVuqSnEdBh
ufm1wjPqLLwnE0+rEey/d1GlE9wMq5lcdyRmIxENEK8cU7AEXoFjwVbL2EmAz7V8wOq8ET1ZrX3q
fFb54veX7FEadvaVa9w4qf6YkVhBNTJQ942dTkVQVkM3cMk3D1BMK8Jy8h2LgialeaY/rVMQv0B/
LChDZ1PByo6GQQN5V0Mv28MsUQNPzfxtSiXC+w0SpXgPKXHMbAYF/y9l2ffJMCtTWsNMlSZbDJnH
JCLd+dy0JnzKZV3VtZl/qYeuDfEkbjmRC+p/xWDEfUuXoUW1Xp3GsoSpPZ6NUyRi/AL6rlJoV76v
0ek3UimSFqNBC30zMnwgDfSVuAZsXqzoQRoUBP39PDSv62U2eqkBTqsaUopf1hX2tz328UcITuJ8
x1eUMRZSTf86hZbItpkUSPjbsVOR0kxbbZRWItGToOVgm6torSAzMSm+sSjw3qQ/psvpojY/qC28
Tk3WdFinmO68wBRa36HduI+Pxg0IiYJlgttzEUCvb247L5R29lbI2ZPbHGyCqkQcCi3IvSaOQ2gy
aQSfIWxKxfikHDT8P/Uv0vRBop/npQXu0NYrPQ8EeFuQ9Nbg/0RM2Kq/qK4MrnpxvUZVhtvYxdU0
gJBa7d8tPWY5Qia1v5Xs2AP4Io1M5Hs+4Uz/os9rEeDQMEUTQtn+dQd3FaFXWXJwBbyjQrIS9Q+M
Hl4W+MxoG4mL+tJmCX/N6JnwpekKiaJwyH3bOXO9nHXW8upS1kPVolK0qDTTuUt9om1EB0J32rfK
/Sgjnxv7MqHQg2DEfugd7zu8wRbMe2GhyzLlKFLiEWPHVlqtjNmwLZWFpLfvmie0LqT3oVyB6g3N
+uC/6vAqqK3hgqdA6dj2LE36xSrVScXaMhc/y+144nEJBiPyD4FrHZsbPnoEOPBJ/TJlKKmM+LBk
vxwpJMoMLu/b2if0mCEQ6lfgZVHoo69VfqsATf5Wl1ttZaDxrMTQX3XD/cuS69ZlweL6LZUofjHG
ZNqbn8vg2yvhgjXcj1iiQjMKKwR/1F6YVsmA5Gg2NMGpIkcngzjg9LEzYhmYZX1fe72r95JAxjB+
44YML6369GOW7givrfsR+LhRYrQZWYON0qQkgSd7DiQav2oQAjag/1qa1DirbbenCnu+FGU+01E5
wZhi+cCBDzO/oQSPILiLzEFaHnAJUONCevlTQnJImWxxeiZONpxqnw2h2oeL/etprGLMw00mu+b+
hPnU/TtTV+xybFCEd/MCZLNxWH9Do7BPqltgba/T3TP7Rfhsgh47QqSm4IILefrcmZnyAtJztvI+
hoZ8oZpPL7b7ndODHB2ldFxFwD4YYd9gEZEjP0lRewkU4Gl5Y/uBB1QWnmWqNfi/CamXEUHg/6ZX
fbGrWq2aUJ2DYmrPh1/8E4i3UdfRnLb26Ks3StNoJ3pE+ZZRgyihHalthdyvYGV0t3nyiQIUTQBh
Pv5KaGAMAkOi5q+sDrtMPrsSyKfMQ0/qEMllAyg7l/JOx2HXgR5hlNYfTHD6UcuqRAWuJat9Ossc
RGhfG9srhumyapDl/Xo4MQGUU4IOufPd9eHZ7I77H6wQphpXkFrn8MTx9qe8gvHQdNDbrBPA8c3I
SYD2DIz7pIfES+Rt7H9SIBRk+iMI+YlnmYbml/Z/HOoMahLA4p4/+R5h3Yvc+bx5dKzbLQfgHTrW
Rhxl1s2mResXrYa19wuQS/pwkB7mf7NNUqv2Vey1H3coqyp406F1CVppKQJkjjwW84x1srwGixjr
/pdbVyKeS/LMaZ7jf2NWA6sYKx/QlnYKrlsDbkdFECXZe/WZe8VNMI6wK6Dhta5MEccFlLg2vQjo
8W04Jxka9g1AJbefPYdRmlMClmKE6Wd9D6//A3OrBxKWD4WeFnYMI1ZAZlQGrGpMCKn9XRkh6yW6
TRKE00XPFr2bAhZtwuf1KDeHjBWiStIuZuCONhlwQelyqLwUVxINm+09cIT8gd3UCXOSKrn+KJby
ogFa+jskIIzHqngBbJhNwwPIuIOwDFQlHH43z9AAepi4QKWsJtJDm+Eh7fKIKrl48DGLj7aIIdIO
T+HrFAwsAcby7cutrej1zwbiO9UPw/8eSP53Vwx9T/5hwX+fIkOmmN5Bz3Q90nM7g8kyQ5PpTwuD
AfTQIwo3KONiuT3du2rhBoxC0EUsWM3gnCJN5ROuBs0w17x5CE1guny8g6JG+Azr9gQ2aJF5rPqU
FrV8WUKctbPA9OphmSr1kdIaIurP7FZRTrcItmlMGClZXNF3R8eef795pdj2hxsFvDwzlDUbpBhI
oTEzY3TwQ9ocEONowlRPlim3FrmQmQNZdW49ZhlFB99MVnZgRK14eKcJyDhNo6t4+evDPRqDuW0A
nbJeo37QyWeR3yLpATo0E5C8wJyqKqz+8BYqJt7KkDb10NFx4m/OWU96D65iGBHlzD9JqtzgWlJq
QMcqxLQeHskZs05bhsAGyDSBjY5OBkPlpmJ9J4qNZ6uF6F9ujY/pt6X4eaMGH5CC8hf13nVwa2hD
IUdFOgfMWilcXv0hfw6vvX5DQ6Qdr53HsezrTKhAjydAQCM2BzPH4LjRGWYBtSYqgYLZ34jx5Gxd
1J+gGM3TaIoYntgjt8b9ft8ny/H+RAyjC7bxMA+I+4kSfKIuaBVye6FKbisksZLa+pAGPNfXISjC
8H2e8adxBH60b1+D3vH9oMqpcuwNbpAnpilpSqLjdoHfi9Pmk/NN5XigMjCOrjhpBksYushMd92O
6pNFJtJeZmAkszkEfDfmkmZlp7iSi2nMjdtWZmqTPnJreiFLHSrKZbmIgzJX4K0zQT8uYdrDjGfp
TosE1pB78L5HoEJeAzwX3nJG3jXwzxRIKYElXfSzS4/aE7QtzKApB++UAWweE7s+NtLI++Zjr8Uy
VlI7vw0ysJK9ZXaW+nJfGcJmNYKvY68ciQMMSBpedvp+zIyjaI0KAI8LhqezILQtGLYDviIqGypx
eMsl6WIJKMmR1aH2sPuXRv9rdSiNoU6LieCazDUtaNrM6P0gxJh1NxscgPMh+GkT2gfT4mpAmUHR
SkH+wVE0MMCYdpvRXVfX+82yL4a4gXtHVtOwN1nWyyvJ2OWC1yKbBNxIBsyQAfFR82S+EzTD+jSl
WTUEa7gN8lDyOmMN37UsHaFAYdd2nBPpEmtPI00J3LQApyydJryy+9N212LeKqigdap0awIUHFRY
72qwVPhoKcIEKUxPOIDNrSzaeUukz8xlqB+/8+FQ5W3M0XWWODTA7nN8+AgwB4+nFxK1S0jrQrWk
eBW+ECsiCXAP9YVq4KhrlqcIIJVnMrRtli+RsgO4TOQVQBL3VREV0IP9OShIB1963c2KIEFKEKDY
ZR2/QcRbjaItUvBjDlSM4JYCf5EZssUWgtn4Of+X/D1I7ifxoUz9PM+kOvMH5a0AgJRa4ooLSI5Y
3BepgqxZxcGxhNxSrvBEWFvyc9QnPOrzZsQW1qcFNnwBU4sRG8WsiYJXSFysgG0+CumH2zuBssh8
rZBxTKtf1EfcR5/pAua4uyJz1hL62WfRwy/mqLguaVzKwnSJyehyFLentpIBgnSwZrCsUoFz3/Vk
1tQpFeYFGCcVDkMsgomtdeTEA+9iOr0rDaohuHHyEalV5H0cOfZelDCbDcVfF61uXtfcLHzckTc/
UqaG76yWSB2cg6Pq6gAwroyG8O3j0UzsNUYMZXp0EXJ6Z/U5iU7F7IyuaAemdJLx92zQDfgJUHNg
cWndkL8pPVAZF9f6Xe1G2pt8/Yk7hLqaIb9tdfDuescFIapOeinbCPIvpityQYHiX9WO3qDquuNr
+6tWsmaVDc2glJdg5Qy3aiZz2ty1saAfzFM/c0zyDxoTcHm2AEqyoq0xRWbYKBD60r8YzADiyfoU
3CsS5R3Fq1hiXnZJ/C9nJjNJaAlhFVBJBG7Ooac2p4bfnV+Y4Tujstji+UCO5U8NX92FLn7OQsye
cDho4d6Y5ziTmskEE2+QR3EAPzeKcECSw5VYVkg2euseKeWzIAisCxdUMjtmunqojXPDq0/gOw+C
XUnrJt26q45IEF6nkoeJ0TcWgObiscQO3dW89fkDj4SSpnQmnI2No/W0AbGALq/YE2LVAkYRkLSF
W/8Ab5zz5Cl4fdWroBBpN3FxC3ptZpxZ7LQHEXaar1y4Iwj8S+w02DTNVZ5aBvZTkk2maTYfJnhB
10dmeAUef4Oofsr6HQ9RwkdT3Pp55uoblZm3JBtR6XMfoh0xokhu6xn7IlPE8cl+sfN6rtO/3cim
pcopLj1f404tARyVQOArkzhV02+2tUaB7lFBMJcmFDcppxZl1fUeRn7p+Or8wAaIeBq6s2EHUbJJ
wzj50p+m9gpFyC0EfEQPcIp60ezlnvuSTYQ+zj3BVou7MvuQtBRgs0A5s1f93J2xgJ55fwBQcD2f
eJbUiqfpYUuxdEwqUo8mEUPGVVEEmp5m2wS0EDk0lwUN1Z0xQdnVI1PDNpigfEWzZqF/ukYdTRc+
4lXy85BMzCUXOkqvAQOqJVHmCBeKvHeyYcZG0fNA8WZTWOaatO+FR2nGR7uywIXfHRAEO1K3v6fC
FwQolrCsUnEUJVXJ06hqiuEnymRixBskFaddxMqJcPjR8rtixtTNq3u6nkhqTUJmJv0B97zaaeKK
8henco3v8yLXmlNSwQWFpH4IwgUgnF05PBXhQEShsH/WSl8BylHdhfaMgqhDPOIZ07yv8ABOe3Px
XAMczCwlhRHJvkb9P/N/7418sBz4hoyCFbD/HRdJxE7mKO4qgGJs6Wjt6uQOG4EJKSMAVwykYftU
XQgZ1wOgceZ/1jvUewGWo3G5EcThfxi3CaX1/1lLemTRruxKfEn/ug9tFjkz31349W8sxuh91JTr
yfLclgwhgXdgUgIuqJLjTa/HFXYcXPKnz7UR7Weg3F4nL4NPWqzwQjLr1EWfA7cT2CULTf0z0iT5
Wzoy2mLajZ26Y/ozCxUW9bKpFV5SnrDZx2k2NATN724DXGypb0+tVxR/HzRXFyae+6XQd/FeNvnf
NaJXzKDM98K4XR7KDwvyFw1S3EeVTaPvhHR3QRn+Vjag/Bk2fLvegZQP+foXhLo2FdCajkJMvJ2m
VfXVT0zA5ClRXBZ17Mtu3mLEacSJMNnyqAsmiymQBwlK2kz7bPB0FDDZLcp3b51Mj9SBCAAz6/Sy
3ezaZ1nO31VC59nwhypUF4NfEmxPEwEauquNki+aWsnIfd8mlFdbx8SBdxNWqzQCQp7vVxoTFg+V
FXYoPwQ6TEpmH+tPRuX1ZpUk0OUsOUtbGoWokoufsBsn3X6oN+rdC4q5ksbP7j/Zgj2q9ogTkxlc
oOiqwzBV53Hv2WEO0U2ZkALtugvbY4bpo86xGoxt+3GNXgspGQVIi8FZCzT55LZXd5fF1rQRLvb2
rk9HeHOhJhOSErA8pmfxhqZPonai1ooFxGBfTPfMi6ua7oHkWAtoQbg/NKzwYoi6keHPXuQZHhOE
6mO8fJ+eAI9TInyAfB5xhfpty3xwmUAia1zKT6b4fhvcVSMLZF48QmuSopjjyFyQvekBAcKw15/7
C5MPyrqOiXwPUXuNk8zYn7XHAML7FDsKGeuC/g0TG/y2jggyYsUwpB2R2UqYU+5BrsJ5Kcz8iUNJ
ZAu/QZiYrFrclgXJCJbFtnUu2/GsMvchvyXtlndgjYJeOahfnln7thqiSe1lAd93KEE8+QdKeHza
HR9yntXzhdzWBeEg5SKqCP+BgKz07gf7m1l1xz5QIv97Wh07yv/xJwAQWV5W/S25brBeeN+Wy2YC
fcKDR3NMP16XwreNnMBkQ9qj4HEMeCxvS1dQweAbNr+ZbZ/LZsI2TuZJJiOLkiNJ/LP+y/YBYBo6
B2JrXprODQlWt7cwhIifpMeMhGbxowtTueaWAvOZMPQdAi3tey0aAp4375ZVQqu9BuV5qvQLq8vQ
SK/hEDvEDW6c6Z+0EZNx0zLwO+v8/W2R4ZX4NY+HpU4E/yL/4QJz2l8oXFI+4XhZvsyf2hOzrvvx
T96ZHkBN1SzJXxIrAGADzrnq8ztjPRq1zvOTzd1HKxk/gmlwBaRSuST80R90dx6NFln+/d1Kpafh
KNv7n5/qZ/PAaI0tyP/kHXZDON0j2s8/cIR9LOFEhJNfGGQpcLy03G0oBZu7dVNBmBEAA2rY3Xvw
MgZ8mqyltDL6xKWVmiHsCvFxFR1gKcHIKGzfKrRXrNvXe+Fvv1AXJ8F+14N1r/sWgqkJgOvTSOX/
BA+0LOx/QMZAA2j8Oqgfui/So4bM4iCvKJ3irqgh+VI9cKM7sdA9zItIaSrlufvAU/CiwBeIAHkM
8hq6OgZDKcLZJjMaOQnXxBX3GqBkzZ/wtzolYP/ED10GE0s2GlVI9m0FgBr8SzxksKp+xrarCfWV
5PGWbcTAj0wpMdMBjF3FmNEIc/+kcVf/WU6sYypDCeSZ4PEQlNz9GFtxtueYcfur1491h+V9w150
5HN4Sz3c6JZLLeRSkpUu6THAl7aA52dpVnfYlU/Y+m6arquHihByBnmqtEcDeozWl7f+J7N9Yxin
NgWt5RXsdLtmtdeo1t8bVmF6wJRKeXsqE4jy/IO8MasDoM8LGS0qifaS5GGk5qUi5+QtKowzj6fK
lknTCamwV0rmODlcUZ+Ix/cpvvSFuLNMo/UKvIto54+BR6lBQ8zPFDSAyxdLC/hfe80eVMPA9pGl
8V7Z8ojpMwiDyEw5ozClLrdQsDBGrelf6cqT2LGiQwR8tW7rlZrW8bJBkCfNOqnpBLxXcilAA4Ax
019EYTIKzImz2bOasPUgiOWartMmA4S5TD/P8yMbj5SR/W++nnRxdIZ7Fpi8Z2lk0kNBj4t9ZEHD
HuCX99osPfOfm/rrqA8gCl9sAFC0b92wVn99jI9l4yYwdayKe4WL/LrSRx8B+/01b8u/1/3hOKh6
jcYSt3D/dkBndk8aJAK7aBhtbvfLz58F9BEyiW58cV/lLU5zAd9vrX6qWSD2fasFMAy8/SbyxYrh
UADFAIN9NVlZ8PDJ6LOwKbTfyTJkwao/rP+MjhvFYymDm+uVQkC+Ga2jb147D1QY75pIXdA7oQnL
Kcq6IB+q9A8cTdxmS9FC0Fxk8dAFBOFl+OaQH02c2mL/EXoWraHEFlsfpcDXdxTRIBhXL8rKY3I+
s2NIfsbRuifZFHNqPc+3DVWZIkZ7ef85Zji9WUcE7U0gn6fiZmFVd5j+lXGNOpIZXKAHIaYeGcGv
S01nj12fgqwacdJArBItndJ8jOi3msM5OYY/jMbHy6g22aZNGWKW6twQyvMHCf9dXtLVb+DM5UMT
appzWBxX5yBvE12dTKDKVRVaBQnnQEaXJ5NEHHB+dUJbSShazjtj+5at82VS9P088LhbNZxTv9qB
NtbTDNHFuPknag/I37bWHgkI9Thw3SgMd7Rk9VLv2eItrmG9fwe/bbc8Gs6xtq46vVnxLpwEJif+
iWE5waB9JtAwL4QyvEqDorW8zt0EBjYlyC40wANTdQc40T4h2k/YDq6/uFXEBxBb+5JjncpjFmAM
Ssd+wvepIiOr0nB+SH7gMNe6B6U6482xt3+7bpTDXz2fZDAIdvScM9pAN0uqTK5tmQxiqwBmxb2s
xmE44YWiOJ+/nD20ucUm17BkoI+ltDANq/kH/LH9CTpMAHCjmgyS8K3zjHgxa72maZoWSFGobJXU
KbV6VHekz1V3K+bNDUeBZcl5v0FujT+iUpckJBmYfVsG/tqEopSlf1EzzdVKqMGH7zGHt6UT++ZR
GsZWY12WSGpexcAaSbQU7t5hoPjdr2ekKpfhJLi700/bkoy+SaZ4mTI7iB3NkeUFzScLGLG+vreL
qRy8t0CObpZwEst9+neX3qR+RMGKJMT2Q775FM/B3r1nBsi22wMIRKtPPGqdxahYMDQBzxJQu2xM
X+41ikE4XAPtEXPpA25Uxb7bD7Ts4XGhaYOWxeza3H9XALsDtMkwxauNBS6ul+fALHB1RXfG6p+m
B806gor7h336pvBQO+SJGvugPyVNMx97KXu3UEZNJf8YRd5Q3zHPw5dh7Z6GdTqk55kedNOqu89c
fZHFKQ332F6w3LBr8b8Xi2DszpjZiN88ss/Z+tvWc619t5MdD0OBCiC3ST6ZCxKr6GsHqKda6hRq
dUxgas9OJPSSPDMOLq6LSS21SRN2E8+46VK4brp+9FtLP4E4b0fN95j5NUCPIiRUqwU1e68wy757
radA1B1DGy3j3DL3feXDs+mUc04uqrxQPCaWIesRHxbZtM9/5R6wiecJM4k591HUWXi7FdM0nYqD
agpOkrecHfAhDvvhn+m7lcfD3S13qczkrnOOGykoD0PTxO5jfiB+pk2rELsHk0uhrVVKFiLVn1Jh
OVJ/l/Y5RZ6azzw8xMdmEo98X7WSGw3ku5VOfO5rGYNRr/Q3IvF5luIaZ4TdO2FslBk/cF+Cq4VY
l1mi+xU4hhVpyHIQsb0fNIzcAvuqMTZWod3Fwxrc5fKnFUey64GxQVCvCdca/FWsYA4uHTXQnwIO
5sCXPqXFhFEU4EIewHx+OTt2E5wwBcmqsiXJjzf1qCqNItfFo0BesSzas1aZ0nMD4XSw5nrPfB1G
nCi4Uv0YnOOcR6KEFJrguBSgZMnlyd8yQfHip/GoeQL+m1oqJJc5itrpJQnIeVM/xlT84daxJaDo
bBbMLPOuSMTK0bp/Wb0EV/GXEKyfW/wBFGAX+150g4xxoMDAfDFuo7qfpi4TU7O37BTQ8lHDTkal
WpwEb/4IIfy4wXSN1mSlSG1bNzArGqLN7L/sJ1r8TLTLbKmXy4+mtKd4MygC1uAXJt9qkczT8IBp
iwV6QpR01DPf8Z8IqmVF94xJ0qxtu8PU8jemXxeyNKcWGvmk0BvMcaTe7heSP9Y6lQntI0uXUUYi
9xssUUh/TpU3ZDGNzHxgJ5LF72sAtkdhafef/EnCsEUb9Qdc6q/S2i0d68Brbm1iSy8NjhxlSIJt
ddnRhp+vAU9EAKH7AE+KagWoOrUvQGWw+uqLMEmcIqvfO8W/riAX82Xb4ehI2UINheWTK3XWc6iW
sbRxHe0Hjv13LEsJfKtf/KnQtT+QpQjMFZdXILa5IAFUig4hexI4OQafcmrda0m9SwaQNctrRec8
yBBj3rxynTLZfmdCJE4w0DiuF8IICehyGru3ZTgKxE9O7YyPIQIloboRT7gHw9ENLnAtodvUFR3N
uTEMAYs3WnCwTA6tVGlQYmp2rB5ib/enmUGze9TpA6IN8/DTRDkfQHVvpzj58f+PWFRfpNdawBVF
WF+f38CZTscMAyc62+vai8tWlmAuBxXD7lWxqAR9Uu9cQgNNlxDzaLmc8JUtkpaY4HLodFm1EgUd
Uru1yCc3475blcPbAob3AByEi+LvcPTfhyexX6u2kQjkkR5txNv3Zoak1nz8Yq5rUJjP0ERjZP60
MoZOlmEaVZv6U7pAbWN/L6OTn/hTuzZGCC5DMbyZii4N0J1OpG4+Mdhgq+DzmVqFxjM1FWmfCJCg
av+n0M9PIIYrd6ERO1U73DQdxmYIMCdBFe3zoIgSYszoyLBr7bFYJZzJV4O3R+o8CrrfD44u2tzU
guy4Sg46muIh2k+C87lMf/KxkPU2uYVRm7+qFOSHc5YRKwbo2u13b9aoY8EAUuMG783sqo/+4eOA
K61exjFYztRLJae4rcsWL1suQjsz+zbWwUeUpv+o99S4ZOXZmijj+F/Qr8hrAOJEiBcTTcGk9nQ+
xTE0IRXoy1+PKazndseb95DZvQ1uggN8x7DpeGdGSjnMEIpKNDb5SyZp+YLGy/rrTqgfbXPZQm13
s4CPExozh7qMfKyrpG1XI47IIiPioowYdZ/BEbIrHoCJv/a0BCsEesQTDcI2V9U8lX5FO1GJJs2z
mWaYrGLmMtpUDkfqf29c40P/zyXI3lNZY6cNdnviFd5ZGZNim0kwqxEUua1haKJ/hU7ojSogKidg
Lv/zE8F87zqI/hv//NdSIwcYCVCM7RNgmlVxWtBCdcSvBiSNu06M+t+tsfqhtx/5/n9Lp8ajJrbJ
Bl2yJj5YkUCh7bElTVzjQ1BF+Wk+tJpwKmXfX2AUnbYygNtqRia+IjCJ3MvJubOFli5tXp98PClL
TjVHSLZ4JwgZWMwanJnLLLvJ0iJA35wLxHPd40bQl/vDDXrnoHpQfoFm4sEAiUQqgxmEGrE1b/1/
Z/NLPPbDdnxD0VhJ9jpEk9+eEFwi4Ecn4r6+yJbUa5B2+L/8F9gGYlgUXrREXk4yNfyok2YUoaih
QZcA+EuRyReQnBL6bguTuMCPAmPsBRKP++YQOCu0Pa5AvikcP9ysePEFcL6LgUuKQgKwLjK8f/m3
sF/ZVUybXp8uX5xPlQ0FUY/m9Qwcv76zijHYDGiZGQdaMC8xHybuinwog2y5UuZh0m+rYlkkV/wv
TNssBpZJw/z7+XiGMGd3EBZldj7FF23Gm8stih/DOsOlU969Xbh3tA5sAIfKYnqDQFHbivNRT4Mc
mNbS2q/s2DANzZr2zLSUsPA4lDr9LDYUW8ovER3xBhOeNntMhiDPA/nwzaoCJFZj5BR2x6jQYgU4
tc+0Ct7ugBc6BE8025hku73obsn71aWrf7OtaDkkuZpSt2Yf0vpOgSnKSZdluZz57paoOWzQKv6Y
TpLXuKb1u63V85Nscmg5bEIjHmTo25dzmTzCgZ38fH91DKhiCavOjtzliPLrFz75Vp7cWSpxffvb
akyjsNFKQRD+Tjhvh3r+T31n1Ia+5+tnysmt42i0iUEKoe1WwkUSICVsgOSJdlpbv/wSyAxW9RMm
yHvSYZtJV2+0pIgj+rkwWCc0p6g9M3uxUvtWvBOnD6W0NdqWpMeE1VaQou03HoCEJDpyGtJrcp3U
jw72NWB33L2nR6PGaj61vD1QNsOhT9ZowWvcrw80W3GqrU+XA3ei9B1OKFuGW4HfEaPsAARMDIGK
YCKfD38OUCbYjwgq+Dq73WktqSW7lOdSOqE0oE/WZBcSMBZyk1OEpFQhGTKfCBfPu5Cm9iDM/rSS
YUFPEHZlAnYKlKR22bDLvuiY6Gfuxe3TLvbiInI5RiyKtggHYbtfNIbIZQHnmM+xFnf7MWlBfTv3
lKSz0b+aEoOXWMBDhJDcePh+1KSdryoNdal9EQDDEuQWNuFql2gdeJJ94CCJqA1eEhccZ/Hr+hSR
WF76wECidx9ZQQ/4CBYzRdLBFAH6jbeU6cS3Nb85eySeDqhtz+d5o7sxgkrqEJGZXkTS+x8WrtPW
qfHzuccmJhpRBFX7BQl3sU+2nUolPxVnA3Q+4/GBOrwgUs0hpk2/+1w9hbjnRTbo3LP9/jZUopKn
MBnHVNJqLQrIeKD/2IoCx36iR/mhUb+4L4hE/DnKTpgc1sG94GuhnJovtBBJ9riCRxWfe17H868Q
ohMrLJNod9ATHl9Pjs3ajF3pdvQCjUyxJ1oFmuksI1Ankix4oL+bJCJ4WRTaVr3JSrKNZqznlg9L
cMJ6LEkkYosORn6cV5EPG3oSJgTD6NaJAv84mzAzdBnBsD3n5bdIWK5aeRx0QGaq0nB/+OOEfmY2
60BJQ6gvPprN3H87aiKNuIn5QJigCOJaPVfHYoxa/y3ja1IH8AdrMqE8r7v/Rq1D5JfHbOk46eFn
nX1kGLsR1rSXj82vZsoKkuYHJjKQBTr8LR5KxI02OY8UDe9u4LXeEOEjErELqLr5G0LcabO2u/d5
fv7KyQ5a4cmgbkHJI1iFn4zjpBTFNqdLz/bc7dPpagRggUnTaljGTZI6+XLi9qqwZ2UfLeDqE1V2
w4GPSJ9rUWZZSskkpZoMa3AFo8PQbQDCqusj95ZsE8SxV1LzhnOwGfJHC+Rmo3yJ4AE/v+cS6vDx
puAZnGngV4j+lquSwZ+YUSJiMRIrC6ZdkMUiflTf2XfvxQgsd3Av5lZ68+foiaJFN6Xl8R/Z9NiB
bgPvWpwUArVdZOahukx/d6AGlvHjF92OnSupgQ4hUAMSqmiRmhZzuITJ3Y81//dmUVkkJ3XcgPOv
54ZgM0BUehSNqc9FdkKV2F0xwPm9jqwOVjS2TkjVxkEpr1xWT7t0MAuixH3bjObkI1gAt0T/adQN
c42c6lpmYCXMLmWxkm82B7EN2LVSlcF6B+L59jCh9Fwl/cMfLttLjsFzMH74KEvKkttG6ZdnT1VN
Pc+ZmI84ZxXwOh+8wyTMJs9O4dU+4nVjPoAk93FYsYXmG6oA36OMwYABBwg6n7KoHArWvhItx8tB
BRo1mNxLEb84gt79aZog8R2WZxZwTZYoQNmQ+/vfGdEYA7ut9Glx2chcKhPVcCtJEhJS+bUWuIiF
R2nmjyez47bjMiK+AsLvqXAOPV8z+roN7kODNJF1MnuKMmB4Y7QWcyibrrr1gl3xDok7UPUCquFg
nZ9iflZlFnN/RvjlGLQzq8hJ8jL+qKPeeCGtHtDY+peAJF92HTQcIWldE7Jwa8kh7Ye4jKWMABaS
KSfEk4uSMZL33YboW6fjB9kAKaDOR9elI3x0GDLvws6vtm/3kVpCr2E+BHpbVDT7G254mGaN0F8N
4rL93Nn9rcY84fqmWX7UUJnXQUI6Atq/WKltVjyZ+PI5etnvJt+Kp/DDu4aT4n8E89SSHasvhoQg
NweiM7I36+vY4dibeUetKQyHPJsJw+oJQxtkUyVp5/iw1l6JVqurHm7UqkqXoZKg8gZpWuE9FQF7
XPq3iH2v+jt0+Wgl0L/aAYDgBETEOLrkpc3fSZ41yvJKtjeMdyvViYMhoScZRsQiSicxJAlRKqiw
+2gb9GPYhtR+u+s2iOkenpMIpcvhUS2B8+sraXfqWKHUO5lqV6v8C6D1AKrIVjaB66EJ1ig1eTDY
stn9CHBBntG45ozZP3FefC9RKlOBfc6GP2JHzq8wDTaAlGT6/ikXBRPndwlWoPvCpEHiimCnCn+m
MOrT7AsIjydN3MCrDHc4QAvbY+/SLQyj2OZP5tWkf7m+aCy2Kj9rzVh/xsmAU5rDW3g5lL0otcJp
98sTN5ofXga0VFFTaB97AH6WVram5lJErti3IhWHXhZnepVIZn6G5FpNNfBId6TlaEpuekhDxCLf
PHX+TQTKUtdZ5aumOpoPI+TNts2Km1+ZkwWGYtcRcg27r2L1nRtqjDel2nu5YlbkjqwOIryUjRIU
Ru9lGSNCuHlrNjA3MZVrQBAG/b1WVJN9+jEcJASVo91S12Ko8hz5PqfnXSwVn0KlW2RT4E2rNHa6
/5QLUGpj0tHWveLRBENjepyMjznqRZ1SnFAvBJ9WDEXl3Q5N/k0mbJoSPilm3GBOlwiWa2qmJxml
/tnTHquAcAx4eYDsPXtMYRvit9OtIzG7CPvJqFzccNyMztyWHWZWnYNloKJ8oNz0j8/EYwL0YSmV
KLJtEXtoXXo8yn4bfjx7H7oCoXlr1pacnIUkrwvSn3fmVLMEryyp0BpRmLBt44xk3tWb2IQlfnTc
q745s9KJsnNa6DSYGikHTegLAKEAM/k9bRYknzAk4Jilr5BEkg02EsKjnvjPVXXNaWk+/SBKH2nG
iB8eokAn/RgAXLl39QiJJyo/+wPcIy/JOLmPIrIeguh04mBEMGAAetLy+BDdkVGWPHIiblkzXHGY
HeXPEuS5VcPHkopeq9PBpEIwD8abI2K+Ua5X6ChkMDywiSFJCU9A8qUpBjzCFOqtgWRMw/fvhC3D
XQTwVkeRcI4O4PsjvDTFHyagre9shG2OfsxUfyPwmoybgezRIo9Wx7Ao+EbQm49QKuEBKrXdS7eG
4U1NYjAYb364YBxl6QGqLvMakv28X67VOsy3Mn+QRkgWumMQN+zNMnI8DYET9Gfk2e1DDM/LR53+
9H4rFUCVjP13A5KTes78P0orYTuLEDyEDqIcsFL90K3v7c6EHnBJcWk0xmsF5yfKvKOpf2Ad6wr7
bXgokgXEqx0SkmfvwSGrcBYd8sYHQRtY8M2HwOBYs3tC9h7LujTIoYCSyi0VgDsifNaUUw+BvOgG
tw947nrXS3fb5OJ6v8xhMyNR83evz/DeEH+cCsk/mPqBoHX3i9+cW3WBQPAf7dCGionrjkaML8M7
8auQAiP094CQ2auZTWoso0TsXoeDSUMXfdyAQEfXJB0eBwjjZWRjjCKyIvyq1hRLTvtX+nFj03VU
ged0ZwxqlpQQ9IeBdzbXLjf87EkAQMVYHx0zZPfh0tYsXqVq1vFRCCrr5/hCBd/lghUfFoYC3WIF
1tFreiRQcvfgEUVhccgNVKdlQU1HklDSP9p0uwwR6m1VBPh3ZCN1hjMt4X8pGAbOMS82YpvvBQsN
oa4WOhV/NPigqbEh/8g2I3ni8sALAbcVAyrKr0rPijw2ZZQ2cPXf6NiQvpS6cUtnyZ2efjtg9Gcb
pIa6bNrTTrGNjnuCLs4ak6xsMq7RE6uet5X2/scE9hDTYzpHAuKj1y1+gZCIx1AXIB3ijE+Zvg03
of9doEGl3iFx4O8eWA9Vc5njCDI8HTyEbjCIcvJAvXHY6RLDztL6ZxyuE9p/bJI0xD12NXZOV+6O
m/PD2xz27Yn8N6AtZ5ZcG5zQqupj3l6A51kzrozkpx9lVg1MySqd3xlnPjgJpBPkJ9jugXD5qgv0
U7IopxV9IeHFoVxUeAcW6l0X1I5cmizvjgEyx40mG2Mb5yzeeoUWW8wmjYbiLpOMQTz7Kk++zdt2
5URs548vFHEaTcqY6flzPbsaDdOeA7uQHwsHZhm27zh964/Yzg9cYKCGsACDFIa4UAvGP977gfKt
7+UMtgWhPA6+xs0osjRf5kLqYpKv7CLmPePGpP2yMFBxL7AoLU1FhuLrFDnV3l/4MhYDCqedMk+B
0fcG7v2Q4A8jxbeqvDWkuIn4voRGW/DQSMkFkwD2NVYaq2ZtYqWi0Q7LNpzjM1YzYooh9PKJaNgh
LPEiUgmsim76P8mMG6u+SZ5LdM5QmKv/lUqmulapo3BHPZC1K/LCPUNtpT0bdOQtlGMOYQBSswc8
gLbqpc7qwscUGhtya/34zHRy8GmvLeGZljsGfW9kz55zFllAhWVhSWL5Z7peO+ocPmEPwQA+U072
FAnXwEhFVaKMzCtV0eXwrs+pPKoDPezMKehYqhzn5ec96BQtfhJJZTtcUfjgsVEmLA8CkrbkN7iP
xLwnVQNLW5S41CQOwiIaongEUEtm5vFGUa7BuAQ0qpKZERfEGHwGKwR3cGgL5upXw3IYEQnbfXTC
h2YuojSeg+ClbOAy/rhSNdcgL7d9Li2zhmwMz44aLBVJOs0kN4/yPfnV11obe/qTYy2W/tqfcEEU
9vsIXCbpA9F564m7VyR3Uz7uDxuRcH8oxUsJsN3RU32pFfbgXrIFID3kmdwPZvfCstul8g0+Hjny
IR/WS1rs3ds1lYCUZb8CjT1oVhkyi03QAlB2gzvv5IUUaExtbnOUglhp/d5RuiB4uSmXMhkuKdYW
EWrmYGRVcR/i+mdAGCiOiaxETp2U5zN7AnKyxolcA5j0XkKaY59UIFvssQzVVyI2RhNGKQfItmtj
eBh8vhqeQU9vZvkLRV20QinWklkt+2QbDFTJplG9KnT5hFNVbxF1ELL2LiyPi790RimxRF4Z6Ph3
v6WN9LpKaQa3Qh05aC1iQF7vDf0eVVP5jmtlH76NsBr1sibuzhkTWCH9pQ2VhBm7JAHRcYOlrngk
2Iboe2EAcd/ItSLv8PYDoi9JU3ZkBujqD43ZtpvBBEy2qOeV70CjGE89p/PdW6M/VCYA7nKkYK5P
hpPmo4YQ6+xM2Kw063z7DMBLKLIe6cjOsJ+E8yfFUQrO2Z1xsfnN8UE8GyY7pPPPBOB5ZeT87wKA
PDuUx1MVCBxIqTxRXxdkXA0MOvxANIMEMs65Zy68kfSdP8FBqdCmAG6tvaSjlVlgt5kxjQPMNfR4
4YaV+32ewCVsQW4Mn6wfesTVT0VhQi0DYplYlWyGCrRu7SfYOz531Ytec+LtSgg6t0NwWTGcipBD
qClm9R/4EoONmwvH7jUFMqTHmXyO9jThGvGBwbyrt3RuEYPEmSSVKkzcCfet3msHHNwy//3kTBu0
WMAXP6RgYwASkR/BUIQgGZjxzXFl1AxAg/znoTxp8tR/sgzfKmpf7DmNPSxaS4t+KAJSZZ62vh89
1fSgXE99I+vIt9sop3nwLzH52XdWXe3RMgvmf0EcQevJy44r+vl/5bxwUEntOmaeTjslZmKt4H4M
6Vehi0/YXkl+hMu6l2WZTgIyf3OwxdbCMvrXgFOGhwjdahnZTA0Wn48gZ8UWMYYdu70pacFokIJd
JNoD+g3vqHUfGQaUp5NFXliET4RbrmmxPhz9TFjjQQrhLUcuax4oHV7eTsicl4ZH4pzOwG7pfg5S
GO0WoEnB7RSY55+ba010ntRl0l09QmYx9SvOre+vH9FB9ME6Vdgm2lv+WVUiHqiC9Ozd2JNaVw2u
OevizECqup6Q4YBp0TCaJo91jkBpCLPsErzXQKKLFR6jrJNrOvdQtcIQtLE4XQ6GzNf2pHexs5T9
i2C5Z6ATmZegGGW+spOpYdTemh9EoOaX2XuTg88f/YouzMe9jz6Csq+F0q8qRdd3KyFFPsLVgOMC
9goC6TxigksS37fuZU3rlunH9rc7FL7yblYCOhN4sCQ5hlOSTfJ4KGiHX+OpAsXbK+tjQx1npjp1
cgzBn1x+IjP0KJdi7SF3SvGnxCEpSWgKX6xC/uNYEzQCvyLcy4TIHd3+8oBn8GtGWP02BeIPWfkr
SrRaP1lui2WBU+dbLzdlJBLqOkzd0hQHcHxYARzbZe4VMlgginNeg5zxX8rbDOyW0Uhxx/Elc+hA
+0wiiPGXuU0MTq0BLht/8QZyJtX+zIDoQ0kjgs/sfSjffUi+FJz+mjly/lk2qytY4+EODoq9HMyH
7NMpsLN5bgUiUSJiCHtbYRWNm21L1B4lyxgRTo2TGztl87zzBnRwWx9h5eAb7slQS7qyn5xv7o8M
6inJ+T7rU6o5hfPOVw4kRUfdfleA+pI/E6g+TnXpYuzth37FS9ekHtm1fHAI+CRREhP5gY8mqI7u
rfvvwjimQDVAcRzK1wHdxwj3pspTjttRhVpABhXDyPkGaEZualI/GVuKoRm5D9D2pNPay1WqcH4m
+KJ7iiCgMSPL/XsMvUgZ2FrTOINDAdA1kyfrjmC/dCpi01VhCO8khjhk4ww7DcpmOQxWUcsUl/Lw
tu+qSf1PS40JacOoSC8tJJt4N7yGmaTQZ3qt2wGirCBE1Gh+DvfwdEYEHR/zszi+AynvTM86DbjW
muC45iykRJtsP2QALNcwwK2u/YFffLJPlG0hov4Z/fNbUVhEThNHUPTMsiLC0KJTdoMAL/Mt9xH4
tNMT4iowERDZxPHy1p3iKKNkYvYnNoRgA1ZZOpefDDTQpHSyo+gjJL6/11xViMeX0K2rL7qZrSYW
Shj43wsWNJ9rf4IpTLDh125LY689oEWBr3F4+sJu6rG7czAYFok/BZKgCOVnCga1FLNx5+qJReMn
x4fnQlXP7QJCkZbDWbKKbw6xdVWwUJhfUV7+0iPkGMRzI4tCV4BZ5G02sY+c7qwJRWAdIg32n+wJ
hUUmPQ7+HIvlItt4s3bmaS0PufrGSan7hAmtv6HiJAytXu9H1JqMJH+pel/ZjqJwx2bxtYdpKp3r
bAxusNdoTXlwnhI97Qyghid7MtlOT9yeuhhU7fPLC0U0DXv6K1p54SB/QOFAPaunrmOraWtiIq++
SEhyFTo0O7YojQkevPP4JaChxwPv6REgG5SLeZED04cbi8j8BdZwkCj8+Ehv7dJWoTaTVf0Q5YJf
dptOvW1G5XNE7Rs66vSqHre6BsZmiWu4h5GPDyyOzPkXzTfMznBcTZiQmnp8CrExbAsUxfpaIKyY
6nERsoC8pU5bSyz/jQ74SIlUen+j0bfXKQtzgKSHoTBep8DdpgEwCIst+j+TNB9l/QICFu9gkUgN
jLWRHP2Cm2e9hZEG9IoI/94q2ZIl9sw3WUz02v0Bggqml0RdSq6fxbGFBfNIN24EeDZpo9jt6Bow
Hv4z5jLxJUN+tvH/Ooh0n3m9o31aWyQWEOs/iTFSMQs5aph/f9awmVKpElbPq9q1m3c54kZx45Hy
Nth9qnZ2tk8sbOtwlITbvhxTCngHMFwXPrNCNVUkTuOqsIUMaSdCk6tpNXgIO/Qz+nMOhL7SlNka
6SwTkGWpXzip4/qQePIipKDf+jeJ7T4lKoQXvv6Y5u84d3PLctiTrrViZY7+NFifc8cZPpRQH6po
WsCd3cnI+SNxEWmKsoEIzdWvIuQL2JLHe52FVVcT7FOsnwgGvjxfHGnB/uEIWXTVZOfkwOO6Hu8p
+dMac4lz6Lqd/CdYG32JTLXntDbQHMMlZDvOUG6bjYgN0Wy69gP3EddkrO/blrwcVLo+vbdhlXMI
rc7vGugzMQCm9OuUzGsLUNNZzpFGsasCZBKLeA9iWtBY0M8t2enVMUHPMjtdlmXCZrSf6HWAUW7e
YRlEyAHsnmOemEkS9fUFGPda7ADOonUM+hB4fFs7GTsDOnFNZtPv97HTYzGNQ7+wgxt5vvKStmmN
xPCHBFCxAbVgiEYYodgQKX1RatiXQWtIKWBTroqRNze4Szhs72R9HL03WmgsF2I2LZ/Irhg3wzoU
JyNW/yLNQ7SgqWw9znS+5RVHWnl6nrk6ZXAeIDCld4BJ9RHZfhLzz1IzLwXjfudxaJTcnQCk3B8O
6T4AiaX+2IHrv9TWEnnjqsPD9o0XQPmw306qDjRnfuMvJCVzbWj1hRGoarBaJb0Y7eI7cQQBzLA1
LRd/rkQC41jzrjD+A71wIVe6P8gh9rap8mm/b4/yIuYwBzYJrPAnhc/U34gOtxUvAqpD8ZH6udFU
2MYcHBx2JkP+vtRbH7XlHUgdjRfU6sIjp1E3djdfcME3Tx3aj0Ce0J952PZDQ1Xij41gy5QgOR6z
DtowEoaqh63jgm7HXcDem1mJ7YE4xnv7fRPDSprutNhSCuD9e+etSgkiTQcX5Uu4sMOvsgoCD6kL
Bq5tDFwuHW8Zo8549oPTEN+d4Ojszi2OzXmOsDl6qa5+pXuTVM6vY/t6+BTwiQKepK5AouKgFjFw
vXarX/d65qtB445++gpqHfDFaBcTZBTFvgdu9qlaNqmxWEkbYHqWQCLaMRBTj7E5BcYRRHw77s9Q
74MNviEmFRyvaPMOnXUz7Zoo+BFAYbbRszMH4mcMX+FnNBvid4uIRM4d8/RrNqppiggTDEX9CJoq
axaEo0EjNShyAf/7ki4XSTldvXJuxiYgrOfJm0fCW3lYuZqbNrAV8k0G5TjBb25xpu27fkGfoGE5
KG8Qsehm8TC9cKGF+EQNW9k0WkG8g5c0FvCGPpFoi+ixVytuwbKF6Fa/pgkrt/wc0YacTeqgphPZ
hP3QDNRDJ7SJjQXXe42/U4o0WwBTgJzv3krhtkFjVkPZifa8Z7Rip8g4M8MX1QIuZ2IdbxLJiDDF
RfrtTpNEWohtrfuDWMiccrIT5CEaD0SIgwSPRzTKrCcnYnEtMtcCL9mJoyEpgcrdEgYtHV83UURi
e33dyXXoGgmuPvcX7WL7w8TVQqh6hmPZOQBpI7c/VhSPISI4LuVKyUlSZF90/Rn58H6GbgFMfOV6
ZUHUMV5qg+yZFHWJRyRk7PEI3ZMW/KcZPDeiBztCji8WfrwNHabTiITGoemOeQdZWUmLQITTLFUk
H4IjQJLJ7SjsItLFrfT5V8P2/bc4IKH9kC72hTZmR+AagNbkCDliqWGoVb+E45KH9ZRDTSycsca/
yQE4f5D0XE5grQ2t+9hkxAnAr4U3+m420SR2883o3dETbjQ/IdUksxheXQKU2KBKZ84QfhhcxA6L
QBokMS4MUVVdR4xdIiGCwWH2XHxwLXtYawb20p3f3Z++/7NTwXuuQjIAvzhaReqPwloBqocgcvoG
FaULEZ+GElUa+0Dcf0U8oo4OkDeLdi6hrdlTw+cfk8nFf3JDRQSfR/qScXZYEfgMKu9WN1wXML2b
c9BYD9xfCEr0A9DiqHhZp1NTMiFC8f25KeR6nDLIpE0amqvVJ6AroIe3nLKxa0Ei2RJzQttZca11
le8rgKjbZ6ZsU6XTrDxGid/1xzn+lm2FimkDdJpw0uNDV45p6S4Zwx7KPqkihG/PPO3uqVRaMlKL
B7LETOjmD3aORw4gI6eCa70X0et6Yx4fs7OvAxAP9lMUyl5oym3CTi9fwhUdcOwaebWa+anztENy
gBYZ/HmzuBaqZjsWucYZzBnRpCFVp+OqoJWKSKBbUht7awVV+vKAtyL68Z9eKs0s1sWQ6b7swVFE
7DCkoAh9Wu9ixM11fTdkRsbcZbE4b3l+AcWvvPbeKXjoIKAb3KfZF8XhVHA35i+MFvzrvUlr4Nbn
gjP8tZd9z/9aNB3UQc3KQeisILgC85jQnvuW7rWzcpGwgZ5l8tcEJPFmse6ZUCuwQ7GKBU0TaYft
67ExiIxYNJnUe56pD8wfOuM6IhsdEeb5WhAXlgrycrc3d6hQnlDxQXUoDPQtnfiH5O/srSF8KWHq
8ol1eIfPkS4yFJmnmkxqSRQpfRK+St23kml4VWLTb2/g6I32xkW/bs6PGXWGSyBJSIN1BiG2XJDX
umm6sTnsae+d1PTQUe5N3U01IoOlUFBjmGRV+N/+4HL6/zYjSj0S8JQtpbDaYnoSoVc/S16IjD3S
Ejb5yHbChxMBeZf08cxMkxI2xmtOcs5kTpvNeb1MgFVBlOVVgVDIT/CPKlXUj7oJWDcQ3PRcHAeW
siw1HEIQ1D7IUbipp2uChhH7cf51VtObAinMtlu7Q8wNbPS5Ik6LxiTqaYABz7zkagH4pDNBNCYu
Xsp/aSZvcnRzC/6UVij8TOLus8hdayMq3EJT4/mJXpFUpUjL66c5bAZXGdCqNeyGmlFpH/DH0OGV
ICylRK13Lwbm9Kat4tI4giJv4+zeshmqd/C+LaL2aWh2gDFls6CljU42dr5gJunWiP272jIR0t6w
D85z/WDoVWc4iDJcNVPb7ho5t7xJPY5e6G3PVS6Y7nsH89qt7sZLYiHO/frCbIbPMwvojas1+C98
zFNdnPOL4FkvvvE8TUDHk1UD2YQ8KSg1bBJkqpp29Y4wxHEL2pXcxUKfVZ5NOSZWktIwrbRmHeGN
DzGSwBVwp55waBepSSj3abUD9gOC0VNRw8FbbkdUznw2mXmUMBcfubXFZPfApLU6t+93tWOPxBWZ
3uDHVwFnsVIfUYca24tAg0r2aq/TLYofeUGmD+7oxt5WKCV+QCjCSjf1TsJYGQIBj8Agiv/2rnRM
tvNfgRi8OwUqjEX81EUsItuCrDidaxQIx2CpPJE/MAxn0iK/4ZjGO8NZMNTNq8Wyb3uCjiRrrOY3
pJnN+x+/R/7FPvck7krppbMUt1+5rQOT7+TC4+/tlsgOlVTzw7da8MS/VsM+T580XWTPikqHpeXP
a7jn1KIM8+LU8L4fIlCdlhYM9fxDh4zMUWhklJl6CPc6B3EGWLTdGQd30JDzPNSW8RKLJ5dOC7p2
DHQExgbRVMIGOJo36XpGVdk7oz4vR7eJS8Jp5wsFpg35D8pLXwmjvqpJuYOlwJJ5jDy1c1Rfj1yy
/bFBe+tjjWdWyv0k9IFUrW+QqXO1jOc/6BS0URR0VuD9yRpPHM9MhnPhzEUhl+T4olLkU2ABglxH
ndw4GDdUIdeXhs4UXoubhanujrAFEKXFwJxLsh+fgxrP3dD7Teu2gHGiUgxW7ozMU/vrPXDd8Epm
pr54vmWpGDvajDaj8HJLNQXWCSaeBgiCeEuPAo1EwfgnxvslZT9/cmjlX0VwKgNc5yciOyfHqf/T
TyMvqF9Q9JtPrtSgN3xnKCi76UDwA5qTwklBf1cbArSdE90wrsHheTnIQjq+3uQ9vDXDvPK/rG/X
UnJYBPkAJ+XJmAu5RdDZnA6vfNIBW2Npco5q7FPZ5C/WyTvMT1z/x98w+0gQYkF7vOKZJI6N1LZY
hi8nLHqlxtuMPhkjnCRBGouqQEKJk87UlOjjheHC8tHXHNnG4FbySvESuCFajBPpDT8822kaF3uC
W+bUYgWCXapCMp2tBrWzED57Y4hJqNrOXDYoZoE9HjROV901eY1qpShK2C/wMC+5+hwME5d+4Ltx
ewumsfY/veMfCIl/kyKRpbpeXjpnVVF1IfjhVS0KF+KHQFN3jj0pbRzqu8dejYvuyUIfH2BexGh7
CqXGlMgNRA7/SUucMQmq6cPgcVfq4yS/JJFU3jMFBAGJuf1Xh9dFaBZCE1A4mRBD1D3p9aP9Fd9W
Y5V3czhGCMC59Scw6C1lHPJaCcudOIWDsXB3GdZtj2dRLkCWPso4oG+Q1zpgBE0nMvfVD1fAgQph
k4FPeP/V+KHHecP/chASlsElsADi7E6CL+VpJHlOvitRXMM5VdpwUOnfY0aQeih/kwaFHAfswjql
TBcsAbYTeCGNhFjCjf+AYoMCfLlWB1bDFVkX78G3Gl5ulcMGJUI0gb8hM+Jf/BYds/Q9QTTGtNd+
HwYL2uc8X8YA7QsmKz7mxHKYmQ7hLwb0tYsJ/pQB7G9MpMQXefaQ7bw+s1n9NxdblfVcIifsRQF5
XkzIy5I29xdigPQewSC8yOQIeCHV8xQiCVyRGy0UkPtGPiH9vJhUXnX5JJwwvu3gffLywypw/iKf
KS0JV6X4AbMQApz66a+sipKdXnjmJog09Rq098rl5V4cDzf3S4leyFCIwd94ZR9vSNt/OefIGKic
wAbgOmVuN9cH0uXCGlBL+fRuj4r32oGAOyv7wmYETBjCvCMiAfe8MvTbpJAdkA/q9ZQ0b/uyfdxo
HSmC8UYegDETZ5CT+OImuy34n1iibR2CQGR5oGLZMogFNSC1+Lhyxyq13ROjwi2+FZAYlDCcZrri
MDsFNrBHVJccfif9tfZXUGht+5Y9WgGzuvm5qdBIsQKPkp+zuQQSm0N91uqHXS2nNHhD1bO63ijD
BfeM9DPL0hbmen+NHso5c+TQUM+dSdBsvzxGpRGCq+QT7WHpvrc6N89SBM0QmUx3YVT2pTSgroje
IS+ljHm6Kgcf0oGMqRxJW4gkrOZ/Yywuv3FcjXw1MvSio1r3puX1bllScfvUVAkP2A4Bc+VsyDG2
coEZp0BIv2LbDKCMbXwLSFKWt64aNRtDCZKufec8nVu0kZO8uYHryxRT/Ter5yNDfG2vnArPcGs1
JgmNmvg1MVGYyzQfjjxa+dPAUK714v1IFkKaqVO/uxOzbwpidOQNj6SG9RPRFmxSqa3Q478e+jBG
kk26VToHBmq1mnCsH+zupEDz+ZZNBCoVVFze13MviJfzFpPECulF7Mtjfc2VWxkOutoVRAnLzuEV
4nArpErg4TE91oxoIX6LRY1nO8qqqSHgD6+hP0eeAOGE+O7xjbOEgt1uFvo+FDHG/W42LsbORhLR
sZzutNC/8C69KrMotxgxS2Zz7RZF2LTIx9SbbUmVCQa248V/ll4KbrujRiVICLW7rrsTHuvcEuVN
JgRlfn/kMPfEfTEss+sAWqeJSbUzkkZkQT02CSE93RBFmR4g7f2ffscoNXMg33UDWs3ELXxAZ2a2
bPe10ZHOyuUeUtV0aN7OT1r4F7qASCmSHIPCzskZT7NiZcSIYEMUcWrE9mrszHb8P0M9Lj/QX2uj
l9H3F+FdShdIluuExxTqK9vKFKWsJO8G9KEi0o2ytQXYVDwBwhn6AZy41hvMS5ZGCd2S+7WlBO00
PvCjcneV2+BkiePc5fAR37UUR2ZhqmawUSGp6zx12Y2Jqg/ww3zqhgmwQ3BWtcKLAVn4kKON5wKL
SKqQlNgxCrYgNXi0Q3ItlZqR5bmZH70iaUY8MjYhhO5RLNsusrysHraCfYH5WHIPiaLpKL8WcKbv
sr7XpDCiM/cMzFbDPUoauji1DF0Gp5r7WefXq9FxnQDe4gG9+bqVRD04kVVR9vysaFPIS5B9Woyp
raYUA+dNVWZ31Bk/ZgaCr4vv0mbWuXqrSpt1J1NxqCpgSEiDBC6DJPA1zc9gOCPId04DkKrUhOyg
XbS6qXCuid3z4ACpi5dZKAEyR1EBjNPzAgfRHLJoY2WYhCAkF/uAEEzJibJzeXM/KFsz3XJ6Xi4L
S7lhqzTuTlImDU7Ed4QBoDyomYID09FxWlvy4Qy9b96QHi1DlpeIGQcarrh6/g4mkKsj2WV/1mvo
dyUiVUSIkL+pxQj0AJUQwgK7CD324xPP+8UGc1sU19vimr3uXi2WhX2plvK7oUlaPe6xhP1m8He+
8eoz5FbW9SPCfcriQ1rHf7F4hrfQOPfhcNLgw5OQ87BdSJtIMGUXOaXNB8//Hb5CvzkFXqWQ81Fl
mETaR/oCMtex4rgsowS49VNGxfL8e6Ud0NlE4wGXJ4CNOx93OI4b/JAz19KvJknOmJ1wUb2HoWRJ
bqpQq/21Oiz2pfRzoVJWxX4/Fgny1ZB2Ykqz/LzYOGQ9loCCnkcvqx4pWve/2TjGtX+oQEFoTdtK
T2j0a8X17baVrKpke9djU2IruR6Ily9ILC9Ye1P/SKC6JUxuza7BYv1ZkgDXecjw2S0k1NMam5E8
aun3krX6tQCffYgraiaybw0lyYXAuezQeCBBHbFTOqKxzb5np+LUmQ8eHjHTQDm7/aZ1va4gJAAd
Nu0bFAcqVata7O2krnz9XhWjz8ELnh9ZRnedGUQoE+WqM7H3hiZzu5gzDzEVUVMBk4SVG7R0QdDE
xSOb2vRytCHLa8mTa8JEertKm5aBGl+8xffQIdZTHIDidW+mzaGGJSaSFaXyCD7Q/73gbZba2kJQ
fSGG4rM8iG2vLVjqVJcukT3+LuOLJVoAI6h/nv2Tbw/zrF3KfCcoXuoGy2uQ+cxpcwzjRuJQcpAz
cmSD+VdKf9l+H5nj6JmvXU1/31oBatJ7c23u3K4HIbn/KndqHzghBtSoNrrh4VsQAPv/IaJ05bd4
I2MV2CbrpYRaDZSqNWgTyvIPac7YRTAQ8uXb6TdeqrMUp14WtjXCgCZiy7QhRkyHw1rE7tezCWzi
WWLN+xWh6eqvUQPSk0QIH74cn6IhlckzVAdjNIMyvMDwddKbcpKiu9OEoOveeko55kUdv/keVUXu
LvwH93KpgYYbW6I2LEQfNQe5+y63xcdN49ikMwv+IKSqu3x3sGRBgmXCM817JY9wyA60HYDWI43C
NfXPLeX+/Q91pgf1GqmskpnCv44diRFVui/22tELk0evdyyBvCUc4fWtmCNHp9M+iabIQc1mYvXz
eLZ3XnPIpzd+Ew9DPdozZDwcOqOre4tFqSaOe9Z8TXSRrkwpnqpT9esNy/SyvW0cNiVGf6QkdU01
HSl1dEB9VZ44cXltbHNwYS0Ztkb0EiukHlIIheKTEc/FD2WoaLe4Xq4ZUAgkOUEQIySopfPMomU3
ZEMkih8o90u48iVaykUY39YwI4PpPaLB2IoPI0XzMjCEgAMiRdKjU9a8xYcpEH051q9UpfGbceKq
aDHzO7jiXbzuZHTeaySSVqDW2g2qrDRCK4ydfQ9d76SEJ6HMg3FW95SusBwPUfysSoaMwxw1Vmkh
tudD/A2KSeO+/7uUCH/LePK7Gg/ESKZJF/n6YcxLDYm7M7LRZK7AkcoVHWDzMWmLJFDCXHI7qJfN
sxcjfsCgwlrTaCInKuZ24U1tTvADy34K3x+mK/gXiAlS+7/rYX4WIbrsSRqz85PiR4YtFQDpw08r
aG/mB9Ck6wxEMyKSz5qotLFNSqI87wf7VrAYEVTVrsQ81u6l9AKdsOzm/GF2MI9hmQ5loQhA+1yH
HdKyuD+gqqBN1PhSOsJ1RnTYB3EO2EZ5ySgc7ZZ2pYVRUfiqVwJrj/QgiDE8RoKaNjJh6RwBYsZX
ZHMycMhfx5tkFZKfnukFh1AoSsycoA0fuTmeAkyoo3Dt9gGM6EFceL3ahmid6B0G4TBGKY6KquyI
84nmJNhcP82UI4el1y1osAO6W+obl1JlEjazZtog5vd2xNYhCJvA/nigdrDg6tEN7EcZaFvyqIvj
6KBqGu6lKi1Kvj1kHG5mEfPiaHOe5syI/zHd+B472XXJgsqXbjaYCKomZjT2FLxteD7GgQcZ2HTn
+s2Qh1zz4ErgWATxbX4mzdZZ2b3ZUKzZxAk2ai4jMErnNGt0EoljNlZ5MLSjk6QS219qBE2LphFP
6YFoYjszsWv8X7M6rOMLHnBHnWJOo+8s1D5JaiLaoPVOzXKIIbhOdx0tTsO8rFk6EXEjsKydDDJa
lStE+0gaTK17lIzm4AqZGMEVDi7sSwKRmx9H+g6nk8DAtFiwfd99glFcBXsjWCuvI1n+LpMaasLu
5J7iWDdkXYs+k9tESXRUUgXXQ1CjWaZ1MQJXPP7InLrJjFRAUozSF5m9ZGHK1iVygXwYdDFNRDj4
d5XpR0HAilIm2SOfUVbAKZ79aNAAkAJ/L5C+wV0ZGHhLTCld0xxf6xWvnFNNfGkt9W+yMzwthijv
C0UtLGN4Zsv5NP0Kuc0F/J2YinJqQWigWCCwxzyoKp3WM2gWfZNC5GwcjYSPjhp0aBckxQju7ct1
h+PF0JK3zdSyp6rpTDqEY6z6iygLlOa8v1G9XkMbj3TYUPcGvpMXCfcCEK3fpv2J4BnjnDW+VpUI
jPfCtEgewbYGGiPHv0C2qzG+P/2L5yLuUv7Ip5pId3sxdLrY+Q6NdQYRT/rtZP8uWbupvUcPo98d
3hPWZ85P0zM+M1LXvmwXctre4okVcsXtFyjOuGcxlQBVLfheZ7MT0NQzsDl4qCsdyYYk3ToJM4PK
8c6Af427eiXQacLc5vxfWEkHceVChgvw/KJCKBhdkIuByuorDXIsJEwbmMkasy5bUTZx/jMcbVsF
IhWiyK5Nyk+2pa2nK8x5GkqNu/jSs9QsmuvmLvdxGe0J0wRj+LD+JLOuWx8ruz81WN+1gXo6i1lb
Q2YC66wnxp5VCciSGdu1zpTcnuWgw7LMgUWhrEogwcoGItTMX+HzL8YTlUJjiKEKDqMpXQILQB2w
Eg1yDNuAz2TBMfiIpi2IDgJjkn8kcJ2JPMktstrpHhQeSbxEjTkvIbmy2OPChOAtLiNS528UGTTX
r0kA/4eBXaa97KOZldexD1Ml0E0RrArjk5ywNBuW4AMNk7wOi9elOgAyDTQ02oOLLX0d2MWzbnEp
9cIVrJ66/tG6HUktWorsmYkbNRKNx/Jh2cpUjEbcLOcs7/QdMzFSgWaDk9QmSN+KOeIYgVCoywVY
rpToMm2atqz9CzwCDeAHUqHj2bdxNj9GLWQwQXfKAMK0d+nCQQSP25ng8SryhKGAtX1ekrNk2XIE
ro4yz3jXyN7QaH1Jz1wMiTZIxPr4ATQkUGICjjISLQHGkj2eRwBKtKT7k+XJkfTLPwI58ySw+ETT
1hmCPUGyWd/NMw8WeP4egUkKf0bAIhbrwVRxikpPXLGITA9fMJzrywGDWfznMXT/AzDyr+YgwNBG
6SJjwhtYubzqyoAhz4pDDl2+u4zllOHyYZZMEBexgyJqmBKujAaPemfADK+bFNaO2N5KPosjfb10
KMfFYPpQl/muvsdfP72esGrpbAISLh2uGknf0Vs416aEHu2b99VE91K25jD2rbuWeBR9u5XD+JsR
F2xFhqqwdlJcE+21UYXTm3u7I6dzrJ++upULq6VAD//+k9qPx+j7NT0i4HNiKjgnea7Jx9gejAt8
5Q72yukbUZSMvTpZe11sSDE0BcYekM4ym96FjtVSsMZ7XsfDnHkRANk1sEiF7UwAJBkyhLuqg959
+ONRADc5lNhHJpQwAT5Byr80/h/9Pt+h7vYR7pKrKwSStiqHBWUqVyl7PEC8kM9Ugsz7+NCKW/A7
wHFMLzx41IBg1Ac7c+vvRD2O66HLGhES/kYINwkWN4w6eMHUAShS4oPrpABgnYtDZsaYIOEFZpIj
hIaKWbuQB6vEixLUzVmY7TaCSSROeaF3b4Vd9WPTH1TuZdCCDVHriS1z9Z6B54XG4lgcdgR8FtMo
ELmbYp/pbIr3wVxSu96z46Gjf3dvpc/L5zuMAqMXspz9WPuc+eOgDhN7dE3Smu9+wxZPrjr+dX/a
sHmTc0vqSKGYGoeaoV9+cdp5by+W5JtJGuAP988Ev6+IszNCnCy2xObDMa2mqjd8ASv92KownJxT
EJukUT6fkDeKHYLcW9Vg1S7Z6/JfPS98+gOUIZ9BZmtmsXzvUmjddlCV0tMtFMHUsy/OKk8QIUNy
6FvdRVGYa8eXFQDofX0d4jeYDtDTINYs19Rey+LWaQrKdN7X9zHC48+JeTrS4WziFMq6ydIB5EoC
2s1HagYjf3TgeSvNexXUROQI1bxAcGPs99fJPyR0+RUul7q2i1ZHCZigb9YjQGYGTpLlSghIvPvZ
Ak5045ofCifCvXdynpNjlyyBJpR8PCpXlLvNaPdw6dpiQb6xttXPqpVJwgdeROt3E2qUuBvhgSzW
tqd0Z8wNoPodNNTZiP7+QMUlWlmfF2EIhoiQ7caTN0UV48QEtDSxlNPJVuD3nFDa0MWl45yc8kae
99QxUfEgUqXOOuoN+SORASXdmXx6i/oUf2THICoqikc5G2puv3YNQAUT/xo/xCvIdrb9SyMPHss3
I3+89+bFgGgFZnb9MxJC43iJl3WH6qJOyTd0ibGTZS9ydcb7WVJkkqZ39L3GmDusTSuWyXiinX9h
wp/X/rkD4MO8lkqn3y+JN+zMbLPWnjF4ex70zlkaRFSnuHIkkkbEn9u8TxhY/CwB/WTQG2bempWX
KNKBMBteWc2ppzq4VXTpy0G1QQFIK96THykIkH4PyQVO0XCjqIFArFeyXocgJw8yKBFK6Dgjq6C5
6a1n+4gwahpiGqop+h9DzBTjyJKEoVCal5tOIyXc16ncheV798kZZd9fQQ2hZilRLyZRA6Rf39dD
4HY7aJrJZPuesqjwNuHHeBFH+keP7RgbCS5xU5UeXCAvTknn7KaY7n29B8Stn940IbLZGEslrp+m
hqGz0kaG4TrEZ23P+H+jDtScLE493rRwGsOGm9jdgPwq4EiafuCa9Vac5v/HVtZpMlvULW10paJr
YFuacfk5ULFnzQ++8FU1/cZc0oU55BTKcpcBwwKdKPxh7qSPMwhuxyEhRRgiQZuq/k5/EJ5DnI2u
xNpIX1JeTLyClHe2JL9Za0gZgNmUhR6aq1heVH4PYNWPTvBPn0XkR7g6YyH97m7gXwAPPk9b/p0g
uQLUjKcFpICJ+2JFZ2HLaL2I6pwtTMXkuSg9XDv1R85Bj1+3b0zKuzyHqzHKIvGewouM1Vn7QrIP
dBI8mLwHksX9a7SZMoDM1vPAYL7eipkkngwPtPufHsYj9Y6HVdDbpZ5S/HB9/iVMXNhgZgzUMLGb
OgAaax3ibp5JR0R7GUcLj5NrQfPDE0EF1HJGe+2fayFEwTnF5X/Uic7sNwxxRg04snVNK+2XzTjE
bITQVLXiV6Biro9F0t8uLyM/jRDa3PvagJMS+4MibwlxgCiMsJhqs9iVwSjeEbPrueAVTcBmCTYf
ByGLFOMfCRghwLCuccd9rpqxDnbsyf5rdFR5vj3FzwUTpM4AeqpUCO5uYx1BbIRhBCltov5w7/XW
4PXpEKwq6EsIA2xwYkT/wP06du00kZVKMfkadJxPdUwyNiD1C1ygLACcT89JQzTcnRcFTDcl1tE6
naF6dZbTz7vBiNImTx3LsYnhJWg3EhTMOLy/uCxHw7lJArHy2BmJi7vV7wLb1ogGcbbTNr3q8eSL
Zp95bzMqnHyMkLNr2ItjhUek/msw1KtSMQkMRXYWZ2tgdoD9qiG3S4FNTmPio6YqVqXSCbiSYhCk
kVsm60ZVlOfGetj9uDEPwoObpuwhXAwT58Q7vvDN1R58NmutT4J5rNtzl9wRVJJCnc+c30rkRq06
E+3MFUhztVKxPVk7CwoCqe4pUEew6+UYGB7rlR0zf0pV4sKaGLpZmRaFGuvE1lUUkyNjS+X11+eD
O9w6QaDO0i9rlisT17OMrDpFXyDT6nFeCnXYqkOGKal3XaNh/3P1+wsvI+uDk3IdTv5yLBfdkDB6
K5NtZc6AvVoJngRovookJxUoxklHaN5U/81pBArfUTTVdMJCzuyjw7LbhjPzIJrMaQxCzvNSxBZt
Vho8CNrLBtFEFoWN69q9dLZG3wZanxtR7B0IkcSBoT0ti2P2+oJw4IMxgeG1x9QSbuvcB1JkINy4
uwKX4zuriK0YMSf1vobYk7AMUN/KA1SUt4c06NTmCefdO+QFiofZUV7/qOM9C5p8NJkX2cUZOCWo
vB+IP6Q0UX5yjMv2TzJpW4+a7AtMjSh5cLQB/pBQ0uTBUkaVI0sTt8qTV8lKYvO1Y0p+axRUCChr
QzXcK7OeF0iZIS6bX5/AA9z93+ftH6VJtEa0sZ8ZzTzMaFQ1wqGhuJFSgMMaaze3oOBl2guCyG+I
+It8lk4KUkbVFxVx2dGDzUH1jojXCPPSEd4qn3L4wGYSlHNigjVKco1AcE3E7cVOYaCaxl5g6ehF
nNUv27i64w/QLG1opP2wzaLfowIN4Hg0W9uKuXYIgkg/A396GWAxsD68CQv5Qz5xF9dV/c+kYD3S
SzIZIcttN6Nt44wt6v40Wz3LTtgL0JB2z3KKrrod0QDGt5HD26HylItXWqCxNjZjNJOs+6Y1YJlv
vZp6XN9BB2aHK7H8isWD7jmAUqx0Pz5tQTtHD9I96jBmL6E1kjNamnwapvUe5d5VYgplfawSSo4F
kn8ww16FKZlRxedfohNkf71qGZdjzs4K6UaNPD2nfZNd6kXcu9oyGm8mnGgQGOXlYdE99eTwduJi
wvnn0OW2rHIlBFA9DtFczyLhhYIK8p3F4l7ycpnVLYIC/VoVlVxQo10Zxw0Lvurs9YZGh3etgDar
jZIs8Zu3zeBzDJsr+3JpHIQP4ACRzL+SDpvFPEg9udXA+SoVnwUUHmBB1fSfJVT4gyRbj1341ART
xoqBK9iVbh1sornJIS5JFsJlIlqurkwQeV+K0JYZvplqIR12jb7BxasD252l/jMixlXw19fp1BkP
EAFnMySaoH7QVKkH2eWZkIiG+RM88nYt4d0naYd5EJt2RYhk1PGbLBDIByMMgAGZAjBCW3LvnKnw
IRfec9gbWGH8ENKYKVZncZTkgSo6x8Q8F+hEKtrkpyI6ekjUaNzPbrPg8gYckQcbYmLnhtjS/O9D
Xb7tw80qtPFOZHaElJwmf2RuiwPIY+t1dx3k5DuIPmYIrdl24NQfjUiMnZYSujKymTY8sRof7L/W
jpKNTipz/SC/CnNAdO4sTd7JyBwu7h2GOQKHUx5yu+jNfasGqnKBZaoFxxOLsGsdKnMUdYVwmpPV
bcv5MYSy7HtVDZSZq127ZOcb3uTG+1iTQq2splwIXtUoux4EYtEZ+EkbkukJIsi8LMppK8b0Uj0R
s5YvuCvHJmJGiUOb2BX2z36TEf+/UB45vs1v58bO6MAYQ/dR8UTBgjk35zcuXYCLIHYNkJGON7uX
f1Vt7bBvdq8A4KFww1pEK1lka1+ymcdtwlVDUezalLTzADBFvy1pMcJJswaRfrZW4GjVUAkwn288
FyirawECR+ZwKjdaKhBqKQz+PpDdoR5sJ2UkofwcJ+7Ej7BzTgKD1DiPSUpW03MfyBfoRYdZp1X8
Ge58PagwuZR3/LWx3R3sDKXwfiljwAzgG2sT8Qq6oCz6PVG63zGs1VwgM/uoVtO8KUpBeRW1+9nN
5HeLB+PD1QCy8VJu9BUjaK2mGfFIyJh64iNXJVHKCPv39O4Rx5zMXWp8hK5AfIV8G0izH1RM7qr/
Sry6OE+cBGjgPELwcAotYwBHy/14D0Ea0LTEn99mmgAjRq4eMPZsBGaPJvHBiFQ5ySyHVJ6MzG7A
vh1LiUbv/lhWOxunsHLHuvbnrmQexpDxVKiVjhcNdkKWa8efFy47M/+8agR2KTxZQVy6kPpeiJsg
mbV0ZeYBDMPbEKmW9YoiQKIeCAw789MlpvapVhTzU0QdwJs4Up+XOZf3YcQ5CeoKOZlNokO6N4nY
ngA8zqzfZWA5jM9C6ypR5sxxr1jaK7QSU4bp/onGI6sNFhDSifWoGsKQzr5tvHE12kQbBURqHULN
bQwjJwkJ9Iyg3vRoUnkifSIVmIzyF1ZZ9PXV2dENXaUCYMawMsij0bIHHjR+FWZOyKN7x8DhGyH9
AeSrOVHs9sUAKsWmQEgl16sJHiszXti1DU/kpJ3JSnqCGPeMN0K7Xf1NqTFN0byCDHKcZKk9EW6c
N/KwTeC+LylCLQOLw+pnx4ZRA5OPmHW5KYFbkQnVYUgONwn6u3mGyVCkTsmsPhmWuhixkxvg9KNm
xth5UFu1h0FdX9pokgm8IVk3XHIz15cZI2lAc7xKwavXQzhTesK7wVocB6++6haQMwuNCRNPGepH
nVca1VpPqJYsytZYOVhPS5FGPOp7Dslir/dAABFlUTynjyTWARqHEd9ETD88g7UkE7Oj9O8zcszv
Zo4q5yLDBIZwFdLXod513jLtKYOh26ticoslTpUwM8/dnmM64LEf/X4K+NtMha9Ae6C3SjqBrIfS
NqTYj+u+OeUIumsWwOT9hiEOdy+24rZ85dcSoSR3/MRj9NTqDRjFLo9cEZIRWv92iNzzAhgc1SOZ
pMp5jLQha6lab1s1/V0XGq9mbBTb7VAySG6xoGOakCbBwEaBv7C2SrSp0HstRGOs2tlRZvrs+Zqv
kre+1PGmxnDzFyePiqSYkzMKgszZc4k56zEr8gk9X7dn+46xnOfESi+DA0Gngdz0L/R5p6/2Rxwg
OGofwhc8ZpLy1YHE4ZUNslkpsY1WLeLSmtpzerJ9G3AlxQWP3qKIGWtcxHklSRk7rk8Am9FZt0Be
eTZVqo67WFi/hiP9dAoEiadd368rCmH0g31sDKmy3SgHABwNJEe/4P5nkOlMEzh4uPlOf1QQoB/5
lr7ePZEdaOwJDiBFEehPWTcMF9wbJ17LTk1S4jzY7wXdyQbhRfu+lr5Ysk6tV8pk462TTweZpyFy
viAUxtuqe7Gl7pySjGt6AxTZh9u4y6o3HPj35gP+MLH03XCnxvGca5jCZcqrDHX5CKahhMkvSopu
Te/UslLprpLuEgBjDU6NCHHY3KOZxEuH1mBdwOceNY00/QUVOT5kfiWNeAoSixH54LbVgllY9jAy
pTE6ok2AEq649GZ0Y9f8e0XahguC+/kdvHgRKlXE7gbC8z8KOQogyUGATAPTlq0PY22lUXR5s9+I
52GiQ6/8H+5HIvdds60M0genr1QmWhStWfnjp6KGAzg6dNKq2GU9iI6H+qpJgzERa1vmBjzrfCcB
CZbm5LxCCMlfazSd4P6IJFM+4A0DpZxnR4qGenc8b13NOiYWmgwmUpWyQsEXiKG/xj4fYG4xcTfT
m/MEYlM/MWQR+Yk/gKylxJfD8wXOrTfGpRcSQwnvYkpcuewatUWdaKHsyK3sbqOq0KNnkBr1HLCK
LFYEjx/VRvncnVcInv/6KMouT2O+TWKLDnwLSjRro4oQGzO6wB9cnPSWmUFRzFw9kIA/lhNHabGF
PbwwBmnP+WmCXKTaB+HD7XcsLs2Rhj8fP+mO88JyO1yKQsQnaNg72harIrKcPltnJ5fIHsaZTcLW
wEZuTpdqamFVdjD0p6HdS6yqFTA/yIuKW18kw2k2+CYjBRbk8paHkMPiTgi9pTtvyOfr72+77HVf
i+rW2EA7P0gXCN2PekSt8n2ziO91vQKWnSp5X1m1CaK2iXIl8lulGE9JxG43bkmE9rP0smS34D5j
5srAjVHvOgMGosUZKJr+lL9vkW9G4WOxrdV0cdpAuDtKe89D87n1xY4VJTZVS2kLwHEXSD/ZRYSY
1G/P+qWyXhiU+XiteVN7fHMM5I13U1Tem1Vviu4XGxcHXaJXeBm1/g0Tj93ndpGFfHa+4GRJGw/q
tOKT8hJW4ndNUMNSpvi7ajd4nPv2qUUX9vo4zmFs/07annd2BniBnywva00Um0jNEcFwQKNoakdo
5UHkGyTQImh0d6Kga29Zi4nGvdqjauK7jes41d3EbnMu5E2nVCmkxf1X9ccqCEpXt/cF2lGvpvsR
xl3RM6pLj+r7869vXiz3W7BDcA3Q87vm6neqhOmtix9nrx0hrdfeJDIlg6/CKcvGEsSBFsaJERoZ
8nkkRAN6lIxleaN1n9w/YLdXWnb9i+MvzsEIantn/uuxM/w7ZjF/rFSKJKG1/JKs3dDZ0VKYT9cb
3wb2oKgJYJvGVzChIWEUv9eA3zX60vUzaE5WtUL4ci0es5i+dmPQT9fvcy5EvsfXrssG86IkOYW3
m+XO1ydMnYeievPCpaiIIngSUlmno31Iv3yPD1M5fL2H299Ot7yUShFywnLU6eqgzMG8SGjQZsrf
YpCEHwlPiJ+VzghS55qw2WR8SOH3L+NLubcCW58fh7rgrp801sSypBV9o79hQwj3u3KMBL9cZ9LG
gj5wk54oPUFXYn6KVjaI1GNfSpOUv+J3dTNBuGPCpWepmkvb6ElZrVS5eW1uo7T72h7k5+XcuMHx
2Thk2kKGWj0SHuIElX2J6zLwaKJDoAdF4Oxscow6r9r2RwZpaak9fvIYkcO2bIbWOUqiHcTfZp6I
3PkygwGXil9r4WzP/inx3c1WZdPkJ2XeZPebCrDd4eBncQHW7SEIETQMHA1LqcR8Jus6JATisNAv
4OTErfCyZxcwN1fiojDQK/3S19zZZbx09MYvTneO2Q1XDjl3NAbpybHe9LZFQrJwQcL4AQWAX+be
0196OMagtpOJrLV+pxzR1BuZTU+2VJ9+Rj/rSgZUncOowNZksXjr6ZFTmZFzUtyVBvrj/lDgdzuG
R9f+Psn6yNtdu8hskH4IUfRFpqXwXdToABYatjWWKAHaLwvlX1b73Jd+4ayKk8/JWrN/AWwyNEyj
ZLskMdIq1wjA/BaIhqDVNW3dO+SFHnj2LkGCC1pc0BHonjsFxxplIg31MOIcSuvVsdO7VjCm3UQX
8q8XDNrvhhmbZp5dRb9Uw1r+D8eQmwfEnh6f3ll81WNjw/dPLuDUZhZlEemGTiIzvBMO5PFSwE/F
Qq3W8Uu8b6my8actgX3byTOz76plu3yqfwgXEC7v+Y/orwSIOqbXNrUq19pMrffxcqThyRbfTS4q
0qfYQNV5+utr8E/6cghvHhdvMKgpru7J93ul42mhrScAJavGw3Mo2i38Q9o532Ywyu5tYiUEt4CD
AI1JlAzunFZufEM5twasPNmvW33mQPuVc9GTyW4BEzNmUs2Ocb/ozYiJNgib7+PzVYpEmKG0VFmb
ZavTiwwdYmpDvwXGvfAh9lpXoZmieUq3Mxh/W10PLLlPH2+A2+qMltpCFuX2ZhmxZnCcyIX/0kmD
WPcXFoHM8FCD0iPe5AeYvrg77O68H2pn1807UpxRHId3gLi5Qurj7MDbvUY55cpePzz5d2JeXTZu
zV17+RzWrEsB/BPnspovEWchMJ6A5Qb0/BfGnwH2P3ur0cimgwFOx2tUDEFsnMwzHGWkKNTDOoqm
dlAL/UNMmB3+xn5jhnTz8IhzwRFFXRu3Cqx5aSlM8tnkyPLekS4DnkTzKVlP61dofxmf82Ov/tTO
GuGwx+mXtaYnV4k0lQ1jTLvI63d1+s5qvrpUdjBXdBxImDzswNEj/tpg6WEUbJ6qwMMp6Q6caPry
uUF+kXIKpmW4vGss7/zSgWQlPrYzf0CvB+dmkHWHMqQU4Yazop43NONglPX422JADtcKCYjwz5HL
uRxvEnDw9LgHGZZWZdwLkgUH7HZ+Op6oMYa24UHc0xZbB+PKU39oYDUiu6R93Vlub67lo0reHJxH
XNQRvQbqBFRHHcl+oB/Mw0sgBbYT9o9p61vsmJY/h8csSmrS2plXqMTzI7P+TlYfdLy47/hh1bPV
xAqffeDyHxW1Lo3NPwbP87mHn5ihpc9JYxncG54fX+1ir2w1BgfRSCOF7+Xfbdpmi68LKfKaOkPg
DE4IIDa8l9aL/f4VxBIz80TqtmMRwpYLx1SB3cIytLQsSIc+/Xd7QEFYnWBGdxONWN7ZxfXSlNeb
oGvgjDdSUQ9UpfZQJoS0usLRRQp4uYTLBcaXJexxQzrG6Ynkvkrd0+NAvuDwiiVxGVqrDwK8SF8O
6eXVz+oyN/qaoBzfxHIEZyQqTCHFi0blhC/1g4anH+efvYM4xRuFpGds6NjUO3sfTKkCa34FYqCe
LFlxaaHNpxmRlS0W2qbP+4psWD9CmTOR6oVc84gt+SFrstMLDOSjOYiahhpLTEOM3A4OPpUweJBQ
tXyYvPGA+ZYHywTxfgzcZGJ4vAR5jjpoblIzH1Wnvvn6Z50bo+2oWeifD6lZalUBVpSmgOTFgG9L
XH6NZHmAsDSPB8V0ikGos+Fgc5IpxyGIeSbUhMZ/wLe8o4ZfypORZERqsLwD0KecRz13H6rmDF+d
9WcFt9A0NGD3c+20/LNFlOANYxHAppCt+cOsnpFEaO5O6oZ82zGMM4Y65uLCmgV9G32KZ/yDW5cr
wJ7I242loLRKf++d4O8gkgR2bZNfjIdmmOaym7+vl690UxF9nGBfrtTyeVTwrEw5jWZx9cfcruxZ
mrQEw2WKEjpHehP8UD9TCy9eczq7CYEZKcI5ps8dYcXxhfAfuxzeXOeAP7d4VENa4hYPh7J1gF8q
hG+2PLvrTSRRRM/GMY3z5NqBUGyovLgjIe4uG3iDvSVcnQgCT3vkjch/z3JCokON6ijUKwhZFYVV
PDGC7dmPzVwz7RUg4WdR4B3TuBeI7rtxodZvUneWpJmFt+oqR74OlHYxHmhQAqNlPoq7HSxX0sa8
NdnidIn/RUp8t/1wcocE73BGOaU/EnAhtQdtN2FIh53+XPwTktXS0QVwJiA1LQLcpWakG0NAqQFN
OHjeky9bFEwpyGLzp3uT2TrVTO5FPgDoddoJ26Ib25MkSTch9H85QY8WYxuqGYJJStnEmprS5Y0i
KVpQ1w8gte5kwmVqtSBeYFVkOUigJb5Zefko7kEohUdryAq5HTQrxJBt9bX1r1Y8n9+vAFaXAUUL
QvMzbti7u+4O4/qIgPIK42QOAQTSkdTCbYMxqsNpcbNljLA0K+W9KBVuodb6DQSfpEuvS7Gfuw/S
a5qPeyPanYsHDDAqdRqr1Df5zv+8zrM0xgl63JWt9e463OXXpvh8S726Y00V/Nms1CVP5dUVtbyb
VYPGtDZSwRokrJiBwIrP1RlTplnibyYaCbOTzAIgWV25Xe+98hqYzC3/GVbglibzQPpsZJIieBF3
hXYIcB89vkFkb5iNhNoo0gN/E0q+Zl55tdl/QhKoxbCs79SZUq4RPiyutUgabjahTLlreoFGPeL4
9lNyt7K8bn8d7GmrpVZfsomK8MWvjuaja/E056iubNCmAB4XbRfF99MDAtYrkwK9x+Z+VJqU9BT2
YLBGl23KbHshKpIzW+ubdrK1uq3dMoph5xximnGxsW1PzyzPVnh9GEqR0fG4XdHu+tguVpE+aVyx
4w5IGxDmXnvOqvEx5SB+n6AqPuonD+W3Wvj0zx94EoviJr+aEiehSzKOeA+rjWQHNs3Dnr5Zs/8N
EiYve0ubDm4+C0McbdENyshyOacFGyO4KsghyeaO7pL2Ya/1J6eYilXhIa/7bTyzw2zLM2w3zFSN
/cGFIqLFEzJ/eGbG/XucyN3Qh3GdhE/7bbd/PXgxMKkdp2p2n5EtyZ1BiFBOYAZondCJ5jvoo+JY
5/QqAZLYMYHRBjIjYDscQcrT/ZInQ4QZp02BdLcY5Mn6zNx2M/SnpDcy3S9QTigcyhnQrtFpr6vR
kri2GaByqiZYg35l0AwShRFnwyNvRPJIOmuKpo2m8ak+AiCGLcyKmyV45iQk8jpS2yoFZXv1YHBf
/9OfFRlSQIv7NbxFhteQfIOI1As6F3vPAyCVk60il/zNXozgUFCluFyawUiX7T551v5m1k2CJ4VU
QAckJxAskYw95NgkwojXS0ZgBP+cqWUJ7qWPBjhblfGdCoP+sUgICZlzKw4FCTvZBIu/ftytZQOB
4NxEAhpCjMpuyYNNk7yKeZibl0Am4RPvuboD31h+cHbFSfhv9CPn4KXss6H5xuVAVhN+/f3/7KD9
4cylmD1uErzJGTltUXMCQhsU2HvF9Q6TDr1awOu+RmOP4KfmO2W0EdP9lQ1jm/0YfTqhFPzszIPI
et34wOljJ+lOc/ndWHTVqTR/IIouK/TjiikMroBluwNwD1salQzKoGzlzgX/+T2pmZY4/nL9rWAe
kNxQJY9+0N/1gKm7/lZbOvrV+rOQ5CYMFlhfUHEfw07yFBeCgvGVTnzcZ1MenB1FHGsf6D7r2oDc
gtC0QtMlnBNuZYbhM8Ms3Wm0apVL6PTg9ok8BJ1JWhEaU6bNz3dXpxZUaMweuYjMn11dG/KTGwMd
n6aOCsfh3CCHr6F+aqKKeY3BA7MpIL204JNobmDfeFQEBvpQITWRt0GtcRIvkqgfWQIWQTBFcA2t
BLJ0aKuLLWhDmiKuKzYbiTLNeDvu9BWVed+O2fOXfmjwB6kFyYYVjYDj8X6ynNmCih++k9vmQcn5
7+n4VpfYv1C29KoJ5AkAPyA2RZfltw6umUC3k9N7ZENVxaYhPQmbxTNB/+ELVgLzozKD8ss9IWLH
YHxWmwN3+Uk7OyVbc58R6c35iz7tzuSBPDlfu4mbTZdXIMoGcFnzhMT4u9BiVL8cuUaPygA6ykDp
54MjEE0y/Mj8jJJI6u7aLWFnqTUDQIds3q45grms38HdH+QctBOgXfMkr1yCkzedQhygmZW0e+Gm
poFDhMyiAhCJSfgONyvqOlgpu/QFGyOdvGlvi7yDzNUxSCvwi01opy90aTjl5vnB7y/cnOTCKk7g
2cAb3OMHx1G6bY/Vj4R8/zeRNoft43rQAMfsbP/6XczO/2YqzvfJ6Duh/oWqbJBDE4itYpqUXPQj
1xKMR/mwG7XUiq7u81aTsh9iwcuPdFyFs0HA0rtYauKGdVgkpQ0PooHSsa7TQAwWkyOkXZmvkkjH
8mwXjFAJmUOfRg5u5L9KIAho1N5EEdp7nSazhdYLK5+BoEogB1bhLHA6D+rPgppKoKixLM0T9Mjp
gKdQiaJ/Bt977moPRqPsQ4NlphbHqCuu2e+OyUbKkE6PsC4UPOV/+BewStWD5/YX6sdiPX/Xgvv9
rhw6wngH0Kc2Jljpyfv6IMgbfXMDlWc7Axe8AgwaiAzFl5N0qQTRCz0a4lJswI379qqL25uFYBzQ
y/EkNwzx9QqcV8zOwZyThL+IsKm2CD8+Bo7fyolZ8q+8tOcB9x9YrVoh1fGjPeZ0qZ39VHjF2nUU
e48qLgBohM98kX0TLzib0KA/47x92bVuhiIqUeabOxgHPbEpuz0Kosc/Z9xM3wK5HpBSlvXjOIBp
5uZUVrdmnVfzIg4j1kReZmpGLxvE4rCCMH5j88YHDcfcqWSIglrT3u3dAKFgO/T2yHe8MpamzMgk
ykMG8oLed/4DJjIO7as5Y/md5VpcjeU6drCC/QrMJgcCx21nkOZvhuCkIViyaOm5g6rzx98me7bl
+3FK5aRT+fxSSvSuoeQ2SW6sh4RUsC7xI9tE3SkB1G9sCRZQWbvIALcpYIohrIf+4q1IGmmKWelA
eXd/MYkvmh8c9nH4818y3BalD+WFR4ePvp51u/Z1Rnlp9/ZKSUtvmflqgIiNO3rPd7Ka+rtCpnJ1
Mib/Rgc8j6KClJPPz59odgGanezA6VQV7d5zZlzDFIR3SXur6BBx8Qcoiqo6kNNokthWQFQHXfff
NUluen6Fzf9kWpp80yW3f/7uLgkdOdsGSXJ362B02t12lBg7iuZv3qQfSn5rWsfH9eM6+UsarnGn
YKJjqRPDS1fYPl4Pz8bWmx42rWuE19RU2gHdfxPyVpyl6M7s1Wvf4lcCqyOPmKl49xJf4/o+5Oad
Wn/ZC5btvTZ0TT6+tm02aspc8Fw/EjIjSj3Nf8fXAt3haJoEL2uU5HweFkHdkP+XN98zs4DrgbY2
CwaDgQSzgClTKu45KIOQg333L+gYXOlTHTirUOrpfCLDVssrRkTHgOi2VOFCM8hymK/p1x1b6msN
N9uQW7oeerpjxwAAcE0aSl4qG68YVZsjwPa2aUeZ9Pn98KpfukiZJvq1CXctdmPz8z5Knj3Wz2yO
WGV5lzwckYFwxgbNNvlSZ4stxp6PMco6MBIWS8/X3HP7TGbOb+5+JWs5IfUYyEB1K/qodbqDqT8E
B21DjGYtJUhHB6Zst5MxQnbjHGjdxc+4fqmTeDULuT03XLDcdIRR9KJ30fKMeOFsTnLdqwBTyWO7
jy8B7SEZKtDjLDQxeygtwHf4ONqYdaBaU6V1uQ2X4M6aTIJuUYDiTRCHscsmL89vftAT8qPQivrG
+13/awRCoZuD/3GI/x1xOVtA//6xHYv/s4wD4ss2mdoZD+FD7hgD0lBDPaINAGEsw0knFG0+zp9J
rDo1YVeq7rlFhmDNG2O5ikwzJ9t7hr+rxnC4Im+GTpHQqfA3JmxWJD8JGGqLfeds/7EXOnYWNt1y
yzW2MvM2tFeb2/C8F93qPa7N6fZc/7ROWGWp20Sa/klRqVLC16TvcJFf72IHdoWf/Z+Tc7uO94Rf
qCQl3cSScBmjD7D+qghtEjHFb/CN9wIvLj6S75UNkZIPR8V0oqYQpmok4LOgDvj4xgAjuP64Fn9C
Od1H0pzTN3dJxsXg5ZGCKe7a/azQ3qucSka6BKScmFrbJaZXZsuwFJicxo5D76BtBjqi4/7qf292
PD39SSCwLsDGqkG7HZr/J67JnmfIdzcWW9Krhs6f6X9f8yPSkSnJ5xM85wQ+Z+qot7+q2Ey6/a19
YtweQyp8lhhKRuQcPBh37CXnQJJ5+7nbyuSf8AQk82VMEQJLep7VzvehV/ELEK28DmLfpFO7Nvt4
l2C1q0cCiRqdfXEMzKOADADnj8ktOdC4qbMixPNu9WHYuvMpeh8qtct2QSxNZ81BI10+ySXBSdqL
0drlN96Rg3MFmjHBeeXf6als667FJmNHcqOCBizpXON172dyAS075e7ph0LTuRXy++dtm3y50A0l
3qUJ4XirkZQLYxn87vinRFyy2E3VDNndpD8yL1WMVtXuOmuHKIVS+kmvtgAzTcGC9WcieYj3UcO8
Khkryx4bEh4eeQR6iEmHQeADhJm7Gw46IRhZ5P9iS3sx9xXyTUmb+iXiw2raPWBzdN+uVZeMe+He
JKJTkD3V2zEjAxfkY2ExPFxxZc+d9MGSjP0JAnshXFeyAm1t0+4AsGPH8XTrhgKbH2nImVbJTMDQ
clHbtMasEo0q7J4YWGV7H18A9/XG7Aeu9FIokmxoHbIRuQrp04x16k9emnjx7T79NjRtSsdKHuBl
eXI+Ebt2XIX99szbc7Pro707ib2SAL974HLt3xIXvQL50MlGN+sSr7e6h7ilCjremieDiCbMNCUV
bYJlh/ztrlChNb8KP5Qi3R40xAfoMotGsuOKOSizp8w57eoVAiqpb+qbGJZBxEJLzSJ4UhG/Tmv5
YRZ66IEAYUQPeSrSE//AUsz9p8sUMB/iRtpjQF6cqVGwpttKfAF21mUTo+Pogj4oze4vZdcjRUHZ
9NS3Sv4hkNYIMjHEyM8411xFmXVUxqKRH/K4aWVRhF+haPDsUSlCfk5tGdbYO9GfF2rPsYCkkIsF
VWsXtaDzJ83xE7cIZw1Sc/1La5bb5S3xa3JRameyzFi4tQwWbOALjPJzZ8xTC9pKfETQB5bWZYpH
HmF+nfUTgIQRYWvOjq+2J/LRKKW6B4yTzymjBK2Y5D4rMyIV1XgfauXPMWHXpMk/GMLbnFKyH2Yd
8713sNgFAlBgyJKH9CHkIQmxZyo0DxLhZHY+OHHXbWi8MMstPKecsjY5iWdnKtMGZHd75RgBn/f4
QE2tWqMgtUvSWJguj7TbJg8Uzwob5IV1OUV8xKHtMaeBQpSOX3aeXqfN2o30CJ2SHo7x0LEh64Nw
pbgetzooz53tKn8wbvA+lWodvm0fl7PCJtJV413eUmh8locONCNUJPExEuYucu4S9y+S7Obo6ydo
HgLFtcJPmA/cAwgW8vih2aBMY5M3o+fZu6sIytmgThrnmfuzzXZrFmSbNJkVMHN+TY0A/ryJ/1g4
mIFvXj1zMCYzECbZEWr94fTp2CCLAgfBKcrqnj0Z3Vg/HmGvNVyfofoI4ITDFviyS2TGSQGHC2+g
Ru54Wh6UUdn2ySIR6BuP2eS5jRSDpY/WKP0bDQONXY5HfKqoXnfU+SSOSoHsLgKxcly6y10K7+vc
FMzo7UWkk2G+ItdO2Y30JS4nXKSKNpsqNzD90ra5BHF+tpUzFpAcrl+D4FISb+CPTu/D9GZyjq6M
zys/DRMr7uthoTVKjvJj9PDhwGf8TClUWlnx0jzXq9McH8/Tt7ZTfdTjcyfYiV7KdyV1637hA0G6
ttdpJiht14XZ030Q0QvgsAe79S1D+nkVnv8LDN+wUJ6SbU/tCO43DKaeEZI0utldFRi3076p3YpW
3BAKhJf/Lmedzy53UnYB6LKsOh+Rrdqrg+ixbDR9XetXt7044oz/Du4iwPfTwQ19c96Af3PkkQ1l
KcHbGEs+3SEuRr6sxiXz1u4NWtj6Ppf52DdTdcpeLrG6CX+RJux23HhHE4LuQRb5MJVJ+sPRHZlJ
jgC7kWne6xURe6ui32zMx+JOhU5T8uvcZm/JAgiukAG0bvPCNPqhzjcb0XZcOWAzqQRtaHUJXFzA
aI5UQmY/+UGwuwjYDYUfvt9AjFe9Ugjlo+/74IUSBMrEZ1XAlcB1+bROkMOALbmgIcwItyNAVB5z
lKjCNP/s8RuyMzU1i4obn7g1sv4X3/c24EYvWRSQZ6Wqsk5h1RVa7HuYYr3tVwCE/UPUcX57cBny
LIe2vO70UpXwSmaM/715uP+vMFzrT8UmLGwiaLj5KMPxs6qluVfOdYhV1bAK/pBQYMH9mHeQcgd5
xJRV03RgXnwpy8Kyv2vQLFe9q24DmBTUbZ6S/woA/YnquCow16G1UtQd7jQEwfjgIJjD9F2gDjac
TLm3bNs6lqdGIEKyp90FRInUHXeJuGfEjKIr9KteFR8X/9v9bq7dyquxO91zUsg9pTfinhhC0YED
spRde8FgK4Zt2N75Lv2/hHHR84UosET+CP2QlN2zuVGTdjhURYudwwSUVr64620IEeQN4E+qz2vE
raZCuJn0hIVp8pj2gd/ZfEVGyc91Qc8cSv7aIHh6DoL8Q0cw/OYS+S8eSHTPkZYjky7tFjlQhrDM
1J0kVjvogsDXZDsUR/HS0TJSKyyqNCln66xAbkPkuYUjzjwlZo40G98hq6RtXfJc41sGpDuXYQKp
dxhm0mYnYQB+tNddlWQVAjLQ2/EKLb+l8V6HgEq3a58A9Rq+wv0nProB43i1zF8sQStK85pkTIh1
GVV7OgrjYXrLPl7qqAIv0ZIVzPumoAPYWwX+QS09GNKMLy0rg5vOWvGiWKjYFg1wqyH2W9DDqu9W
gHKqQtDTUr5aJTzNdDwbmQMP7OCGBMRq43H69KLadWPmC/sx/aPw9XolroGDeW9fY6oDG3y5jHap
TGxf5lmhJ2XV6EC33zEWexMm8JD4iJDDlwgog6iAOTM8YYDurqVjuiTdPldVH3BxFcSbdA9+jOSj
25Sd4qmgvylmWb1sn7gOte3oRabnbmc+ZQGgfnssTNAnOAlLpjDaflv2wa2sUMgmjRuoo9sVvIAa
SDvMXQlEzAP2gGbSxFhKroTbyTPy1N1UXUJVHcGK5Rs3VhISCR4YFFlbujLPHs+v0NbRllSg5cG+
F9rg+ws/SXUGr6AXpy3wx/udH+1/rP0LOcPN9rH4rIhHaZLQ4hltAjFHe3L1cNQ0vsHDq7hVmp8D
IkNYCY1i+eQgSd0sO+w1HTzfIlyJwu5kOybYh63Zu4dyDYgOI3LWD+kmhuQGLK6chRIInBbDS99Z
uFvOuYyZkL78oQNIOFf2I86gu6RzjEP6BrJKbLRkS57v4ks7sV4wKecamtCKSusESNrHSXo7wt+W
QAvTyii+SV7pFkVDxhmnWiqKGbfWHf7ltCgBJe98OPAAewZ7jEOLHTW/uVg5IVTrBPpwkRcD+D26
NKPHc7Xc10Xc4lydEkS8wzJgnHDNOb70jVxDY2Dv/2z3qWlwDahxVg+dUbJpK8fh9WZBBMbrOB8c
xpTpOv/dqfC4271JFJT1iSWJUkZm/OAqYCaHlvxJ0Ib1s0os1/Y63MF+wfqQsFBIWhlsIPnnasw1
vxyWcN5lIUKosBHjlDWgjIa313tcTEjajqqjy2EtsdkW0nQS3pO3Atro4XYcZqM5uSxyhX98FAml
pwKVXSgXYEsPXi0BPJoFirSMp+ZYsQwer85L+VySL2NNpCjRtFZW8VXS8EB1ROv7fV1OnPAZAcPZ
+iCZLI0wo6Q3GksvkQVXzemzyQFXxybWRewDrMMwgEdXwIbwgu2n9Wn9BLvQGPlNMEbJrSpl3F4W
LNDZNYStEEoDfM7CY/u0QQmwewFMsrbnrVzZEYhzeiPz4bT5kJ6rM3M62L0PHCz6d1KmPb/Ruyz0
In1gE2NP/6FMuks7/950lcVxj824CybB3nvPs7W40AwEFGBhdZ7LX0KYQdQprB12tbBcy8trf9nc
E5F2xFk6OY2n3bVBpSYuYn12Ho8+ai6seQS9+M+pzOL/e3Br9P5awhMhQu3hE3XZWWY2LYLX9Qvs
s2OmMMOs1tAYASgtO2OxgrbtR+3wzb/OO+Ea+nscdtYdlzA6VeM+2Xv1SD7CQIPbE7UYWfGM2Bdz
AfPGBEGuSLkocMAjrqAfXl4lHos8sICyWzzebFbuVam6Dgs30Z3PCxtwinE9phf6jqFI6RVSWKHV
QeiKHz/u6bRSuu7w1e26b3p6DlEzmPEIYwOUMor1sKZkNblsuJ+riM6uMsEgNR7w9IpFiLpJ3dGH
9fSd5AJOnDrVAlcMoh7ZgoDyZAWAJQGd3nc0wh9XnmJ2P76Z1IoAw5sWGqPLnrROwtOFk3sGjKXY
bgNLG4vKffNf7FkkW1e4UY0EcD5fzST00iFsc2t8GgAFclDVRSb+svBQaIh0tCvJBQJxXDCt6uMO
cmDlR+IJoBHt+ctJw7bpL8v64uW8SlWRCIWQ9rFL/OETHp+WK8qy09j0aeXiUrF4kYloNFXJbegP
Bs78xy2QDMQUELPJHCDamLEYCFEDVFDTolTPwdq4djEqTkVFTA980zatuOIgzguMe8aNH5X5meQe
JZJcShSraE8pUGzNJzINUgxt0WAa9ByyzYNH+OUEMYyKBSflP0+1hmB0AKk72on6OrcHn19706FA
FXnZCs1HGbDtKgFDyNd/XPAFAKUuGTDyaRoErpXHpwuHgMRkRCPjOKp8dCmyJABasiBKEESP4Bj5
rI2eOEmygPVEjjq6dOQwOZZ4tK8qv5eQXyqUl2eaIjFIv+E+nx+PxCWlMsJkOpTqp+81nOa0B5K2
FdyIZorF1EA7dZnY63qjC8zEwxAXggxqZgpDmUGOelva7KhlpfY1ilOx9t7/Y56zXIoCaJzbFej4
sF5tOgtB4ru5WS42FTUJGrFZviNZNZkhY6OnLi+07Rxhx01fa/W25kcM1CWDUSVGPZU+2DZle4Qb
wlfqZ5AkL9TTZlHIo8ZVbL64FS0O3D4BxXBcw2kpitWzquMqabm8hf/+Qk5cRwahj1dqb7v8k0gg
rDNWaNCFtVYqtDZX+Ai1ApVtZJFlgV4ZPH5wZwN2V9oVxtZx3MJ9bN+ioMePZGP+GdoJ+XxhGxT6
eFHxqhiNX97PTZa35oF6YFt5nY4zaHvmvkZwNN4o9aL9lcgNqo7EGikJ1LAPot22XlQR6djLGUVY
odYVIniKHZ9gDuUu/rgAoxS3oVFb0UH/oYnc5RASVv158zy3O08tT3i3kHQxWGWKDM3Ep6waruav
fhQYnhtJXj2V3fmIhURj4McpU5Y++z2RRV3UWEhikT/j4ESbydWJ7vTngM84LOTcK7eNxvoClkSe
MCS5ITJTAwFbt+jDptA1RQ7qDI+7RnRwIY1r+DEV48sKIkb9d/ezCPaZubw2G36yKxjyUpos27Sb
YjXFFl8IeG5pgNnDDHN6De4vQedDDa9ye14z/mnTsOZrqQeMYjEUWU/GKj7NkSy9mqo1i+V+EsEa
W7HEw78w3INssEGkQDIhf2t1EATavBvggPoAWegSolLtUHHU46yu/+R6XOdwxJ+qFhAwgtvK8Pzm
zGYB3GQsPyJtMVR3isGQRDhppotMhpjzVLgTgK3zwYuMjZq9FpM0GyIsuVOwkzvcUUVFXww59FMo
zhnzoSiBdw1IxCzaHybKrLxMZ/x0WNQ5ZKi1CFrcNMWS/Gg0kYjLZbXjpdO3O2SXrLNVi9TmquL8
It4P5DKe6drYNocUPQxlqC7VSbDvdfc8KKVeE0p8yr/XvW5SSFlEb+D9TyvxaqL8AfFh5UzDjXYl
eQA82mYNih1F9WIFGOoT2FMvpEOSWQj1O85lvRVqw6ALy/EJFjOvR7Ew8TLo+HgMABNAb8IsuPoD
GxDlHDQVHogKD/9FKjFt6krTXbeEtEsXPX01tqPMSDhZ7G9alVUk0rxSj9Tpp+ZM5SKuOWqXhlDK
QTxLDa1T7dCEfAcOmHc/6Y0ZRVPA/jjwhI34k3PJoW0wQQiNmyCgMEjlBRIz0W8dqb/NXJH+3uBf
NGyMxD2ZQSwnNZTTnFL0vA3YmX1H9Q2SnWBBsNgxUbg0mRTOcrdSifBoj/yP8YX1uNz3tjoUfB2W
ttAk9zhU7FA48NV1ZzksEBMfJSIcd/0g22eIYtnz1mt0D19VjQoVH9Cvz2sSZinh2C9vd9W6P954
oKTwC9VSrY9Ag21vKbj0Bu66TPDspSsJW56KSmKAsJ0yKtUI7l15oxzoGRqwrRFV3ivCNYpqTZqo
rfFClCvD58Pm81/7i0gT7FZKFXgnfCtnPlg0qNzCtfQleSAQCFW9GuZkwXziYpP+yCyt+PixFEPI
AfxJTVsGavybcpfXSQA2yyN7whrjrD0pyMfMhH7Nj4REa7u6IoXwJ9C/Z2EAcZ316XzrTmdBNWV+
+Ab7+hcgYy+v/m8jtPR++1xnth57KBDqu7M6KsmIPHqULbAlnVMWGlZpMiYDL3c9WdwVUT0T5K5H
TdPOVWKhCueBVtdOMm9D57EdxXLTr3qyZnRGDLwCus6eJ0QaqzAQHpUb+fbf+ccV3ytlJXMkNaVC
6if/VfEM3sRQfTxDPlopBdaejXpxwIUfd3wmIkwcIoDN8YDW5SeE4tCXOjpATI65IAGYxZ1PlXjH
l3ZH2x4cRQPAm5aut2e1cvc03OIA4K7H3M+R02TMsGfH4kY7wZWQThXP1pd/q+AyCAce9c9BzPDA
K4peFoBsgnsGlRb0TLdEMl6VaD3EO9TjzimwE6lSNCMoBQW8SRAycivR3cHw2TGbLi/+k90F52CD
l3L+F4piZtH6IAJSXiVul6RXurvyiV63BcZE6F6xaPxqB3u0w5c0XOsW2qZyCCqtpY4BxSpG5naK
RRSb4DlwJlXPG+iQ8//toR0QXdk+2mnnWlFyvtvOvcM0QSyIgLNm7400G6hdE1bNdo7zuOYOOV8h
d0vIlhj/b472gkZ8kemmtJ+Xzli1CIzsiCH04cKtRHbUQl+AS9u9JpsyCPd04j40oSH9vo7Yh9sW
tRouEaIQbaJUn7ixfFm/H+l1yzJjhrPt+WXoMhA8cIKP2c/upo4oVzjSs18oqbIs0p0hBU6Q6XUm
2XCnuXA5aKOBS7AX3HtOrsdkkVi0pA9U9bLJ0YlzX1SW0wmk2xPzZOAvKwKMC+uvsW7hZBemF0aB
oauFieiXV3kmZgm1u1GO/PMV2hH5nSwvK+WnAopfirfKUnaJKviqDDQ2vnJJsSW1sd5UlM3LeYox
y9tAvDAaWYj8LpOmCKiXdU9tFeoaE9TnQAv9mxek29IyCV37PLymq0W9zOFBF7V0Vz++tAHf8Sg8
cQ9Ba5przgcUXu2L/WB1EoXz7ZM2e+jW19O8yTKl0iWRlNm/DftRda/eLRVZVK4hEilmxlT8trTz
eZk2HBCMq73krGlohhX+Ms/QFP3/txiGr03wI7LSARxAEUNNEReCs0mG2ZYmpTJaYwoAj75nsJj9
WJIZ5nueRgxb7frQcfUVoPJpv6HiyC4OuKFkAcqYwn0TEPzMVfSud/Bi+Y9s1eVLc6X/YvVDLkQS
1agVM8vw7GAT66/RqWfkM7Dn9T8uFsniDFwLOLI6AcxiYoYaDmXsgsmlyzGKL0sDf0IwsRGvvltm
GxDueGHvRgXGTts/nEGZHOnI658io4YRhObIS8Gw0DkgNwsuqzalMAdjvSmw0kSY6U4MQHlrmfFA
B8zGvIPspz0+9heA5DuZzd0Nw5H9Sn9HoXD3omtLVreKqyFK5NpgNnDO30rnz4RdXYw2a8fkq5dC
0BIP6ydHDcxGSIliy/oBPKeVP7VD78BXnt0bf4xkbBP4pAo0gcDZ6oC8ai5tnkgwpjU6SfFuy44F
1S276i63Y03WYkgbQ+2HVk3fY08N6ntkQDGoyilyOAjYk7NWTINlSSuaCgb3xyNRmEg8ocuJaqhq
26KtN9kFudE6Qwuc1bgpzMg5pqT29KZhXKFzkdsXXnp1r4zzDMYL4h+nmvxJFooqIkL99iF9IOnb
sWEgENpwoA4BmJcikFLCKZH+w7MlFqRnsXMrTzGhKvUGobJuMfDUFVtxr+ik7MSLcoatVxW5Niia
BzuSTHY+bXN8Z3NLDlbH4L9m7mFEzT/WsrdXK3cJta1lvYApx2B8T2n92YWrqo8Bt8IVvxrfAKY+
a1O/9oWF7krJ9RGHFjumc3gqZnOkyhh0XO3z6IRph3jWfASOC2BhLzMbO6z4515uyCninO0pDqge
Mu5tVYm7FYgO26VH/wDoGJ2Ux3Gu4dqeG2hYa4XCCIczNiNpcUza1Dcj4Eiw89z+H+PjkVOuWlCo
rACq/6QaL3ErNd1ZIriurvGuwwB+xSwGj8mXQ/LUr8hCy1WFKHwOeoVN/ZhQ1kP+6LJk49bg0yeg
//5O2Z7XkG43TPLJQ3Ha+MgFcF89snGC4IzhZvWV6kz8zPebOwAmIrKTa5w5t8eWHi48Z3ytkouP
ZduNYpHGhSHRvHZiTeD7vC6YgcGVhqxhhTyjhJ8thqBjwtJBga+fLYKsiMOXQpL1QdfckqwGc1eh
eQ4m4gtBr+wm4RbYeIEJh8pj6ZSacuMamsLD9NsoPsuv+fBDvU9XHklL2E9WsmPsyv9PXZ7KESit
jDPKX07sjyE2AnqEWcSqbkR6oh8xZta4vmdTV0lE4bMTOBs7N2ozIynnpWuKDwmQQrbloyWhV561
hf914/KuuOCuXc+Wuu8lZSC8lLm2tqyxrOOkJ2tCFOTcY0sFZB02tZQ9QIos9J/RQy/MyB+U0i00
jTAj7CzPTygTOTTDDjcmb3V88AEsf2eMLh07q+ZlV/gSD6icMzk//sdv71gaP+O5ETy2/wFpdlK8
1Ry+IU75mR5YouqmmfX+QxMo4jQa4tsir0wczpAyJ6a/Al6MG3f704bmA/2TL/PF9H8qnCY9hm7A
vK8MV538WlYg2HwOsCbIhBVwcCLM4LUtLQA4og324A/qoZmJQn20UGPZdxnwEz3Cs2+kfq0VBEtw
TbZyPbzwpGmzguNFiA6daDcC74JfftDmDiIA2zIasw+JQxV7msNEebSl6tHKtOYVLaQcZ3/TwN4T
MGm+5H8yM8wgcluVwMabRzrUBykDAf61C/0Oh+Jk58IKckAhgoenzZPmnNQaLqeOgRVr6Um7AtWQ
FkO7RJi60rQsCvK9uYVCnXBHNms6TptoFMVn09oxq9ln6K4/lV2s/EjdbQXlj7Q2pUd8l560+N+R
3A91y9mD4OSI2w7JMfL3YeVXpmkXWFYEBsvD/eMuDCNY5/Ac+WHcCqELyuffOKL2eqgZlRBQ/EkX
h1Fqhgo7arnTeJD0XdIHO3AJ1O7PxIz41sYcDMv6XuEXE8Xv9Jm+m5ii4To8vCXavGJcMGWyJsFx
UzntkUEsEm8Z7CdymK7pGztAJXpgQVSGjacMIhITJSwVHlwLzf8JKpv584fcr2fzEuP3INQrKrHU
spNJLFl3sSRrVbF+/lZBFHfBDfU7RsYfWKcFuy+zgAUnL2mRGi7OC34cydp8cAPcCuxZUaM8kHGR
jDWfWtBnPvxd11+HhOHBLr821FOnf5J/SzMcvkdKI3JAaSR+zOQ+fMBytu/d3/CdwuqM2YMtB6bx
m4XmtmBfgsy5gpPtq7Z8uSTV3HoeaxWm6hTtPC5Ojc38wv59F4xa8fhRQJGtsTL3qqw0m8+JffxN
whHS4TqTFsFKoHUcp5lRAuIkRV//zgpP2eigIlxJH3RYjslB5cAhQSWBR3yESokehRVtsegQHfXt
NRG4fqBv8KKec9IgS0AT6Qi851yURQpvzAnU1/XQ2TQss5IncDXA65hHgx7kzOFiYHt5aba8KsJ3
Nj0cZ2wedxSvbIkcEsxhgNyeUWYgWxBXWxNnc/pZYLl086q8sls2POWAjZSnyoFdVwya4JnMkKLB
0a9CtRtyYl47Ef9Cu3Pn+XhBNB5TI8YmaPL55b5/nsJLv+ZVQnlpRbugeNRs9AlKZcsgFHXRQJlR
7grLWNYhyhx7FzHum3HjHi7m1J4wapW2pf9QS8wyaFOIYB7y0d5n2ZBiO1EH4lXnOuohSuLKqixY
CvG0e6H1dc0052Z9BB+2fL/aCU9FSMB+YMGAWLnzm4Q/9bTTK9rQbL1tGBMUDqJ5S1ivWIdORVBc
vFcr+e+00uzToh5AE1gZ3Z6xITLTE9cYIrbjo7px3Pi4z+RN8K/qz/ZRlwOVXsTTj/fEGZH3Vt4m
bYAcj44KTOGSKe1WPwxNwuVVO971sI27tazOpY4wxGTnLPjQHbZ4NJFvGtgFMRQ1XRbwTggy3X8l
CAcYSgKsohTRfTqC0Wj+4xW8pziSaO/1Jygxusk3pwRDM/V6NSFuEhUXcTrg/v78n+xBIhdYIR3W
aV8ZnhYOrAqwLsZOP7tkAf5DbUqrnX/I9nGEXv6WaWKCoyQysyvkyeZHaMciNbZsMZlmdXnXh0Pp
06m8xmcdA3+GzTLIVakYJBIuliwz7nDGph2s2/PwffR9wMrCoCLoLRMuEHn8P9icSN82PnA1eEGx
Q3oypGAHFSgzh9/a90AJ92k2ov1b6TrgvehW8wNfElA+exSBV7K6ZVpUd5r5wpE8hSolLdjUop9w
FYWWxE4NmbBzVqcPw7DXnSPv72aJHeGyyhUBr+MN39M60qhllHM51JQ4f+PbK/NsCjQUQdn3Cu8I
bZr/xkIoSMPPVwwfnghUwSKavk9iXnQCLbDDK+UpzWCLZ2pEf3oJN0wUVY9ALbxN2jjjwllJCXHC
oywy9iOboaOACApehgt+9pk27FSZ/Kke2zOgdWbevyDdgkPghzdGu/NDBHzQOAqsGFlHSrImalOb
gXScusXnhXt15ETf1sZZdnyNDPUKuE/ntVDxgzzrygJWBNqzPIhLm6eRfGvKSmy/cBbJu8SRX+uM
9mweVomPPR/+G1/gfbzXHjY1m4mIgBUnZfXnRGkzPP5Ap+IHvOGanPbjmTkBJHn9wU8f1tkm3I4i
m2rFsj+vdS0+9jdevUEP2/nfGpMopFn/SoRvgc/dlI9OsIS5LXIIOwBsE9j0fuXovWGiScA8UTvw
rSnog0SYnsHRt1v26iPldOjFOLxEJ6jNW4vltKSoSyN+N9axpE3w5YDbzUNrrAX8XIWYjIF7+46u
wQbTCFMzPabyWEAgTJAq0C3OHzZt+b8Ql+NZ7I/hp/WtuR7P6Y9un+BemxExVHQo0CX6dd3QMvRR
v9ADCyNkJNDesanD35tC5FhEgoVEMmTMSrdRTDDzScoXzYaZHHRjVIS3YKBdYg7cZImaZU73gVnn
IE3HoMbm+vtsBoDRdsP5Jo246gA/sd58ZVz+TJQBfxkQ8M0XcYWKtUx8WAur5Bg1t98t54oi4Ltf
Dycno3bABLRDw4733/2DmroO3XA8aoQBhMs9MFoi9oR/5EV7OQKyW4MYUgnn3MOSDLhLRRvGlcun
MV7jqhCV7KhBOLky+l/XJXQ8uDIB6FKkI6yHJnWMXP7gS4dzNbwKW62DrrZ7hkF9P1MOMpPXch1Y
R4TgJaasYsS3ORcSWqNJYYbsvDwZFFx63gjRBZ/812k11jorGeeAJJhd9moCPKj5VFE+Rp9EawYQ
vH9E9Q1uzkSTQetQoh2mdBlyitxfJ10GKTWZqPnOjvwHUIMFgJBoWc39xZo//aHdSAysZuq5wcFJ
G6ZJxWCPu2bUNkRDwVd91Jg9fELX6iqr+iUddXT4sQNLZ658+lp3L95YFpmVJb+BeP6YV3kGRcEu
aS7N2DyZViQIUcj5v0Nv+hDekMK3lWyJI9v/e/DDDrZKT8mAKn5aGl6PdBGVCnkcjYj6a1qEMAWi
mPA4wj6iQGJzWmr7KYFghk/NqM0I9pCIXh5VDVA4JDWGNMNFu2BDii2FoAo5FYwuLFZgVQPGro7W
ASzqeahaROkAmD76TPgzvs5tIWcdBinU4Z4QfKDiEZWk0b6QzXUDQC7ZC4CjwdXcbI/l58PlHBnS
8Gg7AwHdd8/OxUFxsxHr94bAhid9mhI4DIyBV8niSwtLYF3F32xAFc2POpzj0baHtJts48CqNhPY
euoIQFlkC3zB0Qg5FCZlaQVkHflSWjGAoUDIwdNwJ9WLHFGdCwjwS9xyMpaeDrG90IKN3nx3lYSp
10xaKFn9I4wrppIKtaQA3cClYDWXJ6DH130AWhmVhM729Pmtdprm5k5mFHQVc5sZQtXN0/Qdv+ci
WkRjRaMgy1hy+RFRAL/BCmp0VAUELszOijd6yY9OcvZMYA4VkVuI9FysSBf6WVw7VhYh+28IoWVi
gv6ObVmMQ/hUpjvJ6eJOEgEoAekiGJLsbh+p0XlmTkhXus8/Itom60y+mTOArUKRCZFlSyhLX5y6
/Jq6h0vz9rAPsM8kaASCK6aX34uDn9/2spa2t1zgrr8ro3sS51zH5xbHqWBrnr2JTzkFbiKwpEtM
VOZlw6PAjxETphVJmdSEp8M2yrcvU41N49twEvNlo+I7onO5f3enodS75GbzJ9jkDJbggk2truqg
yOBDZj9d7ClzA76vZf/qoRsRH9IvHme4/C74K8HAQJekEBF0FCkNetqL2Z8YiThLDYSf9XtRDa5p
iqy5gSDZxrLkmp63pcUmwXdTnNnyuEgsu1UvFWt3bhbh18dYbG8f98ZcGrvBIlgnI84AzMnH6U0x
5nBPYG5hFOrzaKfCVasm5wkU8ZcY09JP8A+ALUFSvnAy2KGLEF0hCk8DyGtAVXkNVoUIcjteKPxD
O5EkNIkDU0cgHzvwZ0PV/OHz4/kvfFUZoxeNMhfZ/qFAiKkubMnvexpLNEtF+fXmWZziC4egbI++
6aKWDdnLS5/QNa0n0ylP6uKuRfx4EiiVQMc86j/kV9baD98hBZMp1kij1gHgAUvYpp5xox+kA7wH
oSs2tRiGMWUmdVDhnXOJtK0/RPvsh89phXLJhUu4D8u+Ro8LmYwduSkJqQYchua6/1BLshH++ysi
0mt90G00rnyeK1040Hs3/rSXPXoDfPDCMswFN/RSNmH3l83pCbyj4bYdsv0MZUBPvqF5MG4imK/m
MRcik+h5scirc87FDBxuRvFCVAQ6fWPEUU0a4EpNTa89vGJVjvX7Pu6n6NKEW2Zw4uj5edkhJZi+
5vdl/QlxziiQYzocsc5DmMLfonSZOe7G3csYKaWBIChCme6+4wHQMgNC9EoHfKaVnvnINGvdTk2V
vDLEl1aF3JcfirmYPKVxmvNi9dx0mhL/flJSgWzpkqf0MqxMWFks9uO3GhQBERK+Jx9/AFXRfR+q
nqyIuooKXEPoevr7nnjqYuavQa98yA8dELkfQ2HdodNwkMXkdXjZ75PcvJgZqkV7JKLvDLPSq5UP
806GZi2amH9qom7vcG2mp31t1reI6GCO6rz1D+fq30wxoLkBTXq/FQa1WRuWhifELUFRDEK6GQTc
t+ukeHqRQNv11A7k1wQF/p+Sf7uALXBCMnP+kR8Zxnrfkx5OUNWVgGe8LBXdPCQ8MOiuG2EP3JxB
LyqDuuy1DsS9W61+ZdsQngU/bwq2v/CMAwhTXfq7jOQWCB015GkyN3zLCbYOAdoTNLzChvT9Js8N
s4XT7VK2wZvi/fOeJoglHs3FYUNIdqHNCeCBbqg9Ms0+gWgwQUDzRsKB1Pkooxc8qqF55ph2H6kC
JHAg9N/KZY/LnjYY99q4jobvZcLNisHWa2WKahYGc4U0VhVEpH3Bnv7rXb4NbCpfLLbSHZGkqb9n
YdwlZHv3NgqX8i9Cu05N2JVzAN16MshDUwgiepnEaXUzhu1gqfSfrz3gSCzgg+k6t1QdCDlqbzcM
Bh0BaiAwha+vCTYBy6PhyMDhFU2rdsSGpv4i762CjHb0pjXuHT7M7RIE6EDSie1OguPGU+vw4ile
Vchmsw6YfueKQU3Wcbg707KYRPltTFyLyjwF9BXUcYRIkEkmAcXQML/5Mr0MiRI8SMe6dtoAPOQf
0TUZJXZlVKq8dXRjyohPSsAEIyG4rEoEAnrlcPUimKqM2E9RFcLV4LmG2dFScdZH17TZNfoQ1KE0
4pDBLWzhzrEeAy5tj55iTZY0c9+fqxxAiFanYedNisNANda9TIpM6sUuqHRuoR/xcis/q76l6dfh
SnXI8LiRVOMO/YHCK93CZINs3WqGd0+XeKSuRogvU5u1x8E/imwz8saYNBC1FdOrn9l+tSoAQmwb
wz1T4VXvFefyWK97vMFbMB/2yTsd95fUUz8KIDWeY97Hn/UmO3rWL37mjWymX1vN2hqoAih3hF1B
aMrOX0d9BKBzHovxEKjYDN1yKu11L7LcVQP4h2+ZddeOUeV9PtqlyxmPkpCTaLzPbYebtAYGW2+8
MTz4nkk/MsPLyAS4dcgM84Bnv6TtTPf/dKffyG0qLas7klZS5Eq/OHQ6Pgl8TOKAIVFPmQjgs4gq
5qv8E5KqTiCPct5NguKzFIk9MKIGMg19TtWIzz5IhxtdjxtEwSeST/nw3oIQIyPB5lM+8UJ7HfL6
yGYgEX359S57tqLKVjfnUoQpqbNwBr0xEppy8LftEKf0DT3TiZDWhT70qaoNhegSO+f3dB0Xk1Ab
OymQNfghfXDHm4d2TcQOc/Xz2n8g1Siy4WC2Z9rUorRCLGAHX2HdjKxdBiX6hx41q57O75tizdMa
Ed/lD3/bmSAhXrjKzsROdgJKVPzbveLKn8jEIsdGqyMJ6YGmdD7ptkJrhttz/cpgzHoW8/C0NAVO
3/Yr1KdSIUNOopUnPRrw+4kXjHH5Q3f63YRc7RRpAKhTcMmKnsuO8Dwa9E0jp6ngcnBNMDFOlyLT
f2vzboNC9euXUIKi+TT9WtFwA+dDHiQuSCw08OTceKlIC4Ew4rYHvxGYNJoI3Iojf0mOga4yDVh3
2/Vmfz5PFevB0Asj+xwC4qX9sljD1pEz8qVP24NCwCgZ+kieybw54/esfn2XLnx/v7eY5Eh+YUkj
TQCcWafXNvKN0/UJtlrSzrjnSp8FZpBiCLIvQK+jDmVtgQtS8ehz55M0iUlZEWBX7KyhG00QS5St
NYtevMrNDs01hSJHeuDQcinJZ9qmhYnsXjFBS9s7KHEAXRRd7pIdGrWpX9u02iUTKyeTkXOLfCv2
4ApQE1XNy5iUmP43GV0xtgAnVFp0YuZWVCjeFivjA2IR/GSbWP6HHf5Rh84sl01ycDben/abHrsz
hDLjryugtxyQH/NYy4Htshrlu18EKRMyn8mcwc2ACiLlQDHWsWzyYbR6504TgKLySx7JVayC0QXc
zd7alo1mPLZEIzxNRgDq0SU8Or1uCjyk4POOVTmDvjdrv+mBufFO68bh4PGPFn81TLh5jU5ITni3
3qCl16su1voHfVLMEbTk7kwNXrXJtq+MiYa6/wyXfvYuTdK718Bmll3L7LurC4xSdJvSX/FVk6Mb
+xdG4MNlIVYwBBz/4PaWRqJVXkH6L3gaUVgetFTZAO/4oEmnkd8/WFMyj817qWd6m2zvYU2qWedC
yfv+SulOuGF1iJp9RWjAjS8C5TGWl8OIWaTmB1sHFiPeC2jQU0BoFOJe56Yy4ypCou1fYmeEQE+z
w0RfyWIGApYY6KEMQ0CD/yqCZ1ch4yYH2FbNB9r+qVR6uNYk2YEFlQ0PjjFsGm37lmxGrn7I/Q4V
6hqE9Zd3+984sju5as4MR+Ia2KT8gFhiQczXi4+WYdvqvFuN8f21Jz6D/6RXSebEoPF1h+Takfp3
6DQjS87NxuUwYp3nolNjHE1l39t+KkWbhje1BHFWxXb5FZvoHzGu7JIwyIxmQUR4lsL3S/VLjxGG
VVQ0DtK64xZjWFbdA1tHL2b5UV7NMztJ3BOefl69DraRg/R1LhHIHN55qBgbWOSUyMsittac+Nk+
NSx2sxkOD93LFJBXFIue0uQ6B6I6pVcs/h0GdZJffl31jYRK+cSztsf/iSMsxisnb3flQ3nTZzXz
/zth6WH1ewIdhJ6kQoC9QK0pAbmiilHSIzBuB/U7XfCWoQMThBGQwYClEur32vRBIiT2WdITWVwT
OLAZmJRrrqry7C6MTbcqizL5zaWrmRKGk/RD9i/XHqUQrzEdajEuxmF1wnVJBQBpT+PpS5plejd/
ohwUE3w4JULR2gOzwgC9naq7qTIJIHkRKx9uyK5dW6I85k5C1SfvYQCNNpm2efmVntN/qRtm7KZN
UlHYvT5tJ3hlTDytrGcphnr0GJq6YIJpaoPayGpWpdm1bM4ywNjQ0fw6shHcu3Hsx/dk3GVppUX/
03o1wpY5/XoyUmdxzoAFRzP1PHeuziuFX/bZJxi5fMIm2QaeHRbh9DZDu9kLgpbPxuV8MQ2WGzkK
TcRmDJKBQgWCJJDZEEn1pPMEYtsK4+FEhPsNcz6CdYhkA6x0Bfj0+5b8FQ3ss4jCpkfP7oqISQ/3
p7Px2vv8+OWKwI400sX3rlOPucv0da5+2eoFdSNMIVRnmAtL6owoLV7YudXuX2RvMNMFRx0sKB5/
pGvQXCNbt+MgVgCwmF6bylnQwynn3tr6Qkqqp+V6b/nWuagerUZ+jDvnaBGoh1bkEJNyCr6qNckM
kf6Qmb1KuesJnX4mwRlDrBPYZRHvsAx/mYmmtJlKleLhN9JF4qCAM5uqJOLyaanGRBKfu1S0peMK
72IlGE4lWN+eefIiwlXgUwjMId0CSTmo7G9dhs1uItj4EGvWiKLrete+KBwfqHazkd5ClWTgp960
vvB+/928ptKGEorJU4fE5YeurBjwefV7TYHrVs4izQva62utCk9zgcDM4w05GRMqkLXnFSq/Wg1s
gJ9LapuTo8xGfiYBY41cHFfcE7vrwaKq70ydhcXch+3LDf7hkC0svrBUlRbiSwadTKw7G/peU2OB
OOZwFQRuhyaAhm3HDe/KQ3NQaP+9fBwJrRBn6rsRJil1fHxrfonj2jExJK3wHtAkX45RCTWrbQq0
fVNfSmfZErqHtBfHmBsPH7Lv8y8EC8TUmE0jNNvZxnadbWkDnjfdPD5Rpc/4uYdD4ge/J58dXRH6
6DPIvusrCdf5+f0c7ZQSC8kq29a3fbNpfF+wbtlH9g2F2kLsc/W0brzDNZoRpH7+isBDDZJRXRk9
XlLgbEUj+AnzmSxhzK6EA9/SNvpC2GlAVYRkOLRUJkqAOuTosbXfnH2gNCc3iqSKyvATh+/rqdqd
+ehoMsfrerXux6GKUsnoa8mceVMvdKRbgEh/XFvTQ9FXdGGfJtZzQwcn3BO9MQNt94TIXTioY0CT
CVOFraxmnT7IKQBMQg+SWw3qggotgrTW70SodZzY7p92kZ9JUimzveMKvgTrwzSIgcxmDsNFgTjo
WBL+sjqw2kw1/yvt1P6p4s4kM8yxWigGsMUprZfn8I0ajWveSY7o5x9ZkEqNRMFbx9qIZHzLLHGO
O/0/F0nSnQoVXTqxN9DpVchvySMOXO0YDvD6QidUvHi4mON9h1dCanSC27W134kqlzQfjqnSZZMY
gtnswWtA/t45Xha+VZJE6ZcXL+r2VkDzaqaYmG8FTkUzIwlYI1n8t+qT3X1IZa5U+IfTujBQXm2j
aubbhnRV2eKd21lxRZCIyt+nlFlCGES2d+S8vkEpk4ovLwjPACRsfaISO7UMFSyJ973UXsiFYUR1
iipKMOMfjWgsNG+ihuisMo2wbqTWfdn/qFsvO7on8vLVcHJhDtBgUxnk9jJqWcCaPE9/+/6o0xnb
uwzqft9Lx1uKdgXkOsDNbnC1o2+npI2OQOrcYeyv/s4BWLJn3OH5TKC8E2anZ8SE4woCA+RL0IEx
Y0UpsnhRJBp9Fwfww2/pzTz2dg7a6ZhZPxLl1h7rVyns9osqzH2y1JYvXO5aZUSzpd8rpXgorJdd
0Z6Ueucu34400JQF2LRBbBQEtcqk0n7vNcIqER0Z40aBiuxP+jg95a9VqBqU0KxJO+gE5cb/wSAA
J4IC0GwFQcVZya4NgEnHkr97pFBWaIXabg1bAbY89jK2VhygKCjdy2bH8fpo+hOegNaNo3d7YoAU
oN8V6FM+xZqKnWz36b6e6nTw+y/j4OYYVNUz0J+HG3bRqxWljLQwzFYsw6wL5X+pGGSpHfvF8xUC
7ukRtgvgODB/2XEOqTnT6+uG6rVX9nj+xIf0ww0ln7oRFuXnwcxAYqSUmdKyiyuDEj+EwZiRGVqS
VtgOi6od5ZVg9ecX69KdhsLm8UrxbTUFZ+EYvr0GzHEepcKP9nguFb98srDnAlk0gHw6F9QJTQUB
fpKflnk6bNqPnvWPYxzJLVqXlOjc1x5FoeCyLUSPOur9lslrLcUmVVQiKsCGhaz4uzUEArpjDe1M
5WPANeHfLiWOHpvQd32qKxqHnCCeeD+SQfaOIhA1s44hJtpOgem8kpXgupVOKq0+0hBMLcH0wukt
F3PVTRkDNGc2XnYRt7CMg/U0vRAZmwusgWuwmVqFf+ub/2T2TEZA19PWVKKLv9R8BcG0Abmte8xC
7ssuiNGkBOJ6eyMr1aPM9EZnbvjx8KsehgXQaltHdKqjKw2Jb/vs3e9ZbDUbvs716YHS3oM6r6SS
Q8loVaa/seX/d6yETQnvSUWVpGudCjWbNMF/v+QRPmyAiYTk6qPspfErhDBE7s7FiVbJgfJZIiOW
IK7Ya/nj2Q7kGFvTgby5ipqNOmUxf+KL0xX/jAPrLlbVg9nPZLZsyI07/hCslqIlc3xxHVmoi7Yh
XQgdiaMrNcc7kll6CQAP2oXHeEJd7Cc5L9rZhlGQEM28qbuJY3fIIrL1hNZiLr/qva7XcEtH3Ov8
l6P7Qgc5A2SK7dgHiir95TYFGMe0TkCa6ePayNwu2ky+LCUbACUluxaLgk6Cj4Y1Hvwr/qBb7NOB
nAumZeDbRmr8r5fNQcq2g2gjxD/azURqQFRzWZPlrBFBTY3Ja+CojfCgo3X1iJdV1/je8PPLv3kr
gcwDqUprR2/4sVmSJX7s89RSBRpU1DdZAqHoM1kP9GrfVT3/NEPx7tDhEBLIq+Jgxe7rnf/fhXro
SX5I1dyL5B5pRnCw6+tMS65Vge5byFeDIk5k5zBpECESmnJaNmWCMwgr3UJF+afQXKfmYtyh8B6f
Q55imH4SqJ438d0ajQGWJU8yZu4sKR2RR1FiFhDiuIw2RgQmCRtCf6GYl0GRGOb3itz3CVqcbYCn
O5AYLjRxxBNNWKLwSKxEvjEyjWtBiGy11M1T6IS2FYZZalPzwYu0IJpAUPRZBziV9ARfqgu1e1nX
9+YvF/Aj0Wbvmn297hrzIShrgRLwr9Yo3fVKhmMez0g1erXBQQ3CPd2AIrNstix8bCzUx4lXMr1h
547jdkDwvpEN0ZKfBCbTtMUAAxoV2HU4nFoudnrNCI+H5y5eSnyGACUESYev5qNPeUKa5/GiiWvR
DvPMTHjSEa6ImBuoBuPQTtcGVwxudCsXyWn4JzjHaeI5j8A2n3LP3/bLGV/z1f5P6hsd65evEqXn
vyFqx5FJ9JjPStXNrbwfwMeegBGfoX4lLXjk2v06JSHCP7QYcy0FhKuAEXIoVPumG3COmTFjNQxy
icKWDL3YyZhBJUklr6MoAWAqy9itLh21KxlqdZ04/2u5qI/t4CL65me1gGg40tQAdv+pok4SCwf2
4D2PNvyTVdl8s6NfkWrqbY26HlDg02laezogtvTNDtuqQTfvi5bzmw8Oz+Scyx+dDGQm+0dtvULM
k9ip5rGTOAaIYWCXHnzowt5/x42hW4ZHk6jFkwtpvbSxYqEcbWolMd4nNNC13bqC61gERYrRaUYT
hwLwY0b7KL9D16mIVtywThsxpXExFy1kfxoSQIl3MlYSgFZ6PF/RyT80oytRdylQs5A04/DX3/Gt
YF8s67XG9o9fd+v2ksDaKRzziM5Z3m+ClDXuodO/Bb8BtFVjhHzVzNniCC/+/2zUf8H80hOvqeOK
JFC7Vco7h5Qaw1pWReU3pJmfudbiHp2mXbfFdki/gUGDzYgmO+ypKJ9d4K3/osPAsmKPDlYCVh4c
DAbHdj/cOZhQu5g6/gMAMhf6MLBg9K+VtotWmKolpKb83+Z7JphRCxhsb2sZWWM5T8Fj8LpvovdJ
QeCYyzhV1IxiAk0pOags/frQNUOoi1uu+4wRpzbCgfbTIUKe1M0I/DfHb02yN7ZdeUMbWZ8YRoiz
ZAbICGuq+r5BIw5baTa6d5o1+0YIXqGhGiZ3h/aECE87ITBgThEpaoIw8beAAlvzWRvc49c48aTj
uFAIlAxM+62lx5LBJLv9b7C8w8P349TwHwfYuWJady73JGxrBTVSxQp2izmRSxhiDzIjOpA0m93o
YwPBeRYv/NmGKex0lJosVEMOpqMCxHR4Y+kn0EUYwbxHNOCa2ubLEJ24t6MoQFIAK3rb8V97hiay
lT6a+Xn5XXQKLMCsxrXjGhOHvpoKSRpJ+P6MJBBYqFcS6YqVw8ISxs7kIBqqHLz9MvthkuvUx434
C/gNCIzLISRRBulvAy/c1pASF+lq+TMisdEOLLRZopfYsO1ptxRfLjwB8UrmrmlD92YznZ9lSoVa
CiUeFlnET1pWKepQjSMS7O3a8eGgpGw5qhkNC3B4EHDZIB7Z2ngx2j2no+fwXa0t+FgMbRDUq7zj
YGTVKUZQGy05BbdEqJxv6rfiq5fWrvRTpUDzk9z+9uje4L718sPSsb4xzqDq3nQan9dTLyTILZ4j
vR1bFZLeE1JUpbU/UcQ08+n9EkgpJuA3CG0DOS6d6qz5liNUU/mOXrimBO+JiTCd13fN7IzLn3pb
Sx0kysh4wNJFNR2LL17Qj8n9vG7oKyKXBIlOfDyOarh/lhMD5lCC8GC1nan6rG1qwPe+O8z8nXDn
ji/G3ZSKzxyD8nYPyMxE/3bGe/6RA2uhPw64k9+dMDBqQbQ03xhcGhVSdOQwoCxSLs/qHOVqoV//
FN9cAX0pwY1nJziGM0LSd8wbT8SHRcFNsKyEwiGkZ3bOEpdt15xMjDNxju0fGDoX68yEjFqHWnpK
F5y7gOpq4X+RQcgUOM+kIgRQLx+VkQFUmL/+jOAin9SUERn+p9/ufD31dCSUX/NNPRopuHZta+hy
ZhF6mEO0Z1eHKbZKxQFs0RtnRq0i2HBtvF0fXO2++LFIKrAnQ3YbPddoI6aTRDC0yGYqZQyu1wpr
Vy2IAx4/9BQbnsyKCZRVfOrmIkMa7bDmrTeKUrdoCl97Z/0taqvLqjzN9p5nkxGrGrIDJaxiq778
bva6+GWKkIidaDWO6vA2B0sPg7g8LbUsvkpYq6PJ763sasPMyNs2BHPieAAph0Lhpy4O6XDo4vpI
DU1C/PBxzuroZS3LR02UQYpgZrCcm0xFdu1S4lVKEDpUAL+bzEwaVaXjep2LGRZrxysskiHmcPmx
3LNDx/9cYqFuLAqSH7yyF9YObyvUMl8/U98HlSRnRETqXjT6n/4N945YS9eVpb9+iKt0RtWq7Smo
Et7SzDc5JmK7DaI0WPtAf4M7T1zJbT32zMRN1SKChg8QfWf7dA57E/Lt5TN7/iQEQqU1WpEyCTOL
gi/bQQZLl95LN/DaaHnF58z2Mxn0dCLiUZ+rBHk+tHlQYuOhWWf0u/NFGCQ0a8YRpbf3+nMR4qN7
u0OI0Bhs+YaBD8IN8cZmGsn/xYwARKEx2vlXWFB/qZSsfUDyRMprVpU7X/4B3Ki03DYyHqKdtv91
9goNRhI+5+DGI32Tii5bjYxcD8M+VCCP+C73sNu+w8etv7NLIVgU3hXFI7iFUkgbijclmqdR5A6u
Dhy2czdRbxcj7xIATXaycuDVsDGwqqc9EaPA1MVIcJXXJhzK2dXd3AicTbokgPsaf6SXETLk8pmE
jumf+Nx0zjcO/D2f/tvHtzmvTzros5cNPZwzlGZgG1ZAYGmGRYZojhLLegjKVMRCEwCo3U2EX5Jp
Oy41ZdyACdkJ7pDuWnFS8akKsebuE546VcKlbS2e+xcoVDac6OJpiQtaEQRYQDHz0kIWNb013Fnw
D+2YdvGtmRiS6uBcw2uCN0hQdCZbBMYAlAPsO5F6C6Q8iP9RRbVvg84umMd2AAk2WpZj+qshDrvI
DRIWSK90XA+S6pngG6yv2gg29tdPYewQZaEzxL0aL0p8M4fXOpJaaS4JPhq6I8ZCrAsaYZXDe+Vt
ixvEToIzDFmEbKGspzTr0Xw2g8YBJr7UB6yQDHf5NuLb7LH+GnC2FKSFekNflKZ+DpZ/SBSQOuww
VhWCfoj+T9l+v1wP6sHeRq4vaIpMx1hZdyOFsGt6cw5O03vkfZ8x1WoQCgO6ItgEYYtyx8f9HSWh
49xaX9hvdome4OU5Ax3H4V2T5cHsnUql6FyHkEE1nOZRkOQYI2FQ9wHV/+8OQjnIV4cLXyXd5whu
oUaZZdCDn4I8RX79LyRTRmOEn30oV58heAmokXMsrDBZIFfSoWiO1HK9/Hnb4qx4A6XYoEcrKeRC
uAjDkQQLY2HMUfOQTeSN7EnRm1GTDrW7aygQTUNfbD/FwjT6lni1njGgO3ffZfEEz803O+g8wTP8
FWQQUJ6b5ER/nLA6l0RR0khpFy3Opaxo6XgCQuLVM/ycFqQ15SkkFkTGRiZ/bdxgzSALquq8MZcV
QOh0fIFi6vkpkM797uoAnklXGAcAyvEGKUkRv0xZMxNBSaxOkcpZa0gjL/07NwClf/MJ69WouOI3
ifD0H81sPIdUZtASCL1ewo/8xrmbH7QQput+91Z31fSeia4HlC3lgeu7xlZ/UOLgHtyym7TPmy1I
Mdjt70Mfa7UToRogK1iSFdZttdT9Uj1z67+dz4K5wtQOY90/Jpb8yQAwMeB5EfcbYEncWVHsA71P
f/AUH8CgR8tpqmJbIeRnAX1Q8LpmRnU1Vwp83+7Xybt6NKJfwKDAoQTd2sA7wPI+PogXN+KXv997
xWv55gJQnHOicHj4lxfCGGE8FFNRNmVYxUlUl7h+4fKUWiOpmrP5eEqeFRrR4cGKDDJJcAAJcJjQ
5xRh5W8dB5VDt22zwT5ZR1n9UAHP8NQaJ6ehx2mTtDJE3IuNqNLB20gCA8p+0IrqASCUWnO3TVon
pqTWlF7S4b943CZLHfdkfJPktwcoeurfiSNTODkMZ4oqNrZzfReu06Ur4SpTYg8D+BvpN3ZGGjuw
NEQVUc5DtEz8jDSD8tZMW52s12IW+bTrKBMC8Eo8Tz/bOLtZ4puViSDHfMCbdX9EwBtvG+jKglg1
NB3NAVZ84c6jshAOEawGbLch3m/Lxn/CG5i4SXApfTnNLpuxZprEWrS9mi/xsfa/g9SF0YLCpEIi
OwbH3QRneEAhkK0VAv+eoAAth+10wJaC3h/HXfO1qNZvkwOOY99BmHeeigUkPP8Up5xDvwknIHMZ
m0MAB3fvBhLLmdHhy96o2u1jmrUpkBQrGnyYopuY1rOBdEkeZfetiX1Yu9WLXS2BOJWgGbaspq8X
a4P7slqsTUUb4o+kRlTT+pcYFsxytTgd4uuL0btaKGbfoE14TkJtwtS8Qvk0/Sozg8OEXpYj7+nf
SPl6DJqmhUjv9Ssn9ELB0rG0WBCkRTUVyZXuPlzzgu4I9CQWQN3iA1Ce7fTUXfODgF7jDxRcNTeQ
ZwpfTJvlzyC5Zvc8cssxBWpqwlocbUeOC7Q1ws/nUmm7aKOFIMTFgFAI6l9cTNA18Tivwe1DOpOa
MhIlz9nk+WdFjLqUee6MJd5MqlSahDPX0x1xq1EntogTX3sQVZNQCpU/ms7OPxy5Q/Q6N8ErRIEq
VJkGZdRuT+alx8OPKN2QLWNaxjU9jFL7hC7XJqlGNLLP8Gd20hyED1ZqI5O4l4QJD9K3UN0S3WUB
MLUuVMXP4akyp8tVACFYCRucT5Rx89b4vhK2j5qAuaqi4FBpfvGMuPG/yodkrosKHkd4jUqDisDa
xM2P0N6LhHjCCko+w1cmLgx+eA1CbIvSrdjGURPybtOD31mdcQ3eR6K0+ujR7yd6QrNqV4mDYcv/
4U7riV0WdQ03UQf6LBi1Wo+qnsvbRTI/bRU54HAGp23rDDVh1hmLafL1F92JB56YL7Ozltcne837
bC1+GiKdxh2sBvaGvR8sDXw2vctWmFmFrVgvPwvXWn2ndD9yU5TaTb3QZgHootfztBVCY3ay9oXT
XhDZi5SPFkFyfY0a98RplJIQOaFNUk39eFiGfQeXLUlxhYwZhUA8ewiMe9E3mWJKVi2EpfJs3a9w
LUIdbej4R8b07qJZjHfXb832QxXpwKG7rICGYlH5PhH09DKM1XpIBJo0EUDo9pHmmO01eYycGcBS
IdqEmfniQKl7KSZ4Rk2ffjex4SQncK+LeL2YNx4cMSEiVAqz/kmHmgR5lr6WvSivLY9nphESVTJs
bdkSMJhn6zWsJ/nd4ZZ0pSNjTTWVJiCUgxe9wGeb5V8F4IOhhDM67iusLZ2yGl+0emics4bR4qX+
tX9IfjOuJf6WzUKSv4HuGyGOB49y65BQiMPxD6+Zz/1lhHQB7TbRID9/NZmJH7rGAGYywR+U7kv3
mWxfwn8rkkNvY1Jmbekr5vbU7QojMxAmeKGjxMzVGUFwrK+btE9ZrnTl4oomUmE3oTlBTNJqs726
lTBawcoKd5kXmgnrirNxBSlOZTaFSy3cwHE2cn/1CBgBcivcqCysAeDaK95BsWaSQ91ctR2Ox0j2
qzKLO3B1aLzRKMog3agR79Ku2FKx3BOZv6JFUXaM1faoLd+FAce+MZMrdqvKtlrxK+CwjKwjgB/h
lH+aSt2xilbBjEub/xTIg+SZeKQT+Gn+1gBgP3QbTTVX1ZSWRRx5VBZ6IWrjji411gy3DlDNTPvg
xH1ixLppWqZ4HQ7NctqsIlraNJ3laBKXcozXsICqndMsiwp90siuTjuJiLd1JLsolAvKTu+RvXLI
af4BFGkyLaYSE8oSoKPa70Io9NpttcNq2a20SdjkhTNra0QTYjvLUqI9hcV7Uj+O8T4emT9O/MTO
29Dv4wIVWI7wYcBSK8EGvDMd+zwgHU9cmrbpBJ0HmcblzUtso/F8cgLKdJABScj1grUwLLzZC2eQ
N5oKMKJ3HviXsvEfKdNzeXzoDXw4rXXguscEpnNqIJd2mvuM4Da7814Peigx2rdl4SyHyLvjO0Lc
lRvzdz4LkCyoOqKaXNLzH18KcLivA4X0L4ogEo683aDAFQJMvvWVm6AfuhpgE2TG0n0aJlGeF3MX
sWovstq/TsBfuurPmj9RJXy9GHVNMf0mt9xiNJbMTZAInl7jDLR/oJxk54Vv0X6dCYcHEg86+TRE
172rqMXr9/HgyTfM451D15Dezxy7fk/dyofnNuAB10doPv8tATavFEObXqqiwmz9pd2hIBXkr024
x9eYU4WaTPvKdiAnzVRXZ0kLsfl/nRTc0btxUHN3+vGPadHRk92APkgJVtxEWrjqH68P898xQTdM
Tseh1/83NNpqkhz72z2gZP5UJrBsTXKW1YXe15emWoti72nzSvVSKCq4q4q99+OKkVwgkEnlG5aB
ubZ9khBZxgDhfp92aSiEhmqPNKiqip7AOyMSy4ts6q3a0sm+j9Agi9yydNMTGQ/Qwk1qlAE2OBX2
4PBYzMm83oeyL5piQNO6jrmVNBxGzaP0pVO0WUymwXvVFTQRWUJWX3b+TwAaIHeSbPZWlfiL58QW
vXe44Zib7X4A7vQi7QC7qIeo/SErqPIZoTe+/kE2ARRffc+zmQZxix+zKqe8iPMYHNg523vL0nPG
ZGUJVEaPrDZA5Mmol3nHeaGZeSO/h7SMpX8TFMYJnf8X5PI3FaBBng9yI73rxCE8/B+NkW/gNTOm
QPgXTHeyEaI4yEHdm4kSYg2BeYOrvZ594kN/1+gAAHGJlxONoxp8ECgG7MbOcCyL7VZQWkfdmvY0
GVA2VKSp0LEetqm+OIhAFxuWuDVWHyUmcrtu/XYIVNKk3GwHHG66z+ORiZhHCkD3V99FNaK8ia7M
Q0pY7ulsv/NVJBGWEHmgc1EwnpbF346RdUaV01S/0i0fj7aICPmWmHcNJahRwTcxmvZ/Gb//FQK4
fMKYKsdNSUYZm6+vszlVj2fnp4nyO/Hrjpzb5A+MQhZRGBkk+vyrBavEETuM2ODvSwy3Z5g0dpEq
pcyR2GEDfSIFQW5gEj5tjXKin18Sf8sHQVCw0fJFD9mJ+25TcMk/qclAWk8PEQtb2b+GI8B70bPb
jiz22SLoSrDx+6GeKBWWhJfQ7K84wbxpzY6eLYlXLqcQj8KdpDn0BmWt/NL/KJGlBMSksK7RdtR3
bi7+MpQMPUG7ZBIWZ3kWBx5UuRKhgtOyirTjEiJntxuJybRQRgBFG6dqy1Lk0yKnHFqc67q7gIt3
sbPXlk3zRavWFisUyWu6hxH5LCzRnzDUWK1a80a5qi9R7xwdmkiSCyXhp5StQTew7PIBPjfPuiB9
RnhU05qMQVfFKmBV3T3pLT0o5Dl/yTCAzo56P8str1f592k+hyddFJ/TBcbOO9UNwR2eXC/2tR8h
AMmjiEiWkAgQ9UJmz/heXJSIkQxFlsmfNMav+SaC7HjDbBr97psYm3jM3HERmrjTopmXujK9FlWe
C1QpU8hqMo/kA0B/3FGMUKO2NY9oiyMqCRFspDLuecOpSj40CLFeJBVvsDkI54YchBcgzedeTzPd
GMbyeIyYs6Hp2AWLdVugaiCtEmCEkuH0VfKXIRQMyDI6QLSR7y5aoCAXg4/siCPIOH/6mTJ9rNF0
7Qw2PkpIvLD8VgorPfG0DZFBr1BycgdKpt/rxcRUnpXOOyYuGeCFsxJmYtm+3lR14h3eHLU50S0H
xTsURtaR6Q7JTIIuUykaqc6yA7LOGtqs2NP1gMDbT4R4eYLHW4mJ2mO2C6uAwjHYJYZ/85X8fUSW
LR6jeDTa95av4RJJqNRAZK2mXGYqV+jQomI1HCEtWf55miN49VLT2Zk6k58FxLNuTQ6OJKgfbykZ
LrG1VB31+jAZVVgAbHr2sLzP5erhZK/MbIOBI+nPO0ytp88kxdq8KbwgXcLdMxhcuX/p0yA+pp4l
aGa1A4ROOsVJTSHneIz12myrEueMiwwRP6C/V4kr9KZFhy//YzWucK4lNW4eRZydb4XNVNNpO6Z4
9E91sthm9nLIyEhxVS+4VgTC5ARH0XkT/gkCED6mWo/IbQnP7//kWu3h0V6BR3DCrXs78YkSQdNH
lQLTPqAOJSdcdmzgX1r3RhtM5a3LsBrBvMNvlMRSstwM8RVmO4VLIg5lDqft2QHdfQgf3R572H2n
i/wbepsOjnyjC/fTv6SHDJZECaOrkkBDQyJ+/D5Zo7oBoi8vJZDXC0x8+FEeE36m5rOY0TqCt1Rp
09Ue2r1+sFV43ws2nKr1GXlJrzF99Qg9zpKDEZ1phFJsFdzlcbZFXaxoN0ie4nn0S03JbpDGfnfW
iB6SSV+g2E9x9uoRolOb41c3CsqvzTnv2Jv24Ccqbnx5TVYhPUkWg9LtYldZB1uJtNrN/PjR2s+S
yFWHLu/PrqJ+I4pHFUP3bldMOWg4Cg3KXeNoftUlHrgcWRQEjVZ57HRVT61IQTelClFdhI8i+Y18
T8wu0x006iQ04ExmLn1mS5+1F/lJw+dtdj8zO/thB/sOolx3YWmOrpaK5/nht27+o6jbaBXScMmE
NopWedwW1591oG6p95nrNfJT9+UJ3QaSIbrUP4UT9/XRKBkmU9geLGjGxN8mCrLbIxbvF0KbQdRc
TA9bR9WHZAKn0ECWmx2ybmkFHgOI7nptBWvwZi3dBTzBJfUbhEL1y6c4ds5LSqZDLVexV5i8Dcix
uBwrxVxBH9Q9g5CNC79aKUt5FWYZDbreyKKWF+rFR5QzRcKlvvXO3/N5G9gyrIHvTqbxw7mKoxXh
Vxrsk6wRY+XNTY5hgvO3GtU6vb91zM1S+sbmmJQKA1EHVIB6/PFeDm0BFJ0tBZy3rfYYhUvWNOF2
Mj+eVawFE7HuB6KwMsROz6QTH5tywu9v99uxI/3uQKbBBnKehBU93Se7pT6nisb7gt03X0D3a9Cc
7JnoA6r+hGayZEoCVoborBt0wQltracEZ/OLAOEy8mXcYR91CFcnGWO1c2Z7Pgl2XWhPn9BE0oDo
8nxF4uEt3uA/KXeu7GT09xD13yCOVEL/1O0RnCY/HhDlMRZKMoD8Zvu7SyW95UIKXuRGOSWd8gvT
RPTEQJuoI7C5VaEInfGDjGhOQnRdRTSx416ehF8OAEBiY7VezHFNmGhZTmK8PT3CGUJu+bVh601a
oF7nKePbbUa2xxnREQLh3zBoW+gg8zTfgG0lEmQXav8X1qdsBydUEFWLTR3o2PF83wKfRX85z4BR
+s9CgP1l4B09CPHR72P4Po2XTRnjwpmpGAo8cNO5+nsKmLTzsJjzWyhHF818bqqrDna9z2hPyjXr
iT4GFlw84GPr62+rsWWbelAl/hjK4BP7taUrtM7WHiG1mYF0Y3kHxb3FzMRMQhiZiJKGg9ITXKFp
E2exulJnYkrJfYio6qd5Rt0vfKxGO00aV5tm+iEDH9RmrfVV+Hv6IcbWquyIHYe0iDu8M5r3O6C1
uwexmlzuSRAOYkgaif22VsXYyCKOoO6l4KR898yKcRXpPgPbGwpFHsoyx5zhO8xxu6k2AXv/3UzS
MngthF7Wlo3kgGDW/xJqjYrkJJ1IFyCPIAVELtpnb12UVSQ5K9fal9sNfFNF8EPhe5CZl9fz5BP+
o4lHF1AZh71X+ZAMGrBdSbEdmXCw8ybA/87td0yfh/Dh5Ks/LheYGThDoRc8qRLhEarSDqPo8KP/
jWFhmmvGGVf0LA+Gf+TIJJPo+jzerFzimSnet1MQSGZTe2WqpTHtu76dWxG6IEVZ+zduxFHpY512
66e3YhLcmP3R4yAXbo7hEl48jHEfItrZD6ItBp9TxTdkzHsEIaUTiUH/jD4U5F8Gu00hWD3C8hwB
/NCGfbB9gsr0HzngkLVCm66KJLinBErv7v/sz4hWMa2ipI222RgFFNPTnbEIYnEkNrmWwjk7JkUp
n6MVwWQL7hUHHfT6SWmWnNpapmpsWBGNvnf8YIzVYkOXSe6EbzDZqJZBdgfoeB6NTIPjkXy//9OL
GX8T9oDMniRBDDEu42Zyj/GbA0ZVSYjGVZsdlFnHyeiY3D6sVP1xME95TnsbKRKpQIgq80GVfPxT
fuy4bwRYeL+cBGY61f3an29vT1wQdUaYRZQ20pqwXkBxXLuI9fR72kMQ/nQ4OQ8ZIvWZXNFlU/Vn
hPUvXrbGFM2mBpkNc2WZ2wFxgIxfJAXU74kzQh3qz+crvqY80De4mPFvkaRqQHS2r+r8U32G2EHW
MoQBIyI0sypKOpRtWOKxiC9fS0Ah1CHiodapFUxuxaLJDTF7iy7FmmghxcVycwYvrOOf8d/YEZX/
ZEZrTEuINPuOu1DslGgASknkEKiE71R3DnWI6/zOscKepE3ECMwKLwQmysjdOASqzu5DaStZEplX
DwBEtk2HuQnoB+L6gech78U/NSy3YG9ZcYZZ4hCSynRty6aabFUpeQL1BbKeHP1O7jIx59fHNkUl
URFCr/X26oMC5ylD/vF7xkfU0BNk6Bj6FXtVB+F3JL5TDAzyQ3b4i3wkAbUj0IT6OUX0wqOUHddo
vGzLb4+jvTWOi93QMXmC91C+YhSWvHABPwM69msnuaXoF+uh1manI41tVaq00vKp+vOG6lpw89Q+
WaZoa2sJ9f2cWKaahCFFHFshgnokIszGUWR6pSzn52Ii6boC8jYiEw9U7/iu3/bIGY41RVB7C5Jc
kBmfZXOMUseJbAxA0u7xpBUJ1dC72UL648pLLmftKtASxtUldplFlxhs0rHgkZvtzasPVazMsMH+
nUNrZoUr5F/kknpJAgsGmAq9ckgP80UzNY9ARv0GiRCNtti3Cb84sf+cAp3wsFh4C1QGOhxnUc/W
dleF6cQwpdoKeG4PDqA1l5KsLBxZCdbHakYRI9lyOpJYnOtegWGSkvRgLPdZ019liHf7J5zZGiV0
vZjtLSVCX1w6Qz8/fNBoWIKT6YAmX0UTbmGtvgaasfMggnR+ob2z0zBs4+eKlz0NVuZNj960i+wc
HXqu5XsYCo0paqC6OpUBF7CBhUsaVqURRJsS/RYZi2jELkLt8AjawerQOq3++FukmuykDcFqlQoh
BC/R51GZnnDUjkTdLErheln9+gA8RPe1TJC3F4M36/ezekMP0X5TFqAPHwtJeMcUyYSCeX4r9g+N
YFPpCp+krAr63RCn4TmYmlAlg3qX78m/U766bAGYHokx3N1MQoEItHZEat1/51Uu5pu3XfjiVGCj
f8F+zNNiaDBbC8dp17bLKkT2BMspmV3C4cFpeRTSuDW7tnRu+NVb1bzDnNzbeMfYpuCL/l8ifRfQ
5l4nvLh+i89yy1P//GufeA5rjWr9W8032fBEEXnZTgZbhLOEk6O1S4QcYA24CIOfb7OgpKimmCPg
GjLYI+vva1V4DB3lkLbP7rNR7d335YmUVsQypISLp177CRznlVD1NTrG08cvzlZPr8BOjfuq9/sU
QeXOtb90Vv49YJoPWjDGnVsKQ0H7O0pb0jeVIxH9nW/e2aevMKE8AH4UWez8aGt3eZrZ5riFp8ZB
qtT6fIr5cUOpreeKFRXH4X6XHCV8E7vWhdHqJrE2lJYGD8kf1rNXzgoyaUYwDpaLY6FsXRG7cZ8s
R0gZ+Yyx8xRl10K+rusesExwv6qqrOx86tj5R2oAZ9IIWqd5z0pricLBMV2PnthLqZlttNzPiS5V
RI5X3GVuLUBRdrNRQJ1YniRpXYimGgshdDJf3BGgKgRRIFzmA0Asc/8afIFyD5SsGyanSSmZOn0W
enBcTscaZ2ZdqDmfJjCTtOPhF3K23AtixIegIOekfBn8NQ8Tpw1/EVQR/SjJPPaeT26qEEvshGjf
X7h0+KaYHQuyMIfp8Y1BDnYe8L/CW19168OYRO6gqt0HZX7mNIWOl199Y+LSkXg2E5fIoidXEUqr
GB9Oh3FDrKTjZ99DXVHAkq2ljGdajmCviaWAeyrm4W6MAtOmpX7JHXDWCnchSc/pPdmJ/eqWZW/Y
H1cWj0XMDEXNfCrw0JqHB/+nmKLCZR0hqoIuq4OLX8VuHo8XKIBv3q139poW77AEsjexNLIOma0j
XIKp0EN0CJWMDAMauecCBgSFkZNfbq2XVDmF1niw6jlnOvHRqCWHf4hIYb7fqNnIi6wZZyLOr6Pa
WylyPiXwDtci5byjCvET4x0AF7y+N6k6GHSFhDaaTzP3MkXJ9cOADHTL9GRCtk8u4JhAitFvdFkn
9Tyao/RuydDHjAt7eIOgZoTWzVGcoN+ewyh1pDw4qrY2roXfCqQ/S636q3GItBpKP021fVhReZNQ
VejfdavWbsUzWIsa121Dssmt4Hh1JZhdhZGeJibbtZHUewL2zuVsffi5tzAsW22qsXJM5SKjL3GI
rtZhm52vElnyvf/vg+gMjQylj2LXFSfC0fxK6fylMZqgrJVHf9D/BXXOGuMt0VB2fOu/r+8gaIJd
6lfTQjO1HRFk/4RULmmEt+/gXY8cKobU9SXiMBtSpAEOrtQ/cK4H5rur7Z4YX9SZC9m2Y3pR2iLP
zMi+6LTOK4m+rT5FJcXs3ctXcXLXDa0guoactEt+jfOuP7P0wS+ysLphzEGueP59RVfNYLUXf2IA
NTNixfsl1r+Flvx+6QH2zDieyYC+N4mWFK7jFkXgIR9GV5GA/7YlQ2KGpuIJoF83uCZMdGwqHINe
3Ag+vuQKi02Xf2u/+Vz4gGbNB14jwjitmuK4KgwUW3qJbYdTvPoAnV1yom2+kMnh8YLKYoBwbykv
S26JofLlKxnyH22Ya+RGMC+zvhicOMftYLytk3Xl7SZNIjRqNVK6eFZHIw9kvcUqTZlZchWFExWW
Y7/9HAYvSZjYGF/XHFTLjJo6amfDtdoIPqEgpam79KDPF4OeRcsfqbkz6nJSmKTEo41j4Yu5SeIF
j5UUXdcvq6ElxtECS7bGpxdNNz3FhgCvttI9qvumPPXNZsmLWCPhJfU0DYHNdkeX/xtHMKvz8Na0
Smt4Is+waBubdexzo+XVr90v+zuG+QIf7WQLrwjvwDvKuIkHh5gsPrENG8Od4hB2HYF0uvJnzDMf
XaYrPUbpu5zlaAiieVGzCPdSYheHF3tbWowDRvpvGr8eLv60EJbMvB50j9mB0dBIxM2kfzFWnOZ3
8PndR9CP5brUI+ZWsUt/owJ2BKok1q8BWBAZD8lsN+cuw063ZZlSQK1h3YkFN6uDxMmdIebinmQV
bkYsy/lwftSwVu9rOimqy8YSQKC3H5hV4DQPstKmi6mQ3tbyUx8iuQAlZRnlMi4RPJHMZlfFZz6v
9VcpB48h0OjwWC96F51HNeYWbAsqd7PZPCYX51j9ita5x22Doa4HE/ct9r23VWPiNSwjpdrsR7Mz
NsHBrL/UL0hz7CCh7ZoA49KoWow1KXh7L0Pt60RSFE3vmDtY7M9AXK/d5z5908jUFzfUm+AMbNr8
PNDD+EhBIZScN6jSTYsXI5PFpp7p4TNtjdM1uuHzQNwLmymuJHNXiSn/pZOVhjmneF1lZReNPqM8
0CRP0bnDjnNIOEXPxwgaZ8HmJGfMHDhrGqDBlqizzMYxtkR0ivwGjoqzere4CoGAxAF5W5TmbUwa
wOXl49zxApXA2GXWfJGD+SyNCPwXJhbYgiNC26PBZN6g0cHwB/7juaJh7Oxq4UnVc1dTBJSiKFLK
gRIZV19tKWRy5ZtF73OR4fWlbZ9X66j5vRU1PngfSYFHgS/C0No5lqAqw/FxF3Hj0hZ73yVm//kq
2zdj8Fk8SU120TRMMW0NXaPyuTLlqvxjEd/+autStDy2unDVu3tCMqUIahHWjnJmNpLPCi4FITDz
DD9kjvHS3SNQQ8AHUjXgrOPWq3lRkMQcXGeNLFLKZbSf/UdP+SO4awlN9jny2mpKyh7VgC2MN8Bx
gd0HujYbMxGsvkScdAEGu7rQmjkWpbv6wG+HWG+D4bVyygsGPasVL3jWP1ewGKbamBEz4neoqfYZ
6QOwjyrYdNPAoqusQlDgfY57MkVEIArFMUhCBv+6632R+bQ/2+2cWwN9XeEdAzfv/eN9v3K0/f2l
ZfvsFnypkO5trJxPHY21H9S5nq4/S2MehTehg63poz/+ekQKAnyZ+5RW/zVkZb8AuF95FQWrsPZ3
1r+ObnxtEDiLD6fX0EwkKEe9EwYE7XlV4Cv7RoM/prlCYrYYtbY9JBqi14d4teEyeUJqfUkeFldg
v9H9dupv1ZYMLGXcT5S12TRV9JFFMAdQcIf+kxENeRm7SC192EtZlW6NY+jMgNqf5JB+rIQSBGO/
ZNNF0N8bhzDGcw8zwzKfEQOqM8c8z1Xx2MpUdeeVCYPGysAyc9h7QZE9BNzpJLoW6AbT6qsYnr6N
BO6rH66VcivwnNvnm3G3bD9VrFEntkYUQmcppiJoNBBSerevFuYz+lcSH3AeS4YmNVmEQpngn/iL
Aioa9gbb8fwBCp8ae8gBTr+mri7FPp1OBOW1S5+PzXDQZRBNhsEJRoZfzQZSP6x6n1EmxzE9pQj8
Rms7kWE2ocjDj+UydD2hBwwZ3fJ+xPZ/ZNDABYdVhs6j/FMqsb4TqysMPoP4HfJ9IDURihysV09i
7zjZzyQz9L2XtBsAp+xFXqo0i2i5ObkswjizCroOCqt1M8fidqeLEQFuBLgzg88cxogZnH5KEAQm
mJS/41S3Wx81fMnN4uXn8VqbO0CA9zCQ85hespTCpqBrMtNAhZKH4XQKWRYB4ggD6jYahboVcM7B
bVFG5LObLG98Svjdc9RuJmFiUs08WUgt+UxArGzCQ3NmOjKfanBKfYmsv2OvLyU9uNjAWWjwq1dx
w44Cw8BzRBGETJn+PWsb8yBXFUT5BvCq3+Yzy7+bWV8hrBfy5Uz3tNiHnCELscx7WsdLSRtBKltD
DLX24bSnJGz2JD1iNzwHHoCsHMIdusyTmqud3CBUnWOsKm0lcyr9Hk3hYR5AtHxkGH3cLDq4kcSH
ESBDHGeYs4Snu3BmIgy1RgOKN8fo6m+ONZZ7YNXWmo8zQBWb6o+IqSDDJ1rLl6NNHw9IRsb15CPD
bXrTR5+PyBhwEjmh3K/xR2bclkAzdzzw6xAJld7tOI9ahEYjOPxYmQRnIfOTFhCnJkIPqZpXwXZc
1YS4oDEfuWg4pJNjE9RR82yxKt6yTH8mXgY4WHGv2bmGb3IZXh9nghO2oQOtwnf0luvriHWIA7br
5JMzkiFae6zK5gNHrOHSzuGKd1Qfw+H3irZW3FV4hoWMliYYb8JC5PuQ5wru8fmgWrQVuu/P+tiS
FqsOAVkj5MbQgfVVOLWsSLHC+PBBjCipR0mx+LVRgVo0tq9WHF31co416vcmOSsSANatUJPEJlXy
W+TgCl3D1yZP6bQnh60xfG8CxPeuID0Vf3nkzO7nXkrNdFX4uB8BBnrSPu/IrwURuhwQyHSnmuM7
U7RdFJYjr2snWiBCgDzr8VlPpDKw6/Z12N30SepNYnNXa72vUsumuAOmBlz2ndXEXj2sYO830M6Y
38GPlQZg+fy+kYI0emjz1gUbcD4ogRTCvh59+civAzCgy919AHkgybbZyJvmZBxOjM23J7u82FEw
HPgLvgFuZrTFkQ23MMyMgLRS2Kk6qWM11+Ip5KIugD2PMqXwUREJBpmdaXKuYmUW6M6m8cj/wUHh
lYTNx12FQ/37ZVIhqVEh1T9w98YAbhH4B3kZZO0N03q7YBs/W9ATH7LCKRPR7cXJDPH3h6S+xf7R
PrQgk5Zduq9OJzfuUx0ws0RP+6ZxpOv4zvHMGIethxcSdZhBLyHFgMTXIEGqIHytSLVlh9twgt/y
zhmkBhJV0wh9Pg4B+7Dc9HzTskkftPCbW1UNig22Jp20n7wWsUyWaRmEGQT7BRY/TyGKHPO2ocJT
9e7jB/Ot45qiqbvsjKk3uGsAIuwGBFoUqwAx/NFpYnxiXrF5zbJ/haHWoqXmgXuqu15uGHOySMyU
8iYKxdieSYg+PQfoVBq5G8bI5/EuI68PUWIjbKnEsETaTWeZjSD1SMawdE7WzB1SbRCcszOYHcrH
RaNFEdNnkcgyv/SviNB0GTAr36EU9tx918awYFIdPOtKlgKM/6uV+Ac+StjFbDbBUSzOkDhA/PHL
S7UrkRTCkcNaMmheWzxDQEC3vpHr3Xi84faFVlgeV7WN/5Te/khf7bJHbP1GiVg+R2YL/Xjd5wvE
fEOudkHxaSE0jxCBfnHuoFCMr34nkZp4KKJhWsLVfyzRxUEO0RLsb/bdazNL55pcDx0L60hgtONR
zvwMG1ZJebqpby6N93DoAIirsymFoZRonORaOni5AxF2duckQ+kJ17gOHfpnECG5Tfqm2e8d44oR
6XQH78iSl4XFX5xSGrYoCfMmdhMRDluoUeQc4x8CjxC6YfyDLe4N3A38qiqHKdiGGmaTPdGzslMT
xWjjxVAT66WdUiQ/Nn9uR6qAFv3KZjXYwhB2GR8x6uLTSt2iGe7hhaux4k85upWCK7qfE/srQXEI
ptwIVRenmyrk1RSypEZGTn80HGBHUIHJh/K/njmyAbD0+XBiXgaHiq3qVzAGwkk4Smdj2+SyqbE1
Vwl+ltknFnN1YYn+dNeRbIfhiwb/fiPS6ijxkUcRbAhJBUoBpiOKkn44NfPVHC5xg1qenD2KT7eG
3Xu1mKwRgwehK7xSH4eTBNupOQ3ewlpb/J7oZjWc04pvraYyRn6dR5p0UnuCOj+HRosTRCceCdbx
NbBWO0sRMdPrOiK+23xi6Eua1J1eytOR6S6g30wfM+5l92ThaFVT43qIpHqstnsw5qXYiP/h1zbO
DnbCNQ6HxHpApi6Et/OMtyT8Lnwdt5es0tazB6U7o6DwFb85wC3l0yk6yhqoU8OzV0y7tpmI+TBw
AHvtc4HAL1j6sI7PDrCg+sjGddTRGB1q0zp/W1YuSSyOggF184lKcftKK90NL4qO7hoFvRQPQIAH
jOP25lnAaXlJCZ2Dd7b18p3zvZF7ta1NkWj7dkmFWyCc40cDH5TwMK506FI8Asquq87eAxV/VeQq
qF4m+6WMdWvnOvJCZCKzqE9RnhYjdKVnKHAmMaElwDdLfK2Xb40eh8+SXcZTAEs2ZcHVqf7SRGjC
1gR53rNFQy9xP6CpofJ5TSA9jmuKbQBTeZ3AFC+ipaWH6wvIP5w34darEersySWyOoXyRKHBgD76
ZOtbV7QEy9M6fOLwjMBXoUNZhBvynLhfJ1eoQczrMPVdVQmFWPa3dIXHLlpuWIp7LGRhQorWVoeK
eq5Lh1DIILyw4NnnqhHD13+qdvlVjLV+JVnY9oBr+mlXq6elkW1CoffvGfRKuggT8PWi0HK6vm8s
/4oMD3K8W4L2BW0V+YsGNW6VRmOc58e3Zu+9CY5rnuRJlsY8PFAbfVqFOMNF7VemGAlSSGaU2+tA
UH9aQFxAkR2tsKDG4WBxR475ZbwN50KB2YDD/whODurMtb+DZzopPpwKsGj9e67G/N7lxXcPGPej
/k7uKdltgDHw5v50+c5kOx7KnFcb0yA8/1Gj5XGIwS3kb3V3yTRjgLRlOxvaorinkOtfagFIeCBE
ul5HG78ga46xGGy5Fk08TOjomLN22GyYiDmCYiqnbq8OhtNmF3nMvJddMgcRo7ea+om23/m40NxM
+ShR5qzPVhWUYXNVjlFBKlfASTCYi4ZP4gle8RRMSewkSwfL4tZOmBt+e/yTltwLzoTc3ETCUe1Q
P3kVcfrOioxU+sRxpuWzdsWGRZfJhdxIo+gMfzfQGOnISRmpjAucejWOeDSW/MCnWdXpilCqpPLx
4ob304ntW82tXQB4J+8gmldUmJw+ytcMkE/aIykIIkwUea5VADK7fHguesg/bSMz/EcjCFi6HEQx
6zwT8D7DN/FFNPTGFIKUx3MfUO4JgUI7rqCqh9T7kaZLQVZPY3Hd77BQdqW2reHPfTqxB6twRUsk
lLeG9xoFEcp7YDJEt+1K4Ut01/1VX2NLLD0yXy/4h8C1n2Wmw4y5OzBJsuwYUP5xLCtwLo4ZAFdO
0ZWYRsIsVy6bA76RBPcpLA5cFXqdQxv2Ktiva1zCOpQ0M6XPZrtwcXfeKtTlDVagJj2/+C6feezf
AyYS1K+IjzuC9b9ZUumGVqtbcnTcq5wc71eMf/pHFAogsnCXgn+503Ekez/Dmb7EJ5YWGw/lybq3
bZBvf2U/4pNL8mqagHpmDEzSSuNZ04bkAGl+xb0w1kTfGpb9D1UIIOZAbCv6R6aMuA4/4qH5d70+
UGRlj7ut+0JDNrqeJmybYmcsRlR8qOjHlcBvG3BzXkmAy38D8bA3iOjw6dMPwW8t9IT5NvTFwlNr
2aJ/oSA7xPF3f2Uv/TyvJf9LUQXD0JpOasSYBBjriAGDO6xtBfvvtfZK6+juBdbuGxDBj+eWrxo0
XhuQtV9K5BfI8RFwyN2RnvjpOX0S5qA57gmd5vcxG/0VLBqfftOKy7Vy4RkGOSwUYMBHe2EH2P3c
a+i/TU15YHU5rNFStAKFLl0GI3wsEc2UgRQTwTtxKKicY80gTPhzYXwfNefRiO3DTchFU4nqn2+B
C55TnLWW4MbrHdGVjw+6YW8CecmgWjlqb/I7ZFd5QPGsA8W2jwZndcBXlPc6/Eygwh89ip58Gg8L
MXuhUOYhsX4zzB0lu0SefSJc1cD/VVtMiDBPLyZJZwUFwx4Ftq+GplEfiGmTM81dWjoNuds3Xpcf
VXI5oAqZgqOUQG5ZYW5/deKXA/5/ocblzo3tyg04I8OvCVI0RVgVlM3PhxFnMOtY2cKrlG+4PH8z
rinngwwGDw3uSSOBl/ue4Dn7KTd41XmVHCapi9gXK1EVvsMgtd2DHgmldkJbrgYnHPxBQFzkkFQh
4+JDkTRDM/XOaeGfAgphHh5/AyqfyL/vtxNy2qrVeNF/291vyqIGKOBX1s0jJuGHkAqQaV/SgIM2
WFmlCcaJDn38v1NwDKo5KXWXyyBAS8Ly9nNukzeKC44WjXpiOUqLmqAtPahfVNFTUd91EhyBKdoo
+VNvv+yiy2624dnFudsY6/p7HyxbVVYAAP0Bj0YCyYrMGpD65U9n6Vngs3hG3ut6MhCpq2jj/qfB
olzUeu1Qu5VO/8bA1uVQZWXJRV7eVkPDlSbGrM7dwNEfpUgWUk4gNnePJVf/eeLCeGnB4FeTiasz
o8a+ozaI/XQjLFH6b/RSNxQ1xWc3DuDV6b+ynD4dsp5e4aaVBYO/Q13oJ2+g57utiGav2ejT4mgO
aqyNvllopiMZ3mlpTyB2d6klwxwSnmKUfRDm+sgn54A6CovL9FNM9HuzvIFDuJa15QuL1wUNy+Bb
aVWOgO1D1rrb7a6BkHlHGlsR1iAa3Bde9SXLkvpvfUdLTMqCjW5z6qZcN4R+U/sarEl+h/q09PSB
eitz5Wbz9WvusIcD5CuOXTfaU6TERXJrRinn16ICtdGTquukiYzBgRT8cOgE4WQZuhlq6U/aERc+
cbSISW98Su/xY3J1/ZFNBQe+f8XSzPDEKtKKvjzJxZbJfXqAS30v/NW1Q9YPtJhfAKChMxxSWwH5
PTx3PHi+fL2x9MFi3f/2VqQHwxJ+SNnyeugotIEj0bhcqO6OZQyGWoTinfR0rSjCB/vhR58Kqs5R
Iy8MtwGGY/uDyqTFGFC0SHazAA8Zt6VEpzNr4DMpKU+s5vq3DUoGjLmj831sgQ5wRIMzikD0JFNb
36RJI2j+nwGvCvmmIMLqRJpfGbdxwdYUlCcYf7kP47uqlPLmVGVc/AR2goJU8+BsilOJVDNHHTHW
fASjETTcNzWvavSImRyXaAuc2HBS445nX1xLiUQau+Fst9MMMgsk8OvfvpayNrv6fcPIcJJz80Qm
LR2Bh439BiyL+g4Qsp91+fNAsBTr/YDYAUe5scxeuykr4DudAJyJXD00tt+hAoZIY5HASRMVbIlj
PmxuVhhrE0zQWAMfsXX7KKmN2e9DA35wP8AXoyh1aSPOOyMa4Fu82TZJpKwFbf1t4+xM/JDU4snQ
T3ysg7vzcA/MJQGxb1iDNXQbswadQOxGmKDwPX5d4sRfCrXyz2tljuYllGAYQBnYHiUmRI24jd8L
/8w/aRnu82JtF2CPWwKPMNglBfvD6dPNQdSXHjZpZ2K9QOD0jgS36KcyIA5DiI+ND0+eJQJgo2Qw
HnFpPGAdZhf+LVkoa/4KU/rXQKzpsYA/LTCYpFPV7Wu3vCuBO3RBUG9rCKFyYvVNfUPz5qW+jFW5
ZJR86iMqP21Dq2Xr9+a6t5UrVzwXDye+vjYq9XL0O2P7k+J8/RBB0Uh41TSjnjQNNRvpl3xJStV0
ViJxtSNjrknUOrZe8C2Ul7G1wH8am0yHDzbmyMylKbRc44Rmb5EzyBdtPx8hf/nsDhTJQ56niCHf
r1FGeK2yVEXWXV/fr2ui3pLpwodfqpmA8YBXYh+1JBA4FN7hgsQi4xBnTRgvyEP0+hbU1EVUel68
3FEvfWwNpnRWyBx642RgBfYprhxGY2sTKG8qTabkSfCJi365S+DvxVrv4SScTdmMyrmkwl3IO9X9
HsLUSmZhPHdwO5VUvVJk3XOxW2W/QF3uPxclm/s5UN+ziIPNCKXyICE3IRybKtUkub++lVoYRSMb
cF1WxxVoelf16XSKlBI4O3iy/m1TSz+85OyXPbkZ8fXQSXNxmnSy/+EEMa0rTnPvCdtg18MfCYaY
GoUmYc6plF34qukRACws5K0/cfPGaDmeCCT9qNM0RuJncWC6NIA0iAHIXgKtiUje1mrWZqjgczpN
SkFFpuxugbRB0MT6rih+gfvciUq7yU2erE1E/S5TxRkV1X0OGHud64A3OgxdXCMF0B1s+ge6sBGB
IB4Cmb7eeRn8qJvHSYMqQK6FLEC/WK4leJukcquHFv93Rdfv5eF0tcA6nf4dqzL3+DUg/3qP1KEK
jr25qLhLs3GfA/rCFclQ8qV/ND8TFycubDyRFLNIVgZEMlvvwoOv/O2jgCSgNMv7OREEpZJ2MRgh
d+jo8OmztC5izHU+U019rqPLppRRtBv5/WO7gP5kkkwXZAviV/h1QyyLObpIkYSQO1eIOTqeyun+
oKxb9zY3nBie5BEVjHXvVZgv7bUnM+GruycwtYpV411n4iT24wwHfH7CJqHLtX/OmoJ5WyhhUnBB
gefSGZYHFaiDt7nKpTzlmnc+QkATxHr52zlQi7NR+ZHqvYH5aekc5u0to2Vdelur7Df3co3c2Wcx
k9jcLo2L/LMpRZ1M3xaxvniavvlVcgGPyHTEOQ+oJlSfY86p8Hx54GqBvEeJ4p4mRoas+hhnOmAe
t83guCSuNkhmD0D0xM9Tqz+vAGA6Vr8Fctm/twx0SnqpQtuSxG5/zMc6pPWD8Z2ZZGcKjRWoBrWf
1S58TtAMkTqkiNS1zfZb9o2tJmuBkj1A2jdHK9c5f/5EdoHBB7ngbLeRawHSOrGurWRdG3Ld4h0+
AVre4fXpyxfaDv+q2u2Ro/ALUl7WriWVcVWF83jEBaU+pxvQeBPrXdgCF0BRgHiwctpEiRstTeAt
BOzaLfk9kDjbrJ7OsYzHUlWtLwjGWULtkT2kF7ZQzbI5fNFKW0Dvu8jrbN9XautlxGLIdztlSh8p
guxw/QYlQQT1KoVEArADQw88NF9q+i15pClecmA074kQrKo1w53rff2eUT5QukGESXQAF4UQi+pH
y6aldRqYHM/lmPkHLUjJ8XYL08qRp2G/nUe+qefP6rbbq2CylwlPCKU86MLV59YO4VeTMUOAszAy
jaMmdvFjArCoOBZU2wqyRv7ygkHxr68W+DxzRZYYE/8JMgk86od4j9m+NFYEIaT6uSRwV5/a9hmv
w8kMBtSEaOcZIiQnaoA2XzxyX4WQELivqx/qDzCCINat6PgVhbIvwd5Ef4wFZw1SSKrSZgdpDboc
lFq5RY55hBjNEgxdsrBN71BUhJLh6v457hstVUFy0I0x5NxrIQwn8zLYEH7GB6pJa4V3WXukm0/m
K2g2CwV4dDOfseqTSTPb0rovfSZklxsKUGdg38odocT77RbXAcPDbu0HmQHKBsI8JxYg3PzSzwZs
Yust+7uMd/3yzzdaiJISCSf8YcB3Lc9djWSSe44DGRVN29WrcrudMzPzjxMJ7PdVSIXPZVJX5mzR
/PPdPWNELHqmIVzjPNf133zUSZGGh6dQRYnp2ukmSPh39Ifh1WbvI7UG4pzjjdgjaDhZj8rZQhU2
mcUwHKAyIltb9PEmJ6xWXgcb7iAm6Kt6zI5nSfD3NhiOo8NfZa7hNONDm8R9mfp5GDZGQHdzxGN2
y2Xv7/CnTnDZIpF5iskO+jG8LZXg8orEarjyyfA7J4ze4mWFfIIxPKnteynezOW0Qyvl6JWTPM62
uBE+52ZJW/bCG+sGeLtWnKS20BOpyJtDvf9Rf8RwkhcAX1wvMbgr4DFKeb4FunftURaJyBfzaItM
QlmT/+36ajdVMQreIuOMkIbDaIr3hknBcbRLEDkB+/LmGA9xH2wlIbnAFrLU3ZWcnqS52WJ1Ziv+
+PLKjDwZkw5Cq0eyyaBdUMNlsBkLoXqoezKIBCMMlIublppWmKAaw6DRrxHIw6ur/GVCu3OzDVP2
txrxuaCE/GoWTexZwaGNCLdBb39BN1aKCa2wcO0ANs5x7qxi1vEBndG/KNIgdsH2ZSNKITXfWZY2
nd1DAxWEFUB5zBPnGXttTDZ0thSvkptnrB8GLELVzw6t60Ml7I5L/a5kZfvJDj6RayCZQojLXDxO
csfwgY0p0Vvf0j6GuybTAWBM7vZ8Bdm0gPes5azyceYrKwRdvBhDXgYQ7rl9Ix0t6EMjaXwTVy4i
wl3uoQ7Uu8DlHq8ez6hX60Kec1WaOwBrN9ny7XIKLLMwQinSCJx+MuJeTLQcUHgqOdqHjzQE+7VB
m/Ugv+SCml/olMQ527kFJAzghep/i6SeyrC3MYiFIvhI5Rr71C8mFB8+JzoFuQhIffhmklYADqBq
3xnjhsclg2bo+erxo9Q1sB3zY4TTokyloaYaTc7J3WTxJpWFrKc/GnIs946BUjwUNQ61DN2fg8XJ
kAXC0h4/URtMc564iQigrGgen/p9fMcKa5Ku3xgpT44ej2ga+0oLhOC6Avb5AkB1XsWhRwf3ZM1k
/OzFqTWb6v+sb80aAFta44TwP0C2/ng47je+5Qi6bvR/ZH9FmZ6g3xhYK3Wn620sAicvU5YDWAhH
YioGe6PHDFaCSN+dcoIHLlYExek34e5w1Ys/J7SNBxog4qCHkDp3SL2vhKhHDwfiNViZunLK38gD
yhxpTQDRKka2nKpQHLNCBYaHxH3xnv+YXXFG5j53yIqBL0Hauo/Ggv1YIblLaqbjZerj1GLxt4EJ
H6+ktHNBXcYQ7nykVyduPsxZ3vtAq+HAdt04/YlPFrxmq8xqJhDLEqR4MSSMImyQa5KhvPivlIt/
/QeHuFIlP34tAVKmIkm2KAcm2rbFqgga5Xms3JWL73dRZ3ZFKH/H2IjzeGb6M7ZW1r+MzHXu1g1k
cqlRdAba0A/rIllkotTdkm9mkevWGQi8i15TJ2ZJubc4xR/wHRV9IghafwRlcase1heFC9YgFELh
B6ZecWkzDQE4pWNR8RSeORITNfW9lgeTsU+lhthby62PE5Y9YO3J77z1AjTz8KCcQV2UU5YRG+d5
spLymkLTRimQcL9Gm2mpdrszWTkbo8gKyCIo/SyBzGP4XX6Rq8ce/HuLg4I7G5y1BaVUsK/e31Vp
2Rj8oYHaom/AQ4CdcmWL2Q20DQYdpQSRKDsj7cUiJCb48+TzRpmHZvK8/LQuHDZvg+RIMVo/fI6i
PXfWJvKZNMK4AAGLReymryoQdyF2fBlv+XawC09m/bjXQtNT4xNBPaJHqFQpeBwNnsC1l/gw+Plm
CdiBF8Vue9hDI0tHg4676kVz4TRKwaLHDskBE5t7rqsxRhl3tF0A+oDOwB6G7mZCMnJOCEhhQj/y
A+z8G5lMMJfL12QKfXMURZYyxdmPBcLtd91H5d04BMzVsxfahch80T9W2gfTpiFEz+R+iXORR8E5
b3g5Mgk8FJ2svceYtlDjnU/Czgn85OXSyMKVDOsq2zf474TEB7ncwjXbO4v34RgPtZvmqnzh1lZK
O5ngwrlQaOfOHFrtI3xopLB+xfEVyq3aPGytcrCt6RrUQ/eO9pDLHc6qFheTZqSOvGyeALB6Igwk
x/bmG24b0EMsP44iqEoeEPaXsnfdVenkTnUE9+gI9PucgWdbbjqxKqcOnPoKh47WTVDJlpzo29FX
xXxxPH0EkWCzHAxP8xvRJCZBYdsKL8N3J+5AGtmJP+8yJjBYnSt7eKOk0B/OTBtuzBmdZ+B8OG4b
vtE2f21nRLnsNlroG2BXsitJUL1u28TLWZeOeTyoeolCy27XdDJXJKLY+iLjGzzQf8JKP6U3xwZo
QGZmkoVOmRKmwbXy7MsTesqKqLmWwJWEaIcDajHjaJNI3E11nYNLcsBhtKTGf3jpWG3oMkjsstzE
aewR+CnfHaN4DBuBv8f6IjnOEjw44KHND431FgAvtnnh58sFR01FvvM9HvwhLBIe1S5cWJ4lZa8b
ukTpVm5cZcocy2NXBG2dntAol37R97Ept6nKAZW51Ux4lvZp4oMA7Q/m3qkTrhbMqNb9B+q3V06Q
nYGWVwtx0IQDkWXEkjAeVg3HKTeFQD+M9tqnAXIeeQemWpdNNzhq68m948krBCtRCMCWChZs5upM
zZehkJA1TegefQnuH+va4RDjsMwc/06URHxAhMrFbibxmsAKjsaFDRUCu5h6HOtHlvtFJyNhJ5UE
MKRFa8e9Cr5ZL3ad21wj7JygDkSNgeaveKhpEX601hP29PQI8xQvCcAKZ+QzXEuqXOdjb4NYGa1c
ArZQiWebhUFtHzGJIi9P9ddPdqS8HSoPWvmA8A2T4GlzHHfJAcFOeln6UVxNOvDC7i1Q24rxp/Wn
gS+td/sQnBkkzyvtxPMcYRjJbED2mtYl2DDafctm615+IhDkRWs+TNLqWuXRJ3oGLldqrkR+ao9A
rpdKWzEsAtYJg9bMYo3d5IS88Q6G9+BVGq5XHwDHyuLXELH0t41h0csGM0sfk0dsPvvs0IauvhDe
Hec+rJz3tQR73WMlksFP7tP92JSSsLqszB9GcveXxI+6EfQ0FcT5cllE2+LmFjxp3iLbpkwKjfwG
mN5z0Tgpkzq7wA2Oz6ap4EXKFOwhHeS2CO2MTZjCQCJlVr0DI842dluLNs936xKRrVVpBkWSd5rA
l2sWyWrMpN+uOdl4d7wHDd7/uZMD8EmbZ4k3vaudmxypxZi+yNftMpKJz9QfOjqhjVTjyIDFPXcM
Rv/x4fgwdblPliWuUkTJXgKX9TuKE6mxn3ncpt1df+53HYnWmCWYlc8+EtdJAlrYb+EvB6oiPCHm
pYgGqZT+ArJxuTvgh7Ext6gs9vL6ebVeJRm4JkD8xnMUeNxXO/RGZvlgdzMDwBK2Bx67UWNl6gE/
hZPb14uVLcp8oM8vbKZF8lJEopSQUPWBtLEwEvWnawcl24JGLsyBxOhUt3/OmdXJ4upEGX2y0yL4
CMk5Xi+WYMBEQI/eyyIcOi/Ah7UGU1VbFmpww/rbBovHiJGQwr0+nCXpeU8BaiU4rSbdT9Cp3tUL
HLhOjKJ7lS/MZYvKR7TvLuFWGNpz+so+epe+DddJs9DcLX//jvYzOCcdFfKFDc3ip6mJQ3V6Y4th
0C0XBQActpHozCRxZ7oRdchFkxW3d8fS9H9RSvfaJmUMw/SoYlHIf2dbqQ8u83MPcoB9nmQFgRS1
laVKOptvbM/3czrk06bbcPUmB9/1UVyUq9A0ftix7RdX5utad7rAreTipcX/JUixTTDQwDiXFtbp
jnhnDrkQUEgQxEZ3EKlzOhv9welfTd/VfDH3IcUPK+jBJFZrf3k0XBaOd2vDl8syAgXUr9Iz8nxn
lNkvrN3VKPzbEW5LQXb+C661/ApSlxTAXQMmAdWVlQtrbWqlalcuwCC2KuZ/5fJzoh36u8XEUDXW
Wpvwnowb6nBvBrky1BUvgmLCYvUebct4jXGyhIrvTIYN9qgOlrR6d+DV3CVXYa/xQvqtYG/BpSX2
/hVSPNpP56gK+TFQqnYWq23E3967ZcHEvNXZDR9NfHfVEBlixlQASzhPXvh2np+XhdYv5096Z55D
an4GSICmvFr3cAQbQwJ1c30dotUOvNcI+Nsr0shw+KC+SrfAFgy8yaH7yEBON0sRsoCcbKbzaqBs
w4w8PE/OMdxNiIp8UjHs4yJ2DRVREPmkPZ2YB8MYvNi3rdccHAmjClg0DUMEIIQmkGjbMgdwSB2D
hGJ7V18MEROw4XDPuzMLsxq0C0M4c9EbAnxk2iEbwBpAyAoMLkFovJbcOc6JRDXK6BRW2UgtGrlg
rC06mWsFmJf0Uo+RwewC+QMWdzudCVyrkeWmsoaEQ2n6dBgubENDz5rQsU4IFwPXV1bcpmDlt+7/
UWrQOJKaaUWbcbVkQvKTjDuMU4iFNCQ5KGQExlg+NUb1m4Dch9Av72KIdSuGAIKyEJuHDH4ryEcq
KMybLnbIBbdxq9KfzaZKU5lOVz5WnFdhs7ez7Ml7cx33E6ZYLnszN+xHpBgjUkxPQr7XztRVVwqk
/FksrheLlLQsZInp3ixEFgeCcdwzvRn07YHN7l1+0fVLOHfU6OtpRgJ2V7Mpw3hWb7PhV21RXuOR
61eWuLclsyvdVKuWvnQdtbpbLhY+JweROnzJj3VQtVkJDqraRgGC37aBqnJ+zTHUF6UdQuZG2jEr
EDIQwy7QpS2gWPiH2O6Rpl6S05GmVAgUek23CCskCHyflOkkB5x4jb7MRxIF1B+yr0zPruP147o1
l/cP+HWfl6eQd0B0QjJjZEOEohAThREfHVe4Ur+wk2tJOgPCvc14A7ekbKNhTewfDiKGzrJLYOcW
CmJSidDU/TwVQXj/1WhPn3xwgy99LBaMup6DCcKAp0clhnUR+4Z709GYW1Eb1Of31gBmK+543816
hli9c0++V17X5Rnx+jG3Pqn6Und8NyFSJ1Wnof60fMB6MmLg2/LcTJFE4YO0NpQU1D0NfHj+LMQy
67xOgwFnPf/YKpu+iaFB2ApRxxpqK2l8KEpkNmUraBIcAkh9tUj8wIdctLHZy1BCoQIqMQWvFnDt
JEWPwYlkO9loRaBg51ZMTG9trDb7j+x/keRk7nfBu9qx7pNhi3Q0SFDOqN/Qv2GqfmXGLO0MHhWz
C8xTPshcXEqSiAac4RiNLsTO/gwpf2Ih2kpQ1EqItQ6yv7BO5lOBp2KF4QhEkECg4/CeMCPqIV5B
Z2kJVj2T07dFOK6O8n+9eIJ8ACP3OPDNEyfaD7MjUoNkBA/g/gx2e8UkbigZdpe2iL2j0NrClM7G
F/iyWagkUOcEnFH9SbQvOcJ37sAVL4ULP+eUJVnjv6+u5C+FHVzTiNGj8RhwOLPudlWXbNaD5WvD
ulNh0xwUJM+0LyRJDuhw/qfBrr5oUUOiXGG6M7fIzx4Qrsvq0SyeObUirGldAVQN2K+LumiGJptX
oIJ4p2PVXmTwsJCpyPcAQ/RtruLDer1bpBM7I1vCyIrj/gzaTCQGagvhkcVQbMU7P7dFv48yD+KB
p6tG5+qhPaEKXaNOFEHkumg+P2NG80VK9G51nw29jevOiVoizyLwH9Y8FU/ykiq3WWxfaARufQIq
eubJ/dqj8yXTxBsaQDJi3qF3JRGrNeHwiXJw5si1SQriPO0M4+kUyIKzTDrsjIKF/0b+bE1p/1gq
dxer5voLoZZrvy3zJJ8RxF9oRA8jTLpleYuh/9xP/b71UlC/eN05Z8JUI/zEgLG0iaxA1nCspGKk
7GEwFlVCR+Ufx8KycYInCNYopS/sAa5PGQqmzyLWvkEE77LBZHaraVD4pM0zHwgvrFZ8hljQOaE4
pY28nb6HphTRpU/QCInZtEzE90ib38OWk+ydPzfCiCdCYeqb2TaTXKb9Rc+QXYntNrKUYuHiqO0I
0X1gGu3N94uCif0FJRRrAc7v+rYpjEDZMqNtxdL33nXoQb/8oBUQDhcO6Ax0Fy1YU/qnHUZx9s1c
S6w5b3yOmKeZfsXZzmk5FbQvrWtPJWwGKz2d5BEj8zAwT+ZVowVTNsVxtmUVsVUy+F6r4ZNi7cIL
6qNuhn2k3Fh5eAqxnN+XXMt5RfOzDrfZdn4/BkD6ACYr/XjRCsr9bspYWpLQlepZNww4DDweAfni
jLE39RjCXWH5JrtBIK+26vzkS+RxqfiAg9Osgt1gV6Psswd4wM+z1MIVo/XbiNG9kdtg0ryejMP4
uABmP1ixNLq/OGkzBITG4VEqNhg3ftAp5udCPdfmSZ/qzRWQdAXguEkPPclsSquBsUWGg5JEHH7c
346qVIuiZNhfVX9AfJox+66ATsXbsLzREvoxVBuECy3lk8fJZqFSqxBDAz4+E4qW55J1MqAKGEmA
hYD7VlrgbbH/7w6M62rJ9l51DdA/iD/bKuRJ5thMnRs5tDfYolYSlTbdLEvfKUXVVXSasWsOXfdd
dcEHTSXZnnduMACeu+6JJX1R6X/wlPnOGPJL5pMrFR5XrbUjlElf0DuG/u1JtPIVMAyT1o49xop3
KU3PQKNZu/TebcHX7pfhYYsvq/AUDUVUm+WhjURrXCfttnRwLuguFpITH5UoEiSpv0OebxsKkvMy
w9tB6i8qm4+m5NOxzSeUdG3ywMrtBJxOS2NTjfE0A+GZZalUapuKsS1BdE+5InElkg71Ploty+xL
BzjTA0wtfM1+o4Wk6qH6qJtPCJCJQGzFdRwXwyEy7ZmmsBgBtjO8xIwzm5MubyP1Mn+UZEXS/xLg
95hmyUKBhdOVqi3UiEa5LsFdB8jpnakD835EPiSbynAeRJUWNuEfWWaWajazbf1Ylu2rkhVRvQdW
DWJ+L/DeJhNuHu5F8gr4DRzG8NV0yarOdkjDSLYd/ykLF7B8GSbPCui2E+61NT5pD+ImtKqyqrO2
IrpAV06eawDOMm4cp7CSnMHl+MMi3YS5LhB+ua9yc8CYEJ3/6HA2/F0pTP+2fFMZP95swH4hk5IC
0rtdvaIww7RxgBvWyrFtx6Gk9aWK3byahMY1bmtNXYS7Qa1KfInErIUcOMWJHHUfvZ7uiNay+GWj
w3jGAy/txRiMDq8aTNPFvQtwboVZCoDSqnNzqQOnqu16qEYCPLrp5Ep4mwx9nXkQ9cPgwOaAgwWB
8UBofk+OonuVSgwH4IrMZ0wK4ZnRks8QpUi1mXDW8H+r9cvtVrIpQQsy3GzBPE/vsTCLgf1Ie/N/
aNZQGbSqwu4E2RNP34rqzZ2xme4zKPgzNUbWtSYc8ZypE2zrcj07Lol/N6MVW3xps5HaejBnYIn7
SDzGwZbfObl84zE3frjqiI0+pxiDzkKYUNnQwGCrAN8JBbU3j9Su4KaMng3pE6zakgAwzlNV5Mkc
Ph7rnigqzYYXj+/Xh2w3daPpmMjFJKstSao+dO2PQE/q4UfbdiRqndwg7nh85hdOaRdS0se92BYn
XjXZvE2X9Lgg7BGxjegyPXo4jdm0nMtxOwdLMI4YoLXKm9pxxAJRHQD5xW7lPoOjjdNC/dUfXoYq
9ka7UR62zlzodjqvAQxrcsyDhexer/OTRtQaGxU8OVx6qghu0ypgbEPyi3+EF6vMaATP2JMtrQ+j
QD5mSnC/ofx4nsgVnX9/u4UjU6Q0LtzVeEhRGFYnBtnG8xiVQWYJF5p7Lsr3imFCCM/OB0Mim9Yq
Z054z/o5+gZ2WKhLE7tB9VQLRnZGYni7lSddL2D1HRcNbakzt3OJhodZBXMi/d+4Ng5nYodNGwjN
Det7bu5doznDbd31zEi3bSQVskriid9u0IEr6ZCPq2jkroCrzjG/5tJo7HM10aDFx3Y8WfNEGJW2
xQ32DfzWiBeCfa2fRGN+0KixzGzQPDFfciR8+TUhJP+wnfW0iFq/vyir2zukhh57j+4K24RJsi5N
QWLqdv4fgeUOuXnl93oJ8/FzZ7mRGmoR+sjB+FHDOAtT5Af4d4bIet/YRPTpV4CAagW6QeX5fpMJ
mFda5DIFI1pKHUnET079YMcxZn0b/0fqLFtquV30e8ppEpm4+MXJD0w6E0Vcy95qVRgbKgVJFcIC
eskgHaMOrDsa9195+SWZqKAUCuEZmtSx5tEeGUd/4f8TjIuat8NFq1Dqw9eWwyEv147cbB0Mk1p9
4NJhoYquYmwwPkaz4zg2abyWlQLnrW8qriSeq09U+FuQm5eyubQm/fXqjqvvMU8saWtzBZSnUZtg
uK4APLTVF4AtkZ2eC1ZQFcpK8hF0Y9XCiKUGuWa6bDOD285J7q5pKMVDMEu/LEpFTGYHpGp18NzA
ATwfnNZJ1vpJkFt3JrMOh4A86FcO+pFHGvT0d3iR55P7b6/fWfoaEJ6EaQRkmYCeCSpE2K5QR1LO
nRjofOwIjbgy5g30FHjQuQzdSc+cAsPleX9Jnkz7tTP1L0kTqew5uHbMUD4prmXTGRb49O9+NWws
n9V4SzX1MrJjD+WyW4EMzt52GlvSY5gc4+18SfqaFGFNfqnzQS5DeMODWQDGwEU4OT4gERrTpKSa
YV6mFI+ywHaqz292guMVlRTFMKd3Is/cTwNDudIKWMmoxKgDzMbhZkwS4sl13tDHtsqLVbrOmwq8
Bm9HovSssQMYHaSASY1iFtCew38gNfIKIa2VyjgeM3p01NdvE0vV0/g6uUQdsTNKKdn+JIJujuKt
/DgIJjxqPg2cKjVmVi+eKzKmbGl/IMiTR8NUxubJ1x6PFFb5VYxzStfaP6JVb7iv7cwcktSLTLAh
lOyCrcgjxAGZTW3zgrSTMlLm4WVJQi+rOWQD9zkK/1m7k9stOnpZTU6WZJXpe6NzY9AOBpAfIlTu
UPt5d1GGNTxC3yIOZuTU3QlYOdUUlXj2Ne0loPCb/C7IwnURqMdVoLL4tM5WIuBZSuaLn2OdVbCV
R0wb9BTg5Duo08tGD0Ehi0B/VTN2s1nXvX3dy17+o1F/ErDE/1ojZz3x91ZHt53RLyVpSrfffN71
TrL2uL1GAfklYsqq8DRW540FhtLR5DwgvyEF8eMM94hmbZKaNABWe8fRTsEyHj1BV+XAdGOws3ZY
rMOZxBcQTxDzE+qoaHgrVqiQ6uHXklAZNLtV3H/+bhrO7Y1Ucti1ehITR+AJtB65xncMOQ4sMl2F
0X+nbK2b3USt2rmfT2TY9Bymk+E7omJRKoOMbjPVNZRse8Z599xckKHzTzF96/BKiRMrVm0n4Sg2
vcc/fE54ZJYPdRJ3US4xkggdcuxQtVvcYI7+FnfUUx+XASG1TMliMcZeqLIxIDHkkYODt3YHK2aq
QSfRnTARac5WO22AA2wt4P1mRCa0EKfgfyrNFDB9eZ2jFgdAoEYzAguotCOzSoaXXDBcQJP6ZT+g
MkTgBQyg9D3qfrzDpjj0v3Oob8ePe8ppW+MUIAolbVL6Bu866CLqRDDVEXvSS6MIoVlZUoEMiPLF
ah5A2BFmsU4pqimlCpunAjQC9ceycl/Tt6zAaz8LIVuMmsg5tPAYgnSjAPeSDLWKVAOCG7t0BwEP
5yz9DUsT4SpoJ5UoyTDlyrCgEa2VAXFJ+TNMByONGppE90cs90K/HPON0+NG/sdQdmB5WVZeb7CP
iW9Lo5vVzIxv5Xwqvwylfec7rtc46VapmeBYIUNODXAJ0APVVbn+Y4zR9zCwPdiHnoOWBW+MRaMx
HZUfkKiWk+BNIOx4LovzEnlNrpEXYkN6ORJH0IVlHHSbUGOjVg+KVW8qJ/4raRXtodkea7dqxAS4
2AERIKQPto8w0Mg+CTV5suc8r8MeuOwcsmmAoJvJKTgwgYitF9Vr/UpIeCGydwqzI62V0O9E8b6c
F1AYu2uX7qhIpkWGMZR9QDfvq5dFDwHSfO7XhsVC0TIC3v44FsSOdgYa5/ZEuiCjc3NHI6t7skne
cpNCjm1PIgsCw24rnmx78XdMN8mZAwpIYhVFA55Od1d2VRKIw3ybeghkzsf+an1ZU/+mdxW7H/jQ
pYAYojvN3P6Oo3vFNvFFeLJ2XYCUMlAVwQr5CMGukQ+gkB99BotzT9kfXeuPTsLXKBBglnqmRAuN
Ldg8bFAZUMsBkFdnuA3YSHNMPE7MwtIng69bOszgRLiuRj0mRuSk0MneS3Tga8q05HH4CtU+8rU5
BVQjPQUb3H19R3pLQpZ66m5n+XIx43KwARoqlONcYRVzOzxdsuyT7f0+NLsiOsqT7GpzgltoEP+u
lNglSxqpuNfDdToWj/J8LZTrhGMC7ok002w8Xo1sPA/HfZYm3vG/ElKm5VrOYkaUOFomzYtpHY1C
CAnrnaAPXoeBju8jrO7SqrgAzR05pD11fR/M9aWx35E7Rr9kLR4egodFdJIrJUx+rLAdYDDBAFr9
zwn6yvxSljuPj6NRRNONrApJFXM1ffS9so7kjeNzSc42gnNsi012mZqhHv4KIqGcE1zMOtkNZ4Ss
v68KXdJyQUme2zA6ijLbHjH2Hc0/vAPkm3P+O0aSijNEYCXdT3b8krra9u1y/a1fErIQV4AE29WG
12gO8EAI2CzDhFMRVCM4QnmKVsNQds4Ha/dCSCWuuKPIqz/58xIl49aqssuyuvnmwxyO7AFnvq+9
rV5U3IZt94TLcVBTAitwpVlCYYhds8XEqeyVnwe81I39hNxQgzviSxi4LytIojKfrEmV0CZrg+oN
LpZUECuu6HX2aGZmJwuPxNq6jlgjOny4cmy4XdzF4JS8oKxUzOVEr3CmDOhyGtHcLD8BqEpia8yk
d596xOaSQDqbztMlHmP95GPExcbNFy82n1NQVdmUpKU8iyirY3GHiL3mtvhWfxNzkB2OHHZWy048
mUCR7TeRGtmG0lQD3xeH+h4TfbIQKP3kF1brHgqtpWGbVnaK9waX2gWJ+iOGwPHIlTlGaAgrZzA6
MZiUKHU22vRYHHWO8XPHFrTgYne3NMDJi2Lzrvi6Pnp3xEnunfo4OlV5MgSmEi8jhERaioU7CnZg
wq7njh3FDA/LoAXVCfTzFTyVP6eTNgGtWmynKaDYE08T4cWLy8MbrQJBadc6PhYsskBu5OSWqTAe
8SfFMwSrRVaFE+T3Kcq6/HwZkQz74GbCx6XfM2FjSivaekfbSo61xWG0VoNoWhmIYoaBJOzw40h/
EG0Bcm8XOXa6YvZ0TrhnrVP0e4prVARYDmUIADvXnPrTLA+/H8ul2oUbiw6TiJzKXFl1Zsgp9z0v
r5l6Au/n+e1KLcRR1o5/wdPbSTphB8K4JZFRE6iSjRAt5CUdauhkgCMg8KVFsOzU9YeGb4Kr9vSY
DSKWUVAYkIAbCUJGJwWtMU1fZgs+cTseKNUCMAbDOKli5bi9dukozY1iYAh7mNbs9OzIcMuaj2RZ
0AO5XYXe2cijBN1aEHin1YBMFoYgCTdoUm2dCYAAUx6+rIN97v5VBnYIAQiDuUdU7G1pNlGsAk3g
sKOTwbHVSlBn5EuewbATjJAns6xJQyRyas7yRxqe+Y4uWzW7bQK4WS+cDHdRaZ0EXUBRNs5lYXZZ
LAwKxqT8sHKS7I1nAQI/LuMdA5/U6H4LDpq18oKAxFByBfGtXBsUKJoh35J3FXMkGzcMCXFJMkE/
GFjqc175Xp0R8YFGgtI4HB4kNsK9RpaLwCEdskI3wo1xBNoXrOz5Euxl4HkERdpsXFWdZk9/6wuY
WCt7O3B0cqQio4TKBrIlHeozvBNQNVUljCB1d/uTWaCupIfLhwUkgE7BbeJw1SWunTFygFGHnrjB
VtdAsXxOnPov5bvIyehFhEgocfzRHchOkvziZCj3Q9c68sZUXcImaslQlNzxF/Z2yjMRFNyFCqCf
gcj/l8EKLu3tQHv/sEN4H9ofgivUfW8rk+iNgegUHBozgal2F7thAajG48xUm3iOYweli1xqEONt
GyTm4H5CULNJXl4ExtWmbP/SzQNQGVaYghuGYnMZgwvsnVtSmJBLZp3vqS7tbgUfxCKhnZO2OQlx
vMItZ3Mi0WSo3q0gqbgemxLSA9lgES7rMX5oUdJ94KAbQzspz4cU+rOcPz/Ssp5ljhoMD9CjWkw+
qhHRUHdXxgsXzRYd2obqddjcVip8iJBvSzkiI7VN8DY02nf98S1kylBYoadx0XGjV+Wxn/709CJ3
hoIfdpl7PKwrxvhjwmgMC+GmuMz60yo+TKF+HL6EXH0eHLz+hUt8elyKiyU+Oah5HrgMGoMlISim
PyP3oMhbkOKMcnWtHQVKqgjdXSvEevLIvDqto1CFE3Qtm5k6pn/E3QrP/cUl3LPFTU6P0JCsnXYX
r+l+fscftIuTO+3tUjvqkN8Vdz80zdczWypKhv9/gk3AzSDP23nh13A9S5nC7/5l4SDMletsAYSi
Q+4QXPqDHDH60Ipe0zIKSXyhueV/fkOGB37Ik1HmYyxu2GZNJb73RidIkiedGwbsiG346JK8wBVJ
Ozfpz/U6RipsW3Srk9jU2gQSHNyBYe/DfjN+pXl+aINRzF0zFCXNq+/ro9RX4kB60hcLiB2mDWU2
WDgpYxuxnd9qiRKxZYd+kezqCmPIY+/DkQMQXOMi2zJLIkpEulNAhXkio0WWasjNl9MISjh3AG6g
LmO8r6dINJdUnxzd+jugy4FT2MsLEOKNL+FAOFSuBoRPF9N41AWObCH46BPyUmXY1DCkzdSk+/84
avPFMhVJ8U0c1PR7ofUZq9wsf2PNRXYscqPtmtuFn25AmH9M2j+AzdyP/tSyGnmVC8YV2DNQ2OjW
6NilREXYt/C4InRyP6piRYhXtQdAzBQ6VVskKV/rbXaZLWkxvLCQi4EYxFwvTZWdH3xGejtZWBOm
Z2YQ91ZnlDnpUfdisFaFqJF2Lz2l17s2Gyqh8gYtBVKZXTyso7uekaks/uty8UiWXdETcxNGDie7
Uxd9FHk4kxviXHWxsekmp03SKVz4UJ8TqdnhWfXCZCHpKLAdRGNEmdurOF+umFIb17xZQGM/gdiZ
L0Y9qiMUcJaYNoFCsaBNBo/2tESzuHJhBsb6S/BnRRYdrv660F3gkEw4dE9wuUKFKe2XPC4Eg1oa
f2QaC7swL627VxpIt3oQLhxRLhvPgzhARJB+gbyfel2GNYHBub546i7lX5Yxm4O2SWr2QyLIN+Uj
V4b8BKHOL0h5DxCNKmWD7Abt7taD76farTpjEUUh9nghhMogkgbB3cJwtE2atY8B5f7FmAWrbdhF
UDDyh/LrAcY3Og5bCSAdDJLIoiHYBH01CzYXdzcmIHkqP2v8+8wJ5fuzt+Rq/pExxD+8GP2TTVTI
F/045YOx+Z9HhyN3zmWKn6xRIwR9+UKxdDMWf3hdKUZL4W9xYYSZ5jtXq3cHBug6OKahNeBxhUSy
CMJ1hzsGEIv1PM40/wfYIywLBQ3cSJ8T1D5XPp+uCtWSS2NxG4oMPGyPfWI4qz9ZaP9YkJufinsc
MhhclISX6f9XalyrujfgORvlspZ2QgebZId15EPFcaHvrQUtbb+ei7Az98qF7QHny/v0YM5Cybdj
7giMz6CDw/b58rvJJfy+YdezdfdVvw7dQnrlWQhTFjKc1kTNWuvX9O7I4fZGozOiiz65f56sRjZF
w/QTXJOHCM1AaEUHZ4l9N4T/cWH/guFQ6CERr8P/7ruIIbG/CXLNV3Jsei/aHFKKz1W04p300vfV
rJUbt7Qm8sqTfC75VebhnZmqGEVi4H7xqNtMZjkky01Oqyrmq6eEeB3GXZh9cguoLEI9vUoYS6T2
RzUWUdu4jV/KyMof4hFOLZ6gT0PGIq+0HvNJFNZGy8JG9vdkOKgb7Om+D230ya5RUSvbrgF9a+VC
ECatalLhbngGY1CtAH4N9ko89Y9majsZGsfUY9OXCOh9EEftWEJ3uSsOYdb+sneIO0h7lE799r5i
9Iri9u8gdjiW0n95w40nKCUIDBis/T2fdo5vFaGevFdGvZx0B7nWdh3gka6StVQ4C0cNuk8dH+j/
rsE2XzOWI9StXZPtVnCLE9LAIjcTWOG708Wlta5vd6J4PcdYq/HxKffAj/40p9TApUqTXcqnReZl
RqMkyFQhE2EBWVeo2AgATEOm8jbB5F3t5Bwfg/hWTiC+WOCPDb/WAbzMl3F6pQV8sXh04UdkxL3e
1VxoX+BUNEc5RWW3MET+hnC1l23JSqYoEN7AkTercCMJQdDOZ72VnKGXYJhF+aqGXTMlZPYs8YY6
axHrIrvxirnr8XTnvbvL+WPtCFEi31XZZcBUmMpxJMpEaleG0b7fwnTkUBXof3gN5ea4ElrmtzHS
LAZKGz/fW7BykctrJlSXLHN5kf7TCmcVjsS5xqQCKzQxvFRX0FrNO/PN5kBBSTa7e/cxjLvwqpEM
W6xZlp+6LckeGw23XxNh9SyCTv5xL39eEiTKRq0Zc3fPH6BdzCW7Cha0815QEc298bSYtkyAtqcM
cdP+kl/zQ88BtWnFXfZF54KrJroUlFCD8UAkQtwcbW4FaVaPmvgW3VYJmHA6vh5+vkzDJOpLjVa8
nHFdYgc2SPyEJ+NpyG8y7MzcXK8EoaEmMlRTM587F8xh8dY9AyCULdrPlYX3+qiufbuYdYttZjfi
0Qyk9oadS/FgZyk0GHVs/tABj7XIVoJN5rQ8BftPQmdgNCe6sC6QCXe5xCpyzVpJ/LOTbFzLvFsu
Oq7EnFziaaVJK21CyHRGrm234K6OHfnM+6TI1B0rEZGk2ugMpOE5UqkZaty3xGKZfWyV+A5Qb2nk
Zox8XTe3THIzrX0ZfWYTBGEPtlWFVJEQax8SmiENB+A2FEmY/NssMwCltJjk4FJSx674mtL/EXqO
mGCmZKnYGnJ6K83+luRZxJgskYZYPnx0NO2v91AEzQa2v8R/JjIhhgYLVP5TJtORbxQN7/D6uII8
Neu/EmCD7Mk1EUQcBNoXRrln+nHn4aQYs/CgOv1WSV0hvX5ycfuiquDWaW8XgjObaoxCoBAQpzk/
sYZjz6lnmkTf01bfZZs2p4pOZIrJEZjjHAD40Hpu8LCWAx3NIMjAepaLRfppEGHNPPIwKHM99KUe
PATSvEiooTZgcbHhR3SkwFIgPW5leOzugoSi7XY+8cTjg/ZGPLiDJSeZbHJTnC4fASO9xW7yH8ZP
61EBa4zCLfOLVP6ggjeGf0IcPjdiNSFA2om2RgWOIIzheLEWO64T6SSuo6+MMZeIJVKWI97vrvJe
ywE3S0/oprps5W4PZ60IDvXmikt8WgugVPeN/WdrLd8JRObw3U88BCaNMBpG8E+4aYxXlGiC+1c6
lEjO5/3TRBLwS/njNyyHJXge/eEfjskpwJxKDTZtIZKV9RFkrv+1/j5OC8F7WBJVsf1I2SbZiIXA
BiNDS4u84MLPwg/IMtlXG0WiO/GwkdgAln/x9YXuraxOt5CgKFLiVM6lZynyFNXah9Z7FnHCl5aR
K1dDBuZxgbaWbcLiWm/Zj6yfJ0mruk90FFY+KInHyEdm3ZOFdVBAWQD7lxKanqKeUy8HqwD41FbR
nrp0j+IFb7xx6ymceel4entoFYbd/zNDLqdyiTTn9SU9n3OJKVeao5d9Yio1YeStxJgbdT8G0h4F
ymyNzPkf0Mgy4jbj9oJgwuLLKHe9ywPoFlYTQUH6/I0yw/AsYslLnwON+5IsfjqRKldx3AHj+EzG
UWkAnQeqqXH3Z5QprT0N7ShaA/J0F5nphn9Y6Afz8sIfqChelHBEhGGXs/z5s8IBUKl4UUve9RrL
QiAzvxTvv+KkBnvjRlG30xc4iADO7taXrD/WQkj9ytfhx4lHALmKD/wWGQ+MjczF/ixgfCXhTjMv
Gcre4LlJa3V5iIA9Cb3AKgvAfoKx0hMpDL12l0z/ZVEVwPdEfSbgIpj1G2XQdnR1CrWyGE0KO7O1
kgPrXsMDu8lihlRE9bGbjuYi0ElmfOTl6UBWvi/g3McYI7hnO8jsM5ZqD2YuxhhPJqvEabHdDpvb
CPO6YWvLBXEC6cE97ZSKcyDwG8PsDPYo2zPi4sfOtT+3zX9rq/44iXZhlZn6bontsnl13DF9eXkL
jGSQlk7M82Dx7BKkHRfKE527pZdCpChDJWMapSJ6R5EM7G9NRSp7qTCHGmkvafREUQHhiTrYzlLD
uwAto1qndDe6FeMr+m78VWp6B/hr5DiSoJMrkTx4S38jQphCXWw+YWQAnoEOa4iGynqfoMIJR5jE
SxrhbYWo/k0ORDT0WrAdYeWlgHAaCI0BH/6WhDkNu91GvEDQ9HUTz5BJa42K303cFBAnnve3cocT
XyJLGSfRVwqgoHhDCdQoN7Er876OKuRU8LwcjkF0GGkunsYecUp7bTmLuKR1UwsIRHB6BBYA7/N7
xiY5MqvIYx9RtGiBIJ2TAkynriggE7Y37Oh/JofFWIcJHfpKssYt+s9fDCco/2bgU6I0RcgLul/g
1UZrVnfUyJfVNI+AJc+/tsS25OMnGVGM/hGZXm4TfU8BjL8sX2YMWeGoEwAWZU/2D67Y7oCXaMKd
qTZiwl3flXVVxtyctOFwVRLnfhyTXDomaecnWrWBSwLVHaaCx2H0J7lAnpl37hfmivptpmxzznU4
hAnpmmJy/VW8GyKjjPbifdJ/N+kTdp7fIbk9ThTw34+c69P7VG9lnR0rojUlXoqW8Evk7We6LDNt
1E0N2GTs+RI3Aw2NK2MPoYtWM4ShxotaJUONMm/WFuRvIqnRNhr9zed25HK0Ab+sMta5ynNa8Ptq
XIigA4sto00BNF4c55ThjC/ULresbp3ZxrAG2z+NEGxufNtitWypYTWbkP1oYdERuModtWxs3SJa
ahnrPUuJQxxwgQ5ABnqU25Yi59lQq/tDoagZvxsbSleUPqAXLKDkZdgj/Cx3qOMlCuG3gZrS1n4w
5dWDcb+U9Dqx3qRl+wh1rCaXMGIFKBS51SUgQrtrW2mX7jo8q1XfC2DL8Duu7x8bLTjzKIwZYbGc
KDvyMDwl892vL7ikm1B5ywUpPFJgr4Qei6Z2S7wtCs4sgJ3odEftRlidZDaxFmub4r9Ja974dz1w
dAh4NE4LRSHH2wK2aP9YKsGJj4yQ8Noim9cavSXrGIs2iGlityph0gxT+PliwsUdm/lno6gxinuH
ZAJzfwuS3Dzh+Hp0l0qBITGKVqNSJFfgLuCpaKGxJQoXgZcxVvDUbKZ+cR2d0yg4GxwD4KNMvjtI
tRCaE13WKVUnsf6QxxZoP/xG8ln+R1ayCoZ5jkR0SkErX14yqEvAcb8opMFKysYBvkcojfAkh6nF
xaXEMj/DLqud7dVwlmQ2tP5Rjdoc0TlaDRGOvmUfwyuIdkQM5BXEt8Ye9kgRan3z1SrGVoU0zCLq
AgfS00y2fl//MnqkeKXBHM4ucPDPw3Q741kOiWyhY2FkuIgWMoxMVgzRGAJjYoNEuTnllu/hAbKY
nZ7YPbOv83Dwj2htPeY0GWFrMJe/XlinJTZbF2ZMy/GvxfZ42zmzoYPjtg/cUK1i20DkL6SGWQYv
KTe5ioAdh06Euhawx9yt5RikCjbkZXhW9vKfxW7i/OVTYPWYIPytka0kU9e8T/7/CtrX2Vz7AdNZ
H30cxj3gF/ZVKgr51zFSYt50TPasfrTI2bO5FCZ2G8Wr5N75MkFIC6KRBmgd2Sj1ZvCuUy9CR/SV
64QbBHE5AIUGubd3nW0Pary8RCPlF86ujUiq3mk6pezv4E+DaOql9Y5EqXIWjD+z8uKoc6D4tmZX
oW4PgpQiRWMSOVMIfpBZHJGOSh/tM+Iwcc6M/o6UFtdpT8XVX84iXDYOi9V5jSe8pSsPSfUB+09v
yJ3qXsjrbrJZTl70mau15S+qm3IWHhwYLTGKJh2HDK6yQX1Y6d1k+8PcGbOCHTtEHvVxq5UzqkUJ
FIbf0leI2FogPYq5IsnfNiGwNkSE+BEpG9AUlG3ZKxM9cFXaSVvMp6d+cyTH9m+NrYtFzWMULPyu
dEJl7sYD7GGKTVIeJkLfrLPR4Bd7dDOrPEB0zt8IMgn4RSJRK5aTIQSVefJXvP1rxgUWbwxojRs3
EiROLMcPcFBPIO8LLcHbkJAbP5HUtOQg1foAyVF2byGsSCZG/STgRILIXPwbYItYjFLSyX/ePuRv
0+xfFSeVbNHIh6MHLSD2YY2xfPPaeNlquiC3nLPaBLDv8fIeSkYv04QnqTvT/OPdiPxuVLEY4kKq
RyQehbTyulDzg+jRF5mxXa8uwpMsDkqEQqb369o/Bambm4BrcX6j8X3kqJyNq0hGyn+8ozoFGY/K
KbWdpADIjEJlConSmZv78epKJ5feEpQTvVgweFjt3G0qdMrimy92Sv965Xi6TXVF3SmMNMoq8bb4
08ZQ85r95qmKbQJzYVwZmJB2lj8YvHo2py75N0Wy4eJUv5CDvi9eV7KbAJEDUreS2VLrVUHVLBd4
hEjQz9qzhqjQkyes8643krlvKBtQgWvZ1QnPLwNeYCkLk6A/QQNVLMxDo1zEBZgWK4KObkY9YZoT
/bhDOsQrVHjenES5sLE9H8X/DHy5t6ygsav8ixVyeAJ0Osd+MGHebHRLVJheHusUnhePIZfD8Oyd
72JrkN2YPvLWo8SSJnkUESVHWTCXLNQJcS/tGIGK/1iWl+8sD9icnlRAt+m98qs8VOwK+S6Ixjdn
VhS5tihJEBRZJf2tXFznN7ghgxu6r3uvdJTzMYvd4IALTF9jzjmiZ/VSd5qf/g7F+4KcUGi/Rqaq
hI9O5XT3MSRBsxkPJBSSp2tHaG7XjWtZ5/+Uc+AqKO9su3dqlkbVGlv2Sj0JbYk3nTPkL1DtULMr
ZyPtjC3n45UYdxGnseMuJTo3qtaglTWh5MMBXb+wB1UM2bDeXO9I645PU6ofKv7EmB3sTzlAu509
Ljv5nlyiSbeOYKnRxXCWQuH9RrWP+hPNaXUxi41rzlmRoOWtCfPw5zPdaBuHjStRFwcNxX9CyC3Y
g0KjGvDMebhpm5QTqe/UMAvXPNWf8pZIthtAnfAHQ9BiWF8QGNVxM9XqmI66PIpMB1MpzdoLw/wx
qzOCjJLqniRXP8isMHdbwHXkjDdCMmvQRTdKml2RGLBv/UIT+JNjSZ9KQCRs8/fYlCBsnN8ZcTbT
Shte7W7Occ0ECeLdoKT0KCz7yozxQVu/M9g+SwkO/q2cUy7rwURMZiiPZW4bXPyXCHGpZxRIGA9U
gXm/3pKuwK/MMZlMomhc6qqFzBGdSoNq63dWGyeCBjxNk2/tGH5LcxhIWsBvShdAJExkMpgxX6l8
cHbJiwdRBtRxSeZAzvuppsOsSPsIgMKGOmyAXOuJVKUdGTxHpfRdQXLoNLSwZIzpvpDjy0YIvm8K
Hs4vJHrrOdwI7DeueZqhGJSKT45mWxm8eJdW/GWsJgVaol7u5DXNFUF3XG95wXnfzvp3n2AZ3vim
KsD86+2MOq041XgzDeTw3Y8K7JKD5zEAYsNC2QoRTglrnjk8qtD+MoPoazsLey2jfYefTCN6lR3c
pFelS9rV3tTXWRU6S0DJBqLh19KJhJbSpIIFc+1z4cpHiM/fIlqSRGgKCg71ks4b51JWuSJZ6z8H
YHc454JUCQccbCv8pcdDKGBw2fjOd5hD18wW37L7QBDQ2T1TLYdpmNrpK2Kw9/03KcA6bBgLNhFo
KXoY1Oh9L9Ndx8eWx0w6NtKkG46WKAHL7ITCuTxuEPKJteYBlYvyy8N+WsLjGDDDfSufjcePd7y1
1fqe+dQn+tNeQdozHHUQG1aGs76VAV3alEoPFfszCzh+9WhILaWuzjm5zmhGcepan8iytjiAJ/Xs
m8E3dP1M8UjWSwJWHWIXzRPohMLnQDVU0zh5XXMd9TXy3PCVKeHXpix99KEk3gFVxol5emPZP7se
HJE7lLv5hpM21ZqpDoouyuyaRruHBQzLrJ9TOMdq4FajDnNDLRTfAecMaMxnXlqqBNMSV6XaVE+l
1Zm1RLrSJna76XsyQLtjcppzndYvWJBgHskj0apZ2NZhcNwboyQ3PYs34Vs/1O8NW/jOQg1lDLLL
Bt+HA5hbF3hXDHhUz81ev/fMoZ/G06bn/AnCwfi7QqqSJVr8sGIqXpt3JLiCeRO7Cqws+NjkiJBD
ox8s9CBwaQ2OIwUa6Vt9TnzkKx+8HuPm/r1VgvxgMvj+FP0M1b3RwQtnPOLAFzmxYMWPFbwqAu99
FBQi2dLVg6Zgtt1VMnI2F9djZbEofig0kK1sImwxR7UccoWZV2Yq199X5pNCI/kYcl8JCLE1Ybnd
rrCpSue+TYO5A61O3uQvuFXKkHMMAkHr/iiXy25lI4ZxoFBDnSLYSnQ4igfz9UBq4qS47pDmhb4w
Y46Rp+IAPG8F1Bnb626RJbRwtMfy5WMHZ/AcB8I5Cr8EJS3leXTsbOdBRy2u73G929JqcWcG2k2F
kVtCTXJHoX4hFstE1cVJwBEV770/aIRUdfQqZAdoV4SgHLKrdW3ZKTc8hmH7ARH6f36pR5nJBN6b
9G55EeSFwlOUm6GvthWRgDwZ7bCeb/1obM7/RRUsLfLB38dT7A2iFD2PlIik5auYNFYsQHICe42F
D/YSACoVLonTWk4AE7uQ081wwpchYX1rL6kV1KnTchSGx19SMhkuIHi69FLaOBrYq686PiiF0vDn
mhLw/L4ITbhUDjHIlmpI09e7YsDhx15Ec01tnb/TxawxleebZs+UAHHMqDjz0JtI+lAvicOz4u+z
5SQjwuwJ576Q49XfbzZX+Dc+OW5MhkV0YZvQhzcj2FOuWvnIClStp66QqsGI284sXvssMgBCt+zF
GO6ssuwmNQf1wL7PKvzfVHdW0AcZ+GN3Mx99y3HXQ5dVoiyyin1yr8E/WPBKC3RlEmMB26vt0Tvl
//aoVnZ4+2JgrfmJRZ0t8R4Ym12mgPqYeznnbGrUaMwzYpsnmz+60MOiEjkI2YOqNtiS6cl+XEVN
L+mUMp+hIpQQsGH/IE/AAinNOU5ESerLQ/PIJo6dZ8WepkZE6/vpiP6jaJjkXvfN8w/y3cIdAdoO
GaesggeyLHP6CrgW6SY+eC5JmXaGI3ky5ladQA9Wb/eV45/aiJ1uA+TIbgQZVty4oSFiAJQdHd3S
5wvDEnt3cezblOcHK1JZeXHtPlobHffEMPd8fbTIncbXC9hxzsAp3mPSl7ygtg7Wk1PEIlMJfupl
tpz1hP9iuYli68x+eM/hMsR4dAP1G9UEPQw/WjP4hLD62mgVC3ZbEAhtFL+s3j8cWu3DjOOlHjdw
vXO6rcR/+TyDQH1V2lGptAngWKhIA/QrbdZd9czLW67JfbwxN0IILTHUzGa9avepm8FWzCz4Ii3h
QHPpNFVjlVaRmYRfB7ZG0deBOmhtDtglnEVO40o9n57MkHPcrT9qYGj5kTf3ex0LP9IDZ8jk61D9
lns7uJriwxQl6ojy749uu1fwoY+ag5aseFk56Hd5qDKi8RFPd5+K5OaHmuioLixzr0B2PEn509UT
+MrFZiuZKjlTkMcxwa2VRc4ItHh8cUKskXR5PDC3W8Zje3Ii3T9K7A6/VGeRCoa6K/Mf5RImPdL0
aLHVD+196rqgwoeSMIxIi3pohm2BzUpHwfg1wamt6UN1/+b01RPwuYYFXPLPp7c/Hz7GAQia/hp+
EEMEJBWamecKyIepcXvRo0naFGFHLQs8FPho5eDZKdhFY+KmiM9UhqHkZfzHCLzylldR5rpSajGg
8352AmGxNDBz/U9ahb2L1TlsseCTclvOEBhN5sNkJJ68kUmHdchQUCNj+5ZaVZKpIPPKWKYxNUWB
q71jlPN3Ibc/p//xxlF1STWS3LUiwTZmIqqSVJQRjeTYH9Nfq1caqypABVwHPhQPJsnSiHBRX3HN
Zli4NF2CJnSzjYn5afhl1CnLpdQ6AWn6LX65EKCCtjLwzybw0bcVpfGXaFlpfsW1Z73JQa5NO9Wk
hcnuz+dd7N6f9QOEmVSB2WBzrgHX8WAf0sbE/Q98gWZVc6mpSi0KseoffGMvh/Fj988tXA6aYtX9
rCCoGxJh8FC10Xs9K7rEKCTCPrriZX3d2t1OAhtsxfkvjfayVG/PdLADymu3PmSNDsnzCS/oWWfm
eidAITCbPSyB7ZX7Ae76eXr82SSxo/GCsNJ54Za6XxNpijWFDAFIxohPBSkLGY5dHZeYTj0po7b4
FlJO2Zx5mOgi/F0dxpjioNa5vfKddb4iJ+XdIa6mi+jxKSdG8u6bMac6wq3DtnOLRRF99rZu+Szm
0D4VxJ+7uCjg71JlyleZVMNNB+35YmbURLLjVCjchrVFwaZXzuxXhoINCEBlE1nuTCOfcOlmdUuf
ZdRieDDgD90snO74rRy3QI9mIf6T859JJpr79btsWSC8vq09/iiXFLZjTXymiGrCMZMVchi4CxLj
pl+i7BZt8HccE3sNU4ZASSwvjc7SiABVd8iRloRTaXh6Nilnhx/FelM8FZV/Uz7bTjPnipDlw8wB
oqpvH1DT/xXLblRxAxkSoD8u88S0Vjbp6ZMRwIwYZFJOoAPStBw3JUq4L0esNJiPi1160pS6ZT2s
AG2iUdcKKtq+PY5sHoeyecNODtvH6xjrOyX2Fn0K9+vYBRYLS2g+73NmPXmmUxPWRflDcFMJWQG5
+QV8wjqEngjT2emJSZ+EmU/IRmvZZamJePWEevg3a8COPb9nb1lxrfv3LA2mTsDdlKX6S14mQ614
hkWWue1tbK3TdBpknIDcn45G3k+JjcY5pJSqX5YGPeWo3Ni25LWcLaK3oFOZaAT9p7isRr1cSADA
9irJU3SfSOgiWyX9ZJ3wCWtvqXVM3HRuLMklmet3EKcIvovD4RKXKSGRo8LUoefRe3vhA3w/nYdR
/0XzRYNnWhdDTfFGGQ6Q4uBfuso2OKK+uZXrLtL2ccL3mDOI/qNT4+26Z9mNxp42WKrrEyLkS+FQ
AxCIS6UU0NLePHD3vsXhFlB4wf6IzscupRaxai5pZUkny0Sv95XbBE6MO6pYCQx4orGjTtszfuUT
W4SChak83il0MfjrlD7s+vwfsgITRR/tCTKj5Qt4euk2L0sH7rWWRukbKJUex/riKWB2S5o5562C
O5q7BZSB45/oouscSFJcCn3jpzMAAaKU4J1rL3hhePtybe6mLNOlDnvxvLhS5JyIj/+y8qWm8i2h
dgwCwVPT1sOxx1rghxF6Atwurb1q0+Z+M19JYvW7p8C7gWo7H7E0kgxD4ZQEbLzm9MoGUkL4HgPk
vTszjAhIfjv/1MTgAMvsm8l1h8Sr3c0hpwGnFw8vge4vWVjgLMwjq9yQlz5H824Bn301WadPCxBA
CQebU5GZNygSDsX32mZ2l3JNUYzrFPe9BWbqET3Bh4zdtLcTTxSufu7vGZHiSh6IuhVvDyJAu/zS
aY1I/Eq7pwryK5piFuZRYIyUwH5qgOKn0WcJ9Elmu8v+tVIAc1tndOPK3v15l+T2UCNMN4bVnoxc
QT4ShYWNBK+gEEXdqLjrU6JxXRecakCxdKMDSO1kVoG4ojFhocHX2+s/Ut4RUBA9Mz1+dqYeezkX
oBNDphohMW6dudvN2fqxm7c+FWeXcTDxI5yz3s14zrfBaVyRJIdFMXSg3GXBk8cccE/i6a9aB7UA
5XViLRFKcxRn+LU8XZFihxa8XptsnOQPflRYmd08BCtkxC+JTbq8pszQtH+kD8TnUh2NfeyYKPei
cXeaoj9aELAGsAv/IZ2Jv4p4Rszrg1dXtgtnvuCe9t1O/B/EeDR7peBEK+Yn9CbSH2iOMPj0xQ6M
S6vRs4J4qUT2+rX0MYFSg5EByplD31TS6muldcONajz2e3TbLnSw0WCxhLLzwuVuql1dDiahmmsS
rRzZziAH/+vtNJUW8+4hh/KGCMzNZR4QRNtrUqkkfYx7PM1q0cO0xaNXq8b0lqer4Fplt+zG/o3Z
Y0MVin5E0vMw+yJ9hHWuwxPwhdIR2h7fSfVfQcgCZRXi6M9cnHBhVHo1TIQcUun0y3s/k8NbyMY9
JplOqoMUWJJd7OadkhzhgEXVK5nu/bm4SHkEToaEpftiCtBowoaShT6Ffj2Gk06iPO2bz0wsvEva
4Ezi+iWocxHjSxG7iuh5+I9gk0fzweapMfaAWGi4/TQf9VFM/dhBqNI3GZyqljvT2a7Ouig4CKVW
Yvt0kRFf3ifnE4cIl3MNf29Ab90+HNJk4Au1tdwbhFyQcHGb6d79F5MWBRDh+I72feL0DTvIvZHz
F5nh9qismJ06OTgF3si64d7k0R6L1gsRH6QSm7LdLO8Tpig7BoHn6aq5Eh1runZg+vCykklaEbL3
BTsQ3gxMNUHNnnrurY+RGEaKtPwqEtyFheg8efKVEfgjVSVd3/flFbeq6ZVt20x7Z64PGFZDQKO9
BhKRfApzAgilTvlZSSXPZIxjCHFm9OxdFZY5Ie+nUNl419rMZv1Ydqr2PkyjgwU8FB29eRvUsGVE
do5YGCTR+2wzOKpqnEF9VQaheqSNWMxxjgVr8jj83PnfBaginrRyzYZ7pJtl/Lr+P410WC/xolqh
i4Nj9Go8p+Hak4pxTf4hG9R0LpfnYARHlYy42IQVk9LpZUt4a0Iv684oU4UsDzWD0dAwWZpYsTyl
6nPGCg2rl0uv9K+4Agr0n/EmUm6fzQSNd7awzcdpFz/Nsfn1R7KR9Zc3B5YjZud6OUOcXthABOQj
pykcf57nmld7fqvEplsuOO1EDp5YNnUx/pBtfv3vZv1D1jJ5fkdKcXM7Lv9Jq4ilZdkJoH4xCuu+
A5wNDd1A4KQQDDZNPFpXL0ia6p71bPwy+Et/QbOQHndaBRrTi5krroPPgF9FuxHYEz57ypyMxpBn
QsQn7s2Ne5zTZh2ymCarhL4DFt+6CHJsE+75DEMwrvDX1X7372KWzle+B7DnYonlWMgutyJ5F5DW
kJAR5HX+lNC4IKWYZb9J+MsCN7xM5AzKV8pYNPAuvx5kyqlzf7g9aDeFkOV4F8EUbUjofhjlwv1i
ZffE9NlTYiavx1jO3ljr+h80S+CVnoKoMUPp5Yj9Ry+VG1hXDEHkmk1nNdNxqSubV/oUOl+2hUEd
mvqvWb5Vc0MneM1h9DTL5lUhdQv6qEedjs1jOU6iUboWt/2VNCVX33qSvRJuxlgOJOuvugB1jj+4
dsKsGf8RlzNjbyuFZP83mcO/7piz9dFr+mRhxGicHkRjxcR0QHM8Is2Ys6uNgUL07f6X1F7w4axt
0lwGu25rNe9SfW8zp2Raju9bPtkwtyfrAEmG6Kk5z2X/L58lr0yTj0z9Ki8usXgNxvj/D4NZOS+R
iU6HIaXpenY5kEvr4fjtsOhJqziSYgl2U4D+jPVIBOZ2gCuCBaoqT6mBQSVbS0OV90BMab296ugc
CE6kk+QqjTa61sPcgiaSMj79YScr8iY4UlXcROVQcDv27cnicu4xGGHQlOrycPX4CgXEWBCBvK7d
paCYSDuookI7v3D7TeSp8XYt84WSHN7dobrwdeByq4pkb5gYXfVaq6KMz+QUX6dxOPbk1qnvSMAj
Mfw9HAYrzTFBdBUzaM/nBBXNA45hkiXiTjYNI7Dr4Q3cOz34jXuztDGaVP6SDjVmStSLUN2RMD1Q
MTjwEtTb4xgjkL4YU48ArJ/Y2GtIFyGbktNsvJ3GQsdxsmPkWJs94jpwLLyl1+7poXUMI7tBIJQ7
9t6z5qFwHQvm17XgSTdNrvLa5EkbOtY4SOaO2ZlkaDx4E7RYkd4/oTg4pL8fwKmG4KF/DP35pkpX
VMHWw+OmiiRsdnnyPK1Jtx2v5sxR/pQYxzOuk5R76xnHRxhJQcEeeWtFqhpqNhoh/9tiw6vz2vH1
4BfACpXGvQjk0Bp/kewPW8d5Wu7Sj/RcQEcRS88HpSXg7LfgaJnPP94ItLz/z/yT1SOtulg+DRkB
whtdcooeoTkUXX0i5nBSw/1z/JLf+HvF7xhkDJE9P9cIcS67CbqJ1sYo9t6YxThVeKginMK5xpbG
/TxvsIuDOQWEoMa/v2xFKy9aah4sYOj8ZVSRis3s28rX0cEAxGyKTc1Ta38rGnA/HuyfK91W56L/
m6wEcbxd5Iepnw9nXaADqLXUAHZLkVX7p7CfO5uTXifZtfzNSKvTGUbDIRPsUdvG1rmMVCsb1Kqm
fEx1Ltg+wfrp+LO91DXL/Nl9Qm6+8yVBAfOP+ZqwtrIej+DL4t2NaLATRtlPrBFmAMGdodvKtJFO
VN9kQuXNTrQZHhVl1RiGBcEbazandKUCg85yx5B2Ih5jSGGJfSRaZ+YCjDwIpu/kvLxCPjr9kfsh
a7tr1k/5/uRJX/y49RzK9Dx5ANfFm1yvo0G/DpqRnRRpeJgHGxkHEcV7NUkzVcdm0C294orqis9j
9PyEdhUSGmqEdkY/ZWtjDsr1FQrm35gocWrhjpZeRnXvlbq5Y1aY6Rcbcb3GRi5irlC451w/9mQD
6Z+nqbC4wrlbZV2lMTIqKlqSdrl1EkQ5FzNxfUERIRQu6V8Etd4VRSwibpMz/aHgU6kBqmU9iTFP
vYmi+gTwipbpGXAbfmmw64nhxh0L0Zi9VLi7olV9Lbi31YwDDIWT7GExjLctKgSlPYFGfdyZbGdU
+iBuIJHatpvquPcWcjIxm1umocHYdsRFMNUedUdZMoxKgOHLYMychSX4l/iiFGrXGeC6tWtRwo/I
PtF9aX8Wt9B5h+cuC7musjm2HuY74FCm04wQpKLPK2zwpfWGUiqgTFjIITQW4YGcs3NOfCdpI8ck
Od01T4tQ8GMXx9CHE13mE9OORFhQtjbP6/64W5w2AhPvUXl6JljE9bnT7PaAReGftVjwyB8vcxk6
aAJPttEUtG5bTiJmOSZ+yRQeTZFXGSYNgIGUPOERILyFC6LPY7Fj/t/QzBece1XR1xGhXDQtuXcO
suCEuSrU6VC57Gg6/Wvpc4ZkFAJtsc7uqK7o2Atcejfra7mZhgfVc9xTMQJA96mh0U3gvzEWBlvN
PEwGErA4Dnld1xBs8Wk+ePzxhlDBCbqZOeJXlrj5xI70V/uukUqBDauZFj4O3bQRpufoZhNO4SSI
SH1drydjjPmDL3eRPfpxETJs4AOL5UD1M8fITNCLKp79B25FMli/0rOpUwfnTOEMsbOPr00ANulO
EXmShDY+kxSAAng8/tBM3CleQ2K0biT5EIkQPDyRm5Lj2VBp8vf7rbXbDzt/cJuFtnELe27GcJ96
NWsVGBWbl5PmPdGw4zaR6ewKpGXThOC+UaKy9oV3uGf5sgeBqAmUhTDt3Zap9sFs7JGYEVY13kzE
ERy4mqKNkVMNbdqI6LphGVC1YqOz4hz1QRP2RVYzDQIot2t8pnOnGwhGe5d7TzyQySMLyryqN1EB
lApFSD7u5Gv0W/w4IuSENiTkMMTO4iKuBFg/eu2fnQpNYSc3UygTltOSyWKvwz0BWdgzhem0Y13T
3kO3R2CrArpdASjaS/NaoxdEv85qGvmIq1iV9DMWo1onkXS7b39FpnGNyTfJQci8GXIspiK6cQ2z
hAthqZ6qKPJ45K+470Jw/Kqvio5ZeuYCjnF15JwTBz4zeWPEp8qLrNG03EQTGWXPv59pTOkOzG1S
Pmj5pb+ry3S+SRYN7jVH36sb8MTn/Pyqag5dK+heisTW9Mt2Fu0fh3bUs3h7JbNCMO17Iu2ppz0G
0gvIP0H9NMD/WZiGZY3IMfjMiCyo4WSCJVTaiInE3JX8tng2R7BEO5/7ZmihmULblM2MQG6wUrim
p3R1TaWRQM+Yb5U/9oqLAnwSal3RnAntw3pKJvWK7CuNlgJ3XwzwZYDyQpsrX+3FovyAWWuf93P2
k/N81XQjJZ4Tbx3WfdPGk5yyk2Yyjwr33J1BtuVfnIFjbiahY+HwfQJAR44ohMZfXqkTCb+SDqhI
C9Z52CjXePSdw+ieyr0rGOsIHEwGZ4IrGnCHF+sk+JkDCwhwJ5XyxAcixBBjSbJGgPPF/W2eoAFr
57Awruq3XC3QRxFVJMC8oANW5Iy6SWFHb3A1TLaYCxI5a0XnPSptWIJMaYMm1HlJcxh+GocxZmgj
2vo34xxEiC1NEGPi8Mk7Azd1r/JoYY5MaiaED1v82VIg5/L1eqmKvQa15rhGCFpD0VVcN2H2rBah
4gJLL84+IR3cHkAr1RwOkf+fiaTEYGBGu9RR4QW3BGd/kb0hi2dvW4u3ek1FVeqLqED5BW1Bxh8p
vKlruH8iXld6zKXZiPf/BjyfYTARDNOZQm5fa60p/BWTcP24yRIAoIECDUKcXmlnHKmd/6vh4TuJ
T/QiGDvLMOkcKMYqgxkJsWqHHAzQOGeIZbozaZPlPUw99Fx9nfZYfnPviB+uXAPhbO+dNqxO/kz2
1r+H3b5WF751rH4Xmq1rT9d9jtR++qTP4mSxPsAatg7JSmiT+NRlB/bOLHuXcAllnGe+GeNYhkPH
mvYMICPl1ACOMcQpUCOMcnjYvnCpeAYvKQeJpTwFXzfLftfRmylLU1BbDAC2kWlCTqvr0uu9c0lB
XRUf7ll8eOnWiwuRUfzscaqLVRe0Vpm6L1noYk+l50a1H7SITydgQrlJu6SUO1vYv9DPFZIwQiHE
h2z7rv68Wqmn6DioPERHUcIdcOaLohikhw336UyzkF1UdedL4W2Khuh34231LVmWYbjtTnMKk8zt
Q7lUFpVPkrmILMwFNVxh3xtZIpwPlEaB+CpbScD3kKjpU0Sy+GNcETaEGbmf5Pkgkzpya1p5Ib8n
NR5Muc0M+e8dHjztj6mU+a54tI40myX00VEwMRvnSC51jg4HEALK68DYPyi80M7vt6qajdSNRtO1
07QMls262CQ5SCITzbcekWExMsra3VGzLJgXf+U6T7t9aL4dTfJMk5LjtBkAElsBs8Lq31ltppDJ
gq4AqxHZmLxqxsXJYjrSaxCwPSmVqTmOQ+KGYb8R/zBwWReiz84Os+QJwx3wqnuztFHToHVFDP++
I4dBKNCpFt1HzKtH++sKc06OLNYEBCZJq+F76lFUqEWkkZefemvh2Y6O8fxywIxIO6qeP1NkhGGg
Wevb1/IE3oojJghXTW/OIViG8kmgJMf32fOlvhPj0uIwGXpRAq8ZiYvGEeexGXnSlKY/rkvbvI5o
COAkZxJY6RwIUu9SXcYOZYsm5395rEtNWJHRgl//pDZEOxWZIjNbDK6KjC4BZ/R7j46HWHaMj5eE
kPFRfW7YSSGl0DTn1aTJkxNzYvdv3yB+cENfo94cx53dBmLzM441dfGaZ4wOwgexT9b6u8aRxopO
BYLlyTdqk0ZYvrcM68rgoJkjQIsC8YESwPY9YlBHAEQLFU6/Vwy8PsK2cj4ZGikHArnyhhcJHjGG
SEPW1eH8L5+8i+F8bLRIHuAR4WGTr/HCifvAN1WltYMAQ53HV9lBgymHyhQfMdXaB6leT8Pi1v65
GMadq+Mm7+ttMvM588aYVFNgPSJ9Iax9saI4vt31SyRCnQ5Wa3QlSloDbpnRaqDC6SFsdlFfBM0X
v5lbQdeihqn6SyTbvjZO3P8XCrW/W97zYWXaapl8m5giNlC6Fm2eRPtFlCCdFfJrFtZgXvRPZ0n9
KW1JSC4f62ctlPmuR3y59wm0pa9MzijswSbkFw2dqcAUOJpox2TZIlHWtXLZ11fHquUUTl5QKjws
PcuANYbGni2UOKJxTP2gzB4avi8Uni8hF7JiHcCwdVN9Jst9onBFztWumKINaVsYPbJoqxzylW3X
60ndsamToy7OebX/ble/IfYVcckGKdfNQ1rMtJ1BWHet0mXN80QaGy3G4+56Pi5hRiKC4fFw0T0P
hKOA8TOR21DY4Da81Jvljnp8nLnOpnmBl6mQhCzU0hFH7IGyn2bgAqDxOGCAXhyMKAQizjGcpomL
QbYLFF7M0dA9jGZVPM5/tJEPkkb2lpMC4VeZfolx5cI0kKQR5zSTr/KriaAH0yRjfuTuoKiRzyfS
GkKQEfDaebczlX40fj/0f+GGpHGJSsMa+j6/graRdcwTOW+SO03orKuWkF/V3WiccmxChSerdqW1
S916QTQ0MA/ms4HKXxvvXpLMDA8ozYx+RaIMRDPP3YDSWD2EaSdYwrjeg/0BZ6velMQ5uRbsatXR
s5x46lQYOI2pSR44AkKZ8FaLPp5V2RqhRBYzUkd4fV5mr1IVCvfJ9dptU/xuxzXnpkt8NN+6ycQI
sS58Bh+xPll//P+D0JgiLfvSZefHwyLYw8Hqg93qxa7dEdMV0k643BCkY8unNjq8gcrEw1epx2lp
ehWeqWQU+iozsu+HKNFR3XmXmg+lVL/DbadWBELi6O3PGW4KyXgqJli/Pzxogv3i0V1woPjBa5Mk
hGbFb0LpgI8LUl/uT1jnqX2TcfFbMTzHaqFO7T+0yK1tPSo/pQhpPeqtnsdOZx81X4kjevY6E8aR
SdbtsD5pqpi8qD5j22DEj0cBsHmrvgKidvJ2ukbEKvpgci+WY//Tgj/gx+fQ06JMyh7d0S4IQRay
OD3e8R8pub2g53XnmT8a67xdmk4Y7eZWNoVRzVDQk7iZulKYJanC9dnIIeIWebGUPNaGWCYGrjXd
sDY/kMHhtebnriBfkquyLyRCnmHW1mmrJTSrgixgMO3BU5Q5Og6ohRALH5zr1aHCgZ1gd/x+1Eh4
Lq1jvzVeB7ghIgFH3ly6nmopILq5kMMyKSGE3VN4G2mV8TmEubKNds45vl3jcdH5Be5c/Jr4S1MW
zNkfMKMT3y2/omLLKxPjocL2spUo2kQKIV6uJdSpO+BfEfKhU2egA579dk02SD0+NyZZPxpKUKwV
lQwFfzLS1QoprXncYeIuP0JVrcyqTADM8QzP4Ah0hdiukhhd9EZ7MEOT2ddSwLy/tM19LhvZhwE8
4TQRx693bUbRpGmSbFNFwkY/M6z32SipbOMUhokppmQd2PCvkm8TI7CapeOqobP5gpUxysdqbaUM
YM2+ssH5bjvXDyKnm+9K8UOi2B3plVkTWqq8atefslBfLjZk6S63mGrA8ltMPuaErP6Uv/1yV2jN
61XnctFj2jp1fm+amNAJz18zYj2N0l7BXCmt/y0grbf7au8Hnlel6VwEj61OrN9l6Zr8JDCu7thH
hhYHMlxHX6WM+qo72CCFTxINjpZnny8QRfrSywh0JBdmVlv2WO8t6wvD/T/sN2SMfJPI/0gmCaAj
lsveh4K72Q8zYcgmUxOKgmhcDK76eWFw59SbPHLR0hGOgjHnmZ4pnlJLTy3AVTKl2okQwvzdmks7
OStBUKrs8JCcCZ9lqTz1Qn9qjdsZjUcdAK9rU+EMMnBXWTpQWe/Ya3SKO5UhtnSYDuhuw/eoiREU
cZE54yMvQBp4+3VgewzYnzf/pqVW2kO9e/KLYyywN4CFL+7EL8pLAVszN3AtXDo1RXBNamzeEQSU
HNrHDJMVVfrS1O6qG7kXVuz7Jy1+zDGaHBWhQirKEZcc70D/UUs2FLaczvBhKWbGLq8EHQh+4Rkd
g8Eu3Y4cnpabfikGBecC9I8YvgjJvenHPYYFxzCbSS/HL2o/gWgh22xXDCyMdGNyONIDgV8HjR4v
KPcKVAO7rns2QboOCmU9lgU/bFdP3ZvhuT7GlmFCxRCb/+IP8sokslv8QYmffpLJiPUQ13otmtZ2
ldxRr/grxB0Kt5vxERHf/6U9ydeDxnb7j7AmMBUG3pDYhvUXaJfppc1/T0x18VSubvDZktBeYFel
5rU8gRxeDInlroxdCJOwQSEjm4dlthJ6psHGJPzrLEGyVp/TYMtIfhXppnoWvSVOgBKrMgTVLRsx
b1bixPUzFpxOMwy5+pbpj8+ycwKcc+feRsURdYEVuY0FdeYeslUqlxW7dxW72t0TeqthC0iPTork
yknw8d8d9VXv9faj6HA7RhtijnmJ8jK4/pLsbJaeZwW+o9iDVqAKGQf7qkRIOwXsvn92hyis36Xy
hhn7w6QlnF2ETcLIFDthK/ABGYxmfTeOPfhBHty9wXQGkP15KqgpXxTYE7iu+PHOAJCQ6tfuUbb1
nZi9X7OCHbyk+g6bVrL7/xsmlmcnkLVg9v4LFK83Q7z9FgYndd+uK7eylRhNFeG2HFbkfKXgE/0K
/sj0G/C5aG/EuoTFXYjsHW4e+KXrK7JbVMTnKvKZXPsCyZMvC9GxNNpRIFMW9viW906+KNbfgmbU
c9VT3uO6D8uBC4hDAnhz+FpbjBzPP39xuFqvPChviZY5WSiKA4dm5XBOwIhGmy3KbqdX+FnlN9/F
0KTHmAk4gPln203XOm2TV84SnJ4eUH0J1uJhjUOTgHOozLnGu42Fkty6qNg0zts67iO23UjjZiWy
GRMoenjEGwZDKUGaLVWInUH2ube2FEspjYwtAto4ktMjvwp984oCTf4I+5gIpCxlyN+doNEmyTnj
p8qA/XSfxAU8NOdY3kZaFdgueX3bYiQaYv+F3B6KvUsCE7KBZdv51cm7jVjKx6CBuLe6OxAFbt5K
QfEor8CscP4S2MOUSQwnQeU7Xx2WcuGhZXyuTB/CsHHbAYvpaIHGTtfMCsbh8hvowOfCGI/WPQ/e
tSQKCR1FFeL0ObWnJ+UZ6h4tM8XHFszuXScWasYxH2ZhNRbLg1+r1KLbe+2FNZpza1vQQ4dqYEDc
ia1vq0pKiQ204jhSPL5o/zyTl3M8amjGv7OJehxzad2TqT8K4hNt9gq9SjIXs6smlb+zadI2qxqo
ZMX96zImDVIwFYg60jJwr6uq/8OcEve1CEN3H+ihkGdpXlgnzaKFAEIT/fxhmL1k4hMDDljL5Ome
gnjTpd+Zs9OWQrjEcj7cCORzhWX87v0f6g/JWVXvMsOhmSJ67UOgFxkfdxFzSYqXXNIk8S8bITxj
vJb93ghnep/PfgL8hYmzLGtjdvbj3mKhcGcD6evm4pDc1M32iUswyb7nAOzuiWGbTVUPJa+y3TQY
QyR1SAFRF5ZQtoicxfQyz0w3AqQE1tNtUYxOU6qCuHJH4Pto0Jl166liVUq/F7q7VKJI0DJdDzrx
ZtV9mnxn72gy89S/dBQBGceLMWJEvh57i0P63Yuu5kCABFa4OeBuKm43Nl3W6cf6adXmU52TIioK
nf3utKEwyJOVbLPVmygccR4Gfe6uijVwUjpLW4q6Ht+U6oGANIazvhowe5HLOo37ynGM4Gr5Yf7s
ti11KOWNq4fSA/VRVw/8dYqEckfPpHB5Jel0BgRZQv+fNCUj7+lBKLMyTcpduV3C1zTMr92R470y
Bx7LY4IPxHqxePnu03hAFpf3ucG2U2BfJw8jHUjZAK3a/5+XnFOezG3b7KWl53goC42ZOLmBJJ5q
OR4jtaXm9P3dGmUFQrZRCDaGIteozaxWDt5LGJ9MZM1ltvohtZNeir+sk+GdRpCSyG5Qac5ny5Fm
79aYfurcD37h4QBuMHXmeDbBW4VGKVBoKzfbHjsiePGdCGrT9Pm4Rpm5BornMcvDHajEHD7gfDhX
Jiiz6DFSO900l/v8wz2RhrdDFF06neooEIglxlJgr8UkWTbG8zPtPaG2f+YWX+mzMgeLr70OnFGm
CxsWrtoeuL70slqlMsbKRJUKkIWCb8+cuAi96h1ur50QOCYc1qHjBbIpRj6niBdLgEl9qLJH8z5u
Ub2e+9mazlPWFqaz32YbJXS+WdXy2wPhEzN8/bLA8PTjdlnTfn5YsEUJJmvhJcZ3v/0h5zFrgrh9
Vg2m0cVE5zSnBfK2bFj/EI3dwWt0VGjzj+gocru+/qGwY+EOZSaC697XSK1GG/R0XMw2SkAWf7ZD
H8B0cxBW79jHcj+DbqFPuzOufpTyBTyohHXoTG6UK8yGv/QjGk5BHImay1teT5tE4OZOFd3xn4lu
91V3eGYXJLBi3dqdy6EiT0YFNqy1++gOzk2n+HRGxwqvBQzoXcDxAxwthsIAOe58jT5svguOCfxq
G+zwFRn/MvKMMyplB1iya/VTSe7KVXJqK4ZeVRh3q+t6ilL+6GYMe0MrgqUGMNqqWaig9jISIm4z
YaBxdwj7AemJBPfA//suufB0HMa+z4XMRvy3YGd1td7mwueZBdFoTJAXD8KDuRhPTgcFJ1kgeaUy
+DZQdE7Ip3qcbuja0mJEI6/UL6KeiWRCFJgcMibggcxifnfx12i9fjOCQnauMHEadkhQ0xDwXM0R
R6xulq3xRC7e+MFVZRH2Tppr57GThiYBwLjuo6/rlUIXG03xcT2TTaA1fj5EvZOqoOaSnVIMkSah
hfo/1QhL0zI/litjkETczfgnoPeLUUW39qq1gfd0j/u5nweq2n+aDvISaK+CGBl5u3a/vrP+Nsum
sz3w9bv87zWdv8nOi7gSpmwUP2f7Z7naylCtr2YExQ/RDQVbDwx3YISYsaeUPzHwlx8i93avkyvR
pdfae4n47Ho81SuJiF8227wml7rc4zYf96lmCS5Znxqac+G6eWXBv4Mx9Kq3ZpdmJj2lohnLggNL
wEIszNIB36YRXuL9Ai11nCJUh8wl4kMKgwet5MLI+7fSQ8K7K53O0xNZgCRZZgVzp2CdcbD8MZYq
0zIiggnYesl4gyZI1QHqB3NXNO0RbK75+g7rMTZBVOEgLSVbO256LF93UzD1PmU4uU1MirxxJnUr
9i2L0v+YQ4mOMKqXIB3XZVhrFq+mie7OoEQ211e3SVKqoyyAVDHgY2eM2AO8BX+FETfu4ukAsden
Xct5pzFxi0d/+Ne/q/E80oruDd2eLhU13hsKdhQQhag6wenDH1PMXX2IaxsPna/3I2bX3ubHqovj
6Rwtaj2856eTlvPUER4DfcgesvD3u8hIZijCvUCh1Ho6aEPpMXqj1KEHQTm6OmATlJmHwbnDReIS
nWleQQbvO3R0wH7lzGlklFfh8bCbLdqvJCJBQeVEYzD8vpI8OMpHR+Jpwi65d2iJd4n+y7fTn5tO
wXAfenDB2RcpKczfsLBJihQ66Los8pwA4H1HGzUSFwzqAH1sxl3vu6hKQISz65YrzZwJMTk643Am
eCZY9WBNnCB0a6XaEsM3Vq2OgCEnhPIWbTTK10FNeQweSoIKeRtXhC1HHW8qw0NHNCYnSDDz2TPr
VJ+gW32I3aCn+VdSk3Gz0DEIvoTZpSpMshw5WCkgpUKvBUKVsqRziNwXOvZNJzt22eB0NeXZZp4n
ipHqX7UKJGEQxOWsJ7JpnvPQRcKaau5yDtXSk79/SrkeO5YC7E6en/Hm47SFVUPuLwex+3yHDW/R
mV7iWKDEYvpqSU50clLVCWfklJE2PmDU8e3wRdaC1d/L3PM+3HR0GbIXQZvKl6FhCKhTH9HCo2SV
rNfqUTggtBWjNqjJLS9RTJur2lE23Ghc3g11dOQbuZXB3eVBvLRLmLl29Qb6jtrQ4dBoFvTfr53r
UZx8LcG5B6Lwp3ApsfYGgR3rokfKCxnOqx5bKeRXf2CAKlL3etyWTWE/Hnc6JwgyEc+9gX/MCvIn
SiwOTVIeVfnJtv8dNMTDqEagB60q0CSRvPSleAhalozFL4HzqyNBDo0P9cvOVZ9WJUx3Mv9rO4IN
bRrYqcl7weTNM+G9vPKOSi6I8rVpFez+j9ZXCSalmEuqh7TchZGkKFccnRkpqLpcrVWxCLUDgHHJ
8MO7AIRKH6w+EPPeD90wIp4/vQzoAfK1zVzdTSTcnLBoIq9QL9BrKVSDXLYdrDXlfbEO+pA7XyJZ
kHyvortGIkh+shu2aDxNIGxQAIyCCdgOZaN5e1igcIgl2W3clGAtrxml7ZPQYnNLRk7cS4nfc4fZ
W2N8McYLpUMb+p6d/Wp8YVOgpKZoAy/WEgrPbGr0a4c5kfMswRHFkz4LJsZLUmuvHPDI+e5WvmJY
adFt05V2uAGAvrrQtLWMVRmZF67Uep4YFEunIsvMqEY28cMr6jH+VtCRI1irr2Kf+kMX6NZaXLNH
a09a5pbOTaVg89IAGNQoNw3VXqailpFVowvxtd8X276qwjvfYDU5axWgVklwk4EQd2FK4PZ+0zc0
Y3BA4LepD7vjCjmGDxOXMz+cDK5Zn6KHtUDk12I685Pa4OrVPojsxsU30ZXKAqrtZ2CYRViHhQIb
HCEkJiABO2kEU/e5IGAd6zvdu3H3R51Uuq33JocUp7WQ6MJ+lCBHHNiOlov4W/jVmrXIyXOpQt1n
G37BBvM8eEdcsoRLHFgtnX4a4UMqxU7uxLBvnN8ffz6bm3a/jAoRjs4iDdpss0Iw87qIJzUgn7ie
8XPp5DqBy3ivHCFID2w7zYom2DhRVhrOkfcp4RV5xXjoeTQP1rY2KWPrPF7inATGa6T4hFoMZf3y
UVfn4+qtxp2gGRz815Ap8g6nhfmcU0dfkxemgKhQ9rzzqhGwPAwRpNVHJMxrCb9GZUy9hN4Nmmg7
99b4gwKMVC7qoPHvprdnYH6lg5h+vRrJ6jndQQNX9CMK2oSNyUgPG4CyMiBUSj/CkV530KK3/Gqs
EIfvaSc57JagAkiBkScx6Wq2bzSksZIv4Hl2W4F9cmRgo+19e1ZU4l5YJiSiHuhErsDHZwFO4ALR
/9ZucoyHLkKrVDMi0dol7k/CJOVKvRlOeytpEtdbCOIqZ/EUFomQDmEzRhmnT5W/WsPt7H64tU0J
DBTMX4gutAvlKAugZ16uIkXhqzlR9cUnJ9/vLQfEeKW94s5EGIlJg8tzc0LXoku6R8Ut7WcJBpkk
7/3ad2puSfRKR4gi/Q7xy2jjJNj3URP2egiK6mAKIcVTiVy6fjAe7HELE12wnbtU+gw4BNqzGtgS
SfamUTm6ea3nivPAs/FLb6j0wWhXnr7lkcrx39AI/jOIkzzxShEO6l0YyY8ats1gd6cdtkYvy3Sh
m3UdM+sGO56FoVmfUW3LrJUb6mddzEGoBxXw7KXVassiIT05+oUZSmPjeQkRuZ50baNfivtf03Dm
kvDDeDwibgtKcGOK+qBvvjPX3swMAnfhEqjFQdApPCp9812eUTMMJ1mHJ6kxJC41nwq767qc7Mh0
x+VzruDa9ILild6FpMlnJUJT3P9OcqIeD4Mt4zOalwDWI5ACNfoBYzYO4yUuk+Vs+jcghrLBWmyd
NxxZsE23PFVC3DkVNefoz/e+mhFquHUqKku1U1qqbFAw/jNGhjUq+6fHmi+DeqNX4RTbIzVxX5Hv
xmXr8qs0Wh4dVN8pQXf6ucn1jvCaa3GKt1NL6Z2rbx0FlxRMbMx3gwIjvVXQrq//rZAY3u+RdvYr
h/CE9gY+BhA1GogowoaIxoyyZvpt6SJEW5/bOZE/YOXKIPBPDpqYmSkIK6u/YqcQlUY9umO8ruiF
soDWI/EGqB3+pQTttKzflk8lNBgvEm+581Tp3F6AXdWOqxdnD1ugAKwaFQfc9bk8Opp/K4zLNqrV
4fzmIPuQdsHOPwToB1Q/dvAIpAx+rsFK23NWYT9w/yi9DMWdCdlSYkgmtTg4SnLDuL31CnFyt3pH
rxQKChMDo6bSCo3jeCIxhjLPH00+h5Rb2dXAlz6yZbflHRu9xL/kpQ7Age/zBc73uoBmFduy5XBG
mqdFO8mHv5OYL/Pd31WOeuSSTwcvUVeQs/FTN34aMB1tKHwGTx3cm5nXo1csNBFrPFJaYHnH56lM
NVXpWeN35zMiMTPHG8mqsW1DU9PbfoJDFYdGNpM7Nla/FDDkUVu/A8kF2N3OgvRUKXjA6FNN8GEt
TetI/BZdRiBgHXvtgqyW+74BdpWX34LS40/ev9rlzs+NoPKCxuFycHMUpXGCzKsJEfOkjh2qpo6M
kuOZhWnIRZ/ZphwyvzWveOXMTV3U5UXStXtRRLhAcfbcsXwvPddmF0Q0FOIZUNo8jd3lT76AMzeT
ndR37ambii5+VoBCXvsSa5/dBZRPDrzzKra6mKK4AGY7ts4eRh049o8jZug7ydNbEZaf3TTQuq2D
J3Mu3G8geOO0onBzKhZvMrFpzz8vVjZ/gLc8KzxOOVyUV4V0sFdWx0W6iB304EKyIu/QXgeDIMhU
NWtO5tQeVk1H8o7ct5o0ehgu3uccqP9qiNKeipwek2VPq725IZASrGa5Fk6iJcpOdECOr296AqcJ
Z1wxkE8R6pvldWfX133ni8qBfwzD4lEIEz1xkf/9ucinWlzIMuaKv3arRu+ZfAvLNpWZKkbxx2mh
H/Dchi7gze2EklXgblu0Yv4fur3U4Sr2w97+pqDdGw1/BMhfLDxCOTokGzhHr/pl0D428koT1Wxe
bOtI76CFBBqHOvPRmWOq+nmTUc3kaTf9xwktXKAFqq8HNKE1GVIonJfFSdNtJK+D4HIEwcAgsckx
zqY7vZpQmQU9mv5p4w2RzKiDO2C4M2CBTGrByzJKqj8zYqhOxsxRXmL27Af/wORAQZErzItDSGJR
XehNy5EoQ9CcgBVKSAvQDxM/C5T+KTUpQ9vqE2MNM8VCtn3wuajPaF5+ZWUZ1mxbvAotDfnYz9Rl
YE2BAY4ZrosaFLsdXyFgWxMX4wV2YrNRLppzqakm3S2GwHj6dCKQ4dkLHbMahNv20br6jBe7Oa2E
Dew4T3cNaAGNnZFb9/RbyJL+N0f8ZGD2cwkleJWk8nrilKbviMPcrOxpgDtoUJ8KJQ+HURTkcPdo
NejGPEGamdcZbicFyX/JlAC4RSD4HTmcV7S5TxMpgmoC54Pqo7x+uS52+hcI4Yk76AJ3GfOUrKAT
zxohpmYShpAObYUWv1b3r4I56W8CNP6ml1aOcd0w+/7xHOj9eXhv8rVV5RWWqJ3yJzzUWzRrWJsS
XB+ckB9wRAQsnumVMUfanw/1Rx6beGBQwWIzLAmqKQsTlTtT6Zdx7J/bqN+2KtGQUnd5JhKKMGDS
jwL6YaxM8R0hdL8h1F+HmmPKtUg4nM45RJdGhmag+Avuo3NAwtTuh2F+4+evnqMaj1VrDUkdIiOM
KCJN66s4fg3F/F6ovbjhbgaYmACJLtucG4CfABA61SFZmWIFYhVqNX4BRNJKThFbAWMy2JkXUqid
7Lgiwi6lTSCrHwqCYpKyWC10Ucb/4MLMNAVYlL7bDCE7xOaIbGlmDMSFRvRuNUdt/ET6Cp3BqOY6
LxT/hIj8icT5Y6sdGms1mp91ILp9T4NhtQbtEGjP/qQ09obiv6Bw9mCjum3ecuRz155pLjNN4RGA
wmkj7BfFBSbx2u+AcyafU1Al4/aFfiBNnCic9YrkSDKPpwWBhzPmodb+ZGsffDoJ1git7oI2ILXR
eLw5PvdSjNM54r8SLrtTM/uxWNMn1WQh37Y7UfuaQVj5Fm9MrCRdmNKT4Ic8IkYazeSUcnH11zVe
XPGIcgL6k9riLGwT8QPn3gsehQcAEgZNAh69Enh8oB1Q7ao2RE6OnAV9dob3kS9pbgqAjOkK+oma
NbRPEkZsWljKRcGn6p82jcRl4udT6PNtHj4zNDh7t8kfrho7bsDcQrPrhS+WkEsdWZOSPkPhbr/3
+XWitVDWRrUkTWx1E5wlN6+vRMMmzCqtnW6pbGC3BUnGzIO8KjXB6k3CH7f6HZkqgHQLKv2EMBVW
l0MA753s+WRJQX3NWNKeSwBptnCnkXxth4GLURHWHt5IX0omErrXtV/r3Kkujz6gOeo2+TH3UrDg
/AMnJy8hU+sfCol1MMr8Q030ghPefx29YonCVR9gsc/kevpNsc+4PCCVOwwaNCjBeE7IFlWcmiL5
8zbNyN0x45ys0A2Q2m9TC5w1gtfcEM2iPW8ifpJoRC6fXk7OhQCyeWcUMWd3pNvVULy8E2OP1P/f
V9dewKKKfRhvobOVu0AMrsn0Lohut4UpKOzTBhYIGA8EMkcEXSf+0KfRH+E+bVt6ay4+vvD4Nk1m
cecxNtBJgKNKvxQ3tLQkZ2b+yxgEce6ytxyhcW7m1cPe8QgsRXd592TjIepFhTehTtll45iP/+bw
0vDUvtUdBD0RR/BcxrGGryk3TGe50xR8oPCJ5cFS3I5Jlf7CCUhI3v+8k9yT6gUX5eVgzL9zqoSQ
u5eBaT3DPTCI0gtmfrYGQZSauDRHT2uy0VV7gKu7xPNepwuiEL0ecjwv16dRsL5qe7uX7kw8GCa1
OgPIu0gQBXz+JUcROAaC/o7Em/k2Xhjl816ThbtcKAVqvqa/rQncDTTVg3zpnDsSFNbnuc1I1HxI
5bhpLCbuknjSxPGFgSYu/yspwZv9ZD0EPJcq/w5eVNydpjghU+ETtP0gx3adb/yrNBV50Pk+lO8s
qtcOBdjXYKm0JYSU6B+fKtG9e1ohIxiJ6SSi/bNlhEqK677t/75jnSndObzFG1cqAnFx5dRMbLsB
UdMNe0LQAiMF2pBvOhx8MhWEFHYj0oPxLNaJOGayva/Iagem+S9AcdZldQ5icCbnwq6O25ANWp98
c5povI2uLauBQCyr56cGyNgaD1WkK4i9kZNEaKlDSIEdr1wJnbJMN3EZb0wS2Rnd23oDW+RWsBn/
dF1ZQGfGHWPIcwHJX4uWl/ayPCda1FVCx4Ck99xG97/52LpHVB3/YHOi/YwrE8RdkK3iavO4RXuP
gfy+sNy9mFl8ixnpzC9u0PnpDExgB60SDs7c0AKPQWir3XCGyIvXgz6YzwnH0WPBwcNuVRYSJvd4
7cku5+tLnSSDUNw2lI9pKKcsjoIZb01HCkk0/Ipjoq4ve0nNgVHXaczdr/LoYv3L0q/BkNBAU+je
7cuuIEMD+ABVfcDyfrfwfXL0Hooy9EKs83+3fElypJ9NmPLuQTsgiy6krdjJlQe2Ev++EPJKmC8I
MRhW0APFuw/AwlceYdIMexuZERqhvnJoRyOrjRWe8/v+F8A0zs0eIrNpPKH+v1qlD0f8ec0r5yTp
33ojQVmRAUXiNoSDA0zHnGiCcYDwOcnwqgD/TwegFeAo8hqpTBEvUi13Hto3tynyT8FaPqj6Yzi9
70m3XHIsY/su1CGUUcdzcXZyorgfPAbI++cRzCFCdMh3P/q0r7BOBoh/YTYNZU4VTZS0nzY+lBV9
ZSQznV7OqVif1V1tNvit9xkk8VhVNmLTnPvTetddReQIJJH3eG8Zu05PQl0YWUnyJ5aXV/BFzuAq
dqrIs1oXTvC7XdkGq5JHAXPGbU+O9SapX3f0OgG08n9AoMWNfTNx/KxUxKFhJg261E3sBgcYcGNl
PxNcgRKuZFIbkDjJs+V0EA0b1GAtyJn310Lud/GKvPYnd9fBkfDjglkyiWSkfLRgVZZgZGem6Mjy
ylMsPKaoVvyuHgdY+gUOwNBEMysNkUeQB7B1WmtBvN32utFTSthXp5qC4K6N9Rronbq3RVWyfEwu
jKVI7zzuDnLGzylPASD27oOLFSU6QwmkIOEA5RxL0XCfNk/mnAb3IV5Qh/kMYF0oQhQjUbSF7+JI
A6FCvEq152xD2KY+ChvMe4uBmohLdRFHqRvY5HPE8Oe327JHmp3kK7XmbfsHVOmxYl27bvCl4Mbc
9K4rPLWSnW927vjWUygI4DaRH8BCjm32fYB1z436vvJiZehR52heVSYY3uoBn6kxYvqtQe6X+lY9
bk/DBPF3+kWsgC0opBKD+AA12CBfvU4I+jdngj9Qva8wHZ8odyh0rHoKHJyJA5qDnVem9op69DBW
1Q1lsfsniQIEeh+z1gK50cTAS0uvCJlUY7fd+tBCpSAY47Wf0NyWx4eioR5RcOAZ9fZs3+vrvR83
Whw6AmVouQHsmra/FUZNbnVX6YfOb6TLikJ8dV3NPzSnfNHWkDUw47XrF6HwOHU9tM6PlgVbxTLM
BymBVx6Xzdl3RVaO1wOlBRYpk3PPWE46NyCsr1OpZ7KONpGle+Nu6t40W/0f9DLu6cACuzc1X4wy
AleL3tha0PUnbiDNcBsyci7uYqUMBqcffU+h70hgMtjly6/OYCnCd8wbtxX9OvksvOpDSk0iqAXo
l7a0Mqkr3fpahaIis5/ns38fjF+ibyKwp5xAsMe5MsVPFHcJGvgPUbEPT3vvAyv+cLJeb7Jmyzxt
8WxT7Lf/w+gvSYqhVZ3vdwC8xLblOpprb7WfBILcaQC1aYR8yGhKCwDbeSPWiGlAAYlWhbqquBhW
kGBQ76Fd6cg3/xvlVrhbmN7TzaVtm5Oq6jLwvpH3uzwgXpy53F/RukAr+8C8ok7czoPnDvRgfUkT
tZhss6xe3sTBxHCg5ehseraD75ROlxltugUMRXIEEyO6SBNGjjiQi7R9IfmetYiTXffITYYDKrsy
npndqQLep2nzhdoZxHGcY9rov1m49AMHsBs0GkyoYm122RWa01uHzQN9iMUqwDp5BpO3u1rYV3QI
1PDkAZNx6nzX07h/h12IsosHpf14czyXcrP5mc5CxYP7oxzpowfNIcD06HNYYduumURU//zicDCD
a7BIEfFFUe1qTf/jh3nJp0n7352IUGM/1h2BcH2xHrxOLtzPChNQzfVU4Vel7J1r/XNPkpooqe7E
vD0dWqUtrwAwbLMg8TZUlMp0QTvYh5pGPabQUW8mfBo51RXJqbHzvi0uacj2BPTblaYb6yeEtZkP
Uu2/OWSSfqb347cyz9e8aFEsbrPlwCu8fEqGrkHYjzuP1Tw9M9MF+GcoqXOU8GiziZUs94BvjQ05
IQvvlE3p+2ZY0wLCjBIPRWW1TxY9PccTLwvA1Kyophk6JR0li/nWrvQ7NV/XxRZRPXUPaJoEldjb
lY3V7UHQ+x+nsT8oIt+MZKrfxw2gNuK3XK6XILSq2Rc/sZ37CxzqRQSfdA0sgMmEQaPI2mAIMrH8
it6EdUdpeICwaAEhxrZVdo+l7ciEpjKwYFtMScM4M3hhMjK1TjMFZgUXMF/NI2y+F1ZmD6jNsZDY
z9MLshZJ17ch/JOiEHYn9n/0E2W2nUK7WPjKqoSfcF4Y8p7EUQkwUhNE6uHMhclLbt5JbaBOC97u
4uD7NxUWIv+Vnw3zk6kzq30L/3N9j07ZurZIPO22JNQU8XTSbNW8f6LY6LpztLX+mBwTjtxcksiX
vBNxFxfi2ugpCGdka/S0/oeoQUI6R8bq3hWN4CY7Yf0/Equw1RRhef7X7YlaSs7Galf5GN/A3bxp
ExhEn6nODGV4hE6+fIxDDreejCa5s2B1vjjxjWgl21YF1rdoIMu2wnrNNiCnvMKIgwBXCFR0B+8S
iv6raRjZOyCG126wa+vqzelyyVolzF6OAV4259P+ODeSIRQ2PCPN2yG704xuCLYbNDKHMgLc+dn9
nnWbOp5l8LO55cVRstqzdhwKMWywk5Q2fXkfRTp7Rmu0898gggl254uC1Dcd0mmwzsRzVMaccPrt
RaBwEnX5FDis+VA85ZjI4W4t+S906tBDeXFDaiSrZhnPeLLo/6Okpk1DNrL+mAjcr7J2BByaVIXp
qTaQ+dm2/vuDGLvFAEJaiXcLKg3QLE/eITR9YEYI3ctmt1TDpXqba1MO3gpcP4rq+cy6Zbdq4Bma
XfZgBjlIppp11z+D3WG2eiF3RRflZKUP1N8Q1KA9mr8c0vB2AGX9aIDN7AyA3CsRJrvoqOjhfzG3
FIllwUinH2YOup/rCnCcggMJ+6GXKhoCSewV2AQtwAlOLVcdIBPnUbEN6TAVxA2meL4EuRMuKjuM
FwFMwNyCHMDfF1KTQD1VTxEvB0fgatpXnTdKI4/1prxCdClw4CNPGJSXAHCc3nBGOXRrzbQr8V7H
pzehBA8Y/rr5XInRnpu8mChWs90uYb/t9s0X2/x2XdWVtWpOcTvi6s/W1AVcRXGQ2InKKS/ED75E
9LNZO+beM+SAz92McS6d6BivuAkzNL9onCGk7ckmzYlGHDN4gG8XYdt4elNeCsCsOmOd6i6Rcsf9
sNVuJpjAvvdiTGc4mMruU+lRp3FC3hIyPKjVAmk/1VIL+YOilEs4R6r60VQQpNhDQ5q+IlSxG6LW
EhbJGqnYL0ztx63iftvRyy22N/9RDRY1wl89K++/O+fFFX900eqdxz98BddlqI/kbVR4WAW2JQOz
ioq+D9eAJOvUCMu3QL/RBH7I9RvVWNxlqfw3nXEKtE8hOlWOaKqL0QbhyxFJdsGQdTbNjxRRuzR4
7uoWOj/MVPqEctR3oMAceuH4kzIUYu0W5Kco6qL/oOZCeurfaFcig5fOklRm4YBEwWG7GLhWycd0
0nKbmqMMxC0IaiBl7RnzZgkX3KN4yqnSDTU8GrrjUMIO2G1Frfzx/Hn0OAPowPA2wUa0kN+wz4XU
lrGJUQULMB72gatSlS1uaYfFUiau3HzkjE9crJiM8KcDPGL13aTrZFPRW7bWRxZACFS9YE5kkOKX
dqAhrdjW8yjWo9butUOcC78/Ijut4kFFrd9DYFUWlaLl8zNguVsMKvyKYVpLhXIhMStNerW0RG2I
prCFtJxNKRPYHmiXQaDB08fUg0pxj5NNY0IGDLcvwQ2iEtLKRG5NKIPRj5b7/OA9ecJi1ecvzA6E
O6NFpZMnVOOFlBB1dLPydh0M/LroLjFzEAsfWz0N68DqSBMsBTobzdYVOngQR4gzk80xJMLfjkaF
8oRDeRxoIpx8glmuArw1LESLlK02jS5pLGBzb3sFQ1VwJzaSupeQQr3SXIrlhjRuT/kW0V1Iiv30
VEhkebJzXFQYT/xf57k8mYyU0uPbauBKh67thZ48huDGqB53icZDI14RArurUdC/4Szc3TDRhI2F
8SmFfTgEnl3gR9g2xkNofT/D3qBnNLEarvsR9FQtTMd1FY0bNxDkq6GOc2cnbM4WaWnuqhw6LMkW
w9t8vNK16s1mpxuV41aPr5p44CkBzmAPaMk9zdNGYXN63IZR9tfFM1CEmV0iyfvGP3b/xmJqApcg
iFS3Gwk84X+TnPM1d771rsA/BBbyn1VgovlUPbqsdmZbFGDvjpC/VDuAkIOv/rWM4kH2bj98xoyU
BMFfxRLeJ/hFVe8vqAptIKVDKknjl4PogagenUDOcK7SndQqCcFEgCyp8BDr38a97x3UaE8xSgOe
AXaOPrD8wtmrqm5MncSVuo/BTar09OsO4RSkNRol8u0j1DhuXAl0F8GcEy0OZx5toDyEKe1nP2U+
a6fA+iEq5pcjjuvjR1FUvoSbEvN+yGk9XxnrwuIFEsZ8brPF8rAkMVnplVATgsIrgpfgP2LsxLIl
gS5eG42iGNIfWVypcRJrejYcBg7J3hcryAzW0rBNGFeMAqm6zne3l37nGRn3jXXJecru94QmDvXZ
UTJx7D2Fv1dOw4sFPPsLcE0HEA6o3/JdldoRPCJ04GDmuAbxQ0iPWtqJTiR+3YPDRAMcWgx8FGm9
4WYsdNc8WPsuer+vlnWmfeaU2gJRuIClfI6LC6gFFuTXEVJBouIqrTKnPzZfVAIcLJhgUJdi7Ovl
fMD3MGqf0Sdplvd0vrQnqZrkzICil2QnhZ7zBBgz4MeWRIiSaaN80zITxmAf9VnQMu/g4zTTKHJ1
Gx6z1kjLIhMvHN8aUpmofukTTgvbfmr3FwCwNnHmK+DBRV4hte67dPGtzY/Secai5DCJVvkxMhOX
R2COnysCzkGQXbYDya4SRSED4MnP2xYpIs9OA3S+iqZGih/LCnUH/pN7v1lJNQ1RAsnZ7qdGkz06
FBVIfTaueESkv8poAs7352n/moiVQjAomCxN6aMto8UMJFNqcTPaEAn8ZkphZsQqj7kE4/IiEkdx
dHV6rqjfsZLG4izpc6u0XdwAG/zeCqT+h86LjTApT9PH0JnEugTGYU6HpcuOClRRHno/09DuL809
3s7PlUfz5tfBJXN9MC5zUCQ3IrxojR42TqfU9mYSDzRHbGQc+F0ln/Fs0VDrOB+8tJh9Us903AVD
B4k1vZBuHFWZeTqpsh4TpeukurYWe+TuL7GEDZ64Hm1jvqsqNLEc4g4M5dhgQElF8F6EGxpRmg4G
EAmILI02zwlNrGVrxxBhThFlrFbtKrX+8eg6wEKsDFGeivVX+pm8aaF3eESBBE680IH8Xusu92DR
jxdf5DCaiPi5mpH1fvjXD4/u+L1EXXPiHCfsX2XV4xm73YcZD13qDbl9Y/D7ad7cCQ7XtrQnTtrA
NiZs4h19ZKjx00LYDF/dWEI1QD3STpFTC7EoyE3KdeJAhyYSaxQtvemHDwlaFEpDacYsmKZveFbD
TWKzP5BAHOBsfMJFM9zZ7nyvEGofgaUWhjn6NBIIrMX5Do9LHOUxYd64NVPpt78h3i28DLxW/U3t
mJGppUrFVcyW+GqHFbtcr7DqBJerxYUhWrbF8th5Fa69eJnX/4nwgdhHZAhSRRD4Z65viUFMC7UM
PGikAXHLqPCbgrMJdoPYmvKDm492Jl/oyOgK+JkhoiVy3Kym1IbNwjhvNd5qNzD03HRUziRPQ9SM
dIzmOTgCwXEoXVBIS9FJ9F6MM4uqLqoUbHiDEY29t11BGFt+CEa3vp8s0DLBC2ZFXl1mOr+nhuXW
qBwRYqiQfwjNs3roeIk+2DGwi5Xq1yRwbd/603Q4erST253vZRUwq/+KxrW221IAJRSsbOFFfe5/
Okc1OW3VMWWAsdHFRTlIMeGzhW9fm1ePk/Wsg2jBqP0OWZKhm4lBYzXDcAw4CKRX+hbY61gbs+uT
14d+tRC97TTHshHmHyHNjCjXS4jOutxrYqfUxXF404CY7ziWM3F8Gnn+qCBcx+xFnqWyuFRfltkG
rWzweTqobeykbm8tPxeJZKoEDhrQStNCz0FlPYl3oYSfZPkNQLYxj2bezy4OOXcwMQc3XDQOJu0N
wD/IZOjUlPsl9W039PzK3u2V5McSDjEXr8VcX1nxJvj0Bg2ziTYkiVYoldSuTlw9/3Y9ltzhxNKT
7/Mq5u4mYI3sQimoRdW3PPd93CXN2bW2q5EG4/6OJ2/jcCz6DoXx5TitFm2fXXWFRigKQMlB7hUn
ymE4A9uo4D2fcsdHaLPyspOy414mE+zuPSK2ZL208blJFzd3kGzmwPkmXvgdy6kHEF9ex7vS3D2e
VCQA5cyHq3CR5Dm9tXtF5b7YOUoeGIPz9PMwpqOJMUNKYOl/dCYcb/wte7YyiFSPe982zzIL8xWU
xRjfK2CDFEYJq5fm34uw9MNdZx6aM/+T3xrPqxht2v9xPc/B/fdcXebv0wUMGXH7ctf1Szq/k771
6v6Gc9az/u24BJ6XHHttIorxy8IST6nPgby/xk8vxWOuvYeCMy0B+FUslVHch8BTWHzgGiGiVQe5
lP7EDLKcmowdGJMTLLdakDd8WVSJKiXmpNAoKpq/rQvGgrn1vsDR3oF3C02n09oYILoWZzgvNj2q
b9xqm3zrAckaqZTcYh9BntlQTtQN/6iDWPjiHE1ojFKPYdHGUR6QzHSM/FCvmrhk1Bmhy4unGcO7
cXeupSOuGlJHkPIcA8srY6hkDrKd75Yb5JZHqXncYAJsfFvGZcpbNvDaEoY/eyB97yvVrDmY+NNG
v+FXXckMLUzDC+l929Jr87Fks5+kWYoUV3FmQ+LvYq0x9yi8xNO7NrvL1zbXhNpmXrXZ69Kpd8UP
jQ4nc2c3znCaSQw6wqoQu3dERD5T2SgpUbSqIkfvMiBUpQfCbjrUy0IxZjfaCt4vnuEDqKSocw4C
4dH0QdDprBJNmjgt3VbN/+i5nWjXGCIdXaZrVnuAzWfATEwO7NjVUtDDabzgTbxSCeRzUpOjaw9l
YDvWJDAfPPpOYK2ClEb2aeG0kcREeuQVlZften2zNL0VIJd0W9SEy4E9ruwINq9fMMQkbayPp70U
rVbTksb2g0520Ponf7rzAgXfb+RAvtCSi4/LKp1VQ6jRWzcYTad1AXRRCe+F7AMdqHa//SqVKxpc
p7tqxQsGUHuTsUNc4+9XS1WBUwS+QIUwZuCPBJCPB5ietfeSeLm9HH/g9CPpzNmIaOMECKzM4wfj
DfUxpMEM0BR7vSiBC1gtRvWk7TD8cnm25fIL9m4J8fvVi2rOJSu7e2og3EWTwr4a0MlxpS9Wwc0c
A9DrKbi1vtM+6JjXTUGW9nn9MwRTSMKOfd1Ivfzi8rrBrEo3ltzn4PnArPr26qUiG/2aTrATEjX3
8Zv5ZYec89VUP+f+7kzfdtsJGoz6d9QN8cZ4VKH8hOWmPDwkO66lhWybVNjpBPcInHSs2JvvXfgs
Gh/BDQI1r+YQLKsWTuAHr/HCC5dotkGvybQ/Ac+SIUtGYGPiunCZfCQGHx1tmOaAci9qLf5VG1kZ
sXjHmBNZaeSl8hfBZqKhwgXWv1ZGaK9opmUasXEam0twpdoYXjPgEwqnWroMeCaG74zR1RqhPI17
JtSjuMbp5Adw5rOjOZD3dmEgfnd3QpoGy+ytWxX3gWSdIy83Noc8EkCh43r3OCy/6FT7kO+QUEoy
atYLRWRbNpx9JPRU1XYZbVQIu8iWMjm+DiXVMdKqPje50J8UauU8a9ohiU2P3KPC2PHtbBRGaW5l
UmcWk6Pwn+Yp6J/5GzAvOLKt/XWBtJCz8dNEMkfYlpkZpbrQA3Zz+KLrhKb6F4wv2Dfcb9yRdLWk
K0+NzheBzgthqkcPeVxbXyvJgzCiDGX9dIu7pD+pq0yai9PmMwMhh4GEf0ZEIfY206LIjQv100qr
gOGNZl1dpL9FJM5Adtr195vihIvOI5co5Z6XVdVXJ11PxocS92sWPiL5vS7SDeOdZqXMQ3VZAnuJ
jQ7jH6eniKQx6AAZXnauJhnWT8Ix7+zlP+CGDdc3tTubmZ4By4o0tzl4zmhMEyRjWG2MZ/hSiNAt
gqrLf4V1AJWWYykWqkuubykqUnLvIgGP7PJeMfy4tv13Rl4oU8k1Su2RRLVTF2NrIavcBJ2swd4Q
/ERz4DXNJ1caWSUhzWyXpKfN+LX/4nIsG1tN6b7TwNIpr7lu3BB+6LsfMQ5d4wesqHdg4K86xC0r
XQmgJdTMOABqj3D1+YUkQUd7I/Cr8pccSJbK1cHr4Yh2Byy2QzotLQhYl9GDeA8R3g8YpW+s74FO
fHA5aFRRFK9VYBd6E+c0jK19PAaUuVNzSrp1qqHyq4UdtxBxhVyKv1+q/fKi8W/+8DjXOs8Dh+wj
zqBF/ZOcEFzUgJnUzL0/Yg+DET0GSjTb7Mt9peGVlBQs9RgZaleSMy0r1t/gbEQSpUR+xH6GNEXE
ZmM1c16dyB30CjquSzd3a8ENfmjDqnMV/Kd60XCoFnI6rsoD3biRuSyaO5i1i/oIOBKjJr3XRETs
YEQkVP4qsdy5lyUFQ0gMoE6V2xn1JDC1cg+fLakIeMvKv3yvgMY7MdiCwuVp15319zMRPGzZgSkj
FTfe7FFF3xn+J2F3FxrFSZ2tMYQUhSee2RRhrYIRmVWwqKHwcc9cQpbiWDAF2XRBAg77VerZ7t2g
8twdGl5fBhTWJoQRGsXU8GiqOfmz8TfKQ2evxaWSRCZsCsdmpN5Ava1tP5agApw4oUhJ45AR5bvt
Mk6cnt0UaiXCtnKGD/7czG43vuXRU2xPgvK1tCeP7CNf16Kpi0EmFKDxg3CpSFZBX1kuvPEyOc+c
Hr4FSBP0GlQknotFafF5EWXvfei/K7bt9UVA8HG0U3AwY+p2hWIrgfrcYBDoRwcDSkJTwlk1xL1m
9Lq1vChJudpR1XSM5/cThy38+6md/q3Vr8HiWWe3GS3tjR12YMb1xFPLa0+ZXADjDkDq9fTgd3f5
WU58+IlhwADNj+oSYV6f38CPK7+bPIo69JbsQn1r6ghEwVNe8jNVKjqtW4ObSUS6jaPJ7mMGxXhi
jAvsLJCQL+JBBhbmnVpRgvuFAa6kbFGQ19X6inWjZNzDlRR3bPqfTnkcL5ATO2Zga6XDqgSPkqaU
QCplxk8ZDrhToNPaZJPkpkoIIeWx9svJM5unxhbZ6sPbrDwe4HF1TVh6Rxu3GgrEcERTEhTIeido
FHzJWC+MBqeWaO50SNMo6Q9b9QJJKYZuMxW6dos0mTNH85KCj00E+r1V+C5VjJ8uuvcAmML0jnMn
uo4SD/Md3J24hBA9cT24OakFWwdslIO4QHP+SkConpLRzhpS6NROzeWoWtP+A5grT2VG3TLZOfMN
0yU7B6A2BtHe00uSPANnk/ABgrUxZVtvqHDDaC6FSz95/pjW3EZPE4lxsqtSse1wC11UqyxadZG/
EVJ33pMm9n2h7ELCrT4o5ul3yyS5ASorBm4OlePXf6lGQ+0p92QcM71+10MKKhGmIC31nvH6tYjs
Zf2vrCqfLPi5QZGgjmPi3T4ehePlMtSz7r9nNECjKXAge9EuLgghSk4H0OYKMqv9u5r9o+jS3kTY
KzyCsrWI8lUjQ9PDMtwlJaSjQ7gtTGF5bn1MCpmyNZ+SFjDTVQUSrc8mCRaU1bUgECkMWl24yKKs
Kdf+NHxTJjvHyf3EotPKY7cVK3QCOfsnUMxl+vuKdo3geIaZrNleC0w7D/HODXQZdaUttQTc4V62
BA7T5hkCKijPo90bMZtFs+2I9YUpNAHYtEdXJUfHS/ib855d6xU0gM0rGo3qIYWNfXO030LV4s63
7lWpB7eOqzQA3MwLFdinL7WOGq4wTNvfdxeeY1/OjGC56PQAXybj3wnEjDxofySj+IR3qT3dAokD
IhmlgmoayiB6SJM8evH3gmuSb+oUknHkyxvV2n+URAOZFzE6KWbSgpR/N3NSOPYVa+KU/2afV/K4
IXtttfLiWtzcaP3glWdcZ9S+qmcaDBVMBRtUugDdoRr0SyclNriBd4N6aZwmEmZieeX7dqNSbdj/
nqlguMcg+UXHL9b6YCOGEdwPlT0ABc0H62r3mqi9bdQazcw0rBoFYR2UODCroZjbTg8wJgC8wfFQ
t5tqopOY+W+7Y/u1fEaA7/sCrZibaiPZHr8oOKIvl9CxXx1/lMKU4CqmiDs0/eKXJIe+XKCy5MSN
TX2MgfdQslXoTjom4rsglPI9byD60CCR/xA4VsW9MzfACgykr9EugBG6WeHHjN1OlZ9q/uVIDR1Z
830nhcM4iTwip/Pdap9vK7QtLgJ2CjFqKnOc5Hn7PBKW2ImfK3sAJU5LSNT42bF+fAGWASuSwBmq
Svn2mhuL6DfYXtfCXSfTplmd7VADFp/9NNtn21B+0RRJcuZ4fuq/ShVdOlzdkJ9aRwp7K89sLc5e
ZBpqed3+Jc8ZSh2API/p4tj6n2YwyjMVgs/bLK8n2R+j5zEWa+3p7wCMph23452CBtVxS6cHU+y/
zNp5AXgM+Of0CLyQOCvXRsXfZFjg7+0r0JOeaH/TqQM+J1NJKL61xj0YIFTjV7lARAE/MWyBtpBn
20hD4ZgXA/+OqrAgSZzQIo7uzu/K1TlyiO9NFNSqtewfLzA2LppHjPZSYofdqf2AxfKOAO3OTJLV
ZxPO3P/xygcDajuIfAwCG3S6w6Kou8VnSqsGrcwYhXDuN7LdzfgGp2QXqoif8GT/ure1dwpv0bFq
L8QJQm0uOIrCLpzdcrLNZdNUmKBvPMBQH+pE8d1areHy0lgMabKbmK8pBdVJNJE5TALMsLoDNfPK
INUhqtxYgSWN+081IDXNxaRIFi8ACW5V11JQX9mKHiYfJ/0OZWESgPyMP0qTCB0/Oy5JaCPFyzmk
xVE9qnhHmxKaW/q62Dsk2fm0MhFQC+bWleCH0qBT2Ut2N0uGkjHLwl4WGCP5Espzab3iA5h52ZoC
OeMHahn14pwjoTmsbUwcr8HgfwC++m8ivuqZIyhE8/2AO4LFG7vqGup+lL89xmz4O/3WfSFGCW+d
Z8k3H0wSmtl9ipDzo7cc413XpNvdcSUQRT5dRfXlRkTyawlFRA2uSFIGwmXbRX6fJxCvEPjFzUlN
dbqcSEnb2mnmowQGsHAZ/6VZO1bKvO6R5G1wv6nFCfmeK4kXZOE5JITNW97gt+MV14auRgUWf4Fa
P7vSLQkOcpUDkyYIjHvYNF0GqZTDg+gb7Gv8rbabyiC/Wzvx99mTjZ57tXMTaGEDBKYMUabbFhnt
Bb2exDiwaDpMUAodhpGzB7OVPjsJolFS5CpmByqNhVeYKT9Inat2KjfjYWjvp/ryI8yhQGpm+OIt
PVyZUEUH7mWwxTCft9QHHdgoyRniTO1oLVqg8ZTaZ0NYAWtPyLacJ6Lm15VdWl4rEMl7rM2Rs3xH
+nmoZxrpDThjtobvLJz6sXkY2dBFnj3ak4fuj+xlN4nuc0SmEBwTLAbziVfA5kthvBWu3448o628
nnOdbJbs2ZQbWz8wn9h7ZBomgn5kMVwfl0k3ImKLB3qymk1CbVdfVUaCbvBkU+9Ddbxapo2LJ+z2
I7wa/fvtz6OHvPn9TKPEX78U0rXfInHFKm/m9SLhaSB9zDMaYxsW1kOdGs3SSRRGZ/YMUq/ztXYK
J74AtjDHdp7JRhegAXkTdLwDz/cUNNbWWgx8zDP9h3A5khvuCWtGoZZ9i3tPZsNp+vA8+k0Z3d1l
k8wT5Jshtw5Uioec8qmMwUpL6KaeHtmrKGvr/qRtk1oOMX8MPpevMZYm/LJwiEyVuXdoVQMMy12d
k62iFBC8NTva2SruvAXvsMUzfI0LZtEjLdwmafTsruFYfIV1NlJuHM2YG//xbHHsSK+07OLDe2zm
IT+sRoz5h/UxLqsESeLYC8+MzFsrrg2orGFnsjPEp4+rkWWaZsQhEfUtbvq4mwGogkaGX3Ak9uqd
KaDYEQFmELKWtmM654N/Ttc0QIFe9Ll/7FxCP0sHCUVkxEfN5aPfPgP6MwsRxlV0OUV774qpdo6W
RLpd0nt07jIxagzYoAv2xc10c/xCJtxELl+yhJuABtzCGoM1gns0CDzOkcFklt8RbeNvidvzUUst
YP93gm3WssbWTtnRq5+BDLaHSM/BzWx+IUWDr6pvQt2bPju709B8afrAa8xTxQMlV1YEfGd2tHxg
sADOMKdX7gzW9Pv9kwgl3MAGpewLhQsXjyfGL65+5+RSx5fByfjYGbis5vlUd1fMUWUy5gixZ6sc
M5wsjOPgY2EeEGtJhqc4Y5hz8XpA/gyC9nbY0HzTKdq2R8A56EoZI51ZpzHVPbRtmYnyK2O4WiTH
172cMF4gUogmy1rboFvBSfEfJN8NiHJuzlOPc+BFB6hazzvsixWnoPUguLit/3w//1pqqQD6XHGd
B5a4XUzzz2haoTFuKoq5uWvQPPtTigTlHmhjneupVBCyzB1r8B8VoOYN8XNsI1fhALpXYLcjn1fy
ZIyJG3AfcJJwLWtTB6STRYpx2ejkvsfWBJ+THoT8n5MzdgxwH01SUFw7M+ooiVxjRTEBt6uIlDvJ
QAf2PECjSErn77j34j6bIKL6peSvtKjnEtkiL/rQG5DNhG6ki6Uodg5wTXkxaHDtclH7NWaRvOjY
RBmcQtmWApmHoQm99sU74eEmF+6BX0pb17WtIOIGdoTCWWnlye/tyg0wbQBrqumqeNWMBBD2/DQB
vN0ZzB1cbJJyE94XKh8c3CGe9DE/ZswvIelxs1+ni84zy2hcN/ITaFQ1dW0EEPqPfDnDBYhomdiB
932uTG4gSiHF2wSAb0Pyl+ALFbX3mZHgdy08A3kPi0NZvHTiqLKC5p+nuhSUjFc90iEO9gAdm/DD
yMmuAz9GkR+qwiJhQcQKWlAbzOtZnH6QVnEsHqiMDyczrWdyOvc88VmzaSptAe8M3KYfAAKUu+X+
C9b4YdTqYneLCNoig+8lzlxHPm6uXaHl5eAyS4Y8L474zpQ+le9BGs3KYb4np3uZsDz3ExIoN+L2
WnQY+0EEfCaCZNPNupscRu5tRXOZWb12MK70hlaeCwP6PPukbbkCM7PhOPmWGUs1gT0xDNv7lekM
sP/baaslIYlU46tNOu1er9l0t3pqIqmerm9masdSj8DiVpEkliNpDRP8jd16eGZXQs4a+bRAY/b/
/6GfeU2+Qj6H7Uosy6CQDjnMnWLm0cVBL8lycbyNo0fi8Ctvc7/KZ1KyLVEaZ0whtxaDMK43UgLT
K2eYt+HkUqzxsyyGo2TtKhPHhLh4/D4CIt1ItkdzXPf8JRwbj+sq8AVgJLUy7aJODPOJkBmEyn0Q
wOrMD80wkmWOT399nNKIbB00aIrsW0UDI6NHOieXk9AgbK3rImVNCq96cJHr1Czpj8UD2i2hRfY3
Bw9EFgGBDXdSXo+68E1By5icrQvgWPMcSkPv2lCezbC/QupVr7f5NOaB9FCHuMFona3yhUIkJglH
pPKK8U18D9DmO+2FjIJGLrcN6KTiYCNgcdPrdzgJpaHKyJ6+0sdXfbrAYcGI8LGtR+z6fapDFjqD
o2GB0MVu4DFtR7P46qnwZpxaqOPCKlqu0Jsni+1UzIhYrSSNqHmgeAAv7qdXIIrtNIhLsKAj4ByV
twNA6sdHp4HfWLp8rwEirp6aQJ2FJm2Qa2MFkNzkAaQ0dexPP5yNaxp0TYe23Gxq7yqCdxXZMxXC
di4uc9D1JD4GYABathgNtbWXzDzl7p78osC44CvpUlo2XHvHQw+6l/TRR6nkRK1s1CehAfwnXRvs
tfyD1WG7dxKBzm4y4oDUBDyg/rVm8nXkwuS8yxCGyW8oAsexpWfMepUx8SU4fYcU0wHnds9tymvb
gj72w22AQ2rJSwEz/CkVO0E/ymmi/QjIYF+4blZpV0T7/gAN7qaBIqiVtYaFRj+uR/stasAF8rUb
H7vZf1qUXOahNNGH2fkxW/Sm2YwwncBmz8adeAYqaQcZcdpxTxiPEKk9i+S+f4twXBqEqkkZrguy
d4RqeH7o6mskdSO5ROO/FXHrXs2eSipgz8znCD4J9i8EukYsxl5d8wLPwZXg3p/BnZuM2PwL1o0E
ACmDbBpyetyN0H0BWjQD4LD7sVFWP1Qtr2VHIe6khaNG6Sc27dhsfEd+QQM49FTsSLW4e5RNwGYo
OB5zKmzoDMXcNIBwCzM3S/p0XozjS22WWrSLEWwMVz4rSGGH1IA8nt4B/aO1lo71d49EBW/krhHq
mrjWBJo1Sf7ZD9YYfHHlTs9umpJXcAqcGoWtg6KWqTgfFvcyrtvRfky/RlHv8+hDgL4cJ2Gt8S2P
Tp1CkBFFh29/3Dm6YsJ++GEH48U7NWTr8w8EBDfys9rZxD2u9x85pUvD4nykTpwG0mTBrY6WbDtW
Lp01U73ZewwwaKlA120Q/J3pCrJzhsxuS6wtstG3WX/w7x3Fcou3ELXukCoafFa2qrLtUwfAVmmD
lpaql6ENvbA37PXHfh09ia2vlzivlUk3fMbfU2pD6kepgaV4QA5jRZvPUd0aYjirNa2dWLQRVkhC
KLzAuKsQ/C0x9zqyz3jzXPqc/wssu5tX8P6cAzBOwJwCGM4RaC/aF6gy/TRgwJHD9dNDg35mUk1T
UMOr4/lal5l/ATIdvEXoT95+2dNq46Y8vJxeWivcxItCvjbn0pPb0+yr4x1D8ikyRBVmEuflxqZg
/cDW4bB+74MmKvxnD5FdbhCgmDbRUedTKX8thj7W20G2rUv0kF4+GaKudGORRzWAVUMNULPPEMk5
ZfscqIaXdlHqt67pdW5/SmJXe4bP87ryUab26yfolSQljzRc6HTJ3O3RV1eO9OwN/3UcJqzB+6Ec
1L745J849l3ILJnI4y0uQJAHInfQ+5p03CyQfbK9cSY5ypVL4iZA2GCR0lRSosQJgSkTVW8crvoQ
yzCeiBKUWhx2G+6vMyUrvn8JdtXoCHAYoIXBz9P3m1lAyFYcWDwxLMusWGfCEnCTQC2wi0/o3nVR
OTP9iWn21yqyv/JgQP/FNKJvFLbkGNg9Jz8AvgjVP8a7/MLNmv27VMnsAVv7z9Fgu5Hrb50xj2H1
KnVf2ivJdVA8G73RSRpPZeHga07AYTXOgCugbiszEz9LV0DY1vhfPu3SyJqniRySl0nNMs/Ggd4H
LFqfygp7qd5QxP5gEyqU3/JVFObezDMxcpBPbzuJl6rAiaseirw3Ktv2/+cZ3irIoIEzaKhdjcWO
i7t7py/S8IUF5+AjVpj/Kf69gzB1cG7WFGfWjbud5iACptmczx1tt3tUaSMlH4dDOfBZSOhOhmSr
2LmzbLW/sjq2DGAV5HpYGNILRee7UkMrTC0D5k7eKvej5L4O61zLjoVr5MvpNPhR6xtqTZ21Syc/
6xp3nS/xOYwheabigsjSdtCJbLfFAppcFjqYsGFL3D1o6unskSSyFExpTcedyNPSVFmPvF0UnC2c
O13J2EqtBV44jzc535PVxpjJGMUZVhw8cNTf03janM5ck5fb7czWWHqlrr4ybCqzDb9X9cGjXl5p
JX8dSqCsVOVwitz1DK5Wm5hkdx+hXpT4jDUpxbMUgI1ADGELtPZFXMiTveFwRdCGp0pWNmUhbsGI
BvoZTU006b2anZSEET3yJ96vqDpTVySdcmLUVinAw9oxiT3RId9Xq+pwqVmRiB2PsD+UKhO1vLli
e5shdufUvXRCtUFILrx3Z8wtoNUSIFdW6Xr+UQBWptASFwT5Xw/HhWTaHKmnD7YJKIo3xTqX82Br
GyYfy5POENXgUz+1V4sIKNOx9zv2QWTTp3bozI9P16PWZsJAoriE9N9z28ZLvglmEOY3+jt/rxov
p1GrHnD/88RY12d7K/BtPcLJnsHDXfU+DgrMU0axNmmS8tJSFH2YPudgKqVdXI+AfBAcPoq7gVsa
CG4oQlxDrTcT95bQxMF1cEZ970f7678FyA10yfj9Bu/AQGJfIsy+IHUVaRu+bpSUz0v0sWLjI/rm
XrJmNM6AsKBqaZG/zD2w0qgSzh+tbXZMuoeQW6Y0AhDWXVP+DajWgvP54+GvA+f18O6nzcZBr7Jr
OnVpZvI6Sudqbhq5se3xonbtgahipyyhlzjh8Crv/9Dzvk0tLVMdKlvEm2rnQDH3GJkPOTLyMeat
ty2OowrHLKKpH2/MKs7p1Bqj6fhdZUdWSGS2fmnAXVqVI4cJWjkhw4tS9rPkTQOuOhMQD2h0CXCn
79fRiiX9wJ5QSj04EHFJmAHBSt3UTWihKi/WhqD9ICjeExaQy7JZYhPCjwsYnhPngwx5qtFx7j7m
UnVEzkXWLBLOd+SMyPVEnMImtvh2WF1IXe4SkHDMs+VzUVKLjiSNQxAaDLu9jnqP1jQGQUn6CdHl
n203jmpABbC3Q1TtWgEMHf9HOgpB0G7dn0vvPvzDXUBV0vbJWmSLi20mzAYBNdSkeVI9Cpa7Fx8q
iqR1cuSEQ3jy6ttEbQ2C4oQp0xihAgS/sg0eyEXYKkuO8pJDjYGTt1s3EWE1dmz4MnAYVIwoGCqs
gpVucKf52jlABibi5JEteeVJHBYHVgVVwZn1+vsGxORC/i+CLof4sQNXA6SUDsF4SFFSkpwWbFVG
KoWZlv3Vh9ROtjiYLt5Wf2aUgidsvJWLNYZnafFN6s1rAkjw/ktgGYWZgnr4okAxfiqGLwXtEGoF
Hp/WE7bjPWAG08qBNuTb5xCbqmrWQUWV6lBahv80AtCF0tOE/sso/20p5N2OboqnDzAL+inrd5IL
xOKj6+qT+3/fo7TTIDOqoAO/PLXvg/szWFptqzj4hG05LmEgYP+RNRVGhecBlSF+1h9HVFWFXVln
p0sKydhK+C2dSEyKj8fIDCrXBFZRLyYnZAdkcUqofPZN8Cm61hh9wJjQy3nNWkdPfPAuIK7YC/1x
kqv7UWszb21rW2vFQIa3P9Qa7xG/CHxUlim25BuojEKZ8X8rY/NVcLCFRjkgHYCIiNJk+6pCAVlI
TV4TxSUmBNL8vR0z4HeC7sr50tsoH62sGL4sae3N/cznXed5Jcrc2ADIaavAHDinoFBIjxzthZx2
9EKzA1UPQpf33m5G2+Wflxet33Cg6jrDmAvozq4x2TB9raDwsHtkpjL9HMPChcVM8ydn2t4Bdz9a
ZrT9Ab3B4Q9VUfDoC0DvDInhdroUMRPRQMuz5c4c5e1risywF+M1y9Fjo436NNafygi7GSst6RYJ
UCVLAXPxpSEBbp7YyZK2cz+ouiD92KqShLs5Xu5/sK16qOM8W9VUQu47q06G4zaz4Ktyp3d5/FwP
FeRc0XN1KRarGrFUsQ2iYb6XDLtIwljZOWLdLT3adGPn1HA/8vy64NmrNkgcfSkhkTkNwELxRZza
uq1rpmh5Kt+RScdOpQM39YBVeu2pWHaOYkWQXzyQq+L+aioYlzd5w9YDtlP2w+WQZIHmyvGyEUFB
7AL2m6/uuUVFm1Pzblrnge7wEfwyWmbl97DiCmY6mL5rrah6KHAOllinYPvfmgxXwnxAQ4piVaMm
BUwQsxgqIV+5oHSde350BfcNP9OTISvOPEj+XRh/7+oCWCEazgfDq+qayE5CBQJIiyql/omIzba5
1RWu2VhmTOD/nHNcUvxzH8cgJ+LqYc03jzw8Jnl0kv6rzY4tBkeD4THE2TrZEhEP5um7YmAmEYCN
4aqS29Tz3aXn3ZIEhODnLU96qmRoob5qne4gyGbRyu57uVCI7ESgYTMF3y5x2LrwDWfLaCdbuV5o
TQu9+pQ2MTg32FB1pqNWlkqPG329642QIrKARK4cyFs6TQhchCFeuiCxS7m3Rg6eNAw5P5t6NxOb
sGfUjMxPQdQMFumXHBCpsQetPJvbh76Agqitv1DinkPkrIwoaUZvOwL+s8DBotbM3EJzELte9otn
m+rir4ndkh0SBgd53u/gflrCbagL7mnui5z8smoL4C5arOhPiyrY9vjTO8fLv3saSs2Kdh42nJAD
45oP/SVDa7LjjXx8zPjqVKnGyEWRGSfxEHAuCQhh2XMOnzkBFkhgS7g6ciauQf3Y3I7JIOU6En/l
0WXSucTajvbB4xzW89c7xyLoUF4oHA/nPTKGd0QgqaYbCyNPktsE9odcqOIWCG0J9WbGEVrWn3Aq
iH9SKZ4hsh7B+8Giz2mPfKmpA8bPw4hUHcLI93cPu81mHeDj1kf3gFUgO0uotpkOmJNIoMqOG6aX
763VdvFKhk5vRDTN2rp+MJvXDbaOjQ0yMZhR9oyG4bQ+tFXB2JwKacEB991zq/IlleoKquP6vgMn
1h+uLlYXP2Wthw6j2W97Ybn4h2FDgenlEb9ajOKtqPbSO5XSFvOi+ZWf/aKZU2C6wldgcVlYnWBn
2B7yx6EY+PNp4AIgiV3jMXGrc69czh3NrhKww9zKuSmIEtjM3gZ2u90f97v153U+hAhWom8B0/b0
/LcwWwdWHX2BVvGi4BYtCg79WOEWAKc8A8wK21VH8aKzuLwmvxbAkbLtfJhrtng/9Mp6Yqzs+gqZ
UEoyNFI/aclb7HO9zNoGjzmEDt4eTX/qbQXkRPZRFupRmnBIHFNoUOyt20ofY+XRD9Ld6aGyuh9+
uR/82EGdai05djRGTfTphdGxbN5nhpirnAe8pyUv7JY3XRPJMXwZ8WSy1HpEf/wmL3tIFbx45zPO
b5/H3MjwlD26/wMmzbcgY6B4RWL0uQkcZOnOwlZMTXMOcde2IvYwRmKsnvGRqLfbpfrDXvxWnZC9
X4vmWN61PXjiaOs4JhDZYpzfDpNF8BdW8zzwkgqPF3LHy4POKsF9y31xBTUV4XZMch7lIjVLoP7e
XMSp4Wmh0B7raexc6PsetrB+uYUQNR51To2vBTeeQyjtHV25+nq3d/QpOYWxRICOd4ByKzI6v8tV
C+vBL7OzsANCSXfmRSZC3uJK0oFr95uL4LXWlMaqdu5FLoWfBJe8XFnq0BY583IBnFSbWidlDt22
6GM1EORBvTuKJVLM7FFUTE0BT+qhg4BV7F2Rz3M+u+V0o6JbEVxjxJnyvhJxEvvI5ciwDG4HnvjO
fqjatlfu9fWPrZispJl0mgjNCcc58ZRG/swbtl3gqwfU13DPnhqcESJAXoaRHSfI0ypFJzVMhC7a
Y3tL0ZDn1Im6qW40fmb0nJRPUPV/pIBOKtGCEOolvUls/7W5BVnYbDxojHozwlDxZkeW/d7WrHkp
0BrZi5fFSaWclMCS2XoWd229X+Au2EVI4uLd5zijBnZ62gpENgG+xtbRgu9aJ/vQhMsV+l/8nR/x
xBF1QyUviTRFE2EErv/TnyIj/e/caxOIpwjjXQsgUDkjxVz/eS7xlDZHfH0Irh8M4x8xT2gNXBn0
ieUVWKMugnb7TOUCLEVA28WMKAgLF6mDxjE6WWJ/IktdpblHA6a0p2xUfLgelIQtdeOvhAdJFo0/
shw9TxFxyHOsgvCPSWKgBOS5/tNmZrTZwXdZKAETRyJJVvmzB12yymplUf5+xT1xLht8qubdJu8t
QqlB3SaOwbxqxOu54OtQ5TXVXyblrSV4cq144gRXdszCUQzK6RN6HWT6ZvXnOsLmrYe901227DLj
Q2ZrHPg8GJePqsnt051OYphENJ2d80rt7aLNj1kg/XpkRvF0jBv/oNmjTqMyLoryXyp+CadmwSXU
05oyFIG/2fyfQtgb/3jjNEwDsFhIcokqmMZEeW7IRFuv3Wt9snKS/Ym7aqHYeaqBKAG8xY+EXLvc
QtvKJHzw+qt8IJIsVT1T3rt/xrMbMeYWzfPoog37rAo/L+HPv8x0yrO2wn+rHpPpbVf6xL+STwMZ
p9ttcUNbZ/VYYCKsV+Z6Y8jVXfx8Dr72EcfdWYziK2RDxqYZyuB11uTR9TDihelOsGhmu0eRhO8A
JariIRSGTtQEjPpIb+gPi/+hcaIXWkDPycXdzeh/pwEYK3jEmuuH1tfF/bm5soK/3AdAyk2MwUMp
FO3uRsLg0lmyrqN+mazsGtDlnSL6Ts/Ro0tzJPAzS87CXwVGEYKM5w+j/CAlpWWXvhvhmvHRKucx
FFYPVPMdEsgKN9o9Ecwpp2sl9/q2wHEV4Zno9qdYddf2PrzMjwSm/zk2E0xKkCfmCewBK3G89IBO
VFThumTJQBDkE78ASMRI1F7dF2joPdLdGhu0ZQvBaTuVSpGtLuLu5Xm3DQWvSDrFMhVKQGSz9N2q
g1s7hUv9xbD9pPM9h/TqrpnNqSjZfr6Ob7xkh/I5eScU7YFdI6UW8O+FLWKB4V/jE0Q09fABntOR
/8YrXyWtBzWv9fD4EezBoezubYcdXWmKc/EsVJrd4duOJ99UWGsyvaXyPricdNGDa90QanfF9lCB
Gk4OtzgTtDNVQnyPj5YGp6uw6c9ay4OUt23ZTEoToxLlSqXK7Zm4s/0KyOZsdPLhaOqnHTUyehk+
yJrNR3+BHXI4Ox09eGhE6geCwvzWf/LftIYH4AzJKDk69sU7kImMwlUa9NQQjSpVcFaBD1YNpTvp
/AaP4hisSC5ziRECA4N11EPxkPr2h6HzmOg4bX1z8VQ/LDmYPhALTYSDoLE+yuhnJFLzNzN6+RlQ
oUy7jz0z+/gVDYmVw1ziqqEeavhifrpicJYXXwy+GKGeJKNFgjTzQtSZPJ6Dx71SI5t/FGQ5w5b+
UWFZv19g0KENn9/P6q55Qn6bIU9ioY5Y7XFkB9q8D5PoPEFuiyUEMk8vHgHsi3eFyQmUvEmGwwDL
B8Pziowyas6WnrCCFNRC1CfEY8wAGiZgtCceZGC6Pn5dxdqWevIwibj6fwk15IfU3JVSun+TjkZw
Z4df/K/EblPKeTC5ovZv8L5aAF08AW1g8vadoqaBOSKerPIuK+vudWbQUGxIq4io159/oarqBAJb
nMLqiwc+Qyt1g61Wl+qBDz1XM1KicPLI6itWsUB8SoTeG4xISuFcL3bZwY0bTMq1FQfK8PBPgtW9
zjqTfjkVO5ky6jqWmUEbz2PS3eRwC3by5KDnmrFYKBQOsIYFHPtEMu+HzweKJasImgkvRxLbU+91
M+BTrZdY1ZhsI2Ci/sS7RmelKXAInn57cqzLkkn9Yyr+TSPjqlvXx0RF5T9DLNn69C/goi9A9Ctu
yiiOgf2LvzD9nlgvbYhaAxafwFrKVWNr+licrBFN6A9MjnFUKdxuL3gu1Cx8GwjnC4Njk3Z+Pb01
B66S+WKCS+VOztUbnhqWM63je0H2mt/spwvrk7HuNYpFjuHWl8vjx4vFD2vHJ+GeFHGv2a4g33FQ
vshZPIHbjRjFDBYkfYdGT6k7cRkqEW9NGTgA4fwVDD/HMpXl4FMRSqPi4Yn2LIXsi+E/iZZLWIz+
KoER3p8+IBN9yEy8EPLYoMpf1cgesN6FmoJMXm/fsf7ZDOsaKaa6IEgekPnnWWobS8eqjfAIhLhI
UHcKz1fG63cmsekCK+p8IVrPeR4pUK+iDe2gai7o7Yonyvxk0clUHDcGmVDRWCfqQ3AYncTd2HLV
D++OFNy/lkduxPgHlhHetBV6IxmDB8X+S6smqpemhG3i1+E2mZM5m/AIo7IBZCm4pqh97OH16lXh
FwAJYLkHW7Mz/GfpGk2W6IaDDXceP7eXJ/o562nC3LR3GhQSL1cmx6QP1ZfsNiBNyOJzFZyATWpx
uRnT3F6ojnaMunHXJM7cOSR39NMmi1j82Fz4k9ST48HfA10YzGLIGVzY1VaUnr34yZPSjgwrZ6AA
2PDkmDUfO3XTQoYQyqLEqP0RJLdR/9P+QVqKguOfqmJAGAiUzQPDmLeehIsb21w/TR/3NeQAHOLI
kwZjPdcoP37l45RdRMulXn471YLCM1zsndY5j4/oz+GWHOQNWtpo6rQKUJ79d1etSrshJwjkFiIM
+J90Z3ZH8uFTDAgHKdRSyxSqU0QdDTujIPSkVD9nsx2upbHOrxGY6ZUhKZS0JEtpd92Z8WbJxOHm
/TeV9mPgBSjhdbS4RbPgp2lg43kDkpIdHAJ2CPwtvDwI8z5R0t5DNYaI1RM3maUUrjHBiVGy4iMu
5nD/K35jwuIIIm/EPtVb8Ewui9O/TXPk77WxpetzX0LgL2r+qm9cJNyid4tJJ0wI0MwoTJKKYmRw
bmNG7ZbPzNuxNirpjuPE5M4w+7yU+E9XcVNBUSFu5KJ6c+43P7Lv0FjG0GM5FLus0JrdtnupUTrW
OC5cGGUJMJT5nYv2qSztYpakuM07Ff3W3SmmMn3uRJz9Nr4UG7j27YTnXeEBx43d5iNSB+MtjS9Y
6EFTC9gMNJOOlBARq5+qlziDvizpChdEeOWBCvCoanoDVqBHjkwQt6KR/7XkspGfRQy9AFSStso7
O7f3buldrKbePi/2JrrAEGR3UTuw2x5VT0SnZdH+YfkyYM2DoA7ZkFRdf+43VR+w7ie5zIE+qC/2
Py+tBbX+ZSoYKCADBGWPQTOv4E2Ez8JWAM6xI6oP/Wf2i+do/Msbr/d1EhIs4pVXAkBnC7muN080
+JVLwxIgfnTYKuOgNE64I4s7zWcex0FCe2NVuwKsw+XrqzCodc8iUtH+mCqKT8LxvA+2whekW+lG
ujyjjk149bFC8qRVfQnl7aikemY8QkHTTsJM3/n9VmlG8gmGUvDN/Y77HxVg9cTTtI0AIHFCo7DY
GxT0hfLjC0911raw1F10QyeqWrKB4KZ3vvjkNyzb0GpEHe1D1p9W2DahK/cknJZkeY5RPvHIfqJP
HysZUxcnDo2ngm8odzPk4dN2SFzGJMxUsAqmiY7sWnxqK/TDqZ62vTaV1WqQCkxcp2YYBWoV2l7S
M7k0wLX+H+dKY2pq9kkSwQ93zSTvUcPCD5r1TnZIFet81KqkmlUVehTzyTTiyniM4TCc94l8M7X3
HXNiDEsy3H2wz137NECQfss3CFz7BoqdQ2jOsWLntWTnHnIGG+KKu/HWcUTzvAovNghRf5I2eAg+
8MVpSh2HE7CK2gKuSYDpbDXbk5IiB52Gf81IHhFGB5Sh79ekDrKtF4C8dmQn4ZXQarZxBh+LqYJa
QCTLAHwB76uCV4HZnIlapQG4GHlgOyUWq/n053ceOEM7mipl1QccT8hQw6UjGQGC74DiPtEkq8JN
ZBSZrRKBSf2wz9gAHCZEn0u7CMsIxz+KCGHlEqQCbMCyJVEqpBh4uMIp5KujlJs78vgQBxQ6I2TQ
zxBTBTjH/CvwhXuF+BX2pyaBdkZoKfov2FlmdkmYWrc+UthKY7x51WvMwBSpkwoSrgt1Ug51tCpu
7LGhuOZxiMK5+gdEkIrRLTqdLKvN7WDMphhJ3Oby8PJjkMUxKof8n0Q7Yl8AVvCE7TNrQBikYvBr
/bkgpltSl0z7yhJolLnwVsxJsHxyxwmyG3eeK0wHoNGbSTtlX1YZPYp0GDr7/Gn/0TFFv9TYojb+
m5tc7ha/7fxK2shuxmXwKMKeEZd0uBQ3Rzm7UgT4+VcsRYEAjUAP367/ZVE0xzYOjUSwkS8SBHma
hqVBPNobQEbPU4VaO0wTCP88qDn0gXJ81fdDJD3kYhMUXxOmKHcfGBxSlXSeOHBc6uwY9yP56Zeq
INw5R8ZyqP9fWxHGg3J2orfCc/mtzKG04g1nnnOxj4OIMuubiqIB0rRg1BdAdlIqKi4eEBoE6Tl9
7SFORyydygxwfq7Lr8rBK2HC4/WoN2T+8l8EXsQWUF9mcDoWZiR3/R4LuSzkDcc/3Uh7YS+YY+H/
pgjSzuIApfbtrpIyOKzW74MzYE+fXLIu11MaAWSmflKjFxYHQtpr5yNJdeT/XU5JE66eAEOxAYEd
BK6/X3XnjxpCEfGtH4tj5pX0PCy02xLt6+RN+Ks0wRN1mLFpJSWl22acVeKsn+Xyiv1ijEMG20Im
FHLJGZ0kwGzmg2aJ8kNa0hdzMxDK8bRXmWFoHuDtwuKkQyM3ACcxARngjpf5V8f84VazmfWrXF58
wdr+bSdCEbHeyjFDj6SiiKA6vlcfOTN4krM+c3nNdSha28jlZBMESTgui+IOedh4urYE0KZYfpz6
jbrfBZKRG42ZZMifYeDLuvu2yNeFEJ18tBC33yDdLCQcryxxdJVYmCv8paNS9g3ecHxEc8uzbIsh
Y9Ir5WqwM1WePNXzBVYOk9BiXGsbcLNKJG7NyeI7sZxtFhP4V1VyfvMMwLDL0XDflvkVSpL0lJej
VL2DwR8N2wdfTqPefx3f3x8Y3qZLUMYOhVZ1fWRtLYtPq/w+7ilbhkt2LVQECcbSVXzwU0GZ6tRr
0Ss41PjU+e6AQQxb03jp1WVhdyBnz3sfaFELDtZJJ51sR+XE5S02lJ6gI3onJsTqMbnGQAvEyAsk
gJQ9KaecSo8Ny+xnyyjCBrVZ9cANBd88tlUTSkWSg/QMw7GSkpeGr2xzZ6p8/JWwr/NOKK1DkMBq
GPM5trHz3LP5Afu4RsJ+QtOseyCyO6jX+NGJXfQV4Rv0GqwcumZd7ZrSWba31DbolHHJrnyCk5nW
r3k7WfAyq4fEr4wv68GLYxan11eVWw/U9rYeuTlWE4MQTLdP59o8B35EQk02VYqyrAlA/JgAaw1g
5P8F/MQnkMhXbmsxaml7ybNEH5LOOd3k7NtuHM4bDhCzvCLf00hBIZmoQ5tBQpggGqkfqe5nhykT
dtgMqLBiuA+ijgCsL06aG1DFzple3CxBknvA26upquyCJXJp9/cN13co7RYgeqciKAOAvaYdHnrf
1c8UrE6XWA9wOa6TIL/R4xrVxS3S0hswGOxmbdv9oMGVdBfoI6gAwr6q4bfNIMlWZy0sVJp3Bha9
qDAs3NNqTEbEWcg0LZk8qgrnfFnkTvdgcZjmTvkC+nb71NsDKl0W89QP5SWFS9I3Hi6UjNsZmcBF
Y1zX/NccjiwZiftgjtOeAmzNt+Nqm6ehdZYbPmygQ8/zC3bYGxQR3LNiIqWAtO9ZE0U1VEHOBS/c
m+tB0cR0MEk8Y/NL00cGIndSVak0FfuyA1IOVIgr5T9MGGrKUyl6f8OE9LYMGgF53hCXQEjPZPAA
LojRNiv8oIbWTKmYDIj+Trlp5EeP7OYVljJWJqU6kodrVUbJwEvQ+FwJCSCuGMSfdZ66mbeLOjIY
FEsTLTZhSuk7xTcJCcipI9qlpR43j9eEWAmv9QVBvVVKULKXVxJpnVUtcf2Kk1Jf4L0YunHMs0E3
CjLxArtKXqyPiHRdF4yK+FUqeF3IU4nK+hw6nZUZZrgfaqRqT2XGbZLTJKo05JlNfTyaAzwBdpyn
gORYAtBEngkE3puyNfIqEo60M0s5WoDXn2I8MHgNs9tZliiwLkNnb92hRzKnGFe3L3akvHwxpf0T
0dzhYR0sHSfwAkCMC82jqbteO4Br4ru680y1vUdzEHyA+cEGZ6aUUYny2MLzv7VCHsYGmx/isnVW
F1zHpEvuWgTp4KtXtGzjGPJGEA23adzEsTmi0aa9OT2QRnbP1oeBlETfZiHfIWpnobjPpGw9tsoi
IAiOb7FBlm6q7PaNou4ohqcsDcZbuDBooVBeq0qKV+NQ5Yha6ay2YCEu9ok7BenZSBuOdC8U5q5z
4P9ZKYF5kbe2e3/tR5DPKK9fnYtvzn5j4jjsuIpS/rstJydyut7fBs/z8kUijCnUM0/QaQy2OhXL
BBJHw6nFBLgbYkCJ6RNsc5O8AwS2rAz+kFtYNfZMtkgkbCCwTEVX/45R8mtBTCz1WkJOyVpRhKfd
VqUperFfwRtp2G6eSygviHhmRSTID0jHA2XY9T5/puh9Umg92KpEvRquGV8UFBoVUT4k1tinKsMV
pF23Yl5F1cMATxlcoHAErLibrNYKgb6gbehQxzI0lBhoWHi+amEcFsN4Ng4Ukzem25MeRvKGinJY
UaNxTELbBCe3gC8FhE5aZHHkq1B3hqVMaNbzY7S260yU+IdF3mMVFAz55bnn9DSWjRL/kKARLO5p
GBD48pthM59AJBgD/p28l5rRZNxFjCz8PfJxoRJou001cGrjsp+l5sT1c5cf3sjT8bY4eX+Pco8x
Tk12WQmp0ELKEyM/nD9CZsNbMcSHTe/sfNMBO3aNuqHT9M9pc8S2k1+rC4rScHRsx5NIbQZl8ocI
KhS3VyVBXLn56JQCHcCs71vN9L9GlRS0ERpMQBJJ9T5ewspQWp+GLPYgDxrWjLNH6E0fYhOYM84p
bUXN/ou0ZZj2orMiUimr9+bvhg+uYLQyBIxBze3IQ6W/G0NrQJPNRP6HcSkW3mgUncXgFLFFPp2h
eK16THJKEfKD4dE4Pg302nvY5hBGquPSCFVQH1aQ/4a+Po3sWrr3fpGuRJAipruAaytp06lCtoaq
Z9oR2jOTXbwlQYf1d6AT2oWcgReqFrFnP7ZzKDSdqff71T2U4pp4VP4JzlkwpoUeyrD/3l7y3rLb
xWFBaXZG0Rs6w2haWOKW/IAhaedIzRrwL5QA7y10BW2Hq3HXLNYofcE+KCdWL8W48B9kKRjBR0um
a+pYMb36aHH11zdWYFN+h2sTwgDg9/NFszLqv0+YqIyfUw3fOMG/Kb+6Ode8dZXBkKYWDv90reEn
gocD6guQRxKZ9tqmhP8KpimDWAdAI7tHo1Vh3ouc01gpErKxsU8yv6EhDCJ4T9GRDw6hhiRVXqSR
sW323m/lF3s0RK1oUERE/+7hqNHPu0EmpUsaZbDMTho3LFyiM6+iENK+OlO8IkuQ+adFBNk/ApLm
gfn4a9QdDZyUp1/aIQUrvxLksm3FChIrPUhAl6bg8unV1PC9A785Wx9tENP8kGiXvmvtM//Lxb/5
uw714Sc0p7K4phXZXr8FVShCJxTH98LufgxfMSbG8HhQYM2oA/yOlWWROmLVbLJUxjGJ+3gP0VT/
3dKpxiUXoFAuC+avhTgyyAmAPwSSxkADSarYc48cbw8/hr556COcQueEMSBb4faE9xYZYj7oBp0C
kIqXnsqVMhCfKR8byATYdPp++8hxm/mzxXBCZIwtCYIT2vlzVEhRKQZe/gj+LGdsbM+jsXeLELq/
/GAc3wui+ia40a5lJE6hfzaIaUoVagOoQ0qnvrX5+PSm7BrdswiOb8+T+x9mVAMYxpCg3HETdpoh
O+eWc6Fr3VqyFiECEpe0L5ri9fDm3QUgKyvU5Z6hOSnwbPXaxl+DxOuBOvCjagxGYkF4JPsXblPm
Fckbm/5cI2YN7HJg4E11jktVisB0ox6+uf3WmuHuNW3angUTloJKSjTgRuDFoTnSnRftu5VZw7HS
kU+bmtlbLIPr30mPojFwiCnuhwc08wHdNtBcGm56OGo50njlqIkOjdkxlrVKxqEDPV2Kslyl8974
6HrnthqHmjh9eP9zMxgnZd3LAvQQLMGtPnLvXRxxyVxzR8HUDg5YmApCFUVlX1S+p74DFplwlPug
hfgoXw0HsPpN1mmgYZG9UvtjsxBjbT6W06e+Q1rpI7OdvAzZcWMgkVwM0IPibQh7bBAFt/ZruPH4
D0ZABYzcxqprwU5NyMlLfugeZ51Ohy7Q3GjZTTLLxVIJwdB9bfprs6+LZjOnN5NdQkKzwF4ISibX
Kz7mX2tU9KSmO6XtrHax5e8/TqAtmF/1D9mwoWpvgGBkB8V7jxSIrq3Slx8jw937IBZLhr2XbLP9
XuiGWb88ZqWyyApTdd02o8AbVzvZz+sFzo6Gbmywx6iPwQQ3OBaH6GtWXkhj0vDNluGfq9HfsTVO
CN7nEn6oXhX3vJ0f5m+ctmKVGjCTRT98JZlDumWJO3P8hucBguPp8ayLeNUkwzUPJA3IDIdU+Ptu
ohHXsUZn65befY9htbgD4KozVE6hM0zU01KDCsWv8xPKPxVguxyIY79GDUBflAxoY+CeP+0b0Kh2
bO/35cb6A74K8rfZgavw7YSEIjbEmK/iIwRGaj3IEbwe/rYfVMtzdEjvxzIpBExV/IJQFcaHMzY1
OXFJ5ZQdRAurdOnp9XqmSjd/LDryqRsrzRs9GsonRSyaxbKNCQhJzuebXHY37O2pxNX65t0/H1Ok
Lr17pHQNDu3z/FmeVVjkSdEmu8LGiKeP6BRzlVk8kmNB1ay8L2yCQvrQ5/p87MBsx+vP3dLvPKca
7ikVqgV5pvSgfyhwTXcROtib3BLQPrJDctawH30fjJnCL7Xjss7JdsH9QXQ42makuLH0T/4qb237
VmO9I4GizNmfQjZC9MZs9mI/c4tpwObbuEAFGftMw0RBM03tN8+cJ4PPF4WVlQpiVb2xYuWxAjgl
kotjvaROdwqJ8Vb0gUKyH5RaUnY4K6xTTYT0pJrX/pktmMdfODuOA1xofDcl/aG9TYS+jmwAA9e/
243tABzqDHAZoH8ltywRyf7BEZivVRVzT2yEBUhi+zF6Om2hh5M5sFaFF2k/SNEgMYgggkvkrD8o
f0uPkJiz17+vFdbVwDiRwwTkHwczDbq5uuREluT+EHkoiGD6E0DeROkTi81tpCbKCNewHpgg+DMZ
vtOsKRfp4nUNpP6xHC4u4O0N74C6IGl3e0aaw8D+w/NreVSSPirx06Bz06AfPy3cI7I1oZkv8BMu
9pFGnns1TzBTRwvvpBTiQVhDxyofR3Hq/WXT1Wge5xp24QAFGrlsWyTyKEXLeAEutJzkHyCVGlZL
avjf58WiIO7jvQ9QhhsJus5hnN41XqlgOnpwoba3lyyC4bgYwiooysdyJZhsIvB4+JUkZ3jBZipW
9qOSpjzGv3miDSRQmShKzVu9XR354noNoX46XNeLImPAZKgdanQLlNd53WJc9EYlefSqGMIR+M+R
M6wudrJsUQeZhEopYEh2Vo8po/eQrjFOg1X+mkdwT+XVXbUN/sKBmeqADJZ+wcaEgFJG0qkQtYU2
LoakC1ixP7xbLUpIu+9fih0BcxTysd/tOBoHMnaf5O1TNs1vDDNzy9PwvanQZrzOq2DGrXCfB2Rp
yT5jShn6NX+ia5CxAVVwk4KNB87MX19+CrkacE0cAQ2BcmKIukWxtm7VdFOtDgVbZuUg5FtWWWcC
h3pSoFA4EUY+g6+dYh46jb+28GwIgr1FQ7sqRmJEGRJ43Od0kNmkXCRAG9a6eQhf++IXrDFE1bLX
dSvWIC+xx+C4JWR0/hxzjjtYvG0X5sk/fsGe3cOCMheJkAt1B3wIFidTMOCIXbVsj6Qx27E7Oyl4
eDMOgZkkJbrw2WSew0WFwOqYUsxiKyopQU+T3EILQ9W+6kW2ZaCPOeQQ356jWg8g2g0RrFlnq7f0
q0MQ/alJujvrFH9G6PmRyYci+4OBnrjrqc4AMs5Syq4DDsbC1pJVQs4NX4XnKiNPi6LbxGhCBUBO
uNvzLpeQ7FxTOM8vLLRyPKbTdTeIQ6H8o0N/TSHktLB5IEnkeQuwatyRq2kZVJj5Yrjp78w87iTn
t1riU3wgfglpaK7FD/c+nV8uzrzzwPxTt4dg/ORzC7zNNXr7DeCclyFwnNliKaLe+vewfRuGDfMQ
hyIz7rxJHoHtA9QjRC9inNAcWxLiAD11EnloLGo4IH4vthv9mteJqG4/xk505Tv2jRDRoahj5iEl
VixJz2NXp/SdTBHvU+jeytO7Yb9T8yA7eDDRVxPWxP9fcCC6f0iVMgB0Pqvfj3Xu7nGnBunIYBXC
RCpvJZLnyWumMHCbP51qM2CaKvIVp2qevcppISGkXI64VmfVPdGSjxg/tzZJMKtNdr+rZmh5JwX9
ftHV5pYzME1W0wyzJdzoucphJNqeffp5EkHN2m1nBnf8V8KNgJYlndLgciquYrJ1Yo/Otq1YNvz9
nmNmvO2+vIXWD324q7KnfdEAO95sV0UOwJ0MyKCkAZGx32EhYdV7DodoWheuAKOMEZ63K1BK3hki
Sa5Mmz6K6pfItyqptcBc4njOwye/gl/kAmpVTnJsB/hx0nehH71wLGc3GRUpDGN7VMYRv8B39zzA
HKeT09oOOaA6Ip5f2qUKYp6cEsKUknc8SqDNyKp/5YqdFCT22j9u5y1E8acohikJVqJ2KV+ngwAR
aor9f9ARxTJcTmVxeTWsc4qG7IgQxTTh6mX5vFgST3MRZO0wnht9hfvmlqMoGPQilRmmyI0sKpdH
8Csr8cIFCeNGT0hpSVT4hfOTWI+xD5dXRKbM+YOnc+vKwPEc4ZG7NPYrjGPYy6D7pSM8q3fpEV2C
Gspv13tlyiCeLdOShWNC+5kk+jbV7fwh3Av5+L5iw2WejXS7nkXUCQpqHGyqgRw3AzxdAIFVjI/F
u8dNgIfT+jBnM5cMxSmkoR3/gJ/nV2U029JTpwSTTcMyJz9UGwgmexhveK654JtV7QJCgk8T/a10
IxnYDwsVhsEAt23FfWGLOxffR1TilmeDV/k8EAMKh4MOjE+rpp0SYGNkDZkKtnhCVwjyPMkbQghT
ZaV1qaRjJ/Rgwq91veAbvYFo02U0Nn8pvmNowgWhBG5m+JTgcbG09lFYxyiKF+f4hsG+S0CQdFXI
wczSBngNxKOSGkXIcskFEbtoFASzRuc6f5rg1rMGoG2LCijU5FNK0t50ViQPQ67lPKuL2eY6POes
UnMPfUfLqydDQ5yPVXv5dKbwFvmUX21OEJ/QMxaFBU5OwFqIisNIF6dGM0wThRuGSAR25HMSGyfi
PFkYIKUdv0zjnOlHpHirkfli+HlzlG+d7XmkBVcU2HOoYbxACin4CgH4XDz/4LLSg3Xb6OD8mD4Z
01mJF9yGutqgPzKpK2fa8Ctox5eOoPIuiNEkDIDE6ER1pvxWXMEHaZk1H4wlXlNtUW/h9eHH5Z+a
xdt1MEvew7BtYOqshKU9EHP9xuzgdoKpV0EBRzcEwpf6mHRawRO/VY354981KGCgAWobWQzV2pBS
awLPLGQLpADFmW8/0XH3pKmVJa7/ZKQqIIq294veKIqU7Je0BpddzbVNYGBfz6WGzxTwbmTB+9aj
rHbXqwAl5IBCKMU4iV14tcTwcQb6LK2PZElR5OYAn/AvjdKwyiurxtzLmHCLpdnWXZ6V6piQaoWs
FcnSq90qd4tQc9Af/ZjqpsAxTGL4BuUAqXd3rG2QmFHVmBMD+T2dzIJgZgG+piSEz5GiJOX4n/CG
pfJN65tJgYheHH7jRZXv1I66cVE2Ufej7YlDcp3f6h9wvp1xckSjxuU36SVZ9bNyv1pMtoPkEN9m
ibp7nI6aQynoP0nKWsV0bbhWloRzWUMsRnmzOPaq2MUhuGnCx3fgvuCgC29Y0cm/hDg6OmVZCU8o
KRlAMvxDrpWNUPxdAG5biKccOhjEuL/94yohCad6ZyzcSLuScp8L9+7LWFZBh61CerZHeHBS0f70
47LSSJyVmE6E+fuSP71gDGsFxLa+cT7ppqJIWzkPiLXaI3mukhoBqBFpkycwsf9KmU6lRuho1N2R
FNtFuzAXxnKKp/9hz1Vbjm/M2nGLIJ9gmgwXIbZqFmnl0/y+yM9UV4ivZ5+oZ7FZe2tvMTyXtm0k
RbQbvgd6WeZQxUiGd3qP0eALMYhcOnlrukouB/p+5V+WPomh6lc6rlSUAGb8EhzEFhuNQSavymLx
lEM7zUOo78RJOfGgzTdXq/J7xgN889vTsK8d2Kv+Tl7bBtb3LmZZFW9oWrX6Y4nFFYro95eT7DIY
0I/Zh/PZ120cIY/h/ujBf9JX2dIqtx9Zs/Dyns/mENP0CMgk4v466dECpQYz1bI9VZQA8nlXzkyH
RXhy0bXUYUDV1zggfRADxSEqhEJ1RVEAroOHx5PvHXp5TrysyBYea6xiZKaZtNIZL4DhJK0JUjX5
X4DHyxjnb5AXNc7YA2sVi3+4Eb+8DQzCawcH+x/nZ4qhUrwbhqfW5dwxWO8Lz/3SbeteIznFiqvB
u0e+tYJdlsSZOYSczif450NS9yJb2ckemSUrhyr6VtUUBZw6WbyLI4wU85q7cOT7DPahSPrYCN2N
gHFfdctWw4Txeuigb5L6pWbDjB/K1QDOS0pAMA4BcI8eiS1Uk+qAhCd0z/jqE5nx9swLNtcB+Oot
EcaY21JIdGfXQdMKwXR3LWEiVU07CqqT42bhjT1AVbSFJfytW5KEMAm3RTjM8y0WEYEscuFhlt65
UPrPliIKstPunkZ81SX0XURLFSKr7lr9PfNQgaqik8BpFmkN7ddSNcObDPuT03cPd+d3oQ764Gs6
cJ0SdV1AmTOF8Z+zkAsaY2GCbhFYpqHvph26+28U39r60Kow1+cFZTEgKY4eYoGlQVbRDXm/mzvy
Re2cqSIahigzjFlcxcUdYtG+OLDOWEKL7H9RtXmJGgim6lMQ+cKveyJVibxkkQAH7jQYHEpYpM8U
xC6Aeov/eKtz4j4RKf2y+IxfWOEufU5Za5qHNSOOc/XTSqmY2KaIT0A3AGOcgsjqHPmxRmhO3ype
U4ZRulIDoai3iN8Hls5a6BC0C1RMvrYNlXWrQ/VqFoq0daVjLrk9sIQz9WhZsEl56YHJr8e/MQPZ
0krYhbiEPEjQg533AAtqWCHAz6vW+3dRkczyob9IlMuY5JW91OWiKITAwSNtaYoEtPef1NEulcPF
GN8XR6iUoe+gfZenqi4kihCouC14KAdF4TL+BpPuVBegNvlTtTcL8P8qR89udW0oL9K8URLU644C
D+8kj8tuKshJZ81fkV6bxUKazNpuNY7zBViHKw2kLwUGCPVepXfcRi0/7QX/iy7dXml5zABxZbHE
0xXOTcCr6bKBM5f6Lln/ufR9GqAACS9oKmqw4DL3RjZV0nEzQKxJmoyHjaB0RLiYQz8oZ2FI/DFz
i0+Nh9RoDQKSdKFhozm0W3IDQcgNrsy816Hb+dB5urc6g0aQUUtwdIn5xc4giKMnfsZYIuFR5w4/
VvlvYXhEAxXQeRyTRNPLPJqKVvVGM9+5dHbEKwa3+/JrQvABmVnKyvLtBrHjq3puZCASq24iNx1N
LNeuz4BJ1SgAIoDBdZHLAnq9pPlQogp8pxvaqbSlvN11ILEcI7pzcZLtTXRdiNlJWCb6BMofigWm
EKwxjT3DJpnTU+uX842XMCeP3uk8WLNtTJ7UIxRxeofQ8zHwdfRJy3JaxJQ5XFi/QRjyFcb8eXMe
KNNrg9rc9axkDfkvG+JOtYzI01IVxPX83mU7ygqBOOyK6BjUYXOkjTnzybhdOYSPB666J0jqY9iM
HDQAkxuSGGYxxlikMHFibnjb7Rw+Kq4Q0Q3pcBxxIqamVwwp3yE0sR6kjZtvbDVi+cL2MDGa+RC3
B9PLOgl2xSOVPYEzR/Gry7vqMzZfZmaSUt+tNFTFH5X3hLNG8nh9bYjYZjG15xEbAhp7fU6wQsjA
E8OuwYmRT5tj00y/WCRmZTcEVo3bDttsjf+OeP8Xf4vo2co37J2rXzP/hfAkaqxgHhROJhUfAoI5
uWqzml56437GFb6tJnaY8gFW6DdnwL3Yq4KoNGBBBMYIMT56nLQspGmnY9f4ceio6yEh67f50f4K
HPq+tE8TYV3PSaJtY42+YaNc6N3Oiyolr78ly3ZQCJMToXPwgkdUrqpdzVvuennioyu5DrhuhV+v
kMrmUTu5SwTa8Ocrx0nOH7Dp8rAF5KWLyQC36caa3SfDh/nPHdwwk/T3zY6YHGZs3PYZMIrD89qY
NkTHX0gmkdpE3JnB50KzTyMR9BMbD5j2vhIQGbke7f0z3XZhMQp0HscmfbqrpgJ84AzZYNQqIzP9
oYuzhCUcUDBTNA/a2gGwrmfr0pcENAuMYiB0izcS+aBU6YA0SqmlYAKAEHhF75syTJadP4+/+tZv
Ic4hXWHZI27OXmZ9yWf4+cJsRt8rnH6PFakD7Ne9fgILzeKa7n/6dhK/cv7wE8+RCZY5AN6MYkKw
N1NDJgf4h1ybypyAtL98aTlq6JHdNqmC91kBqcEeDG+k1p9mcpn2ABvTFs5eto/C7aVBenSPXsTt
a18fKDrgAFf1cugdicmWzFRyHV50cyCwd7MbtSHc8iEQCpWstgoyHMlYrHaIssqq7+Nl1SfZ2Qhn
DMwTJDL4A0owBG2z8de7N8Pwp2j6Ld/78C10rbUmfZf9Iunr7/w9gXDxbYMnrL8ZyKJhhDRVRyyl
TLbEtD+YFbo+Er7c/UYxO+nkDP8ICDvAH075T6xnc2TyWo+CWUB73E38I6yXOe+nj1W3Tf3KE0oz
/Z33eUj1b71JcBTePj5BIFVlSGB9IvGCH+qovw5WkDcbrS855nHSX6dlu8dTCNqYfKORzz/Nuvr+
j0np3ofSZcszmTV6pANDkMnby9PoXe1KzSiIyu2OrjYxOC9u5urwvw+LliQkg/j6e+hzxD5VW18E
xVkftBXifcBIUtp2G2jWA4bYXGTSwXY2DtXim41ZD1oXFsUKNGhzU7Y4Q9mzzKrM6JHDVDh0aumu
D93tExlS/ykYaSHDsV2d0weVkFMfEZPOl3EC4QJ1TOVcK0HgqkahN7ZRXjZKwBqv4Jg0zNEUjwK+
M3vYhbviErOyzUHGV1vurEK1ArsNWZGxBUaQYdMaC3eM/GpkQKeJvEHeQbC0lUiWUckslAF/cTY0
e5qtUBthvbAs4EZLdcfn6i9QF9DJEHpQ589y12sIQwRkqUBSwzjnh2y9cu84519Y5hmOsg5qrTok
0uKg0XPxADKWM0gMzQnC0yRzLOAOpJZVPizet1k/ddtdajr7LYaitfTdJsSLnk/MxWpu+HMejaj6
WxVGVBNDrcTGHA+gRwt3pvbq5aUesy/Gb7BSt3/ZG3YeW/2IEqFI7++cpQ4fLtlZXNh8tlUCXDyl
uUnTjfdYYoWmhoRuc2zfo3erBOdBjMbi0h4Uw5TWyGdjwjEqyK7fyjJkF81/SaixA8QXltFKoaZS
OlZmW8SVcJ3BW6SX2WS7dkR9oSgD2wHm1BYlybhnieGtc3oxi/XbRjjDuCEbk2k77N1X7hABzdHM
JQOCD2WAmF5t0RBoEIGxMjqFqe7z9IxTdiPEqDPr9Ay/9J4lgvnZqdwCT5oonL3YqEaakQswohf5
FEbew4dF5ZQZ0kcKVvFKzCulxhJudKvLDy/ohDgiYSX5qRCCt+BAsZVMDAHjVanbMkh0rJSd+au8
kyfr1nT2KoYxsggwO5ED5TFr3f2g9ocOIHd6gnjvGEjK5ZZ31h+Sa16Ov4sd/ER5NPy4T2x4aQdx
LLJZeta+pZVAIwFpEYj1ADx43IR/TEmckxJkkX2Q2PWH3bHcQe7PvpZvLyGBq427HhCi0tOJ/Gg8
YCotlyAuILrG1OJXqxAB/GFXmXPL5bLzvlWVnYKMWMOxjdf0dMvNm1yVn5f9H7fn6cTzLM717LEz
SvM0xB7SsqM8A9c6y5GrP5TLzPCgm9nWuMaaeBHZYMuimPBn0jzd3ermZNJ+oyaJx1AeCwhGx3hP
DRotucrAJwUIGqxTnhamPnsQWBCBkLlO7W3qit/8RAS3X9L82LpaokOHxqv2zV45+lW6kjWOCGDR
SKj05sOu8Ckg98jMnMMv6rEBJ5hO19CiE5qbyF5TWsJvme70tEY0QBcn3uq5sOXIlPyJp2xMBDjr
Nn4Za7ABZ2SRsmZWnuT3paQqSHQRQSpvE6llOi2/pEB7FufLWf9WqeYcUtpBOFRgwD8L9nFDwpay
B1qfrHPbsnFAwx54ZaoAyYQuCDp4E8mI9sor17DjDmrECShWq9cAcysTKF7TRlKFsbodq9MmJt0V
EjbpJ7FBivPJy+fz0GNjFd/leKZ6q3fBgxKW4E555uLP7tT2VLbX+EprNWVN3dzgcLmb2BZrk/73
g47Ddm4CZ01UfNCWRhD+ZRC9Dsby9vAbDnHYBqnNPqmNY7T31IPZIimujfKgeg895ut9j+ksi3vc
DERdw+xoxSimFA9hNIZN51txjiHpfhldNZ2FoNc+lP1DXOSYXQGau6KVxXohGXnWmKShEaKPFhDt
awdmvHa6XdE/xnDUA+QAnQduDsVEmRbNDieCLZ4gN6iu1ip+qsfAlq8C4tmvp1RX8U4yNL01xFwV
a4y5x72cTezgu8dB0BIBnJMuXYbgjj0BXzEUn1HEzSm8Dot/+BHd2RH4SHwCJmtodFZDJPmbLSie
fA8b+TwfwXbXWXHrJWm9pA0+/6e/BI7rcSf+8koyqBv1YYtJeQEzkOnQXNwYQRaJJvf9FWDW+/KF
aqYrRHaxHao1BYI6gCmXNwcOzQ0Z2OYzCLZwqM5R77UZzZ1lH+g74xcbL5wagW0ATic6CYL7pUVh
0omgxfe7H+yz0tzPPiHojWi5lITFcoJwyWyppLM5Ehai98O60SorU0csQ0Oiq/I6BEihZcu4WEcj
ubQDtR29Gp3nyfM0Zj/tVG8J+Eh/dVwNo4vfqm2fHf12ibuBX0fSQNCRcCrbi6lhpWCpSAoQ8S44
jJaQr8/AtwF4KRDtT+QktIMOO6LZ4YQYrpuONJKdirLzdX4+AMcw6BbexQuNk1XMgVjbEK3wW/Zw
79wnV0ihNadMb5W+r9OzuzkDM/2X+FNWgdiKudaycAn5gPSbct3x3eMnYmMmmo/nybznCO/b8Ul3
xZXxb7T7SAeWMuoUsgeJIutgilBJJKsOOLaIzZDNnzmVp9TfWBZMoSUj8+qToQM9+S8T8HAJUMxm
OSy6mME0BhPw4K6JHf+0zPFpzoq4joSnwOgCIKxne8lDu7RQYko3lGCe2S3F/NgQFD13UhdalrOH
0B4JjxhQZ8wqe9DM/Tn8TgEUOU6CvRQKVZyW5yJZMUdt78EKqg2z+G6oR8RrzXnLXOuACPX1hsTC
TU54afb/r8p4UbW8/MnGnw47KXcDHnCIlVqbjyNJrslxhOfKbAAHNskBmUnIBQaO7iGZjjdr5H9D
euuMJ94ATX8ZIhxo0huF+SjWjTLN+VVtfewaik1atwBBmiFpsIqDhctMX6d7SAFEXdmI+Y82b/vB
wgk1OMh3cplpJ15bl1xE9rUjq/qTsSIM5f8m/nS71f/8i9eCtWQkEKG4upxSV7SAsCtgTmc2L2Ib
3gJyZHA5O5dBirDYzRJ92KY+rjgqx9kjelmZCUBjgb8Z53lV6aph/MQptnoDOYWyeD8PN+Q80mhx
Jt82U+7b9StO6yTxyoA4uXR9ITCdeZAc2TVpykf3qc/7SWI3nfeQx9iZy+s7rT2mIKlOYgVjfvdh
O0Z1am2cxsAbl6Mr8OpvEJSe7o2q+mUH41XJ1JhjXxq3NqhS/KXoXSRNiINGynBRzvRMPlMEDBtS
ENF1deqsOpwzBETb4lfq19MywNTQdKd199mFSjj4HT5rQ3gCZOCWBEaBBGUpNuWXR1H5GMSuNThM
ehjyaQljCvRuTNlDoL9e2DAYKK0PTXKY/2vU0IRc4dHfych09yc4kYk2GaL24djfUgyIDi7nfS79
VsU4wIvx/NNZVR8R+kl7l1tJSx5+U8PwXs05vk9mQDiiTUcIc4UA669+1w7LY6fWqxwIVNKoMTgu
+aOgvKC9Y+a2qX0BfBfAgXdWwCCJZnz/ItprpqA/FeMR15n1MSgCzuhedLwq9vEpXNT+6aJB7SdR
t49xCG1eCJdGmd66HyiiDOcJhTWe3esDp63UAtajteg3eMaZOtdE6dLauXQ+PRMDgE6fErAya5kw
KynPV9KIZB3L16vfIBA1WUVCZ5JsEFcpEfSn33YvMiSS5yIGDD7bhZRkztDk/DlOlibG6s+uWcju
whvT0WknOjD+fpoG4KVoMULEF55uaE9EFlZ6XOSdxNGafqWOPUnuyimpyCq9SY1cLZsK/DaXAXAo
yYQYw/Qs/SWSNVJ92SR1q1J9kPlLNMnx/1Gip4IpYc6C60e8d8Ub4Wsh8HSIQpRjtb8KF/xIQ0Ed
Xdf5bCAhgkazN5nctu/nbH81wDS8xnWCChd57kLjYQI3uJbD3BOs4nejrNyw3vHBlBhjBJPNPvUG
Vw0eGZUd6+RpZ8hltPPDc6HXYw0/yumpY6jkj6D1Np8N2knXHjR30NszbjO2fQ47vmn4ZJ3WxVkL
r7dER5eiW2fB9TZOm7faJ5/gShdipIxJRrFJJ8ehEJv5+g4mausaxAs5CXpykOg3r7Wj9k9YcgBi
ViHdu+KOFUv1zpWnaGLHHtOsz/zmwfnHEeOhRKDJj0e/DccaUpbZnD7/UrsGdSutWcMagQimVSjz
6m/fW1+GGVEsRhtMG2OGHInFDg6/R1IXZ3B5iFfOKM4CROC6MZyxPGcit1liHyCwPid90tjr3JvM
vyBvDtaQdKKCgy+cZ7CF1+oFlFmYtHw+iBstnso0TbdChoGKSmVEk0abT2MN8hpb/u2mHG3EO3Bo
ym58bgVxTfyineu36otnDri5YEUwJ1qxK3wcJMeUL8cXwCGkwfgwTLi4YlkZWXtcltNPBUHjrKmf
fxiDtqa1baxYmAW/4MECmRjPVCYKKJC7c1UVQImjC+XivWGyoMHL3TrrKkjx4BUuXlhHGqPXUvfD
M2wSGVuuVqASsHeeX00mBJrEsLJdpVelB9gqtbjRg/0ZrYe/6QTSp5+jnGBKOQapkdOdl8Nvy1HC
mARQ5lMvu8GxbK+8PNF+X+0HewzLdRMDxdfYfGvQAatdvl8hyAWdHovhuNavFXe8tDKu+uvxHb1b
HT7cy+eKLOpOJ7xUbItcFKekFtERJ7RzRwViEYWRfKYbC9HCeuOjHqYmeD526RjuhIUoYR5jRNqH
zVnT33VMLSEvYZllpLao2rfkxtXOzpihmQMapeop5DQebbBw+egg8sWR8KthELjvn5qtuhLJGfhR
bNfR5vQcMHx2kvB/MbU/eZxYmG+1soJAfAj7i7ZCFvgn2fvcbsuKFtWdnL7nw9At1NrnS1PGwjPZ
2W8WyeRTyW3ZNQn1KdTCX5wWdGPN0Uv4zEr6jMBQrH4RKkKGBkgllVdgkMELR45q1XXa8IZBa0o6
SY+V6uZzOflaJy689UyT0SdaoZ0vOyf9KCaH2y7AuX7xUb9gMHbkHXTx7FbLcccfYL6YYuDc71KZ
/WjXiAU3QQH0QCIXmsBNWP456ovAzUe3AE7NhdF0i3PWt1CPVwDuRm+MG3Ngn/5106uBhCXlEUuY
/t2ZpsZxWlsHaoorK7T9VWr9LJrM96cRQx+i19/VCNyldY6lwESsBcVRHead54bmE9CLkf/Muojq
dDFY9TSRg7njBpXl6dLQjO+OZwwWYRyrAFbLrkjlbX7cmrL9yBXRL3REnovjgW9K7pExsU/cVLto
h+3shMRAwfyDvnhy9PbWLNxo6phq/mRLYoD2eGL+7Fr6514QX7NYoyvu/afFvX21bu+4betX2ROw
aILNHiEZK1RTPg6NGTBKdUhIUW6BtoYlRrPpLq1E2t3JOAbu9DURh5xfLclaHIDZXnlzRMN3owHz
6bVFMY5bkayvKvfG0rbHyo03G8M/qA9RCxg4/lSg9hcfI/K0Y+jHWeeBtdKYWH6YgUplDPmqaYh6
RaSu/Y67ki8r8oeneYo4xQzlNEo7uYeJfL9aTjL6dW0rjGg+HKbelmR6mNIeKl/seWr3zk/mYES7
EeFIKJHCUPOkN5TZ3FGIxm2r4/6MIzsnJ3/BIkwh9xBaW8LZBcj7xuMTzQ88WqeEXXI29eqcLPZR
K/8nX0XtN+FIgCAOOvQjEEnpyPEw6uBLGw/FTokg2EWwCaY/8ywspCxpbcLxykz7sJM9nVFtywX9
4ti+LCZKavhvObQynqAIzHxdvpbMEE8UZ4X+FYnF8JBT0EF2thEbsbgQ1NanW9tVh6cJxJNQOpCR
1mTeV7Povh7HtgkQowp4eNPzkaDx6H6v2t9WipkSPIwCWd3JPudpPAuFu4DMMAhGhXDlCv23y3na
b3HIz9lV+xZmnhyFcrRZhGTs/bQ+/+C/u5VkSX30keqOB+iU+Ndnfntl+UuWzl2RmCIokYiLCKHq
0tlE3WPq/pgdnNLTnjUzvLFsWQ11ASSK2rW2YhsKJyOfg3QhV1ccp8KA35islZ6Ps8vmuylAUm8M
I7xea/EraYKGGmDaJ5Xh8A0zwzFZm7GvsTEwKUfod1+91QGA02kniFKc1f8nqyUFtHHqTWAQdFz5
DeaGbwCkzM4fWymiGkQ0SlqSYrVzYArrs3hA1WZphLH96AzFlusyOwpCq/go/xNLDhwykwxT2ewD
MHB/YPlk9C/5/RNnd5rwlR0ty/B05sV/CQscEBdJhS2ziqijCmHmTrmN27ls9CjjersSC8z4h5v2
DfSkGiN0ZI4TXL/OL3v3MgD2Psa4ZYFdzlOeDpmMhd3rAsdHsU6yYhftxWwQepuAbWSd6hOwEV46
DKVa3RFidz5oGBwADFPOEkzbIyJOxcfwODlwmQFFneJmzDPnwPyIOnr72j/k+d49QkU4oWOE1Zyj
9AFLpiXzpiO2IeZZwXWlJF3L7oA03kB7V9l7dZ6xYY9ByrJF+9uKleV2W9pi2ru4ONuUHd4iTkrh
QrOJkWttsiMW/IWYH8FwbM02F2KfNe+2fvHGYRNh01sLDu5zmPf2gXoyPyZT05KOXSNM2Df9oYK3
nz3aWUN82Jxa+oGrBDMMvuLZW33vnuP9s4xfZWAKk7kAnguFd9/AIyi4I7P1bbsSVDAH30K7kEWL
VSGwt89eLQrvIgNsgHfj+tJ3VV/NTMr/vSxXC5nB+8EYIYA3c3Pgz8w+wES5fgwBYoYaLXlmWvtU
ffzZ5m7bCCHiCpVWvhWd7y+Jm21Ox3+8qfpD9AqgRKOlHt7e8rog1sBzwZnUcUiysCiRfeEidpVT
AqXMbX6f2xBrBW7+bgzrHpQx/qbPllvuWNJsePuZ1R4OjobN6YUpMRx49w2LIWKZsEpGwic9Iimc
HlZbmY8JT3tHRij6OIQVvCq2OQJikb0mfg7GxqHex4J+J0seVXuvGCwvMjuDTeTQfvPsNGhzu1XW
LdD7dmAXHCGM5NdkFZtsXG1DRkjE+WgTA4v8VUUw/FZ8I3klTkBgYoAtgHyQd4CYWISqZV/yaG7m
N1BwPMGRgG4hUBZpj5XYW02pE17hIzAuRDrjymnU1n50UuvvREtrRM0chHCjH6s1ysLLIjB7CZiS
+Kskfljb/8K8RsLqhnFdibY5djHuDLEAitjJdko7/LsegKb6hCUJlbo6wat8iP3vZ5VUkXfqiGXC
VEEj+th6s2FhBaZA30kNKmNKh06Y3XrZy5YzcO3Jb0QzscdMpMGUisnbiuzjxhiA07aEiDVxfgGj
FzdZxCFOGg9pgbUB40KHkar23BZgqrrdy/BEDJ4Au9+AxgpzcPmLIzwBHEiw3D4v1qbjvvo2vpEs
5QLOndZGFRGGkTh55h2Ac6xIXAME571jwd74x1bcPMRmB5g0rW9jnXDaGSWvLpkX0Ih+zEZalkVH
kup5h9Oz612/Z9GeYds+nYnZfsghKBfHFY6d/RbInYvDMzwvML8f+cFL1Qit70Xn7sAJYdcVvizy
lmSEUShKCp1OrsPxeQx80lP9CkuP68kwKVye18LK64cgy5pXEmiWdNwIa/MNLQKCNN8SXE3h5yYs
loCn6u8qED9l4hBxSXBBJaFyJUpb7FOsOgxzQaXQecyJ+nRgooqBccaXE9CB1/VqJjOW1iT7z4T+
2RUJzXIVSR2I1qaqUtyElvvecha8sjNxEmVGO1O892COnGQlAsC1sk+exzUosAjvZzI0sEuMEDKV
6Ta6abxTNB9wirXN9c6hNjC1r/zsJSKfKO1YLLdPk8RMM3y6wB69gvND7daESsXiKOJzYsXkwntn
LWJ2ne86b0WtEiy+J1WcXd2sZH8NE+5Q0u2yaZG35RMmarVmpJHizDYc7eG+3Q/deVMjYUWtUEGz
AJKw8/hzYOKz5oFJkvpogHsTRGr/RoFfC32gEQ+1WsMNdoaAOoofw+7ECDDlK1aOJDDaRyXsC9Bw
IPjOlto96vUsuN2NZOOItyYeQkYI6cxeU73BwevxoVqhYoIbiTDDIr/VgXomG0MtOamu40SGTDu0
0Ps7UguSfMGMyXDOxdvU0MHFVfpI2rl/jDDyT+tAKfwr8jyPB3TWdLxh7TeyjrOlQRvSn2TsaH3K
MbHTQHDdsR3mnxi9qMPn/2rGag1Xh4fO9QgQrrjCugpRPLjXLb5FSYEgLucszWb1J302UTpG9Qlc
9JD8wNXh/9Kd1AjKd2t/Jh10rXK+UK9To+LArNAliawyupifjHbJXlslOc500Xr0x7AFHrCvTL4B
LqrWMbxd2YKOhqkpvrfL+DmeKutgggLVoXK/A/CHIaC8Jbm8MLgmnWWszYNH6pPoxuV58VGhLlWH
7nW2y4pB+X8mGGQwByt+MstGop54m0Dk960RVXHf+YAcwmKbE6QiYxWw7BlRmPTRa3K4H2ZxDgY4
UerMpZR2lFSz2IcamWFjl5P8VaGM3DSYhlRAWkjgILAbaxRrNGoyZPiKH2/gM9Q1CzF9YEJ/uW1q
B7ICxHzeQRBD+o0TeBpQm6X5XhEYZHnsmSsa3EIa6MT7VDFZ1AEinhMpE6NMrql1361mQuyw+Jvq
21ahYp5P4AEyGv/c75f8KfF26PfP5UhhO4JqBq+vnjzxxEsR8uk7NuItlyU38U9H19RV7bmxTGOq
n+du/A1nqezOIVnXMLgzXh2PCr4KLJrlg/QwZJJcZzFqBWKCeVkvUThvfv1hfOFiTiKX2IzYN1aS
1EDOaJfNurCfn5L7Eb/KgoywJ/BhguC3AsC4puC9LDUD4lxo3Fi3D+fDyKK5sOpMWH5lE3CIH8AA
WGu4qevm0sC5A4k7HOacOc1YPWkY5BdV76rn7cigrcZVU41bkc0WZUe1ThVaoLd2T4UlT3i56bLx
H2KJC1kRRPWlZcsJCc5DYt1ADfHwQDTPHREBve+LAnPTsDQoFt4igJ78iz3fhwmDD5/mTFikOE1A
NDezTtq62NeG5tQpYGzepRWgGp5kw2ZnD6bqZVWztbUEedUMTYhOD0PtEhSS+6w4Aw6Tpx+E0eqK
RlpF0AT0btfa+V+5mnanfaLO7l8g7ao0nj1JkVkn2xT2nOHtlxKc+2kUWbb1BPDeAoA6TYf6j+X0
O8FbEd/M3mCIj6Ajw4T8aKlB/2TEKipQZD+xGozUgC8TSBxKOW79xwamyPHBEDccqk+kTxRi+jRz
mOFW4VLQuDsw0GX3RHFwBzy7aV1Ld3iYBJX4LZwL3UUdlP4JTXg1c8/jfueJtCL5pvsFiC7NpWcQ
F2f8pnRFihenfU+EkQdhOJU9RqRtvL/die7Em20P7v9l+z60IyGlMbLVLDjJIdTgLijGI4dyuGCc
Ui8FfEIYfL3faJ57s7olxUH2KhjyPwGZwd2jpFwjfWPIq08ijkNwHq6MR5YzQuqikae9MePaF+20
DLQeQduXzGjUFhlL1wHXnHPdT+b6ocwHCm/wq2Dj11xi3QoRqIcgYgZr3glldBOJUC6mCnybGvfc
LdXy8Wa3zyBChKaiz1DGAHId2UsNpQJObHMAYuvXj+pLgkR3AldSDMeKtJeYWmCSxv3mVLononAj
6MIEoz2BopceeQHxytjEEEj3/GWkRm9pfDdlFlU9Y+E1U212JHX9I43C4HPIrgepIN5idR9hE4Wn
3waXhc/Kf3PY5L9uPCsDI+CKSv5vInucdOs7lYoHB5ar8EXUyxpo8LjGy4870MSlgfOotY6SU3ak
pNXaft6PsYvkN4uyRY1bLfBjTb5FN/N0z6U67N2houe+JZmMlslhWwmuh8ua86W1DYKlY9qM5P/F
KZv9c9a82L5o2auGKAsMQrc7XJl/qk8R1vCP8mpaWoy5MM9l/lBCf7A01WE17U6vv0x0h2LLHe7q
MxCLXclCMkObZi/ZQnL+N7dVT6AIpvmLhjRHyaLW/ofCfmrlmSzYwirJXiRbSxZpJhMXIsC5LsbI
zdDNmftrAbX9+FTpz2tBKrBW19NWPK245uZVDKMWBVcKk01z2z2uDO74rQVmnxmWPvh6zfnc0Zmk
TZpMoSHrDu5O8op7wg82NrWcxytUvck/zZRYjK7m5fZ+XJOeUOHRq7JJ3+63seFrQowVUOM+sd7b
Q4tn/m+j+43yAIa9y25Vsim9KAoYMCpbsgaZfhzVYUEw7NC6NDF2YO0LUCSv0M9Ub+NEtLza2dj8
WUTJ4My+rZ2t8sMEIK8FWcIFdj8g/ZMCxKS/SZKp2wYdphPb/63SMm3mb19PsTI7C6k3NwvyoV6C
EdLKw+sLvCPwS9f/uH27CO40Xd4pOSPvF/QB1TWipMvA/4L5eZZBkXKGSUb+Cz1n+1d3pBMMXZnc
LZEia8az1CG7CXczIrNYWwgEwOpD/KezCO+sBTnqo2HUYJdVLEiFybD0RX8Juu51rnpkx5rBfwYn
mHISX18bDMONqr6hoNChxd+fyOCr8eWYxvJNFeXUk0qEji9lIbbJP5V9YIxFP8QzESXT6gtYY7ou
CE/UkBpNqYXtnmBSuxGSJqpIZR1W+9RroPG0H66euh89fUVxhs8Te+tyhmcFEvrf84ZZOqD+VPl4
sSuIY+Lt3snjI0FPJgsDp0/4BJ9YhMt/wt9+0quXweEC29Ys3yG3+MpE5Z50QIm0JWi7WMQ0lBRr
ASGcgh7+PQVPVvBdA2DsifwdEe6uoNCdfLRgqm6a5d3qvIuXe3dj4/0aHThj0DQ5gi+6mJMd6gui
dKtW2u2038Wo2o1KM3Onp66zhiaN6EGzD7wdRLffKsFijVk7MSaRbaKrMa7C2ZuKRE5bkRkHHwMk
oZcJQYXOOTF/TFRhXbSIrxWQ2jpsFtN4vC4FqpI6VdpQ2o1NhK1yDMIsnopM4MAwqC4/pvtgN1uU
hU8uvXyqlCvUzQxr9qs+u3rZl7ld+E8VHIeH74+dlx8dQAgT0KZKb5KOLp3ov7uzmFP/74/uGK6B
+vXzefL3uoYLCieBQdzQnPV9/5eBDZJglXpUVAa4gCAdEK0510m1inVCBcKzufczLZ9YGoUxd35Z
PYQiEO5XJCZvBY24vp++RE7/Z1RlW8CtUrEKavUu3gvs8ruR1bnpLQuM69YdskmCPSX3jNv8osIe
A8+RcRhQYuHGhD3RNEcpjT39Pr6cS3EdMTtmJAU0M/uvHhkN1yWhDygbR0yx+eQvLfPr+KvqDKCO
zdoF4WXe6b4VRjshCPI3jkZLOwhnNXg9aetMG98dUI3Yrjsu5N2TAOEeM//RwYs+jqpMe35Jx/Mr
NinfDMYvq6UV5K63SqUgzePZVF2UKF+JfDMScwSClrJbx6zddteFDmclGwzblH5w2QX0N0j9j5Xk
Vhl4x0DFt7L3bP9lHg35ZGc8OuUXz0T/pTyPOkLGevzMY0JugVVcN80OManRLJlT32vGu1ElV5zU
HEUxhrqBnCq9UQ14zotQ0G64xVa8JeCrfLRde9aB0sfT9Fwk3bUsc5NiN8jQU+jn/Wfb9LdMI7Tz
rE0T6ys0TEjUj7OnjNtCod7RzNLHlxJ4EcUcKhMvOeNJZqty/nU8qnAfXo3wUGhOp48l8Qgf1R/0
7v5YoJA2tLDiwnOEz8Bc43LJkHXWC+wgh4EbGFwZhfgeIRiqOSd/cmbCe59+P8Xr3GHQ9YxtMM3/
8T0i24v3Nkbwk1Eo+hfwlPr5X1NQHjvnPPAaGVfDnhv7iBVyL9kZGP3nRBkb3ylS319A7kAV24ZU
/IxURifRIwv+i1OgP+J9EuG4g1E74PhYkK78nR10bleIu/5cnlxbFNzJu9DGe25BydU8GjZ5R4XR
umTK4jrDrajxGYzum02tFkHRcRqhK5P/zTuqjvNqyF8caqJqlWEjoJWEPb8cbUkdbRgPu14/V+FQ
LogfN5b2yTGkKr5LeISE+kGdujJoRFDbsJX9C9jwClu75P/XrgWFg+dUFh+uHRGaj9tAhHZH6EwV
fRF6RSiL8PLHJow2RyBAkq0YA7BeoZ3fMt+Hh3EQMtHl/BDqPWdvI8IUQtJzEt4A6UhR8xQIFYO6
WGgOD9f10fzkH2WRQhoM2pBjCbQHwdn3Qrx2xZOOUCLhvUeyxWgiaKsi3RkAmVUK9vZowU1ykWbc
Ds4wy/+IcJy0XL2CgaQ6Ek4sHg2zMaywDQ7xkbjBwjtWNT2vGaTqvduxGvHYgSDPOl1z1HiY2ZIK
ZIQQi/f2stgsEHzxsVFdhaH0xY0asnkldig8jCTZgRCkD7QMsenSdz6bRuGNgi2XVg6JvupQvpJm
GLyR5g3XlG9mlruGvRNfUR3QTo/QiK/aHkLfU7V676hRGwqrjkWuKl0gEcy2BSipBV08xSariHB/
v6yrUBqKEG6jMTdF/wgdSyJlSoPnJqRTQu9fBMesmt9FmEIx8vBhAPFg1EIP9dQ40e5y876PRNIa
2HZxN9urNnVbbUyQJyRrbeX+vKxh/D/aTnzxrDguTSYD46BT9KB3DqcVCLhYAUJLoKom+2OjM1a6
5n4d10O8f40nPUpjSxXXGfTctzynX3CNeLPf7m5IOh5ufAlKY0h+HEw/a0Bz0cU04cj0ObATapRG
/CQVsreHcjcopPwF5RpkRwKj31exLA9FSGLDrKZ1Ub+F/FNOtk04DfoJgGoGoIh1eHETUkCx3HNP
uQoiLGzWdKmaUOLPITS1xpCn5XqBXHdW23bNs7li2Ew/GBI7jJVtxFwQLVLxJiuamDtKmVKrEGo/
ZptI8+4hYR5ssjKgRvocD+PWrImpI8MpmJ3aUd43yEPZMQYIVHu4GP3+tuXz+1w2weqazs3/et4f
mg8RgkY6T5DkP35CVGgNgmZuHS+Ca8AC8eNyeTnC460PoWyK6Hgvbal3zuZqiOXt54HwbB4OOSTG
qGbIUpe6D1CeGq1Y47HIkUpBtkt7boefxJtppLdzNbIMvfnFLN3ap4nxB806lbLEdUCmOOsi8tJn
+8QP8x+j9vjr5MM65Ad83xoxSbyG95mABc4ntKMAUeg66emXwCjR0z9/JGhnNDl+f+HHfqaaMO+7
8D1dn7LbN7Ia0P45njuRQ110C2LVbp4phI0cLc0sscAbqaQqkq7FkSe76LVAgPGFKVcvHt7+NyVi
83IglVldoIesj/Yr/WHe7a9odh8l6LainRcXhqsiEuVMp9WF6pbkauphlYv0CnvoQ/9HaWlUPn+t
y4uO/edXb5MFnq6zt3bmjPQJFnsqsS3oMcx3aCdJ5yCdT5mUBx4Us+s4K0/g4diFb3mx7he73ori
17bJEr9wjvqXnjli/uWooRRPEU5QzlkcqR/BwXpVR2pGopMnniSjUAQ3p8dmzz/0KLehgbNIaINL
GWUnc2GbcAXkjU1YSj/Jxkvv+hy8vWVRXv6xeTQzxzGvlBmgJX7MyCSiLYyoh9AfhTqhJ1AopSN2
SmUODf8Esze6kJQxR8fzqzL5Dxg9Co/tZ8wVajZmO3emjXB/hoPZtUeDMDJwGUVWUtPIgjXyUNoi
6msSKdVmIb2ZyyP/mqdQVk/6G5etZ7DSu1TurzbvNFwYqHsEFzkhXigaQGp011gtE1nzVBront89
m4xZCKA7II7gxoU6ZTfIyZT+BNZ6+Ia2d0Jvmp1Z65MLZi3bCKCBLQ7s/Z8+vzIZgauX4hvmfR3S
a8KSN4bT2Ntak7vOQiUFO4yPPXJSmEPtMVhoalUagm7M3yzXRKTpQLg8UeXG8Nx8ptiRVthcGP0c
Qe+XhDc2l85HCeEmn+i0JCgxgkur2Cc9pztzSN06iszjcvRbVrkGDKXq+PbdGskcCoP6qm4QR06f
tZyN3aVwV2C0hmvwhQHY1absU3pXmP0/0oeql5aYZkaubJ+ziVGtoFY+Fd66WLPCcz+4iiSUxhNy
dNWCjTf2DeVPBZBBLmNaDdqMR23lMcDs+5CwDeEw+J9+vY/WSnhrB7lSD8mnDR9sKy1InLVRv1au
jBC/MPZy+wiTggUVVgJci0agPkqxzOQUCeM64VJMfM2l2YHvSbOtj1X/7VFt8sThl4Eixy9+1Akd
XT4M2Y02AFKvp4lIpqd+EBSIOmgsw51Z77ZWNXdOnMmoPT5Mj4J8YyBywDWXH8tyBZtAWp6O4xcV
95FcgMaUTePZHTQj5K6TpUnt7p+Wk6jtn7WXZcHQDfoyRoIbKajq0ow+4Su0VP5YvNG8UWwuZ1jl
Zt9DORPhS0y1sZKaCnOJ3XjJgNoCRuwimcSHy60a12v+8gn/cgO7EZRI9Xau7W7NfYvbpJnGo4RL
4kXZoeY2wdHgMIMxKPeBz6zMCUwsi2mqydTJyBCNYDJTDtHXCltihsMKM9z6XddCcP11Tr8B6zPL
HN5mx69+mTxCax7Hbf+iemnImNkfPXtLYsuiVeV2ZS1/NmEJTG2p/I6+Kx43YFiPfud2eaMMWgVo
6+vgF10rkVbCxHHR7DgodHMezaXVU35ip713/0PbSb8UY2WW5VpDVDWpbu0SSsHVRK8YOFG+eeci
XfN+RzyKXCQneFMNbLCLWQtqJYUzc7Nez1CTjTZAhOHkQiTNyoMuUwJI36Fih109e8owJtAfcK28
UXBou/QNURF7S6sS1C5FyLpr8j3VnbfJ8imODej0B4u/d2L+XnajWIU9XmvgOiqWQMqEt0elI0qT
yg61wGCJFhDJelyQqD08S943qn+fG92qlgjitsg7SJtX97eQdBuog+0mxqhDFw/qdvQNoqoPeCzd
M6XTF2eNxptR76HtYYikMgMVb6L3xNIFwuqzEHWa11Ctrx7fq8t9OEW/SlNbMRxONvgiHhDqHyhN
yRFfVfpNh13w3V4cnlgXd5DpIdDR07eVz96HiqUflR7qOcd+cLXcROyvqI54qoGoAByoCt1yWOZ6
/Xnk2h+LyacYsE1ESRuufVGyonFxp2C1E/F6qifuAJUQuELOyePuUZWBRXbNbGKmIevndBimdGoh
8kcdn+qCVbno9T3Wz1DAWBadvywUbYcJ/wUv37RShcsImqpkvj162YIoZJnwD8dCty/rQre+Km6t
KJMavgzWhTR77san/kByt4htBxHFoBykxVfkxdhzXup7/r+8VkArKzCCicZsL8KeHs4f13hlvQbS
LtkIpAcZlAOJBcK14g07f8LCLME4njyD/PQZ75s/lhrZZY4je3NjtRdX72jwFcsihQBf3VDAYn+i
WhxM4m4v3mgSPNj2j/jNgWNU4lkpGhKrJVD/AlKUZEkYdMOXrmKRWDLqargUZq8/soAig6wkmOid
nEP33zR16/Dm+A8LPSLWYMDnId5mvbUQMyJPoxh1rpIhSp12W52yTBXzC+GCf5lDlBBPQ8TN2cK1
mSKHKaxPorMTFSZIo4ZFIEf8haV+aNnV7zVqiamCMaEYDWovhtVslsdYonPQoSfUwBK2T5rDu9E2
983ZhNee9fG7wqVxqTkgj7lWzRQdN0cBW51aCDX9UhPP67ZcJOy1V2vXnHga/ZiC7Ji/DINzFtWZ
3w6krTK1MQyWzPZhMCX2XcvqkpdxD3rPA6qSUYB/GQhCl0wbwpg23e7yBMRjypgiuweOiZrHKtrb
G/ykaPaddXcVwhUCWiJt43CDjZzYjB8rLcfRJCuCVJo4kAtzI55iYbkrYUz+rCJU6D+XSpz8gL0I
A3TpO5IzfaR+Hvcpb7f3tlgMAGWxIlPhKk7MEP2VxCqXHeUx4/odumg9IIharDKbuuhc0cYD/GvG
vWPUm21LD6ZfdjRUQpdUR5y4t3l17AOON7QfsXbE5jqouuodATUf+4WacWhhP1+p2bv/bIGd79tI
AlcywwtaU89gHg/+fYTfjxng1i8rqnSyuVBEQ0f0CIagp42yHhTwzkE9Z6AUGaI/k7gQp5KSqv++
QBGqpSNqXrkGfuIERjjpxav5pZrdI9vvhucz8KkaJfAdtHnzTaAgrEc2LACY2ovCOrBfAp7spMan
iC4Lj8+C2gbwecA5T/LJ53w55h/ZogtiRholBg2MCQtdin8vVHiFHR8QolK4oI8oMWbV9agNTaAu
2UTPgIjYqCoayZjGAFmwgcw9Dm69mwNR+itmVjv3sh7PNqBhLvHNvhpE085puPzc3j2C0+OY6jFE
ir9Futm0mNXC6dGVf9tASDayewkqUTcaxO1s/tgpTVyZJoShvMw99gC9DXpbJOcevJOEbQs1llUv
SQNPKUR7lzXqIm8s5YDpTcJDxIHrNMRKRepSdo918XyfYo1Q7gB3RJcDchIFFCWqm5bi7tsZzOlW
kbSncsXPTxxnCybnW1w74AorstSMFycQppDAniJ3JoG/unf42guEse5SdNvEtpk0dJGqdnQl/0oP
oDTPN14ymWmYxhJzsHsv4G8zLaLuFuIYRz4FKU35MqnoowbM6x3gF7n2JwXLpQkcLIspVOng61vB
y3fh2f5uBFZGdZsWCTdyQun/aGl9InNA+UAneFLVCFr/TY0Tegt/F9nWIHXqEaswLvStcEQ5Nfyc
373XtzYVyacM5bDcTIQnGjO7Dk0fshidp+WAMp/YTxyOjgu13IdxIL892liSHtdKSMLpgruMBXBh
x/7t3UxZmgI3q02ZdMeKX4JKq6d8MmKEhQeN2QHY6sO5FiEuByYzRLbrUbexAnD8Ihlll8EezABg
sgJCbOoSqJt1m7Ogl/gHmXFrdOlxE6bZQJ3G1YepsBTgNsI2tZaC8/u5WEwtA6Yv25+LIf/Y4X9H
Y9OVWESSmv/StVRK7NhY3cizgsl1EvHFMAdQyMUsFhA9jzy7elBnPklrv/oaGL2K2ip0Lbig8N6v
79Rde0YqnHz14tMzUXqLMU3Prvq4UaK2Lbp/Swq3JZLjZIb0ogNGeq62dvAB8ywnk7OqQEYisSXM
sjvoBW9LFqg+ave2jhPl3CTLgSngtnyYog9UhTzAUtusRYhcxmilLRIpSGs4PHrUvlSVp/JgHC8z
l5N5MQZk0i9uWezqPTSYU5MVqXIdjuFd+c9KfczXIr+Bc1S9YhWniRss4lR48XyMA2Lpc0+sucGl
2A2OfADxhu5ccFo6iab/zkd01YXppPSigy0ZTiaXa+u07FqUs8EFmfROE91W4vFBOt9ftgX50E2U
O1dGIUa9RpMPsATPbAqC1tZ+axPUrKFhDaHMm2EzYG48Mx3OVzUsPhtstXVTpEEoGpliX/3Rzepu
8/jXNstUyJrjasXPpDfjzqHTCdxhJ7xOFFv2nB56/jzYXZa6bMI1j1CF5ed5cMmyeTok4Uizet8E
fCMshT6kCFeW+Cv3c0v/fOyY4Ql4A7whVC+0aY9J6reAEpbr9Iey2zqYhiAWbMabbI6k45RSaSi/
51LymKQ+ap8lDzbzGBHD8p2lTqx0fO8+b5LGe356+UntP+4DhKKxUkycOZDhfVQc8s5B1dp4zTKE
Ph5PY7FByvX6ATMeHWwsgtFVWDvJQaQI7JM5bYXyNPDprQHX0GqpLHTboIrxSwbB+EFlfq06Lu1d
8+l1b7+EARdtfQScX2aXFNpnGyyH518/gmhkE6QZhl9ZfRTmBeat1aR9HgLNONl9H93DpqdonNmx
v2Nu1DBd2AV0kWW49jp5gR3fthaADpirBHyx49nsFcKxAeEeIRcBRoTGZI69WR5W6FzjoVCur3EL
9SE3BHWkuJA/bqu0usdQ3YE31xaEABhCMrMa4kCt95HyXYco7p47csTIIu7ZxNJuJ1VhL0zE+xjU
OBhMvkpVNuZlPEOW3ArJblil9O/X4JwX3PKJJvLY8NQvEljRbhpQaIveoi4JpNWlUadYudalTo6G
SYsT0XS91XTlhprH2F6qSchSEOHZBEJmzfiKJ7bdycCEUnXe0YsXg1pDmNQerAKFCpALrqDjdWaA
yHeNJwMFJBROsoX0bBUk/jwoOliZi1WV0KYDKg/Iq91ScvynQcRAkMiYhd/dw25x48nyVfWoz5PG
xHbKZsCVMverabx5zvgx+8J5x8l/Yr69b78dUpMKwHt8CDJiyCa/l9J8mke7GTpURNT84hK/MP7L
9vmTO2IU+Dk94J4b0I6niMUZzCkVWGnUdUM6W7xkvkzHB1qOImvKVeePHnzyQXdhWqC1khJ3MNTb
kwp1TCQ6uAdSqI1qAaL25X6azioV9BmBBDXjse+pTc0SD/QXw8+fYSZfbbSbEEareqaOFx9bqCyu
gRbQ2nIEVKgR5a3XsKIrST2rRtWnnMLY573MeDQaF5drTmb7ygG+k14qGKPoLHo1UhXZDMV0/8u/
tpKm+KycQAmLEyWJ0PVtCJ5bRoylvu8fnr6LxwOKcwPUxhPcCRCp3YjIexeqGLZ48FdNYEAxzno1
zJzzSDNo4EGG1RVMLnuGugYYEUB/PHq9C8UIvBY7gbO+v5p3vf0g1llqQD6dndxXFtNC9bwy0E3h
nWOlMsN0vu4iaEgRZh8dTuYxwN3KpxVKJ+PbgmStwVff4cKMIWL58cnyNrIfwJm42echbyNjsfdW
kHT91tiCh6iY3iic4NebyUWhmihbY/DQpPhUGxQW1LM2U+/cQMzNz4x0VA/FJiDdyZ6IObDmDhUM
GWZUYBzTNryy07Ej8KHcAi52VuvKpQM1QRXOnktcdnbtxIXzFJpCyqFRG9ws422IUOjqOMRLKjg0
m2s+mvxUK/eMt36i6GCfStoojRbWgkGVN5sHitRXqmXVVgJkX48EzFEJ3XoVukUOJtF6bBSceYMA
slZs4cPrTj9lj9d24QUFY6LJgaoGSmuzqs2Hiy1AcImSLaWI4Ia0aBytGGNz0xiTeVJ0z+F6K6tt
krvE5gEqXo8p1kKC9mQHRDiK/MjD/Aix2Eh7I+NeKihbITBMZDTkfRgWpu7Fmhx4uh+EZa8zthhf
Q5W+LoCMF+jogIpZn69BotV2I0p+jj1zFT0bCqjUjTZiBPD6BHItEYenTnqRox9+mAiYJvG0hbm6
K/RDmXElBlbhIPOrQbTokIU7iAYSsTP1bTgixF9w2t1HjtQYBEtYLQOh8y4TonuannoKRWJ+DWxO
JSD/OByyPw+PeXHBs5KvbsZbOPm6392eODpSmCQTCppe2L1UvLBexmDDm0QtvPEZ7XS5LJBF1uqi
5Yz7eMj/wC/8gtUdO+KVzEjAxTgAtj1slXLqIegcwiYefms6NKAYtJ68KF2WdoldardvxdS+2hrz
S0CzANTIDQ12vBY7VQmDpVaOlQY5fsIPvlvlEiCPAm/q8O6wRBH5NmUklWrSeX97PD00tzkHsQDn
kBxz0Ys7eJ0xsoQF880BnjUzlr0H/zo9HhFV63wn9IZiCrabuF89EC/02Si4ZnqzQ1P0m3FzwdON
U4vqOUD8gvrygIRRdzU37B8v6R9RNS2a3GtxoW4Z6emUPXarr7PUrv1yX53IDvdGitnwqgqEKbg1
fE7OcnA1RWQBWUxrBv72ymOZrvYi27nmMi958PUqVAK829vjOg6UanV6t850FjifM2RkU6M+9CM5
brI02/nHUFOxu+RMU7B5mEGWNb1ZJBvMGYsHSWzBXCaMLVmgrOo5u9HR7mmlRkmrpH3+cspT7Jps
jweWgwPEvxlSaiXYoBBEfvuHTZuc3oYBv450kMPeQqVkFQtmfb/Dj3DJVBfEkxlkcIO/IdtVGinR
kMVABSGLRv2sGsxI3TPWxZ5jHd6ShtRYUvkG46kKJkmK+vtPheJIFhO174tn53VoHMhX51I550Y1
QoR91T0i7tEfo/+9GXyd5g7jtO43UKAqDyIWvKoiL2lT0UEcRlVRT4dKa1rCJUYLw0Glolw0QNSh
HgYSjMRfvp0x/nRDLBeCtqhWQRM05Hk7xczTvh0tKuFiGidTGTesp5d+T4hN6DnBqSa+tBB2UhZP
gASrCZojLmYsJgHX3Yaqs4g+WWi1RqQuUtrkpxiYOd+CjJNEvtm/d7OdN8Xye5nEzFc4R9G9wbvM
6l4IQcYGoHaS7CwKz5DiFYrJAcwmYS6WPW2uVUl5H1e7rbKi8WIGpM7LwtEBX9OkD0hLRhkEKgBU
S/6FGtD58/YWXEyZyKlvhy/LoFYNDKeaiC+puq+cVJCGOFliq1WDhGSrvU3DrvOdBKdgfIYpbiLu
5Ps/Swf9UuNgtOt4vadYxoQx7ZE3MSyW+q5qqZaiwZMJwe9ra/3FbT/0MWTtJhRq7PGRtn/EoDwI
KUCSlgLEfGLZci+y2NNPHdRs2acg5u3mzyMf9GxC1BsXPblSzVpKJilA0aitH2KDlTeYitavhxV6
WUGKzHWWNeLpZlupaVrsuIh021gi6w6zPBlkPenO/pYUmeVrKUosI/cyXtVbgMYrhCmjCowfVDTA
CWQfeyUz1M2E6y/OIdFMGJAO5nRIg4R1mKuLq/wqu+YlFM70heMJfzZ3JR0IU76ln+fHaTIson7N
VJjuZ9Q62ybP9YTfur1m7jbui3JdDLMqIKRgywgBQvUMiUFDvBQogKoK00o6WDcbd4orZIJ5ftX8
VlAx6bC9sq0fQircuVLJZVazJRfot5TwGJSpLw5bA75qT6xcYZmICH21NvI6neO0/PzkR+6sBGfF
VDfGJap9RS3c/ZYfhBRCMa6C/929ewiw89seOQXZF602gKCjPrmS7zB3dlgHPzVZL8fo9CG2/89J
dSfiM65nvAywjVM3MAYhjoZ/fT64+IQ7YEWRhhmyufpXhX2QOCqV8z0+nmYUZGKj7sMrybdkUmjO
0DyXo7sxuZHNd5+oxAlXLx9v1+OvyodVPudBieWXv4Z1rkzwbr6i0ERxhAlrloldef9CsDs5N6pZ
bAt9CEGGpAvPp/SgJY1mRIv7mu5jb/VA3jHozSFHHEfnT1H4GuJWb83MP+Xa9dSeYUYMI5xsoKeM
RR/6w/CsADzgvax0S/rElcEDZnevojbKpLolaVW/equrmf8H4ubQgMz6TbWFxQa2m4ewC07O45At
kFdgxL7hr5Cdg8LRTu5Fru1Hu5Ui4QkThQE2+efX5AwpX0Z09qtmewJThrlWjG51TfWL+yQaybzB
FpShBYRjBv+mPQOY1X6A4c+W6CO+h1k07xVvapA9aJtdYWHboe1ReRC4whzDo7VMhDM76R6NZscE
DH8RsUSaWlslszKNZSkda77nUiwaFRD1e187bkueKv13vkhGdt62cB7VPFGlRyCgdVrq7lYq9uvy
JXMmOAACb4JCp5lrH3c29hLwRG3WYNAl6uApnSQwKedGZi+/1uGmnX60qqKFPN03/2IYJmAhaxoE
fL+YJlrq5dDPj1scSORQbCEmh6gS5hVwDK7QcUPKgoGSiReUP9Cjff0T6ilQKdN7avPstn4tbd9t
PMotO3KsFqoAg2FuZwCMab1N2/JY++rNMYu+4qHNGdYNC1lXQozik/QzRevnY+uHyJJpZ1H72GJC
pT4SUCcaL4y+PIVLgZs3inEQH9NCNMlyitedUXWZ8CnsoK8O2g4kiAYlTez1NRKfusXi9GSYZ36B
dBGYHo8KBUp++4BAzXL90nMpzTea3XNdIZesSAg1VQ3u6c43dkgCdF9MhDPhFQltnxtyOgGKt7ft
rgJb0sWyr9MuO/MuSh/IlafUPgD53PRezRDXCb2sF24AKrpaa+BOmYPvCq1BdmQEGvVz+rdRAbbD
JHOaIcQdMzhG3CmbmFK9rEMDKJDyOnRRKwfXYu46fHjBgekJDSzSm2vQa7UR5sajJpmlMnevY5cr
FO9foNqmBrLCnExXyViZ2sjThITq1yE5deHJxsoeVcWcysRVEq0sAk3ql97fnPltJauvoqeiHeG8
uY90zCnNUWLm2/MzU4iLZpYP71xyXEYJWfhFeAhRds/LW9qKscO+VrtdSebgozPtKJgFXqYCCBDX
0ECy824WMS/MpPylMMkG0BkYKg/G7XNTMiE91Bk1auJ6YaaOtHzISN5JFI/m4t3xEEVm2qj20HZw
yVXUXa+bbVBl6Nm0j9hGd+SuLXZKLk/ykaX9mofg25qFR5SzGZ7mfQ+5HuhRGc2blrXvVdQUfDCP
S7pIAAEk4E5677f9nQsLQQgbg6spIFhyCSjPbtLJOaWYm14hVpWlhvsT1DmByoHSAoxmRsCu+vKQ
HjE6lD5t/P3tvuwDzTJxHDoz7lyT7GKeFgRK3Iz/UazZHhpm9BjNggfrTb7k+MpGbB4z+qJDzHRk
WMU/OwypZTOc3ySlnUEkJG8Mi5O68/209ZOUik/hhnDh1Y630FM4IU1bGjACsbxztNqf8fMzDXgI
xI9ckWKsK76agcshXXGFuMQmciWcS30gX4ulGnf5ZtJZhcLLXRYPj3oA2DY5Nem6E6eB74shmUqk
RQSxXUbGMTiEKvLOSisitDXoNJjzVDrWcYRUQtumE42RxwriIuyKKxWvQIRMWiDjfJYDTCGuLLhN
dVbhD+QncHm+Q8louqcHQD2MD2iYtwk26s9CbktvJ2A2AE4stFLEucGXkjiQyWGR2gShRVkJhuEK
e1V+4ZuchNs1qhegOJwFOCTAKFNNZXrzldeVSp7SkAwB08A3rRzjL24XSYBuJqJLKu2MX5jQJuc+
o1RFCStkUV0Xaxr4ncnvB5cVpYdWc7jBoG3X6jTWzNydB6n6Jm2SlgN6j3a+t1393Eu/zfA1D/B8
1DYEayOFiMyy65/OGIO68S9aqQVaajusLQYcyhLkVTTlFQgCDdWYJwAW6aud5RCVgWhy+cjlYIXU
NC+odEt6h8zkSFVLL4X/ghTQ05lxBxJ4kKwVddGhsOe508Uq1YsV1OB+lrpkS/HRC1ePIP+exKCn
sOIBEcL/XxwBoi/7WR1I/dXSW0euKrZiR2GFxZNNmosq0VpphZP1oPErNaiUESyKY/Dl0aBcm+E7
PoLSOXSd0olwlcD5NhYcLb2S/PD7q5UpEozo+yEPI9dIvhc/4Ee7ucA5KMdlYbSMB6Kiq2LJf2+X
AYwK4TsO2dQmDscvgjTK0xGH2KKZ4ZcJXxX6Wq1/ya6Dz4DYzbtoGCeIvNpde3cVlhiavKfTk4WI
8+W4Tcw57DiSRcRYjdC0n47LrlLkurKzfXAAAyefiQyZYMEtvVzV6s6z1RaBYUB9IPuUy34Ryn/s
Mgb5LBrcltv7G3ExETp4aE5HVp9QUrwVCrPm6LFVB8hFU4BtkrNWhEYE1n9wuYQvB99yPRvqoddg
+PdpxNl/WKViOZvinDVErQ9skl5GdUawxejKhjrtVarqJCqAd6UTw7LTfi3k6vXyj5Rfc1FsGUxq
7XJomr8NceQf1DehgelygNAOQbQqImeU9T4EV8UCRwzpSxFi9eofI9/RqwkJvsH8crPp/9TKm9X8
LjWY742iZEEFdFYggNkSG+fVRSv4sUpTfWH4bjxezV6MvM1Iq0gCuqC83hyc/JwWdvk2Du9AiY2p
SIiRVHEEqapb/3WwuTIK8cHcbKXEeL+5j5OtlWUpZEp/BDRDQ6ZTkkYm7WIkHEkyVOpRWEUxbLB8
DT6Q9YNWatFIG62+dOX6Y0+yVZ00Doc+qtdhRviGXGsq7SkAxrIIrGge9tKvuPDXZCDhnBW2fmmx
MebaIpKlFmbg1ZHnW//WV07Cfx6ceX+0hN4NnsX5Ip39HRfXlwMzqvWpGZqnd4kOqZXQNZ12dtG/
SY4LIslV4AdyfDvote1cpm+ohWf92QthT83lJt0oh9Wo2oIjca2xBYMVjVenrUqXB5/dd7ZNzItX
WBuQcDsijavfHVcF9vVV9PC4Hp+Ur1uCBkftabHyiQgmVaoG7q/mLePLY2uMR6RBvXEm28YJ43+3
ku4VALU9VDH3U3hKanoqIZQJnNPorFYF0JJM98IfsNZUCIKpmTjPE/AcegDxaQBHaqNBG0HwPcCP
hWVncevx0wF0yhrPlLl3JZRVgKTH2/ox+xT44LtWvxt4PD2RhCNqWzwfOrJupmy2cal0kj5QTO5i
PJGdRfNqCFc4kjyAM57SxwKdju/t+1EAerI7JFKWVtKM/Oc9SggEt4HuwyCZmB/1Vgl0jdTQWEQn
5WLiO6D4FOLFQwQuXwZVd4KgfbTyrZUDarVETA9v0KfY2Qs9Jdz4BckoTYOPtlkNlAP/eJ5iuBo3
PhfYZES9FEDG+6Bl1b0kqY98He0B7Lw7NxGQugn+RV9bqwuEF1OfKiV9/dA+1fTK/QVidPzQUk+V
AIr8hlSUQBqHtmxke7Jzj6exIV6HvnTwX/fCuMbK+T2rx0g3Nw253b5CNqAI9ZLgutac8YB6E0WJ
pI2LaOs5b1PvalAfee4pe3ig/tEYU/vFeNGNzBzcmFdLwfKYMq1ZUitc0QgcohogRdvjeWgklIEA
vwl8/EJVHLGncAI/sgS/MSJHSI2OwJ/lOlvapPXRYrS4qIpExgBTEpx19HjH5WVJ94GPYCYxaRvs
hO2LkKtxFpX1qNho8XdAcIKI9haX9Asg4udaUnV6QK2A/5MrVepGrX5kZkGXv5KmPRzO34TEIFKj
pHjfJVMd2hvKObja4OnHdKCXd1bILo7mYiW4OjhNFuzWmEuk1XsDCW5kLhWSPuYampc0wSDrDWrV
k6KSuI/1fX21k8ExJddZwS26Qia3GL2NXW8+c6JPA1W6NWRg8vMgKftFYq/r8eITE5UbFLh5uMbH
/BNuc0uhSaTrzr0xLbt5EQVKIVGT0aXUfYwJ9N9hj6u7klfojqR9tjNwgOPn2xudcdYmJprJ1atB
4AxGd2R0ZBxHQE/AE9AZgZ9HjzQMdMnVixF9hupWt+SstDjKwathDf8OXzdZ2WEv4mW+zVtWGWqo
zGCa9neWyFCIYGwfNGAMOvrPvIkQ2Hue8d5MyPns5oxYoKK5wSNCHxXkoNI6kJXKFP04M+M+IeIA
Z/6M+WZisAwkr5xlZBqkr7e4J6oJga99ElG+sU0fNJwpPWIL7iZ/UrJBSxJ5+BGAFgkGO5QEerkn
zgNmoOH8CVrbMs5A3TJlLCCRU69kfsFhMQdHbDvJIIz7A2W33COI7XJ6+mH9wlIqFIIluyemN5og
CTnmTsBDIJOFoFGzDqkG6hYnFfy4uSTfGk3Q5/ln+TLiWuWabUrsXNMyEMupyu/CuDUT75fg0c4B
/Ixn6WejDTIhVvf34eIoMawgkABgUcI9u46b/Gth95qGjXxDxPD8HlpAqZyWEzXHKSiZivh4PDsK
0/1MTZu7k5aFX2y9fAhPiEniSgYEmRSiCs3Rzj71tPMY6eckma59Aq+alwvO29Q/I9bxjjqry5ln
C1qC6aTrZ1PORK8iCvHMgHMP6PxfLr0u1IP6I5DDNOa7kZ6ZsVtcBm1BWuy/Bxewp49dWF0CPkIj
0jwGfxGZ1IyNmiubJinmW7hh4X0FLkkFn+6wOfDACKWuxwGxNMygsX8I60Abi4ymRfS8syyXYrFn
y2OI3kSGA0E/bND+ZOHH5AcNdvJ1JEAqOn0IdYBguiYvBlte+7bM9I0M9pQLkkqVDEJljnVrvAAp
jqA5HV3FSN+MptzLHIdTIypRpvryBiA27BM33OgSKuGW1pBEH+deYUd7rjHm72xdKos3wKhcVvBc
lT8vBvotgyWGP+mDp/HSVwzRnDo9zaZS1r5oQ4s0Bv1LPDD3uWPGhHxeYGSekTz7M0f14UaZUZsp
r+gh1bWaZY38nwRT53PxJRChGwh2gMElOt/jBo9CGMysioSn4qoIMw9UAFJ6HGZkRAXLIcMVDGMY
n6o2ahgV5LMCTKXYe7Sgq+KMldK8yNj6Qc+bvFhHTWwsMn4z6Z4FgbYrbxn1JNxIOL0mCQY0VTzd
SH+px2P58P4AXNjlLjhSnCWN5j+GuViPQ1AdiwM0t635CbKjK5W5AwFNYZhhayrbHdFjeLFZCN7i
xb9UHvKkVV8AHA57bes2/pM4inEfEbbopeb5mnBCv1jExhsyFDpUHoF9nd2q816Ylj2tdwFpcl0Y
Ja11iBpmRTCKyPOKhXT2IOArzwCBFE8+VbqBFKcw0AlTIJAOI5hxfxePoBqtjSemz0TnaKCpuxph
2J8Yc2JmBIblHVWat8NanNj73oHv7Bvhf7o8srcrMwQhcraVT/DAKPrtwioTO5nslRIJIyI+YcIN
0A12XXe8s1pfrHoCEZ042TTHkeLdcOFwJ0/K7Ii9nFTXgSNXl9BrAQiqUjr+ExvdMtwz7e8xn7/t
oDXRm4tYEt0VV2u/q0FR+u8kEI/6JbqwNKCylZbBjLbeeRKzNDpG9KbAlxe388ruC2FQ64FzGnBA
caiZ9YP9FkY6PPSAmyf3kyayelTdr2QW9MV4NrdK6QaGM9tw7Vg//yvQYcInmiYySFIrtR09NGJQ
q/o/e/JhbjYHncbyAfHSHyOjxBEZTUOr/heQXYFXkwo4Au3LvN+JKLdjas6ppXG5BPoFFvH43tbh
HHAUy0JeGCYkv38QWfVPkmZ5qQnyivfTH4n5ilV8oK6dfEOq8H3xaO4hHAaLotmxKw/cOUYq+HtT
cLARXHOoBAL4kZelLXAs90v8YCH0BGizsDRZcCmXDbbzPmYX6gUhqiL2c4JrsgHptbxoyTg9O8LZ
XEeFoKj1JFIAEe7aRoF5m+vX5tOdspMRDkwKALylF31ojBXUtLSK8DtHdrY+TeWJ4g7f0kSHqOS0
gurKgROYukAktVtYzkO9s25Pe9NFT9Iw0sRjUf0NpWmc3xrSF6PQL1ge9CpMw0nvQRKJXQ9OABhQ
TNeGXjAokVz+AVfCDoxXCGCAJlgBIw60AaiNNGLPhU/XQcgwb7t2VuaIdEHYNcEOI8v+CkYGiskD
X+15U93SnLXRCc+aojFIm2vtJQnqnO66vH2gTMkesPQe/CkYsTwyxzSXGQlbEbpmFx8WBDVgd0Og
XmtrtLeOJ39foxxC9IINgBDe1QzAJze8bvOuvWNUSbgdFJzOIlbcldNXbezF65AKfMvSsQmPaTii
MS/DVy6q5ZCYl2UhFwt6SZNx6SBEhxI/S7Q8LC6VRRXYGakzOKMZxrJZV1OeMpTLCWqf/bfHzXu8
un0JVT3+bPU25+SKcKIUZchBTjc5wFiQVAOBJIBGL0kLtBrctPfBGM/YWInrKCym7PlwbUlfBine
AAZ6umtoltvw0rDz1ebztuxEoQQg3seCHrshasVyASyq9vVjGCPpL5j2E9r6ZIZtXnZKvrlrcQoP
ivV3gC8sLzIpVHQVieAxBuQTMeoxuogrH55RQ7+JoxhEk779/N0w4YNoKAf/V1yyEG1HM5NGHReT
H9VrTchQsEaiT7/mGbG+nLORIH9ewY0mdUAItBb0XHznE8jTM76HNYgW+n8AxNuVaayfiff9HiAz
V2ZPn49+rF1SzZ0ryYYd5PHlixofkzTt1xUGcAR9EtK2UZJIMCZGB+97g73KkFv1JZ2J+EIh6dxK
/VFL/Vn2PoFOZYnUm8zSG8Mqn6Zu/xZtDyQci7e2hdMP78at+hzXkyYusX9Z4bpBU3vNUO9ZAJaG
NKvcXGaXUOdrUc18fBkD5KnrEWSHpwWfCjzzQ/9whTwNZI6RTl8yc1V77nWdLe9GBrmdPskvP3FN
FIdEniHUarbTQJ7dW70KtUQluLcYI9fkXmOmXmBY28gk0FStBABrmHbtKgfCl5lQt9c29IpdEMn/
Jj7uUMiTmVuUQLzrMVYI1Rr+l0rRQ4mRzLqEBPFoS1RjESSALnKKP2hEADaolSpNVg87VqwlUcw3
v4b1SYD8vJWiFia6wUkMNkOXSTZytxw70+lPCf8UzvMee5QOI1gUPb2BBADrYVK7QDp3KR9iZOAO
P+8ixm9cX773SRwZ9cNpb6vXMH+y7DX1ReIUxqz9UvRAsNESDuL6xuUkbV/cppcHvKEpv/ea5vF+
nDnHBafkAIQDousghPB6NEn6hCEYJTQ+hs8IGtOnL/x1VjGokk5nuUjjl4rP32OJMfLOUQ0tklB0
oWph5kIVGDCDkrMSIloOrnJZLCqAdDYD9/xgH1zbvemongazwgglygVKDV69DwiYRCkiP+s6m8OQ
OFGoyzTe4UoOJd8RWNeJYs7pKpKqI5p5YkYkiA0338/9Acr1qEt4JRMaRqXoPIiptWDC3z9UXmKb
+l7JgyYOu3ZQNZRt3ESzZsfw7urxgOMkxU8r/Cfgq98dHfLyclL2Klo3TSUq315StxFS1T7/pzTB
84g7BkCD/NSJ4slbsJwVv2ao9wjAQzVb2pH7tXUo59t/IcjKdSmWltW054oH2B9MtWp/TPnxqOHg
xsVo1fnbMU3cH73WzCsXgLgozRB50r//v4nZ76wa1GOPC3FGtqV6bOE2mwQ/0Tx7F0+R1OSk/f8t
RXIC8NHOWvHNfhhxeMou9w4stEXIj7dtF2YDNeOFEujKPgEjUmUbdQMGypEP9RY4ZARrdqGMnlcH
OxLhVvaX7lfNXMURw4XFrza0ZkFEQHRAsge5CkRSGU8aCtnoavHPFA/SlzcKpTMICnnMX5WtcJFN
b2P3MBbW+8cdBulqsEC5mC3/RVNHpLS3qiok5yNgpYHdNro8qfYUMykC1BBvKUWX7n/oeqxMq7Gu
8qIzDlOc6X1NvSjWOJq3h9m2FlMzm+MPwfc4f9aC+UTY4gUm5ufLjZ3DpoMExPAzQ6yqeYMbRIOO
UJCIbyq8lBVAjgQYKaw7f3YjJjnrb3x/CUmKNUYfUp6fuSJAkvpyxEB5QgFf7dONrVroVT/4kAAF
e+oJT8xi3scdXRNUfhYRGT+EIYVGFFCVvxQF453ZTOOai8NfwfLfZ4qfOfEdsD+LvfcfCJnfXvEV
fjmTsb4u/GBGftnqCwQAX1Q5oHi3rLZ5SQH4TlBB2sSg3EdFQK+VzenKdyMv892rf4+jJTYouUno
XjTmEnZG+uZD+fywJ8cWwez6aNHIMtYPCsb/eKjefIDkUlpXe4oZIWwHUt4mwpWLrtaqW7oIumsY
KM7i8u5q1vxV2/ILZZ/geRejacMqOBTZNKeFS8frF3mAvGtrbnG4L1A0Z+FbG4UAE7DGV569Qaj7
iP/7nmsk+Nfp08PaRMFMlL/gnYmv6LlIlee94tWs64JLmIEHnju8k2BDQE74EwVsiLTyBL6gIHgZ
K+OH4n6NvyFIfLHF5Tbmebp5/6CYrGfveHA6VTUdWu1no/J4UqKaoL7yuvoF9myyk7jLh3J/eL3b
VBV5aSN57tLb6Ppx3qyncV+7wTcRNYIB80Vugboru5CBIKSd1VnOYNkQvpVrfOIA20O3c9ltCLGu
gHAP1zZ3Rjp/D6QRQtKzXrXYC3tErvF8Z7zD6YqA1KxdqEggG79gD3G8n7b2Lg+WVwcQwTrbzs12
rdY78Vmm2RXLrzKloNqsASrlnSiI9U90UEni0B5mBdm54cR+7qe7x/PMomGb43CDHGM4mo7Pgg4v
MXdPw5BrRbnW4yjMMS+8DDadVzGjzyY6+sKqCvfzIrtVFc+ygTRdQwf1XmchEINKzfhvg2r8xR3m
I5XfKkLR0NS6aqJMQKSXk47hMIY/YLUeeQZV1j6AWln5PvH7RyFT0fIvqrgduDOIAij/fYjtrn11
FHugyR0d0b3O1Fq+PqGGegnOPb1tkiJ61MEcVO0NAtEIJ8pLxyKVk8W6HQJirkH/Cb8ZnCRiuz4p
d9YVeSi9QrR1MirvUGFN1qnyUWUkFrvB5fSCSN2tIc/iSqg5E+Ab5BQ2mQ+gVIAy8zJps1lp7AaP
O3XJAslbuj2HWb5xzdwpS0UJ0PL3FahleMqM5FFiJ4ywAvdoj1EzRBIn4HNAYXCgNbmk1PN2TVbv
LzZXlyINUiIiU08953a9LD05OtKkh7Z8CyDvV6vICLfA/KhlKq/JD6OxVI0rxOPiKYG1/YBN6GL2
fn55FZukThPlaT6TQzHUTMDMuBWs2VWQaNQeq2tdmRAMrNKwe+MdG2mqwism8Akruz3XqKb0gMBN
uTSghDYaDjK85CIZ5zAAZmUDpI1NhOl/hRhQ7c/2pFecc/+eockJ2qXgLbfdBHEuFbOvACL6coDR
+9UyXNcZUKrvVcg7XG6FgCM/kWs7DEEgqN51cwopG70rN3Z5ellzdo5Sc/4PSvJMAN94Nlej+NlT
vAQNXY4/M4DuiMZyVFCKWnJ5yFKt99c3D+aGxY69cqLZU8Wk15NJjUOg6HNznzYXA69wNNeFfxer
vzBC8lSnwbdc7+OF4uwok2YlqjHF68QRM4En0q8SWwSNYifjW3A8vVn8B9KgQRzN9IbLAskoLsE1
ehsZMgBq6uXmfrCQdSVFsS/h0d/vbI+HaAjSAR1N3b3rSZXe55Ft+aAHFOvOCnaaEfwZSCSx0Kxa
BMoPhqxXnbgKKovv2qYYvX9sj/ImbW7F2vjOZgTE6/Nd77EBp7Gin+iK6XZx8XznohyrJl5WyLHm
+v1lMGMxmvvt2S3Rn/07RqRk226e3ubGkLDlrbc6G9Ai6tZ/9bp1AE2Twf7QWfL+sDvwzC6TH4og
Wf4ZZWeJfC1hqBgeTQM3/phOFf3DdLQMut1SqAkAK30MR40GiCDPbyqVe6EbF0tEAn0dGhAJcYkJ
RyrzDIJM7mE4R4MgDowx41Xo8jaOdzOya0AaNoDpQ4BBoTpkNWf61cvFC2gSTIrYzAJHvwunjvmj
kUrRidiIwESC7vOsxUTL+JB3ugGqpfcCxBI1PoinklpZkAtNp1UXQQpXYLdDra6PO7IaOLcKzBcw
JaUCJSvDWL9P8Fq90FwTcJlv5oELJCxc3t9k84YqK6MBoCuYm4piej2kyI4O/Cgm0vmiP5uIpSUQ
H2qyVFJBXH3qJ7A4BnLQvw7TNlGOqInZd0lmGf6ty0fOvN0tl0GwlneaqO75Ys9byD6t9tp/N8gU
merJ3rFOVMYUdH4HD/XqYyYjCiRwnBFTdyqhzhs51ZmEcJgMo0vqJPpf5qFKC3WllP4gZZCtvqiQ
BKns9MVAK5o3PBNM15YYOL0iDpzLkFcRUgrl8kWCcNsZSMKvm0FZzROS7FnQwdT1UTLdj9sYkixy
YOOj+p75s00Emq1SlieUM2VG/l5eAVD4u2qpMxb6+tSDhkjtOhtVP4qgRbujtgVHJqQLdwLZUJoM
z+zF3GPGhAVpsHeiuVvEW1P5tZQR3QNjdSIx5Xo2jdyRURHBv5eXd/vgsFo0/7tjr0yx1Owwe7ZR
H7dY7P1BDCFHEPte+04UKVZj6BJ+Tw+AmTqloFxJpOmzmoc3j/dOQCsrYSEl31jjWNeYwOJcarpT
YK+FUkiuV/qeF12hFEKQ3+KkZ/cJvNxvi1Z6NpmEZBhOprWN3NfcNIIJTpSCT1fPvOq4vop1ec9V
WIabSoJzo9BHvJr1WGOOUo9F4vY/Q//RFH9EdYTxCxPimJm1winTXOyYtiuXqq1xLi7tzprJrukw
kseFuXVGOZ2qrVIhCPtti8si/QQrJAkRMM7r/GSe01NYsYhRgr400hejeoBNDbm1h5ClYcWvV/ge
sG3InPef9uvgAGkrpkyyxt0kqy2qNsjd1r1VWmBWJmxzWjsD6x9sRKGWZpIRHgbhpD0cJJl+w2Fo
obUbj4z1nI7ank/90/sfcC/5H1QVhOmCza/v91Bfwak7CYYlPf5XL2IUh3YDAY+0Pz55hCbSKQGq
NW3cYEvFhfN34lgXhabeekC2M+dykriqIjw29Ox8utVAuHaoZJ/9+cJU0Jq/lcw7XRs8/CfGgLN/
tdUsTa1d5AdTqrvuBVNZ7209oBiZLZ+++L7/90WAQEzYN2pRUWAPyNU7IOJKkgiGmQmYnVp3T1ng
lKO76CH5U43SPizhOEIog7trCVHQskrpAUGdaGiZ1x4IgS4aDzmHAOq+ygFh7kqneqSipaxS65p9
+JmDEwmrw4vhgt4qetTpuBTI/9zMAvWkBT8aTRwJ5QXKPH20tnrpnhtvxjPTPCL6ilqi5DHd+7+l
AaV0E/+0NG653rUt/CPKWwjcHuGc5fnUvuvPL6Il1M19b4e9ddNIxmGibn/tffoQd5nuLwyCSmvs
H62efk2wIEsmDspL6jyT1MjPelJNjM0KGtjevrbDiFyRUXjObovJfxiZ+TaAuwKyX7IC4Efchq5b
SDueIglqEB4LrGl06V/MXfGeXYuWwAjphvbLzy5HICnSTECHPI2Qx4OKdym+F3/lgn/jo6W+7jq5
y620FPMAMNWP8+mABTmiYEH3NzDVum5TSn8YCtv2wVrUgSb6SIphwygi1hr81vJj4FnaVLR5r1V3
6wveaNHLTF6W13+bWRcOVjAP/N9njGjkUNSZqJ+hzTWiuZqfBCCSFBydbA1IE4Cp6Xyw72x91kdg
gZS/zYdLzUvngyQH7YTySf2Q2U3KR6WCIokUF7/E+lebgf35HO9tzrjQc/0C77DtptK/TZmSFtCt
htEw09cuqJQ3GbdjICHH95rdjZeqDiyb0MWXGhgfay+BwUtwwFyps5SK3BT1yMzA0GSgHMmXd8cS
xC+YYaECGXb9GdMea3G0tuTYYnba1SoK4lBvO3yhC6ENA2cH2rwjAV9Ii7Brom2pEgKA4K8WAGaP
yLofacyN7jmLSYHQCHvhXAFOOIlrA94oixJhIYHVBWus0kf3JWiRe+411/DsFlQHz7nUpiymbdx/
VA7l8vT58omDeizsxX5lXAAb416pLfV2yICdbuuRcOnIJTPB+MWPyspjEYbw3gXYpzHQm/B4IsrF
hmYNc/my5YYXkQ/vAcTZ+yJujkYn4FDa5l8eRDG3kmVHCF90WjvgTHmxeqFKYvwDCANTVaRrCKV0
SXvmR8QKpDSDgF/qjyRgEyy2j7AUxqeZyAf+AE8Xst+JscCewwIfY/zyEgDy4zWdXz7Rw11RJ80B
nkkJmzUhFjLneGVN/RQSN6Pm5O6GrdFiIQJl5XkkIuiPf8xLxf7cRfMwxlwzWjKBA5Dvxk/mfPJQ
mjZvLOpajrE2s6/qNs2VuSU+WK18OaIvpPJPBE1AoPSWd6Chx1+6UwrtCOByZntFQfLjOa36Hfh2
MARnjfkNu/FEZyWD6sW0lwhZuFf23E+UdUDdB6X4Sgp/hK3tCRawLT1Z8VWWuJd7/7sH+U/EUs7R
bah0BVRt02WL+tuVf0PeczAgALuS9Ik/nWC2Y/KcEkLlWzpAVLnDZlcBS8+KMVxINEo2E8t+qdqi
wBUG6frPr+s3UQALNfRq1b56v3Vs2+mJc3IHJzl8zjHtaaLvT21dZWvXAPF6jkX1YZsm04uxYQxE
QCYY2K9a3fXtR5+6sD9qXuBQxU7HMgqgXwDy9wCoQDTXh4NoTLKff3aAAD/tuKMFWeNHLM20+wv7
elLCEMDVIpAZgKXcxU0jbdbF36lr6BABVkMbSQ+cLq+aK2PFxths/LvYbAlj4NuMayFgd8b52k8F
SnELc7xt3dbfxPyWv7k5EPn92D3AW5L8XoWbyb0t7nDHxiL+Cikp9I7uxUl1mHDg06Pv7L9pZKpc
cbky+PBn8jHkSgT2EymdUB4CHgO2J56ge7lcRbVdLyLkwjNQsOFT95M89ymIrvFNsIx+KAelF5Vv
40kC2or9v9ukAe+KKYVySsn3LZYieWwK5VSVvTaSRoftOw9RVWB7sdjq0haaRzta8YfySIc1lnZX
ENkrpK8u1q2XpDvuygnfnw1eW+c1n8R7y3pHV4oVaP2EzTtDCVFeVjxIscw2j6srHUU2ch9n1vjm
3P9fv0mQwjIBfaoalLQeK4N0fJXBPRmZwfvgn9JVwtOTBRTvcBgM/ll7rnikvwoDlSbcQRxVs/wG
W3qLmMj/s75pi/RnW2P/vh9BADfsF8yTjSVguQm7JC/Q50RcKY7GnheIQthkDPZ7crRfe7dqy2MF
zjj/OOLp5r7Gq0wC1EiOE3wOS4lkbdn6U/7Jbz3qZ1JhVw4Fw31iMNARGOqgXV7IleWnhOw367CB
Ltji3hcNyp7AzLsSNpwVwPIj81GUz089srR576CXJJ62Y8nqcPaudqFxCgnikvctiuIqBSDQNl5T
LxMVHPUhnkyAT1Crcp7QDrpv+PPsdHOuvQAv81Vd/aOwDv93wgOzhU6pnWnb4WtTikomBitLvrzZ
8o+QZCz3vyuFw/YCjWyRUd6P2lNT3sVF53QwV0psPlBhVI/ChTI88smjgqRJjAlUGCPJ5PxWV/Vj
hQrGeagGCnkucSZxiuH47Bp8uxwksQEyPlqx66FhIIUZni6asb5zpXeWKI/ErSU4OrGWjEa4xuH/
4YvFCRscHFdfPbZAL74LLfIDkaJ0ZwhOHjO7NT9gwLT3Rcm8WHyuewVRKHy679TP9vzg/mN8V5sC
MbRysw9qrAGDiDq67QB0AFNjapnmcyviIO8+7GUojT7unzIzUaM1jc0dj24UJK4RrhfLs6oSn8ma
3w2d5AbVgeEi8YFo7C6zzgCFR73lMyF+eRGEtStQO0gdcp3PEbXHXF2U5cdwhqIyWlexc0EoksyN
h8D9dd4w2W5UUxssX6X7Jk1QUJouFRDHQn2TCiZRkPaB39bZ7ttQ9qNSeKxTqMkSUPCk3iB1gMpU
2YQPtLvRR1uDepWgPzV3Jg4AewnGgCN8U+gcoliN5vlBdRnQLFCuTaQMaqO+/QIbOIvYACqBNvDg
qo6dHDpzogJrHdlQZ7kSJsCe79Rr8r/CK1+UelQQfcxQ5Pj6G7O9n5hweMBlMDLYHZPKofG1C/Mk
JQluXvhgjcCqMxgo3pW/M9VQFaLnMGnTmcSlk05sVcT1lnuyb3d+QmrRr9UQkXLiC5LHvXXh+JCj
ClF2t0cWDR2nz//+ih17+riWvvEDFpJE2niH7N8lPqh56cZvzych5IG1eYSCYRUluH5G9BKzO1hi
fUntN+dVRKzb+vLqdPOCwP1iRzDWN6BmB3nUc8vl4XJl5MW7MuiakLbvzpA1x4v3K+aC8zBL0rXi
1SeFvNQma5yhUf9QvMEMIKI3Sk6XL4XKUiAfEF+zJSaBR39AqpeFJfKsM1oVQehT9kh9NBKbWWDE
fylcfyPKV9XOl8x1ABbemCCGMjxguUC+DHSQvs3jNVu7sUjK1jcDHAKceygz3f8MrMsJo+mBuoWh
AfCUYNlw2H8krQQeZaBkUrBDkUpJiIpvU/rq5M+ZkoD2SbyW+WfvSjB0M+0MyBXnurXEF75gb7yR
jPPQaIhP/xFc1cVhlnx4kSV4Kz9f+7ElRuvuMERvBrH2ow6fR0hzgPTkFd7x7Pq53mewVC4JuzIz
EHRxgOhKXXb24aWhmR5OM6OdrfX2E/VkoGLVEnododdIhwWUxJAsvXQ5nQyoc8eT1javTAqnGD+D
ik7np186Oy29xo9MjQev/qGvhekRfaAkiFtz/qTdg1V5NcDF8TsNIooCj8/pBQvfTqmqWz77Dpzp
BNFA+PIsy6hpoU69V7AB06wT2EXupuLwk+kY1iC2n9jSIUQrteAFnArRzTjaL22ix+rjd6onmG6H
ZSZEDs8XrfO7CGNLQH608UpuCziUNq690MA/XC78kXhmBXkhn7zza4oNEwSi65BzA1kIjUeK+Xv5
bWhFzKXZ2fyifel2bPcm/Iir30hcePetCDwAnBF7rhBkYi1EksalpEtY9rnkdCOfLf9pp11rUeIA
L6DOx17lsIefbIycSy4Pd8fO3IMamLmImZm1pVErhaqdRI0sh3+e7lkCzrOC/qZIrBGM/BI6QyJU
dj9CW5g2wTZwWdM0IlBFjpW4o9k6qx+g0sVbAG8BDUxVuegoT+EcHF24b/drbLcReLvZL8+JtIf2
S3MNUAyYtCy3ysos30sqnVkstKCyE7HD1/uPz+bD8bT0P79w2gMDXZiKQ9Wjw8+rgwtmcPXKIxH3
PJJ2s+eNGHTlu86QwIuO4ZxJ78vhaViw+FalY5SHoL6lSkYqMsM/Z2iLyFMzM6WiQbicGLivJLne
LUEqbP864KOdiplMzQbpO/NF3G9+jKQep99YmvUUWOB8MQn8Ka3KsOw94O/etLCx1W//7UKoCt9g
f9MTQy85jr/EHZfotNptrbVBYyqHKmw6vCcpoLXcYsWYv8YTggRcNuVMDLbHcMT2wEbxcoDzK81C
OXzAlcAKOXwKpLTRULdUVLzfHphw6p0Q5QjeDf8BM/5b5hZihqkzB2G0ettgLNaVodrVJrHXhKWw
OX439PctsPWNE+DigRdBLVGUa2NcGMHCZOp2D4h3iBDZ6N7Gmk+nyLcDQY1TLo8kpeq+GJuvYWA7
zqW7aVWIrYIgaKe+S8U3dWZRV6/7UeYeKmeEx7WOEDbFKBX55tiEGQhpJAFHho+TulZe7461nXQ8
khihfs9pCDK902Q556G2Kx4308sLVIw9KwID1WEbuLEGNCR46Ri5AFsspnZMrNgpHwcVqZ6EWrOh
AyLHV1+pe7LgTiY/aoHAY17yJlehOPWFMlA7xcU6BWvjDlYsWjLspY4dacpCYxVTKoFqNhrlY5Xv
CQ3zwsB9z/Z8hx3YZmci1hkKc2CXAkcizc22CLfWpFSv3K3QEpvsBqSEKl0l01IaPGmgNhR2YezO
F3oEwWcU+X6regl9iT7vTz54UMGejSw9LMz4yiENsr7FEFk6L5ZGnuiTWipPiZWk2MdSflIR74fw
h+r9RrB8jenMDmPLIzIq7rq1kbkQj3U0W4S++tY+RSCnwZC5QnRH7X+tulu+KzaJNYgcsWFrZfdM
C82rhFtSauKuIQuSSvXf1KNO2fRrjrCghwRTzS/QWHEjnbeDUhkqTVg5und06xRZbOwE4jmtFS/g
wyuYmW+LBXUb1ZlIt5nowSKlRm87MEBwGQ8uaYJm1jz0aR98pTjnoGaMm/3F2AMduuS2eYu7IgEs
xsgZwOCuzniwtWPVc/3Fs2wTU5HbBM1ncw0OylY7Ydw2cyZt0P6zjBYOrDTC9tO87x4QM9hPm5o4
uc36bLqw7Cbl7x39bWeIAjd+SA/8oi5mC/lCOTw5GJ7L+7HF9E1nEn58fILbMciJ8o9iuFylIfv9
2RvU3NpR7sqA7iuTF5MgDjd1cUgWBrHGkLdqlFtllF1vYHbzbW5SBiJrZck696WUTkOmFGLJ1B2D
VSUKkTsy+Lp7qpFGEV4BN8hBdor/6Td8/O/CSSImtqJlZ4vF/Mo097fywI64eZH9sD9mP+3YgHtb
o3NnLbBP+fubRejrTl7fesieIG6Q+OBRvVDYoVd41Wjh3kAyXRfVqwg4coW8NefPWaHLhDgtGzKr
swM97KwB8qepIgbQA8pJ+ooWfQmTQ2HSKMmaPqNB3JMa2icnjRYv7TO40ztR0V8lkSS94DSzt/MH
SK+1n4bFVX5G2NCkQZvbItyHNlC4kLtDHW+Dk4HDwFvvUhgClWVl9NcoJsr+W6TFq11h3HDq8Cjo
rzBgHAzzUIAs3UoMF2fdmMpv6JNmav8MBcxZ/i2ygLL109mIe+gWj4qT/YWzoSLDA8IW3C83vS3Y
CW+jFUFzCG6zzkIGCKDUm92/M4ko/CtQa2rXucpw5lSrspzXw+qUB/Zr1leAnWceuXkt+mCFXbxr
kYNUdaFoTaqnsJV0y+DiPm1Qq7JyFuw4dpV6bi/09CIbSoD9abmLp3wSD6XtYnzx88Qwno8XZVfh
Oac+5syjytkEJ6FV3gbpEt//wh2YQr87zACXy++zb4vBld+Qjt2EGh/tVCF2a/rucHnCzb0M+cFA
Z3FAIDa68Vfl7cDL01Y0MftUgNt5nClsaK/IyVNBydovcw3SGxFMBjo5sYCpNtCgJNouadsP06tq
AalzL30I+NARwAi0ym4TAWHH3GTolUK/xsuW0o9drpgDimDzyXv/kKnp8YcK7EbpsDyvZUEki0Ug
XFO7fy1238wSxUwEiGQExnDiNYjcARkvKAhSbytyejmU7lNGCkCn6BaEn4BkUU/zec8ivw67WfT5
pxWPhHNQsOQGaKW5IzSLLJdXfk6zFndYd9ptVulXIOoYalFBkyaRFnRXtANsT/JY3+VGSC+DcJqV
YdaU4rUD/3WeHKTqWeJpVXhuE4Z+gPQ0GeTcMcvyj7pV2dt2vMW+3LCbhcGGuJ1esDA6kFHBRQNw
Js7JFsrGdpgiOQvshNBBBbBdnOl4MJGPjCOns1W8rLa8btgFG0d5AXbARGq/CerAJ87fDpgD//yS
bBagviM5z62+a8cYO6XELpPJJIBEsPK8S5nSf1pDVpwHLPscWe1Pd3ZZCs5jCfn7XbqhWZJ9IuoT
sTLy2UXCSCIBcUe+XOh87JufZ0pXsqYnJ9TKpsT7/x6IMfGkrDSte3isqM4cjmt4x6ygELPoLUTU
M2og7BsHL/vtOeldgwTkPHRWbjkl2g5NIcaGsolAAHRDBFcgHn2cjym5w/6sw7gpC6vddw4SSwv8
RjR+wdw5MB0NS6kXjl0T9Qil6UuVws/+valoI4B7gnou0m5XfUkh8fHPDQYyM52FuvZKnDCZTIsa
ufDJo+D+Cu3rZxivxUBVMuCUfc2byKFkj9jMkLq2Y5G2snlvb80XPlVLtWkm774KWeokfyr3AmtA
UkO5LIEUgfexily5aOVz0RqnVHKvcHaWXahMqKA2SpNdUTBr/QjoxwRi2ael7f7A/hkfidimaGca
byWNUP4PnQ3t11kaApfxwZcjCCiyUHZqwbFVM/olXdoehuH51TXagjpjCV4DcLwomILIRYFpMELl
BEJKfN2+ma6WmLSXLecjvXk76iwPbDPXtJ+CnzXnr5KWfbZ1DACmYxh8z4LU+s3g249mb6t8LN9V
GuUAKaw2uB83/t44ePub46wHIWpEg5tfg6IXqvotcMmmXDLe5ToTofY61PykYh7I24lU06/He2dB
8soZmvsJu63snt6BC+gKtoESAfxxzS0hrB+akgsi0iOzz/fVFOPuGNUwhCbUlaRm8N8hgkNn/M4G
+IyZHWF5kidlkJKpGRXvd8DhxXIhb2jQGSdMgwmP+6tqVBI0FZORSQ24io0FTjGtNFzm7Di45zmE
JgCts4TbGcMw9pE3fsGg9F6YR1pg/Xw7iofZpRZMbadrChhCoUrNEJQh/w49xM0tm1FAwRRrYKyR
ci2nOdstZSs7hC9Mdgxy/Ji8sCsR2MYZMOQZF4fJP3FQ1fbJOQ/zrBvcnCfymrYLTSzsnQ0QbwWS
pwcTTB2cSUd6toDCtaXHGlBg3fAu5DJvEljLJ1TQQbr/Z/l7ANs4mK9Ifd7mq9f2Klk+aY4NtsFq
PCof5i03DZA9uIw6tq2yhuC8qyQrBnY8ktaFF4Dd3PkWfxya/Jp7L+rIeBR9UTwzrrJhWbUJgACi
CEy0DBQ5SEgl5XEHWGZ/phwtaXYhE29zM3PT0P1xzr5sZgCUWiMmAxnkJLVQTS7RFLKNqP0rRAfL
CuZ/lhBj+2kSXvoRcMaMmnEGW3dqVb8pwANcbZKuIgyGxrKnjn6UcZFqgtgiR6eLIsBrNTqCi3jB
G4UgK1zECoL8PrZMfTDONZD9zd3/nJCl7nzy520Ibyk+dFXfZ31UNXl7guP6fW5H5ql5og/y1pFL
zCfp74t+MXpsZAkxMvu6M3Uc+Bb77wAyn5DAvC/OLB3389VMXsveAQ7yi1lSSTRNhZlIn9vLWI6Q
TaO8BlQD3Py2f92mBk3bv4wJk+SAAiQFWSwSnJlWcs88Zc9T3d+iatYAcm1IYG+dmEd31JG8Ivu6
bNV7yUr3b2FQB3+V+jHwy8B9pH2BAMAZ/bSLpumbm05DR4p+nJ99z/t/IYBHo7G3bFp6K3DyWwkp
oNSG28jJcaHaZzv8Qs4liZPTtNm+mHMdxqEn7hOJJOVGMVJQUPwPB2TCRZ9bXVq0BYY+W48yCI91
u0cr2VE9g2HaeYPEZn1i/7hSxe5GxPK0qRXgmoEqR8ehDoDysaTavYqbdWPc1GB9NLho3oY0WKL/
USoB8W4xwBgYx6kNJzB3eufDX9mr4uYwidnS4ZQCkRxpmMj73gJrWELWRKcmeILyK89kfVKp+Na6
ELWNKS1ufoX0uXm+2+mDh2X3yynCZ0B9OkRwUpSJyCHrgqusYS9/pFScOoexopVgV3oWOwBxh9bb
z7dRFYHXkTMo3MpAFMdyAwnbc/33WR+fVChbTsXNW7Q48kjfWwijv6daKWrjbOizrS/Ng+OKXfKH
gywoe5M508HNBzx9OYIs382JBAFyYSM2h3lCUkNS/4YY73RVSzaExz10jsglZlpBHxSB72z23uN+
urFpQUoF1OEDnKcwg0IdccPQitmeeAKhKdh+akcX2d47XRJfkJFfMdHcEZsQ3ifjWCEIYc2xFms7
9X8N53a5mSlHzAFCXQULv0us4U0Qa3TmUK4ATjpVf0KxLsOr9MK5WhANXSmtw5ntzZq9K3a4w+ey
yPsng2jKM5dec4AewFENH8OyJ4g9PNIziLubZZD2aF2LavuHNkPFcSSM+mPEpUdbyHMQjKfELnA+
YJUvNy6IOGhVwO64HZTE3bV6VjNZidACWYSn5u+gdu0VUk9LqDj/6UmrJmUeWeePoVeiV52J8TbU
19v8Tf9GtN/mcJy3ItWBQAev7RBmC60rz+NL2d3jMnnJyPK9HPi2UxWXge+Lq/wLRaJ1T0rRoqSb
bBUTmz++Hf3fl2nxDFgLKXfVh4s70yl2CVnr6HnNr2agQOYpoq8fMfHbyp/F/+0CHPaLx5yGpJCb
RCrgPB/ru0s7InMpKNOGVnH/hxPGD3Vlf4+xndlihynTeTd0GbxEOeU63cCCLcY9DxRYHf0mBnn7
635/dkxsqlBy0mk5BkAlmkUum1l1t/YjEUGHOebUTH+wiFjyY1BQ2X6uDttllfDF0Lby9sRfWgdI
B2gq1czy5zEP8sbbpI0d8We+mqF/JFhR62YrqKN3yn+G78BjwC4+5t/IP6I0Cou8AnXzoHQDz5+/
axCw7W4NTkivWoOYeqyVpaE2robcO+ZdmCut+EsIG5W/6Ijr6tL/mjHNtug0fMoB9Z4PlOool5rA
eNlnPJ3RRuuvQEAXfjo41QvRR/U8UyPmaAe6fOG7gbCBLT2uGm2EGoi/tUVOlc7tq06J4muSyR5A
PL2mkkR9pSrTFcjgRHrpykegyfXmjraElENyv0fj2Ms2VGDmJC0r7Q3ZNoPVHdJcOzs2LqfokmsT
eR4jjzmn22nzSvwAPRJgsEw+PfcQ0SNKLkeLtXuHvu+QDPE+N3CC6nbKTCVj909dgaL+CYKMMO90
Wh2kvbPfwVuL6nwme15FlVU/zWc13Bi8Gum5PuEpCkCUlvuyk0LbTOq+RNwXflnFosC4o2mURC7W
WQc/GQBBcNofTIv5RjY3zY3nYzXl4j9hAs6AYTfL3v6IfA+P/V9zp++6oUfBQUrqDQWTb6j4jPnW
d/1+M5Zugv0/mLecFb0beTp+n3zdIby0rkzIdMIB1re9cwhLRwR/btlI/p8tbg7pI+EvnpSK1V9n
olK6LokUSr9Z34bSuspWm/EGmDMsvcn34S5UvBHEsM5uzyZUblBZrAaQXmT3q01Oq8Y8CCNGlWuy
Q1Odphazgem7rrFDRk7h6Lp7fk4gjHuvP7nrb/S9bwYAFVikpL9KBLeQ6jw4nXqnryKD1L7IYxGr
wPm93MePr03MsxE81c38Kpp82SaNO7eo6wsrx4g186Gef8DwIbKOFVg+3ZP3n1yqYk82fS/RMjlD
fKupe5tjPhhS4xJlovrDuFcfCy8gtHwrHhWL7e/EK8v53ntOaPGKQx2qZl3zrtTLALbYXfht2uVp
+LQGKgiM1KrtAZ2R7rbK6fHh2I10aEI5ElugyLRndP7tngBOMS1Gn58miWXN2R6a5YZCKIPZDyg+
M3MeRycJPxcn0YmpsM+CumFm5qTJ1qHxq8YB1CXDVpExa4gZvSin1t02IRzM+rLGun81gQ5YRBeX
4mEgbnXslovMoa9cOT/b/kx1419O/I/U22WdphCXyeTJRbCMcvrqvwxTe76OBq+6RXYFnwd9l2o4
FcRnlyqP8jmQREe6SkI9QiQV42PRE5cQURQHMktp28rSnQ6Mjwag+FZP79DzrHQEvbwijULh/naS
BFr7sNVoutHUwlSMWJwKAtdqEoAV3tin3+/o0wvcCSFtmsQYF9pzv1QpiZObKpySMIsbYyiKO0r9
61i8gbVS9v11Ives/UyhyToVzYH7bEFFp7KNMH+7JJCeU/b0umnICmRlWLeZVLHgJnbnCsIdWEXt
+tJp9L0YwYBWHpOGIUgAysxeJtER3JVaiDGKWoGkbtkmOGo1SWMKqWl0b8g009ZMrF6yy59VVT52
07tMG3TgPXiUIFwZTzJybFX8jKlD6R69z9ffaDpH8A2OXY+7ZDkY4mhhIqK6SRU9Y/ZBYoq7b2kh
e3G7RvV9yvZbKDuUQYAzsbrdUBeR588lK4ENzZioDDUPgu4O2fgAME80rnvCKS2NjOSGiB/Spowq
bUGDvYAxFJnA2jcn88OTxStcKv54ZIp9rjPy0XI4SlSV1/3Cg8DUVtB0McN1lwJKNNB4JVv+LLLv
RWlegZlhEkefNJc4FuyIOlHZHirJX1sk0kPhGkZCqpjsH8xEe5X7dugo+np4rVmMwE2eEej11SS5
d34tPKLBYjHE+nzXP4VTZh12RHdLvHOz8OphYI7H0V0x1emFRxtx9H4czBWTNkza9Its0QlguylX
TMt7eiNeY12qGZV7ya5YpLxjDBgj+cD0Omj5OJlcqbJSpCuoBCUyE7Kxv05HwLtcAQ5T1PQDzR1+
vTWy+KlDEI8UhJFdpKK08yCUbMA72M0tr69ErzJcq/Eg8JmicfTcxYm1Bi7YyuFyPlmLNIt8IJW0
Y1fEuENpxEVb8erQg9cEmIzb5U0AMWyOHrjuEyRjBuZJ3O5lG2MIWtx2QBRCau8H9U90LsJJheAK
YNyDq8FVqpUHV1TFDYyFqWSBML78XBJS6sXC/oWc1UDa8Ds32N57tGm+nTpa4NSmqyirfNCJRDkN
YCnIGP5cTrN4aALwXX90PEMeE/nMKUuX+V3IwTIDp7KkxBHW3ysLe89iQdrAh1hOptmgytPD2zSq
8AFdOJY3ifasyPtMSNWoYPlVY4AKm15CRDoZ3MKsrrSq9RvWta6C0vpOTygHoGy/EH89xIeXKw8j
q56O29Ivv82WlTZki8/ve4545UHQrU0GR7o5Z/q9SAzoXq0/Qjp7LHEYv+m0T63hWVIR+lHqQN7e
Q9ONzCr4yPJq7UT/1U3NhTl3G/nZtxC10XMUjvpA4PnsXZK/YskWMoHcAugN8MLiKde1mN8k1igG
PcKcPDmEl4ZzFDj65S3oOY7yYOGSyfm9+uhgIQxTP55+DEaA+YHzXVpud4rxPpsCKrFHI2XwQrid
Nc2KDLDeYRD17IkksLJe6P21gLdYQZPVE1y/TkkHpe8t0sQMUNYqsOEYMrYKeyEdJHSQeLZ+1bBk
YIOP3BCl2EO53aQQAArAwp8mx0TOELcZPz+QNHCkuHtU8DZcquG/lGLafHQjqbWcBb9YPSYnuHlM
3qR2c0w78+7MWPWrjSRwKjJoB+qyrVcnk9YtKZpevQDmwFmrJUPh0YvNW8dw+X+Xiq7jsIMNaAEX
KjUH8IQZG2XJFW8JavmaXYriteECuqKtC/G2jZqjNGQuzrt23bMJGr1h4iz2Mq5ZGRah1tvefWo1
Kg//mmIH29EjzTOFUnngB7jvldf6cDU0dtQKZkbfUCyOyONXZhguDicPP2Yank2QTa0B10t8u9dD
BsFF1bHebcNo3kquPXwiQNIWNLZ/iEYUqSlujRiaoYByJXv7zTg/xIACWSjTkzz8x2WxjWmLPVVm
7LMmQRtgQsPcVKBIk9Qd6yzxTd6ngvmkXMJL5G0lkl9o04lAJv9BYbJDP5m0FcpesYTY2RHJQxwO
nSoJqPBcCphONM7gKY5YOhWPMPz/6EQ4Gm2YshkomG5ajhDYulyH0s0zcq3YBriX1PPqLR8DTZgf
vv8Gril/HgsxCHR1+JhpFsp9H2abZ1BBNYljE+v4rXxdeDo2MoRUkgACj5BfNGKyDZ2HZ0xob20y
youAwpvYrUJFWTCUs5zVSlicwrJuYuRclBbLEaj5YyfRmAV7WyekUwHod8RR62eKgOFFwcl0uTs7
tZ0UnMBe14aT7pktuqKHZwPmEuRHfnfz9r/BeWtXqjGZOi3oewtGIpqwusieT8IrCV8P2tHI8MZk
T6ax740JadcWPXdpn2mIpF72hTxpmj9KmfuLOYqIHsXOoN7U537YGSApk5kedbc7tVzzi5ceLgXH
68Fuu78Ql6R1MUT+iVjns2dIASrPqWKI46LPu7eCzmM8sv8DAjRUBIO6nque+2AWOTcb8XtZfLQp
WfTdXO3+8X7VcgU51xsxU27T7WP+xZmwdiskj0DY0njulN+2Xzj2ew72/UdSZhYbhfBiDaWocSUu
Jlc0GDS6FtiRemzkeqllLDjZBgnWAS4iVeieLMLD0L4wN4R+nP8NdA/2ZOD6HXykWOwost9gb36d
cZSR5bGb9PNluX6BHRgWlEhLU9tBV4AewLHpmD4wMquhj1PwPgmg78+givrDkdfVD1cacZZ/CBob
Rp14KMpu/Bs5AemSWE/t0i1BQWfRsZVczwaz21nVU6s1GL2uZocVkF7kBf+iw70u/lWdQ+c67Rz6
ptcp/or8Dn9OxTG/nrZ75aemf5GS/G+8RRvyeePRb8L17uvxCd6Ka58mkNsM20JT3xNK1ynTFgWd
Ot3d41WMnQ48yt+XNnVndiUatwawYOPkiVIBYbkxP8lGG4cwdWwzxUDqLUyu5F2IlbV3a8uQd2u4
Tqn0SRQEWl+gKPIVikdKfPSASne6cgH8y7S59IiBxelYhR2XoDyegSJ5VrO3e+dr3Jt1RqDa/jJK
aO1eqfP+zrU4195JHCHLTEbdX/dstarD8sKmbCs7BpMcqBgBbYwB5+lSfYoNrnReJNBoVBKjY/7H
QFHOWmyoeqF0lgsy9yhcEG7uuE3QpPT8DymVOC8f1kscPyO0dYtVtKzF1ql1NiWczf6NCesuNYTp
H0ganXv9TOHdYYICpYDfaU2dDXZRNdLN1vvZNz+YtfKdXLrmkhd5cj7Ucqwb4IEwzdz+zMx4/Ss5
RQKmacPP3Pg3TIomhS+HhC5U5+Tlh8OJSjOdtae9F4+xIqsf6KRikDGXqCVEp55eSCmJRQzgNiYr
NSfhamv1UVDamm0r6TacVcfmadV7XSqhCktA65N4bRJ+sSivjdTXbObTvCUUv9cb90jlh/XMbFZR
UKtrvhkxZPJCdiIkIzdNGsJxJBE1jRKRyqDpLBFP+AGHf86uK2jk6Oq8rXGwpZeW32TvBgZtkuEX
Bspmd+urgBnD4Hq3tvJZhRmA6UiYelsNgcDdqvc8x8HDnNTZUC1v8OCpGxvmHNIhnCOvfi9vuqQd
CnrNBmbjUannnX/MupOV01FYvp+gNeQElAWR0KAIAYde4Z8yj+USAJo9Uxm9e6qUlgr5/56gNQ+c
b2qVOo5TbdnX/I7QolDM26OJSkuqzEQSLE83VlX+z528eFNCDlgYuCfkNPkh14/NqO6G5Kupdyfw
sS+SBydnJnp2lFsdL0pyjybXrtHOA4+LgEEM2Q1n/hFpLYbexHzBhYkN43r20J0xWTjbMq6gbj5T
i+ONew1+Pdd3pq6yfSRWjSlshoIxgJKTcLloCwJb45dr95HAWN0gVPmG0mEIfaJJUfxf5Jynl7DM
5pgFOAA4SCFJIp7UXmHYVgepf1Y3AmHUoiM5tP+YoGeWfR1dHpPU9CMDXFQok+XAvVWm4wSWd9pA
bFuu+PHEA0kuZ0lfsPmmGlrFzerFLUiVuv41UUsic4eOTyhyqhKI/2L9PO+88MSutkpUAxTYsc7W
22n+7X6/1TdlQYAky8egIUdmUB393QbYjBHhGqGpaig7SiXeo14d9RNOsdMJa+Kd6UUaqDHZSthc
etyDYiYlLWRwiT/CUanOE7HtsR4f6R+RRLBi93w45pX9v9eX1IzuIO4W4nK2RGlmSaa8YhNn6kGM
lqBnQ5PzYl1MWzhRJCr1qdTg2Wq6LOTFa5R2al4ssARcxDWlufB6ofMFJuLgBXPTOAac4MKv8Xml
IExObIiByVFWP6xyRx0XYo5tuGYTsfRjUeqnqKGubsnVRhHwdtTWpSGmaOS66YFgse+QdIm8otuo
SySJP8LybwuWr5n2g0o/CyVU2W8ZFLE7MWUnruWt81N2JeR7W039VRRRFfVycLV/2zcj7U/t3bVE
UvBoUF8pYPrwr7nkwUaxi2TxArSHjC4uLz8Uv4g2/L5zceLWrt0qb8y0MDAI4YzRdAWM6y9b0jSS
el8+kJ6sIRG+u1jO3E2ajs0YkCsf+iX+36h8xh4kc51DKaFLY+orcVLoi0TOrQ6UcUOuSSX6rg4X
CjQyHJVzVPrLslIorXzV/qtq69uodS9DcLPw144ziqh7laXSJdM0GnUtpdm6COKE4uO53/IO4AS8
fVs27MrnZBmsMvGCjfv6Z1qTvFrZyS6alQxO7Z+1exVcPxiGqzKTE7X8evlFzK07PMGkLj4njoMc
Z9SarO/reCQCOawOoQDXAtn+z6fifn8PgpQ+cxbtxMxit147xDC9IKWXCI4vOOV8a6yYf9wZd8KC
Sa59mq5TXCuTA+xOuduBE4VCkrvtDWWpYLxRUam8pQF26pGL2ypQXJUreaFf6DceaobAh2vXA5bz
KEsgAJRRwetlck813IfSLwOp/vr7sjpPj6xUiRGz7Am0PoGlqMBW/4JSeN7L2BF+lnrmp821Hjk4
bw6eyOm+ss/7qzdNAX8qNwSz9kE9SrqKbkBnTgjVpvk0qe3JptKw2zNcAAzTKjUrdemjvqliLmu1
KAVJ2dcf5qQDA+mSpGbcRSCQ48CkDkmvB5JKO3OW5WuHs2BQs22W2nuG4n1ke7baKD8Wdrf1gr7y
qwiKGE3s+pXz1FinD3A5ll2Emcg0o6NgoBuT7BUEKYjwzwdeYBVOXKM4ioAaO8YDzd1yna3ajn1s
47N5dFgfxFHFFwEi23kCz8Bd8QEuz31JjiwHvm9N+nA2mGMYtcKnSZ80d2w9ozsfr56OAPjVMpNy
/g3ss8RS6cUWJ44bqO+y+7nLvaB0Po9/yCzdEb5RnhlnuQK9Ecf9pTxSkMF1AKx7GuHPtDXpR3lT
rpDAmVZ/SunfpjJzDsr03yVKT9m6y9x5xdXKzR0kZ6MRSxQwDJREzdmDpMXRZui/x8BDUCLov/jH
M8stBZJ9gw9tV0L6a+C+H+c3n1NnDxbagsWG1vYLWpyICi5XXc2ktkbsKdByaun66NJz2ZZ9/AXQ
o1awG6cULvclhTLBvJUvsCV8Qvt+dIYkJ0C7j9wFO9t4oL7/JH8w/QfzB9YOG8XSDu0GKI2BRlNm
Zlt94LlXVxX53xdYr8PF5+lUD31vY9DvNG2pVZlSRsgiRZdJZkw9/TacXCybHrZ21MyvR7lek70m
Hqtqo0P88MhWBTshlJG1VpsmdrHj4eoViNtB/pvB5l4PAuSDSAeeoj+EhWQC9DGQ+ziHew0mkxyH
Jjp9JJ+KjA9J+sA02FG7DoJy6iYRU+wQmV//r43+VmeRqzIlUfQe+cSAUebVShyJv0mv2DBjOG4E
MPv0N6Lw9bcvJuJ1TYp+h1N5+T0CPu6F8ITT1jXV+ny6iE4HBXe+aAp2MsIA5NjcjKxbZ72INCuc
R1xf48bwVw2TPQV+8gwLSvLWJboM2lbpMzuNsW4SzsjSPrVbbxa9E8yi7/oSAG0cFVmndsq/u1K3
PSMhsqlodv/KzyGsCEg8lUStBtizKCNIReKI2Jcz7Oa0pjFJBv2Ork/Dpg5DCN6uF/QXdZfp1QXf
ldRQFBZyUqbgb01h9rjfEVg5VSUZZmlIGxXFPrON5y4NrRiUngFok50j+Os3MersNW8k+v/wAWIx
/J7nNxlXhgjBuNC6/3IcKRIXVK8S433CFxq+lTw+N3r/WCHGylJ3MT4csTcdXgvWOBOldQw2/+Dt
5JhOLPdS4btBNQloK2cGnS1P3OsvgGmmIyI2JmOBRPeogfgGMwFlL1aQIboo9+w2lPtnzWmQe0e/
QKVZh/UN/DFZ8/EIosoN5bf5daW2DsDOXrrLr8f1dHcnqd64lCNALhrZ2txFJK5axRYa/5f+QFlx
DmQ9JR35/lDBScfxqbDSBEfDb/6wMUI8vHYPBkyp7jwam+kSEcZYTDPpQqgge4r3mNNd/0qNqZib
F4M9eykIhpUuunBXv/29FhKFbo/r+W0ldQQzwAZLpkq8KIGf2QtGZ/P8tYFwjtORrXwCiwjFo+SP
JCc5EM7ekv9ZcPMgBJUXy1MHbQLaCOay1/8E2OW977JWuKzVIOv4t/dcStLntRHpfGSLwD4+Hcuc
9rMsCARRwTqV7s9gRbn0kUQxJUgFUxaf7leNSNCqTb6ozkgoXErk68o6dNk+3iWs/QE5uEh4ZJDw
tl1VEGZx+ebzRttdyGFe3tBDsrT1fcBH36VXuU9mdlEgS0mR+ACZEpEXV8nhDQYH+6z8LEUhZ3P6
wZui4rRm2nCowAAu8B9oG/QeXutnLF258UWNyeUVFP3x33GQYRS0aHrauHfO1IOG4HOB9RLseSnw
9PwglQY7830qQEU4MwsGA4KzVfPL5uTMXQbrqhgMN9ixH6nZQb+u6gyOdSCvlkVvSvvFlLFYKaMe
WJ9xSnp8ZTdlFSDeBt7gBRYI7SV0Bq+HViczDm1YRqMyfMO3Aa1oTctM+gD1h5fDZO2A7P2AF0u6
YMrAXxyn/hGe3egyVyeBh7kri2gpnEsXn2uhLgacBL5Yo7tAITE5Wt1eUCiehnJKpGxQ9O0UQkEm
15I+aQCqUT3R2JzXjpAG0zh3Vl/jACgaGmyqfS7RdPme+Mlt4udIJPlrTbuGoA9sycHNnGCRjH41
e26rGNGk0NQkE5fb5RaDxObhJpOzAMNCkEgzRcp1ytWJ4eSxRPmo4G0HqQkqfn2/U8CsADiHDa9H
ZOVmgjravWEg9S7Q9dR1k9Py1BmGg1O9zFwyGGl7GDDUfcr6L0AvGoo2tMuUoEBBBWivzp4so5V/
fYtHLhb99LzwEzjq0HD269DAEeFuGuz1IiKp7SxN0wuSWq2eiW9RS4rEGl8oNUaACK2rOyNbzsoO
Vd6O6SyMXQR5O0VlsACVZ6dkbbofY3GfNf5dhZ6WTAoi7UCvPLLFKwPMlgMTFu9k6S3neuKcKbN6
8PQWSZVChPD0UAKkIBcKjOvh7SowmMAr3IEkCUqs1IHnqAZ2Wud7wqcohwURWsXMj58Slj9LoH1U
yNvzvXnUo3xVbqZJKGZZCibA4Hgc1lQRSsQhgZjf3spG+SC8jLL5vXlNztaSs3OWrVj1xcFyUXah
xrm9UzmxLst0EfXcILUReRpMs2iHUspb0K7UUwpE6+EpcW7nZbghaCPiPaw/U1b4OOy3SXAOjgDQ
cukMOTE2KEteMhA0sKKe3b3EUZpkrI2zEKPFAi2B6cMK5CYjFJCAYbVPBhQ/uETtElgemFffOL7N
cR8Oi+cfrRl1JfocwT9kWTfUek3EMTxnz8Pa3ZujkcJgtrkIaK2uYTsC2I9tJhLmdYqh20KKPSgv
PH/TpwdgDpm/RDiLFEYtMPQcMHRcAh6W52QDBMvVAfup4Nm6gseiHruf6qaZHzaSdfz+ZCyVRnR1
Jl67pQCGQxqd6QabL46O1dByIGzLMk37uNjhBjKlkT/aEK3oMYOBbDMg/cm/cSZ/onMi0EHousuJ
6hfvHTTyx5kL+w25iH09JBCwuNoT8ZwPxIkhF2XljEemclom7v9tvyGJKkSoGhh+ubRlrx0iHhtX
CdSUWf/RzLwfMZ6h9xJ81rW6WVV/W4R+jF/bFGyii5ECEnGvOW2AM5sJf+bmFg1lTJ3Portad+0g
0K/uGLyos8FN/LQisAp3j6a4N+ljgtOT/9kchiuZDcWzE2lp7UqdhKtjVimeIVoHFeso6rEmiPX4
53nOHviMywD/m+YI0rIkw1kQquup7lVzDl1Dwf3wOYQeDNwuG/xaKbgg0MCmammP/9k8e/EE5wq3
7H3iRheY2x0fxbFBk4jO7GloEzhg4Ev4wiFw6fglhfS2vQ037837K98ZDtVNTvxDGM5Nh0vevGaT
4gDqKo9ovkD5eDiOYbRsHqYMXA75l2boTSrrplP3z0RlNksptn+UublG54OpySJ5zTztW3dahm/M
+mln4VSpTSDkQn3Z5K6Y9mZJhIjM+NidpZHfXUP+/omb1GS0Fs5cKZNLj7qWb3nhOVQq+/Xkhcq9
OLCqVw9omcDf6Y/dMrWMg1UdVousePpXLZVnC2bjJwJ+wtdQ8qolyZUthwki6Mwf5/cv1S+GUpCy
LrMbiGJCLMreMVYGd62721yMjx/joeE0a6VUasc/kjgZHmAma+auWnb9k/A8u2SdgFJt51Myg/Wc
w0c4dyWzqv4YWGV5Ea1ybXxmBP1T6pmcgll2oOvaURqvy0c2v0JwZenY+7XjCgs24mA6vhNzcyO2
G78hsdPUaXsz9juXEBmPpIrsXb9/zJVkhrdamWH8LgicxYnfDAVF6ga2UqUYZ1KrARw+DIEs6JHp
hJO2zgO455MEqZHosIwtCAdnqw3OIXgrDf/uX8zJ8VuNRDTPY1rcwr3wzbQ3jdzivIAznigboNTy
FnRjB5LQuVIaWa9c0wNIWV3TCwZdtB7xlJEo4wkih/pPQZSbVIPxyaAzPtJ6XuaBCKuLP170NnZL
stN6oNM1RY587J3UbaQz8n+T6XpwFKJbBKT++gBOgdYh1K45pXiKPQsqNrUOFp3QMfNmWLJ6gpE8
ILb1CGa5QYTFf61yN/dOoq8EpVH2csujNU5gAxExksbQ7Yu2zE0m4iYmX5l6slda+f13WjC+N7gN
kf0vj6nmCYFGlaeSEgqKPuugf6g3yVVP2a0FYoGwwrAXYWwOR9Ngn7jlRlBymAdnihE9fP7BQ7H4
imx5+sdzXxRVwdGxNiEANu47y3FQsrtXP6gEpjjAgoA2yEmyVV3YZEg5grzGjVUkgx5KFbo5CLYv
5f9h9hbJiL7iuSJJHuojwveYE9/qhfPloOKfS8abL4M7wzgKHMS4xiZcIZpc8qvD7ZEFiGol7jsw
zox/hNtJuTLHKMR0v0WSkknK/9BdetSVJTFlujKTJ0+PRs9W3zqDrfq8yGSIF5naEnj5lDyv6dON
Y2v4dTbB7+YChfc9v77asXgg4KGZL4RPozGlSf8SxvqPnJWg3XSAnMZKBWhrdxVzpvrBj02GYV4U
CxlJluE7FFvfoaMTig7ekOx4Saibh/mI39jKg26DLQZ+Bpc0lCAJtYjYpjiTroZsDAyPMPUmDWvn
6Q9bT6S8QyAyFtwVMtTAO1TFQAtFF0MPQrl6loavrHbob1WchGWFxyeD9stsHKceTlT71IoBKNeB
P9VIDtFwEZf5Wyti6J8LhlFqEXJkIGJ0BlEdM2MS56ALr2+vWaHmYkYsR4DhopxZiJqMLM8ZN9IA
L4drG/bdXoIZjiFXdgQCPSdf46wnYo/l+SX3/j8IBFI4aZnemTm1VvyvVu7vYJ46IuykTGBZNVcR
eyTCasr6Pn0efT2qHY5MX1sZVS2t1U+IFcog1TsUY6SwLBd8wiKkkC30hnZENQj+YdTQxCnWDIrv
+ToOWzv9TjNbpAa/p+VjJyWtUgZAuLqeoNOfyptdcNZ3DjUqg0VE22ka2783CIl/AsbcDnQXncYq
qV7uZM0mfUN7UzDnZSX6DB0/nwd2m3eBUryL9FamZWJwxFVSw6kga1zX0Reagm39oxI5cxcKeLeU
h524YVUYCA7MfNeMuSpU5nluXvyH6dfVuUJWKIkIk3qSP0t+P2pE55abZUX09hJpZeOofGFEeX55
m3HrGt6zpDcOtmEBx7BGHXHGIEuwOGpbj+7LJTuuvkd9toVtjV1R8VUDv93mcao5LepRCGfSoHFS
nZRNGSe6Q8VoTzCcwCrEPT9EJ352WXPcHd+gUblpuovF7F836QnBdh7kApygnS+aqdbRA61kMlAF
mXQzMUUhrwz1JzQehHi3BTyhBTdhgLwPhOAzjUHYElnzWBpFCPXlclHlaRp1XZJhVBcTN4giihDd
Bm8vRMqH6RbJY5bamTZ4/cssMhi0zl/+l+0HQPJ5AvHvQPSZXL77EzheJM5lkRklquWAWdQ/x6uG
SznAezM8Jhc/xoq12HFTRp1RbUvwvy3+5gvPfcDOxA+hwsz7aIQXoo9njBqSD0OFz1lMPzJx+DkO
b2NdkkC1Ir/GfLBpJHxBJANxxto48WKq6iP57cmNbxBj+PYFZQJUYeeV6mKEqzr3HhdrCnFQCtx0
RFHVVDJEv+XDActpCkwlxxlLZarmbPLZmltzQsljMLhHOWjhuKWXCYLP/E9Jt8PhJmbfKnl27rIu
xw76qQyVEuQ0cH4G7KyKBaUISK+rLNqz4IJ0+BWUhhROgBgLDAjpwJvrsj6JBHzRdqVPkBNM/TPU
VdeIllo3BNwcyoXxO87YVU7Xf4Nq3OSU/BEZrC6kpFQLDahPqTRXMbppqc+V6DGVfWFNuM22zYqH
Tx/HhIXU9CbRcsLFqCXgcy8YiM8HBBw7nlY7+k1odrkgw16aDr3bk95xtN87yxuKA0WJRWEMQS4+
Igle69dQnvMJQjxj1KAmyKP6sbB/tfLArnjQMXMvh8WouczOpd6gu7IqfaqwTS2qDGKOXV5ZHBSN
jywnXpZNZnWSnvDbbFaNeSuQaaJ/1CpmRFneJyLCPBsUcXnLrNzvsJSiPIS7EnqnhIOB2gNfG41D
dMZNEjzdtQUX1FvLoG1QLgGaJvK15BNr7wF1BD7tfNnUZtvetbv4npZc+GNBdHbOPN96mt5VW0V0
U6oHu3TA3aLCioK6RbshYndic+/PvfRBCOBC0EERedEkr8/xuO28GkssESb/muLKlz8lHkTfsAfL
ZwnrKISr3CFw23T6kKw4riZbC1uyPe5DaMO6GENemG5D1Bgsfl+PitUr/yGoRZi0/gteXeIkHgTz
mICA+R6APj0Ucc9Xzv5B00ILc04yPO4J9Fyn+TQKQCTqcZJkp6wjqXVTNiekTTYAtsiXfmzfQD6o
RSWsRn1p+Ek8250pBk1l5spJsioaD+3z/eQOuyfcrxNkSSu//gaGlMO5/swo5wvxjQaKqybqUKys
qdcBq1rcYEmviIDzqpyvcBe7Y+nDLkm01MHWqTDSF0hSli+ZK6IH99Bn99OSZt8Gef3VgYporvlx
TUBAmnMcfdOkr8jHATApCqrlOlDaS/0EvFpEFvEGp/bpQRSjnv8N7XgBIEFo2TE1FC6zSjnW0H7F
QorgiY5x87ftZff3WIA1gQ7ROSATYt65FYU2WwwtJHqJhpZhCy3ZCAQuVwrflBN8x3RuF97eAeF5
9MuC6Byu5f/nC+vSBKHSYurQkRMCoyl4ru6CvQSuVJe0eUegftireJm0E2M5VAfxQQpYsyxcVo13
ZJliGdZD198SHQuR1q17+AmQOfbCBauGWQPqUm1pPZSm2gOddq1OFbn8B0BWeGG6/I5tZdEyYQMx
8F1UVqMzCYTirHP9TmWqwEKSWeq5cZaU2SZaerVWQlHFO5pGxrMTlTmZCopa2jZ4jqr4YmEYush7
iknWbc7fHNwvyYHeB6tss0sS1oc+xt5Kzg4I1tFPBLG2ASYcYf+IYUlvhxzbIT7lzQ0guveRHQDt
fjm+XN2L0aJ/bC+picW0DC7zADLsh7VAvwaTJEZDFW35gvqavThsPEqbVBltGzx+Isd3rdXH3dGV
JoEYoK5cVnQKu/4pKOUYNVlX1B+d5ZH6MaKGRyfLIAip4BbyYat15nZ7K3CpJSAeJmS+/XBNgyMI
rRbZrWcGxNU88eg2iqQbrLu23Gb7GrY4fHszCTymKcXBNqFZOSRtCKqh3/qI6NZQSVC+3O2+0BkU
eIz5Bv7/EoR+s1zsryXfcs10D3+Mbdfeb6ZcTDH1D02ODCASCKxzAe1y7j+xZRhFfGi7Iu0ot6x7
Uebh2eQ+JQXQ3I7QZzejspdXZzpIDGye2fT7xPkvOoOPvBEf2E8DL0UvcUHvtOIo+cfJTWD3WJht
2ML8pdjE6kznLrlcTXhkCTibi1otB+fGEzceDVlPuNnGpzKizN3nWMnY9eGeUuB+cPD20KJwbRtZ
9A80nTY1rLYxKFISi4I9j99MJK+MttSfOA22jSwsUL5lHOGRDgZm3vdICYzxSS5DD2mhrz9gH2Hz
v9B+qyMXAnh+RfEszNhSdbb2/OctngUG9ZuG9XWhajWzHw5IsSADbRfoY/bgkButIRD/kCNUbmo8
TrjRLqljF6UiLOvAsWuL2O1kenZUdu/quNDcJ1Fj+IGxGi5CxbktN6GxhmWZSw966ETJU8rvWL+A
Qmq8YDbXqu8SHwWeHlMklDB+eI8HYyro0SF4OsEmGLsRJd4d/Q+xciEyyKwiselQSYjKhCZFU4o3
l0UQTuGPO9AQqIOu//x5NHclpZz/ks9w3Eeqr9eQGl2LcAOsVyRqOc5woiouWPbOp3lrMmRqFM6R
OEiW6LOvJlJyhJj0vEW31JA0MjuJjLCuPXWe85uxYFTR9RAhwR8NQ3uHMzHhnFDGlJxNO4kScJ1N
CHCLlOpaKPzyzTkHeXV+yJRiwWIv5q5AFe7XHPpVFW20aYAQjdBqzIyAONEZvZaKr3dRm2kygnqs
0XyUMHyQDqj3mRxb55mgeWR3XGuPdYQyewUE+H22Vb/paWhL5GbpRTK5l/wY8tzIKbNMM/M/bEso
KElo6Y9tF+GPM1b0Sy2OfpC3be4pdnA/uU9IpvVmMy1LAvpcf6UgwjOi9loTpIPerWbOhutt9YeK
KZWERUUFGgYedkq4iNvNM31xEUh1eENU+lmWTNpcAb0uSzbnYYpz8K9YWiFpjy8sSVHoxGCzE7On
2UF4TBpwtJ6pjzlaqTz27IHxwjsye/Z96jEiqCKvDRDyQn8/t1BcyA4NYri44g1Lx4BRQZAVzSov
Wsr6FufBkFfZC65xyGqYJSvJ9UH1uE569fjE4H06xb8Syqo6qjQ0d5y1rgQIDt2vSFY2s4YjslHl
BHbfqQXrQ3LIB7igwPloQqBb05Mg0ZO6LJHxwaTWlYbRLoAz36KAwsUnTjcN/S1j18bhwqz6j/nF
49dCJxh2ZS9dkg7eygK/rq8ClzP6X5VnKujysuZQdSG1wKHwbfkkhEr16VYAy7jHDTWOFhunsetL
GrvNluTags940i1JsMyKc1Q4FqChZ587Zy8sGbnPmVneeMhECprdKeWeDwb8M30sNLCbJ/L/Z4cM
WwbTucYxh2uzNipb2oNgxXZgY66MN+LmAUeSUeLZpH2hA0TFNoxT1zhhytCiR8DuOTfN4HiusiM5
D+jVxqH5jO83yuNEYhj4oBg5GObw0a3oUa0aqE71a/a2Vwc/bA5DJ7ZrK70LAHG6KkOB50hL2u3z
BYcckrCdGeDMCCmRObB2HcenEZJK6PVsBi3XVr3STl0H4w7CcIO3v/gYrcsPKoZojvsxrkYfeHeY
Bo/9nQdfKoAeFwX6KZUEhclFs+/vEMJICTFjfSOZWT2XzUL8/etnpAyZB92nW1L3Pk2Voyx1fauj
ZwkSK5CKcUGNXhayQ7JyCNOJBwslg3Kh3W0etrGsCPrZS3g4ZPSkAZxg/5jGErIHWZ2CTMjYioa3
HUdhG7Tf1+I/iQ7ovh56z9MlW52Mp2yH01QQEWex6BU6+B4/rZUoLzq7bhii2x0SUMn7wd1KmL9j
6kyC6TOsUP4MW/gMaT46nt+NszDKVVAiKSr633evAn37IO+sCppznGJIx+3T8/YGCL4RUUSdlVIl
TM5LT/2t3h1rHvWmHAaFWwlRtzvJucl/W3qUKUq1hNnTtHpxwJnBjZsGx+VK/Tn+dxeI8cW2I8Yx
oHTY4+obHiaV+aCyaUMirMIYtmvlB1xzdLOtJlAY83gVlh8vB1+u0gYq3p4sOgmTI6PQ0LaGmYrd
KVpGr1S9kkbl+0YCE9OVJAZjCgr8EezDp9Qupbg31hWsKA4Jo/xEcrTN7o97qW/H8D/BZEp3B3IO
ijx2Re+UiUj1gcH6d9rWuiZ+V+2GePNfSVdn/R2K6a9we8pknv2oQexxlpCDrkxL02v0pJN9Rsdu
H2TYWIeoZ8MiZoSSuhNbCgXZYToaELckhd2BW/5YaJG/V/CUXGvmYYcfNUGvym2V1P24ugaPR2Hk
G+E5EKstJzXV2BP79Jl1REpTmyi9+nllGu8NaSl1AYEuc//Kq7TIirZrrUoJw0fBio2sKPhqkLLg
lTyAqLHC0rOTtoz1IApPVY1qO5rXVeeZAv8wlMJ/xWVCqYp8Jkm90fayaSl8tnjCAPCF4sHTPX1V
zqg9CwwThWwtjVWvuMR+dQn6Unz2ZLG9jvFo92ESv9hwjSwUPe0ryt5kpcphwtfoTN2mpFCUIFU4
Ijzr5o1XI/GUBBQsbNHqbR1EUT1Jj5xZQHe1uDDRtEk7WN6F5q7m/rsCcDfoWIbu62pRwkAA2D7z
/WRgRpqxRG79cIAQmGdFmdPThddYVnur7S0a/x/93N4sgdp6KK+ZwzEIesuUAW4mi7dfwKVBt6u+
kkKDDejWMxVenidEw3hvN2D8BxrL2l5PJwqM0pf8hdxibVoHHH1GHgz5Vt3wdcO65Fw5xxHZMReZ
1XE5RNzsILnKKMJalzv1coLskzibHVdVrXiBLlSr7WIAtXOPWRjGpC28vsL44oNI3XRcFzG/5ESN
mFVZaoiWDNskrcxxnbojA59UDAresTPODKwJj/6asYZ/4xDF1p9Fq9AZzG+7ONTu2AvT40tvmy9y
axBXhHtC26LTHjcq/5WXk3rtDjEsBiu8FGdiaPBgF134ouKDRgbJbrMLVluwN/aMEdQ5KLpDquES
/GGKdGNGgVNMozCUDm4ShLwA5ZLx9pi5d6A8yE4GX5Grn9cfdiAV7FWLk9Z+xEy6l8WInRlb1AlS
0siOcar6smBQDrNFzv4YgB/I01sxLy9Tw3F7euVs7yKmlN+YlYX+VKud8R/MJEHYiXqWBSaiBYj/
zT/sTRNtjCsCRRomTYyZe1K+xJkxOKyY75R32ql7chDJ5c7GwUqUwEccPB3OtUnduwOECm3t6C6P
xmdCRxHjL0KBXghNnBPkHiY+bSjk/liJeSyg/0eIIuws6sf5rG4Cv0s2DX0bTr5Eoz7jdpG6TpTa
qFfR33/Zhm3tX2tFhy6fwZek8yLa5uDvYVFxokB2fdkdZZT/spczDsqfu6HbMw84BiI4EXyq5VcH
I3NT7vQv6cN47GHGWAxGpD+zOMZPb+RddA+lvtCjO3Xqj5l3PGoJHccirjkaUyAI3YOJ0BxsfDnI
ntBxfX5//XGF3pZcIuUYn62T7ToyTR6DYVkfByPvzkTrlUbRuzv70Tk0EqYKiOI1SG7R2ywTB01H
ek6xWqdmwO0kqH/UVfDdZ6pXrUffw7+gSSOPp9F8PzXVsBgFYSR38bRGa9KFXFdaOLPbUhzfxxyt
Yt7Ys2rdoJigb6lRw3hzPAfEEDcB340RUeFpMc583jJpSlC41SrvO1MPJ6f7q54S5Q2smaf/BUdA
5P5fA9llnrWybUTCLdG3FlWXJQeFM8e6EaE3ESKjTtuYokYuUb9GhSKPEqEGJv25QL6ifqUDpsNw
k64eLlwLMHsMKsGkua+0kQQVQd9KOav/C+h7a+AYIVm9rjR4sx/JB8Tl3G8B5EhdAUfNx12/GOL+
pBiZO+HMPTAsDXtHOFK/EMfGuJd9u/357ZioYmkvh/X/P+APZ3sO3MqNILr08ku75f7GAVSikGlT
daGneGNdGnia+QAwverEehiG8EFwxBswQOrE0YY36zHnHHU0kOyt1fnChSc/DaldBPwvS1Za1Awm
DBKObxSAEMgPU5gbZk8+bJ/gr0y+yzWqCbMAqbaqJywfElFjTlden38md5sv0Klvpy79AxVaY7nF
VB3Ku3i+N4ECAdrnDJ5VlgQypkVjjqbUSvMhhNMQwhLE+NzrnWAQGL4pWnIrEq3UccNN5USntt4A
EADg6+g0I5j+7Ext5rNm3utI23scGuGB9e2NUymlcZjUR8yF4xB3n0O9CfFc4aN3ztkXOVIZqkQZ
ZotdOLeOTDPe6onaVhEh8y3DVp9LCfpkJ49gXu2pvk0N6C6Em29YAdmMZo6lmAlu181LrSxxkQ+S
sj+B1EanLkB+N+oObaV+hNqBA5KgXagH6+TaM9zDi20K05oycjr9HzSiv/jPUI5S2/HfsJilJ/8Y
ivdl3Qg9AQRutGOyeEmfSgWoC3mp4Blrj2tLJQhbBFFBsB+kLR9Py/b/vNOfPbuVSLX9JqZEm1yA
6eMKRy7sM2SIeGljvAaKY7n2SGzpDv13phjTtcA2sB/mDMDqH62IRerP3+XNzuX16pU4i5lOUJEg
mFJLH7CEE7BbrlhYFzhDyss9vhCt5z1EQHrX5/hMQE7c0JnmzdYzzaPhAV6MgkYLntvBKOoI9lFj
ufQ9KGLJXv+bNNk6Q5/159FXhdqqrcXKXDucUXFy6cQmupQBGoCQYJ3POUyEqJEsdDPOZ53lBuJ9
tIFac8Hrj60CFUzWZLDVvp4453AQdO9OnuH0FCrnII6BZliomW0Rn8VEIHbHGxAwNB8I5waOD7Pv
9uOd2Dkl24DQJWX4qyvMEicaO3QjW2b9nl8mdKXAz7qMcOTfFlCb2t5JiMt2E+9hLhZkduPdEbY6
7AFHsLxJsU+tPV3ygj69CUALAHQtKemt2X6jev8rzw3nkoaVs6GTzp1HZAK7DiDOaSdea73ZMmUW
nSbvLsJM2zxJzrJcObybua0oW74sCBOqeRK296ZVpDr+3uNHrTomE+7+dGPHXZWVf2zKBuTsDXA2
E002pjvCbNov6fCd+w/yzgDeq6uR6kMNRz5Da4nnmKI/dq0fZNpg8Lf0ryn0i2Rz09k4CUxBH4X9
X1VHHjcP2zYY6oxpuRIDg63Cf09CiMLL5QICpxDad2PfCX1h1I+Dl5FPQWV7rjUYUxF5S51aPza0
x5vprQkmYOwgSlNYhezZvXwVlIF2ZMeUwBjxR0ovT/BRtk1Wp5hbAIRQJSTu/HFFe3AqYUvpTaHy
DUt3ULGhUwb1vxnIqOqgygxKOQc3XsYXa/QTXF3wDvasHU3fm31LWuNN9zCAFoWAQNJ5utXBcwQI
UnmhKer3Xoiz85w5AOj8gLstQrRxAzRxsKDX2PUZhoqY9m3VUnOfrPWEMODbM+dttE29lDAQPjgw
bKrnGWDeWCjnoJ2eeb49ZBBHlhLAKtLLFrpHe+NN2Efh+pOTdld8VUzLOHSyfRWvBuOWg7K3bvT0
3QvrPmrcdDDezNKer2hlXePabqQc8XOLeEdwDMRoKiXxzWlecddd5A2CgamgKUNNejwt0qCadqr4
wRXNh51zXoVaruBp6gPTOf9S9TE7SMUMAnKDUYzHNxU7FHaS5PuzKiNtBOVBLjDvSg5cyVTQR9so
vErVczE2r5a3tsx/000FE/FJr7geOHZLGkvD5mMbRV1V8XNPDkN8X9U6QlDl8B1ccGRhnymwHOwP
KdAQ6mBG4Lw1LY/A/w2kk/eoekaFSaTrBnhw004D+kuwPLnOHIq+pRHYm0zxsRuNwkHTYUYbsc4p
QJKJpMK2hyqmew+wEP9yyOfzRmBlasn3Hgc62/sLwd8+8UaInoJnnd6WJFMyWUEvCplNCmP1pK9n
eX8pGZ8NAbCwxIJNaNL/nYHQ+MeQRhCpCiiU0MEtWWps7Y0jsa571lR8LqVQTZ3Vir1yxR51iJvw
5LS5XsMNe5uAbmtC7oK/1rsWkvLVA0CJSQU0ebQU+4YRwBfJPFNEoS7IWRbcF14SIqSpxPmd53uQ
wYh8DaoGVLL/vwHnxGyF8dbjVDk4+lteK79aZ1JJaO6YEBW2O43jF5HtE5j1iNPlaKiUchT713zo
n5XR0N95O+qDCQcXeQ74SNb3NXUosEiu45uY5UD7a7JV23Rv12Cjd2yvx+aZgE97+ImUWMtEvGeZ
cuhGBcSuJqOsubj+idZdgRIKIgbVzwOrUoDOhAGJifEjycWv2LkAxCKH8Db5ZU6fx5B+Ck+qJIHy
d+KOJ/U2pT1CAg4v/4ecuLfgKoqZ2JJJj0POvI0vQl2ns02DGR+kxUdMZC8IytkSijvZQW19YSaJ
iumaHkbAp7DwT3mauC7QD8mobwWUZNkuT7iwRwASaAV1zLQygiagQJf8ZIza9Z4KLKNKPDJhQrlE
zf8mWCa6CRt6vfcxFBXhuvHwyyuUqgQ7ce62KMeVwwDLO/jGUGOXCdXmfhqLWJ75zINJcX8fsm3S
xPC56xybohTsh7r/6+GNlaJMREVGpMt3fgwL3t6KNb2y5zXL2OgE+fWXrSeQLqTk2+5krIpqgkt6
x8OGNLCis2b4RA4NZVycxXNEqjNfB9jAKd6qoNWhmAq8twa7lUsAPBwllHvf6qF0Q5DOzKtvJSW7
z1lDm2f6Ir8mRH3cF/xBwnPGm/kDK0qidVeLFXRpTZ/dCwxIWbtRDBhgxpii/IgyFjtAUx280lXY
DNj9hoFOtWGgbQoblIIfz4uDYB7VrDTAgSx3rJM+sZBnD56jBFopnQEPrRVyle/YkVNGCm7e2SM2
v6bfgZXeHhw7Yr14AuNZgXXl48JwFXVJAwBQjfIddPb0CXxl/vxWNBFfO0nQP/KITrS6WuVYid3b
w0UfeS7g0+z3wOMsDOlmEDIpZTEvF8wYg3F/mJtiZgRYvtWG8eFFXENtaQxv+25x34okzmlCjnxE
WmnLPvIO0tVOm0dn5we2bNtcogJLzEQt2bFhkuGRupo7iMBcNfuerTQQSxmTnbjYTIOTxF18dF5y
QZU9uHzvHOkjkWU0dOQftbuerSEIjihJ8VgcG/l3shqZxRNC8iHRGsK/P5Io4scuMAeJtVAj2UBh
g/FLYrZqnB1eqhdr+QyZufVD1vuGWomH4UZ5n7MIPDjow0bb/2CeILsXMXnMMMOeDWpXLayEEgJ+
snkpZHWQHwQfdlkqJNUAgeQxIPPqeVJTNi0Vf6zS3iEl6AnJ/g2q2lFhZDJhDuwyi4OtBSiPn/OE
tDOOCbn5OdL0FQtjCtddOhs8UB2gconZ88EV95j5QWRM3DupNpTCg+SbT2sG0PfRz0f+GPPexRDw
Ek3jV/Rbhg6MhLuwL9SAHRgKIz/X/sEoeBvIB7nIeN+KL6M3tTKrxH8mzQFTuZelAzIPTLvWwgkt
xXCUkxScqq9BKd5g2YfFsIvLQDKLB7OgGVB9Qy66rcXmovck2KR8/A5P9BsDVwV1/P/G4uLEYQvs
YoKaYz2wKscw+dsNK2x/Ynz6WTPJFX9vrVE4vNPYrLhFFDp32GlZJyebqI2MSdkOaePdWxShOAHA
brZEetspxRVlcSd5K0bIEnmFTTlnNZrOnwFN0dxEDnkcpKbK/46u9ZP9j3VUQojR9BPnTY76URXw
MfPw2mrnGETYKXphgXs8WsY9zsSLRKYn6bUPXFhrXbgTM8MGBM5HDzButs/We1r9DjXwEd7szrVn
cyVaY+fuNcWolw2WafU6jm1e0+4ZFG5gHwbLYva4vpzTN9ft8yc5pwwMRsk1nRd4yZ/eEFWNaSII
Nz+LIjwmJIRhN7ejay7997mIibHpav0SpQZ3NgSBddYXrCBVN7mT/qCOm+ubR4zdpLOzRldrNrQJ
y89X7D5FwmEwWshx/ljzeteHqI2A8C4zCUWzIm3zCKi7RCNVzUtb0BCc0PHCV72LYKes3QWqQPiG
MD4K77n5O8q4+9MjJi/tCSxiHYaE/bV5nehtBGZ/fwydl5tDyiqF1wrBdPPqgxJYTttFAH+1GTln
Q75bthnZbD6fizS3S3cAScMJdTHEvhCW/HtRkh152uxjbkRaHLjzxkzi9BWWQCmMhyrgqdrwRC/B
WOEAyo0RPzVMp6+tMne1effO6v2kFcQfOeYsfMOQ92uqPyt+IxD4JSDaFDiA2162hxLUJuqyAhZv
K8OmK/FAsHLyvl+iSLG2+1qaJ1bv1FmhDI038uvweRZw0GHsdFgIC+CUtXQyFhXEO5RF2OlaapaN
3KPAmkyA9HkwG1G/k2PIcMN1ZGG+DpkIU58tGHe6bot0PHHIC8V2zQu05lXKab3F6INC8xMWZ2FN
0JqCuOZJQY+zj/cqxZuSWCsPuiT6kVYg63s55FItHbwwTBXQKQ132it7BZb/xVK35+sYZ8I9eKvR
9DAii8Ow8YoZsWAPA/bJFUWMIrQESF8BCGuDVLQWEocOyZGHcJS6+5bYWw23R1Non8OZA3qOrw9r
i/nA7EbsYE5hnHssQWkfrkUDm/JwZKvmJk+/iylKajiamnHBJ6nQM5HjEyNDDdIGlpTB0sQggpg8
n7Ps96ksGylGfu1jFY5arylzMpiSzE/KYB/B9fB72SbsXbSFkTH6jkYsmX+EW/lZ1Mp91ylbuKY1
SYk/7RbG7G9ccy/G4IiXAAXHyWHgfmyN/UEhTNgPystDhCu4yjyR8s4jYQJt9wi52xwVWkKj1jpF
y75uO+Xi1zeUbIejV6mzJnxoNEhaeiYINXVRff1yp4EojuB0FFn84POrEG4Ko5FY3LwJR290r18a
yGwxb9OxV80KOD7sYm5FiRc4tXcmdppZzKsGxy1Xg7o9BTnqdxA7nN48TEvKiUtDXLdHuJnYi3XL
Jjtl+7cbXI94Tu42n41thEcwuwceC8FlWxi+vtONp4LLr2qrR37eAyac52zPu1L6mBYAJ3QDbxs1
llNh4+ZFy9JjlzN2G2iE+agYjB6ZtWzMTsr+/LSc3FiKfoK3JPs3jWvfP3sP4pdGJjVFLVJjj/O9
BEPM7bi7V6PZq3R5oIr5J32uAftegNYH1oJye0nezYk2ClRzir9LooPjtzpNBEI0+hgWiqzLDwai
vKDk8fuGAQA//+KpLtTrgJvxzQnPTvy4Z83ApUeXIN+Iu/69Hnx2aR/d1FioMvcOVxy3PVOrRaq6
aVkXM3ppIEdTLmX7V5Shf6hdtUSCLZ0GR96lKP52XYi6QcUDWkZ8+EBSa+MKK9BIEbcgIB0wAi8C
tECFUQAptmz+Ybwdj1OJQsPn2KfsX86SMbNUYrs6NCjxehD8zyz5Rid3cl4uzrvnRg6CJ5dY1Zxc
SSuafPPYmpYjSEZc2EpAJu2sb/CCyEPrdIs6WLToht0vXcXT+VP10wfC+Do8D7VliYwIgGY6uaBv
WeoEl+ZiaHr4/V+pJTNQuN/U938gC7lPI3oqMCHfNHZrHOZE7UBTLrFyL4BkaTXj9D/r/cCFaOmq
Qk9Wr3+rdRANuI3C0L1Ki9AtKvqtSgxevyHeZopzrhd727cHKKFJkJYJMbqMG5yo6EJ3cZlkbOkk
hRCIZHM8xsmi/IT0VkKB+CwWV9yLmcl4hEwHRjIxye8LLT3nXNJwryt+aehVmXvC+UJcL75JSoVP
OFGfJtC6YB5RewP3DVt4pkCNAKoh9vjz7mhwmCMDhg0oVGS7iXKq06nn9ipaOlGjXwwOVWo8pgFy
blUQryFv9jY5fQnhVCXqZjt3eOqRDExsdOMBB6HrXOBuyOmSPcjx8QWehns4iF5Sh9oNz6KTDBQw
sYcpyAPn6wWjA2A6IOLeXt5hqoWiKeN8V7lDRyLDd29H0/U5l7CJNNjw9y94g+zWBtbAT8a3C6xD
DNc/R9t+K7TyrhNMRVb9oVLujkOQrFIKPdFDEh/xOjDl9FN4JQkEcv7hDATks10bX+om3JyRMds4
xbCHUPtlfdBgTyNdPqCQtuMyx95aGAmiUdimId/byqvE1NQ0uaRCq0HbAQLBh+P8X++PQ0nVkMEi
m85HUWPauf8FRisGIu2qRLiLvP2hVNlI63KZqwuS6dJz7kCG386inxbflNrbla+dbxmHZ1x5DkQC
6ChJIyBaYm92dr0ktq4it/Fw/gbFHAqsmmUD4K8fSSjhglTQ3QoCTFRSjBpLczIeAX7aq0JgIKQS
JirkAjoQqSbnKXzEeqNNyFkKpLNfUAoz20if7w58L+MJC/jOAFVGZxrmep/KEBilH4Tow2IuwaED
R8zkzj5uFx40SCtLRlomCcDOpn7caxM1R0EReEXsAiNRql3DVpjmfLrH1HsqGT52aaL+HYdSpzds
FlJz3h9H14aTzvIyhOQ1gzJfBSKOmrlqmwlUlvytgMaaoJC2uv5N2QsCSxOA83to4/83VRbLtRVc
rFQwlm5Ox29aPUrmRR9FnpHdRifYvRQ3deNoVOP4Iz6ZT5O/D++tlNavYpjhumGL2eWDbDCeRcj8
/Lpc4Y4EozG9Myu5KncWPkhVEH9Fy5K9/2GcZ5d3Ff5O0xGdsBvQZU2dseRRlZMUHzAXhlqQtpih
7amU5VRCK3tLWGgEJFajoP4sPzaH/kWMl19M5VotrWJr6lhz/AtB416KG12SFjXmO6oMoamdiEpM
uM5KpKexbAvnFbU4fUS6I/RZYH3XlsqVgCDbUz/oBNZSt3xvOC+9uy3KzQ1M2mtluEnf9OXO1bEZ
Fzknp9t5znRsEUQCGcDhn7xyLDkiX3sUU/iRVZv/Nv+7sND59gjWs2GXo0bzx1Yl0Tvj+S/tbNRg
J+T174A2aKVjJ3ije+HSRTn1ke0dAnHZCOtPCMFTbs/HOgSb9XsQbwVI1qtqQg4ueVZ1iM3PGGq4
KRUL17HalBrmoN0MFOSCJDxy7g3j5InBcvRqmlk/8V87zzcYdDX1Z18PPvDeJ+kTlM2KVV/N6vas
WR2FAsoZYK4jnWy/65LVWlWz/Vqs7cjlV0TsQko1w2VIUT/JqLYrgIZoGzv9rcQv8Gnts31258C+
i6EmdERJg9iEs581VD9KwyeAqRJY4dFo5ZqE72gZkn79lZcQq4tNHTtpKFEoKczwWyX4j15TvPez
G7RYtGsz3nSkPNUZlobnjC7SddowJNB6jVrz4IcV07WbtWAbCuzznb8QlGo7OjLDTL79Kmh6u6zR
sfciE8WkiWrjIQglWE4Jf/V8oOy+mU89t3RerJSYJ4ddnp1bPQ/Ix57NDIbxBe17Iyd6M4X1Eq1Z
YH0ZWqEK6CSJtQoe1O9T4brLbclDzpwWq5Id1DeSUccOU1B0cwErVPUCvlDYgpHDV3gJJzR3vx9X
FPHsMnNwXsK1oKoRHBY6xE2b2V6BdSv5y/ZqCiY3PF5qcFYs3STWZJzsr4RXH1kEYE/nqSw9DzMz
fXDMU6gwNIq1e7GnoB62N+F2a2Qbz+dg5dibUiiRjQ3MxDkYX+AKZJG4N9piJaoZZv2r7fQQdj2Z
g2nUz7QdyUe69T1ULZHTHURqKmGx4aklKHkwsEDAlD+3PwqY23tx8/HxoElyJiUkepPwVgmz3lyi
dfdMGZUAGB1TiQEABiXnFmmx6EHh49Ui/XLT/IZTp1w1/6w90FUlJ11F3ijGKdyBZZKopuv9gzJM
LGSxH0WQzxsJ5lpNRljo4sZQ5ntgVLMRztW8UZAvMUNGdgf2jOFnqPH5KvszGCWGgsbKMZ9VByBh
MayJ9/nmNbBstUchXGKaRF+u0W+p5VqS83Nellac2Zes316AdTMnXORFUU+Gqv18wHOxFRphnWhs
N4oY+b7V1Z18t2CY34m067wBKNH6FtYqeFT/32bWZiuw2Yb06jzbLkU6JXfG6unFEo8SkIsrEFqv
dweg2g6vMovmrfVqxJBTTzNyGjc3wkRL0kqEabirtjVqYWMJL25AfNiwI8/mtx4WaMrj+GlwQuEd
8FFV/gjaAmF+5XycYJsMJC/10sQ+OBQcjMbvn+rQMKc4SFH1RJEWIYp+AswGw3RQStz6nsfAlm3N
Yz+5ad4BTocz/H78qE2aRi7jU/v3eUUSHToQAOVUt7cHhZ39plRCiJ92l+4rfugACLWoUAaF5LZo
AcZRR41ajMmlBulrnLiyGJ/P0FX5DW1XUtHLav5F4fsDLqVrb8nL1JtLyUtZf5odJj6XPrwDtqP/
fXTArrKcQRNRchlLCCZ3VXggwOCBYHP9hRqyYpk0rnyC0jEP7asXcOPTkJSFNEacPTkz9fxzdpaR
TsnasdpIRkBx5pkPFJzzywTMwDLGWAuH7DtvgNRhJ3rU1tlh1ZuX68vy8Acy2roLkxrbNV6KmCc4
J9n6cALyiZjp4AxaBai4ajfKgBSDB/Uyk7w5Oq8ooYvLlkgq2a8eVf65ca5Pciym0X14JxdZoTdy
ROBBlM+XXq6XRxGsWAqfwkQSFZyygzHUvwFMUNnmm8x3jd9e4iqiUQBEyw8ivO25mMVVlpl4OWRW
XVYAKHsqiS2uV7ESfm67rFLj5O1keTQTiUmm1JWNHCJaGT5brfHoC1xoR/zgrq6ErHpLW8DYqyet
E6HtYADG5vYK1jqm47m2XDKRjXF99WnWezuLu9QjJnsZLnd8J+SUDju2eEBG+qqjAfkUxdaFolvv
LIAg6FGSRy9wLBDjPnrir7QTf1v6ss+CseCa6evKZGy0HAQK+xG/LivsPzq2RUOrzF9N9loqozfo
otpLPNF2BLSmXWpl9KfjF/rVmOUofc++WtrQaGtyBjG6qEl2xqBjwbsJOJH1YyHc07iGVIkWAIOx
xUsvUOKoXgjRc7oZmFZ3TrgRwpDSa8wcftljCmoVK9ytHjxh7chIy2OKkTXRfirnayGXxh9tfq2B
WPcpd2Rtdx64mIdLWqgTA01ommRiAESO2vGA8e/ADqNXIPzZzAWlp+p5uEOIp9j8NyML5+socEwH
mrQkGv5AbzjPM3x7BSLurcozA9Boa6KuMTpXmmi54NIHN/mz1/C2eDfjs2/kRi+PfqnjqPLly/jO
Qkhlvary2qSqoY+uDOUdAgxOVG9SXQWmokZkxVbLQsfJLvcCW1OO24izDUcy/pdPtAgMlI88SzA9
BKIwpyMCLvPAwkke/w2W8U9D7IP6GIfeGIgnx5BURcpIWKIzWFlPntJT4grqKVRG9u4rxjh/0Bks
Wwju7p5BfkGXzj61t+S8DZzTD5s5w3QwgEY7RIM0/ZJAXijK/SQiUjBivE9g0+2oMOM1nTeOn3y2
RlcQYxBs3JZboNTYjxpAtsgvGoZ1Y5fn8aco7rcBZIjvAVNeKetwHKSI4J/kOqrGiI6PDfiPppQ2
F/wlKK10a+0ZsItpU6b3W/c1zVh6UBD2PKX8hSDFmbgI8e1h1cg43tLgJDqBuwHgC61KLIQ+1tTw
Lez6eiGqDQGk2/gH9MB9Q9jfIt6+pBHMruGSDOcDhylrt6a/8mv9nnuG28Yb+3HP+BRuhODXX37M
A1A+ys1qVD+fduZvaIKNOt3FOvlbAy8whS0I0hyDvPwLcPI7H9vp/JRuMELUmC/FiMmKxbnmKybG
YTKwVZLpulPvUVmIu3ElFB4+xY1vtUdoOP/zlB3rRJl0fI1AZ1fDn0n1CJzYMk4ZXA0rXQoqZrDY
S0eLzOEwu0ocXxT6ENQLtGINghgndOBlnekD/XRVdRgkMu2QhPp0nOoSO6H6Dt8R+Eh5CmKvB7o+
GFga0Csk8GeZAqCQKhxsAwGlf6eSWh9P0zlDtEwagkz4mwZOnlTdnIkQzDIGjzzHizhPiIXNHu22
wYwgaFcwPgIdlvtZHzsUWWuJiV9a5IlOu0UKJj+f5wu47YPExSBAF4Vfo1NWUQ0MTtweBqO1PPEm
lt276m/yl5Wn9naAxq3QFA7C1C7cmoN5edVawH10zRbDR/b5TWNzmUvpPcF2uLPiBheBeX7X4GoY
afeWGpLSC7PCv/D36eCQqPLQue+FaEfAudEGUbzUYnod6tDeb767HcoOe+zCjroOqW0GB5FtFdcI
zqrVXNuO9BuVEGOYeNHRqgmiVv0Z8qY4BuDat5+YPCrt+FdxDKH2MKy8f/7LguG9aUVvdmON++io
Q71RiKMv2o+vKBxTwZibruoD6SJK/APx0klcnHmf7xmrkftxCMnlTC7TPGPxoel8YL/VWTSc85LZ
PrPsc1b9sUleo4YRBekQWjiuNDmMGAfqatNmi7X9nTZgJOrpjlWd2acqA+6jcT+NPoRXp1V4eAyn
iOM3lsseVuKwKPGb0fk3LayxfGMK2SJVi6xUyaX5svcR8PWqLnI7qa9/msxpmbw3q4NT+jFiTeX+
BQfSdOMgh2fd3uZ+TTCq7YqdGYsOEv4I6nmPJCTEwc1q9X0uh7oXRPjTRhXxv8z5VH7T/UHbm4s4
hn4uJf4SRkHFnHeE6Wz/tiWGookUebKMyHV1mzh8/6wT830To7He6H/s+WW6AIm3K0JUUTxRBQP1
kzHhTIFfRvO5oPNA5Z/PvmQsbJRMUwTUBWCTSxgsuqJlwktVb+uH55egOFJ/Aj1IYMRQH7tfKugT
pyGB9sZwiyjeU7R524H9Q31s4g6+2RLIAjGfqNWRGYugkp3PekVz1S7kIRuKrayN80wbqHayMfvb
eFBGbSubDgfAW9l+4v2NLoitEYPpdR2+80xxf+qkUd+EGCMXIgiYwvK5avAs9LUgpJejmX9I+/0E
tYiZsxM0Us0KmpDZbPL/uB07pB2+qhDUSyQ29gEfI0o4AKLqgqPM6Y2uJRAL3FILeOh5zU9Ks0TL
ckcZMy9y5L40ijYKZTchJt6OgCEPurw4bAYi+Ki4X7TWCN+pYPE7AgSip7ReLUDOgigxL7E3er6D
Op3rKaeOoDyl8Sh2gtJv+hRBEHLDyK3dgqc1hGIbtpVxUQqkH31vn+LEKTillcKA/8C97j9C/7w5
ZDDc5M3vA866t/vmWWRCubbMvAB23Zv8XunFdgWxFxeB6mZxA7t62Ox4fqgnNZPaIpnfrCA52pzG
um9KsRfcjQb8imE2TLSJU7aFoWmBhAnQoy1ARRoPAvflXXq6YiDa678Tvi7Pln2pZeVR4ldpJtn6
5x+LK1Y36gTrOc/gUMR8LcNFJdmqIiCoE/bq/k8CiSq3J7RaKrqJjDLTY7LwJoCOrDoZfuqBbRGN
5NO1GTWm1G4uUW6oJmc7fnX2q9JFr33Y9ivqrW3rOTsSZnXLDjqoit27jU+zpEWmLSq7WHyLRkdG
GIYWRl03aMrcfYvs2HvbCuknjtTxfxbn9UFFVvfW9IJF8Qcp7LV1qgF6HIh15olU9gNTtyE3uCvT
j5Ta1WQwSOuP2u9hFRzqVyOHyskw6CdpupWbpB1pYobzaYbMz5/TrlmEqp0VvkaKhOhSzSkdPj/W
/35zZhLA+2vnaX48VlgXbTyyihwmSt16oL22Md9vQokrHRvBF162jRV6dSxVvHQ+kETgK7jTZMzY
28f+0m4KishPAr+LnVmwsJk9KIVYKOlsTOltXWYwOZkVHA1CIlDkMMQ2glky1ZlsOBzr3zS+xFRj
UnyMi1P515kJ0NJ+4uZiXfOQLwuuYQG4RYO+U7dbsyVXG24ao8rRYTIYjdXI6UPVQLXYpR51NeTY
soj7EqgvjG2a3dJa7Br7fq/r+F9xSoSeINNNWMDAOQCT4VqTuLs3nQ81aJ5ktnXbAl/7BLQyuT9r
YST7W9J0UmAOBoVIrZZtMbnDW1kVeeJtlk778oL5xg93oVFoBELMfteIeWxuqwR6by+KcZEjSfeu
P2OC/XMT2dzJd5GiGsMvOapR3ZIsOaXBzlVuyxP+7WCipVRubSn7S6vxLcSnfSQqfbMvw4MYXiyE
1LvTHM/zYYoLhJuXYTgaT76VdZg5R4kcJDS01quxcciheDjg5Q0qNz2uO/nfWQlNa2SloESOXb5a
2YQd/+VBt4l7LD318xfV9+LXFTPoQo615Cow1yLVhjjfGrPjdVDxpvH0y02CjEY68VOUjZtWTu4c
KyvN9dlFlBRlvzBvkp9RxHwsd3KI00d/m3fKbpWkr8+Kh/V93XYCRRa5eIseR0LMi0EZ5f1u6Luc
qOgtDoayCZ61YCXLkHMmZ2uVLmMgV2xnivsQK0/dQRzmId8e6fKqNGtK+EQFlaFJXZfs/KfLvH+I
IER37iD+j5U9x2jIWsryFsNRqBx6UZ40+WwfqWYUAFhPE9w8nAPQcPT7jiLyB9tR6htpbsXycJM5
nNv32pEm+aOPR1LZcNZmwdI2IV5u+7ROWdxtkA25KpQOw/vgRn2z3VgpbCQjY+uqOJLbQk3mDGaQ
BNhOWhIF+dIepgnrZtHOsc8iBCfPrEIk1Nl6m+f8DHGOjQuJh9bd1I74wQCwZaQs/jGuh8jDpM0P
md+hXXgADjQL6T8uoIlwBf5vqcEi08G7mQKvrSEHFkKpMbtj5w2CfWdVuiqQVGG2pd9cicwh9snS
YIOYu2Ts0odX0R8HmbOWdHlUxmQEpVMkj+c9gPsCYZHGcP8IqQQiZsh044g2huPJaFNcCZKbcqit
vIMjSiStAnNGpr6Zf4bMsb2lbG0FrqYHqLVXIXYPIUK0cezhLCyfE8RRxMSpyGw6zJ5BujwHUTU4
91hsL6qV8eyswj6WrIRTh/A7E1yQbTCgGr/zWHUZQ5h8NZKrDgVT+I73x/+74KUy9ai50Lc6WIkE
i8nA+bkzIVcg6PM93JYdYTKX5Qvb8kY2MpFVRS0axPGSUnfug6LJmb9IQJrbc4V3p0BRONYYGWV6
UZZHfRGWgZFI95/T8QXRh3hxFRjNp7+oxk5RSpSzYIAAncENpuKXGzBc6zKR0ScKGDX0cmmByfTE
33RLwgtwbUO+ic2DJ4aWeMIeO3q5/pjepqiXKavWmlZfLvT0Pk3P5DkctDSP54HJRL8SldsQ6WIN
MUXUJM62BDlu7lIdAnHPPvLaXoXDegg6DnLi80dJzCrTTlH+9M9YCoVU0j8hgh0wHHKY27sabFgb
7QcukkZrSBvW98dwUy7S1AerMZkqY2AXZctBPbw0sFqNFtfWozvrWscdWeFvYz9arxJWJwX1KjdE
gLi0LHCBcCMWat5BpXX7uOSuqTMM7Fq5ZQdsMHQNivbvu9NbUIVrveBVvAvWdTCPNJfVHfAx9erh
jgqNYcGgaVm4lfNDjoUztgT4uRWyahEzH0EZqaDNcxAWa56wcflbYZrUvgxr7bJvHoNo10CZkGIe
nPeYB2EMAiJmEkfIteDnTSJIltqFAKuAaxdFlf+kEkaXUPXkrw7PgtLqkgii9Ib3FnydTR2Ih0M3
gRwxlqBiqSYF8FIMOi3RF6hnUqUD/a7vEQDtqLOpNvIPc8TMn9nLMbacgi0MA7nv+cdGXXtU1jEe
LmGBwLbP3p4x5w4EEbs05ZrDZ4g/7FfB+1DSeqlu3tpB7CB43OHXvOHGd5zor4k9SNS08ya8cvH2
oOYAEQGSAq8F852OOux1IQxXsVkO2TDjopuimULUL//SJknTiH822FP8h47G4V8qRbPYVW9XhSBB
LhTHisPEkebaqodXZEHZ1PvrngvZ5onBYH6AvjeImbFmcfVwk7xBrGKbVoVz7APtzUHpgPYBznlA
lNDzTPsHdn0N5aL5EjtFRaYQpMEdoIaWdOSRGq0pBHE7iPk3KbBBfgKAHT/kXGy8u6Vj9Sms6oFs
ecNEt2KtuBQscgkrCHXdI1Cb23/L57jL/FTGsUuT5nuNkfrVMp+cc3c4CCFGfjdRuDCwdsJ2xNB5
/mWw8lQA4/ha39uXTnLCHXCrmD/DeHMPmNvf0BSyKpaVpBzyeAOV9XAKbyGmBRkKi0+yETiQeO5x
aLnsfFzlmgY0sgXQq1XXzMvVKFL1wV58LnkxhVY21qCL8vFPr8XpHHK3du6P4Ss+nMEnoAhp7CbF
+72gjZMoY8EwGc56pt5efiW/FbuaSgSH7gv2GOKFQ1+GimAXgPvn+/u2/kyjXGxtZTv0AoETDHKQ
yJg+2IfRYH+6QJClvLDQDf71i6FngZbSPhnZ+t3JDwtPRNMNrb7To4VgeTO1rTwYflnfQCqZ7R8T
3Xay6E/fifG9f4UcQT1YaN+moDQS14oE4Lo0F0MGr0jQQt8SjnYp3LNQfRIMkAiXptSbB8JzOf0e
iiQzdL0iKStZ3ggSxsj+q3fR4ZYQEyE7P5Y673+la1C94ZHfIcFPrXGGzGUkAtdayzkQGaR5YxD6
O/jgI2JwWg55eR+DqjMtrVUbyOtgR37gRB0jl7SzRNmgJQgBYzDx18AuY9fI49lPETIAGl6EYq4N
qzAq7U6LPcXlgwkULN8hLjDSYaIa/eTf1H9z/k1xB00dU8UVkNzS7HAh03HqLSjV27SCj4CMep6R
KSfQnndd442LGWk8qHN0YSW65JQPFhfGuv+W6vf0kkTEbmYE2qRNiycIQT3zqVPcFc2CYBXGwYcB
BU2gAfvMdm7IuYmDnMUD6orSWEjd1GczgZL1POc9lhWCkMbBcXX4haJYWl3WnRTC6bTKLmqrO5na
Ykg0CmMA6X7FPKS/kvWTVfX8Z9VFX6JXRr4Krlb7E+in45juX4SIkoCdCgRnz+SycVYKC6UgNyFX
X0doipy0gw1XoYs/TIQn2nU2skuNiG9phoPK0WeNxo0Sw6z8BIHZWSB6k4K5uQpgXWerc5fmn3VV
hfV2lR5nOUxEBDyxaDBYNU/6yFftyf+pTayq3g6nIq3K2/jACEWaw023/43VQHzbshTXBE9dDkNe
xD2iaaW4RRuD71E2IxZ/0xm/c+IQSL7LklIuKWp9dGyrYZVMEBOxCHbgeJKVsonszeoZroWfAHjF
5DyfLlciLQmBaLaJeclGSSVv2G2Q8A8RjNR++TLzXyKKKBn2ZktiaHf2Ze8McS3H/gF1jgu7l6dv
txipo25AjFkUHAnJqK18NRHx6+ZaxX5PEhSv0Rauahn1xqEp+k6buCOlB3AqyORBfcfoYBysBVZ4
sUCA7v5UnbmZiqIloPoQiJ83NXUKd5jT/VsGTQWyZZH65uEmCYk1GKrLnkZLzjEXsiDYkaqFpEWi
ncFUDVoC2pZA3GU07+RcjDPUNnOVs8Mj41DYjpTyn6LhfbJAYlmd4mTc2092a6xk2ntwhB/9Kntn
bi8S/UWarX538nmlbJvprBbhhcEIvlyTBe7RQ/sEO+WdNvPwWTmIyWHzyrYJU82805qHKSoELzyD
Ea9+oYNiLh8m94h1YXj6ViwFUKsX//TVVjRX9CJiCf7hyptfGpqnvCWGkr2YUbIrYRgWw+tCISSh
hb4BJOr95ziQ58kJXUx7etGbe5KucQGPbd8hHTXTKvn1oUopAXHqRZj5hzH0oRtaGkrqLRFvLe5Z
H4adXpU9inaEB60tmLiWxJn2hxiy2e1wADhpQ4lNDMk0soRCcTl9rcDjEfVZPyu3DGQddi+vzyeI
gaEnApmNz+vZWVHvWBqnn+qQ28lcqpFOJ1bXWyJxhb/ou3IAh7G/Caxl03QitPMddz8zeIXTBSjG
WjJtKg/Z6TGF9MI3jQim3Rm5h+bLAC9IhP19NmZpEedFkrTGFC4rTrajDyix+Zpbu2IOeu5xXef0
xWEryaYgf85aJpgfaUj9lbx5arOGkWHWX5TZA86LHRhSjguz5OrCID0AZ1ijlE2KVComsyeH4dtE
GXimFFexdRgEyCGggp0nYZ2wYjG67/1QzBFghaBtX6r/b1EGN/jJ7dX4glwxpDHGSwmenyaF6PNu
sn1miZdHIPkDhvcehr27PT3N+j9T1NCebEUYTHQR5XpAoj2Xnc8kdigOn4pPXWJVoVxc3zRoDlST
kV5RGLBbVpNZVfPYTsBr5oTFAOvL1fzevfVUlQJXdH2nOenx6nljhuwJP05LhwPCaB3T8zonl/0N
reDkLi/MARdaKkW0vg3qqoKdeflRih14nvOAyfbJYUyHKA6M0QkRMGvIjmQxmJxTFywWwB3auKcA
xR1iszhnAqWenzK/txSuEUy6RGrdf6Bg51+uknMxD0mRirAClUvqeWCJjcfOEQFbSdOJ1KMDOKRH
xSB1f3xYda1dMYlBvmr8crtqD2JGaflq1MVf8ekRmY46FV46b8vKDJ1mEh7fg3ezUMMLP01OkWyV
JRCgN1Lc4xtbBKtq0DfgZn37G2gl9y3U3LZ0sMqq2w8WMnvyPIArC4FJk6Dn5xrUSoBNg961WNdO
7tapaPy12E1kPIx1MYtApRaNaQzrmr29ZjEiEjmv0r+6vV+zyL0jQoBlOIH3DSon5g+sgbb9wr/q
7+bxbc3KSSQTAshFi7xc/SnOjxNfU/zdZ4TYpdw21cU/JUNW0jepfr/1LF7dEAVB45gJ/pKpipOR
f1DBlQNzxX39KD3fJPSpr6KEmHCyaKYqZqkNJ+Mi2ImgUAPelnXMJrroPm+9drVf8ORouqdV5TgK
XgyRF4GZrBz5b/evyftFF+d94eyhY4VA1kbxgeySCjUladCSInmEZxG/nRq3xvLi1Pf//YIcMRMA
c+NxMSZMEUV1DALllbon58jIfRMDYnuCfxf/FjnX5p5n5yr5vCPqT/QAODDv5smecX3GMi+Mn+ii
KTngZ18fRrurmf8JXJburPPETw1HpoInT1DbJsMxR4KVuH9XhE8Lav1QHfvReeMy2LWKd5eLlyBl
2xj/cgNIVlp6YQ0xDY02ZHhxKL++Y34N4NfNqzU8Gy6rLy3q0pJ8Aduf8xCEJbt6DSg4ZRPW7QGO
VKHDEpHG/Ddtb0EOBzJH9Ai0Afa8wSTtsKiuPrLErhdbGVzxFlKQ6oqad9/XbMXctpdAJdSa1a6p
F785V0azXFM1sEqbHuKwcabQVRox1t2D0ImnsteK9aTzNGHSspksuhQXfz9MdSLO1MJx1z8l8Hg7
ZDp1O+842kou/2yiJG5Oz5AzR8gtVqJGw9Ffxcxm3X6VTQpAPniXwyZz43KV7fH68GvAMwmycGgd
Vfx9Mofzowwts55xfPJt6pwEqokKib1Vuws8YGm1TDdrD5uGxguvaLUVjE41iaMfPd/Dg2pLxzei
vQz1wLzjFc7TuPjno4tFCPvSiOP+XZk5EfouaZ81hqUV+i+ehI2RGCC3zW+M7FxZ3grZiT+LwDzs
a0tklCvAX5PtsINXphKW0Gy6v+LFOXG5rSwpG+C4TpvqzcDnkkXuu3Nk4zVWj+jUswMWIW2RExJu
I/Q3BZ6D+m1mNZ8GbUuN5MqKf6d7Uw/v/52hE5Dw0lVRbFHU+qTehgHcQlZsLBE0zp4TfDEPFqg5
xVtiH3XfZCKLtU1QUdGbnvGVMKW9o5+OewU8c67dyXqs+pr/D2zNt7BgWHW2r1cSVJnMfdMYF+Z6
RrdyruLsAzVD8OVSfYnKu1kcDEJChOSAlS1VigmLjhra99Fnt3EGVuyrZcCik7HgPdOZSQVdWPzL
l3TwAwzEPCUWR/iRYEpe8PE4sPIdD9Iy5eqTiBUbc1wf4UB43LQFcYkvqluTnZGDzd5QJ+HhyoJG
6AXJ9ISLcC7HTGAJBh+Ou/C0dvCb8Je43v5+nwJfKZ7tcvhbJ8LE+cUhJWMQ1nENmG5+bIu39W11
8ND323tv7MhZvTOnzZ/KpoDHh1adzURJDluk9ycE67N0m2ONX+Nj3becAycFqS2pqmFDRTuRPA1o
7X35koGyftAQxos2+Fi/VYwfxgzdJUX69e1T919cTj/Gb9SNQu78SyoAmUh2eTe0y+e7e4eYKzMr
fWtYHFBGnb3rcuKqoKx+08+5BMbEV2h+wJypYHA3VqxigzOyeonGka3WWs0HgSBClVlu7JI+/PR3
X6v9CeCrwyp5vhLuLgOqfJQxsqXqHVGYF90FjVPctnnjpb5B6NFNG19a7/Q+D0c3mqBQwzWcLhCa
EmXjFyaKxyD4AReSMGDNpRjxBURsH9JOQ71XrGc8fAEH8BSpUwGn9nnP5k/HiUv2zYO8/u0lE2Jr
FrMBboBgLJllFUk/Up946sk7cKJQ8UV8DCrqP99YE1cDG5c6QOHK5YBakYkW/OqVsyP34Ur1frtC
lSO3oN/1xH6I1p4ug7alXQJ8A0ocSsK6sZrwq7MiigyZU6oRACBzdVzv2dHeUFhStn/MjFiq7Mi7
4GCYHcpi1tsKOa2xpzhw0/kLBWG+aYjfXT4cALeDGLOQMm7KhkflGTVPE7GInWSd0syjt8XAn+Kz
ZdiSAWP6HEcrKLJzDKTuAiH45XNOwxcgzVDTYhwiRJVyMvrMWmxuTNIGDAt2GeeQ1hO+xKJVE5to
shoWGzmHAVLcDnXB9UDoSH3yUz5zzOw1W+PONTIaDV45I+CMAvYcsEytEYqUN0V9y+EtwKe0/4KQ
mvWpLD9KSp2S06XWm1Y5ovIjsvnzRiZEmpmC9XX6oKu79+4EvbfFLmAOCqo3gX9H1vt4VqUwX/rU
FIf6sdE/L/fQl0YQJCjrW5XtmJV58i70pX+vKaUdLrDebo5IIcSSp3B0G6EXbQWFr/pO9EeE2NRp
xW48jrq3zc3+EVjuX9dn42T1HGDcv1zodR7LLf0rZyV78zZgxusZnA4w8QpiGmgu71tp62tKJCfB
FyIrfFCkKILY5dCmCRkLilrG4N9x26ATNlUWEQQDzA+ClZkmzdSigXcTz8CAGZZC/Kmk4HfJz6qx
KlvBwBT/ZAs9HKDnktNP97emR6palhZqtzlqKpLqKD+zcQLD9gln2MxH1PR0sIPdMaPWy57N1gKy
6AkYn2dAHvF4M2DkCMIehuQP1lbBlFpxofRkj/oc3qLo8Ia+rPeh7aDgmL98k19Fp6tbixHVGdss
AKweoQ3iF4qEFFGX0aGbh2Z5b+RUJ1ojLyam4ZYN+ZSmYsn/uQVTVMUudmYwSM7tqK8oq/9wnOUL
mVExTdkybONvIcOV1OVmsS+FlpLmuvzFmFMitVfsoukwxJ1J9J+Ywj+CndqfgdBm3a8E3/PMeNUM
tISRVQ1zRmLg1tFaSOonMGqSB5PF/Sfsro7ykMgrWZNtv9jLg2SHcqEkmjlx3/592aGh7ZmCV/j8
IDOm0uT/NEj7f+OfwuQiYaH0YfSAaMjvdi27gdQSfSYkVsMlHJbVnZ+w9djvNRBr5+JyWsEXxtDJ
9V7FjBh6X0D1OgCrO60i2BPcXKKwjYl8kMHtjtgXpiaowXzxhTb/ffzRZ0PPLVszlz7mMmsMO5Ug
gKXavOdGBCHdy7hZ2AE0dJO3iWMk94WodVUz/BEh1j7TxFOC4kkHgqemZohcJov0Los3gD1aG7UJ
x2S5Pwi+CStAKox1KVS+d8G6bpbfMdQitP/w+1+EMxEqisy9Klg8FrBLUemyTssnIxvATgrmfBtM
DAQer2c1UNde2M+89KmnzBfPfCHx4HY2lvIMKjsQXWV3HHQcI3OYYVYoWKr3m6KqzEaA88YssNHI
Oo2LDW/UKUNkgnMZR26Dis32xLOG7q0RjZDOW8p+8k7rkP6xrKAt/RQNFqyS9h8o7mH+o/4za6ii
+8bDrP6ZRictX++Q8ryVXE93LVjTOBcES8S1RT3gs+DUEjqwGEbSBYQBs+s2TToSTfH3pNjCIDQl
0DczR1vLTVuBjh6jDxiOSTJaJfFz2KNMiKDMFtupgdz+sW6IS0qt2mIE2M/4fihUTKFu//xXw7YP
Q+Us3E8LdOT/NrtQVoznJEdTeQQHnbzy+0L/KFIBwT+XlUOiAKd1nUIEG8GvpSRBnvMeuvfrIC3s
iBecUg5rIRSdIFkrwqkKvGv+0vUI86SDpMFid8N7kQhDav3rGcjrp+wg1D/yGpMKlXhdzKSb0w0E
qTewBBCzCyTKZZ98KQywzj4w7RvDGNT2eRYaJbMm23INM4JYBGgpOBcap4e1Fo46fdZMSDTY21m4
xoIFhmmo/sPV5PhR3Ksnecnc77goAU1t+jQx1ce+O96GZZgUhEU/ZLkTbxsoyPUh4OIsuWChFmvI
YFuesCseXn9RI+Sq9KHpfLhLtQB8Pdbs+nRnzvRpQ6Fq2IE6/CmKUr0U27xtxWT4m8bwlfEUZHrD
vY4nSDRA5yO4uuuM38V5Qu2hKFGI5f7Z1S2Dih8MF+eq8AVzyetGV4SUE9cekQZj2wZyKCbX98T3
Yliul2lZi0ptIFELV7UrDoh/RvZQ9QKNsfSTtJYZiUNYrtjnrm+1EXRzzmK30C6y1TAin1ySm4mA
pA/21QStLeMnl50OVWNiJjvtK2PEOefMbc6kCgdJPgFG30wfcIMa4PdBXXdC4Mow3wk1GD7zrf7N
uGMNDQnFYqIkWOWmUvcOVVcEpnkakOE2mfygY8p0HvScCT9g2jZ6NjdKHQ+5zFl72RaCP2HzJyN7
hnEF7Qza6W/k0OBMyOqxOXaJX8Trpv5Lc+Cdvt6Q4aiEEDRSP95d+dDjjPc2lUry2ETCHLBjqWqb
rw0i574K+6ayzkeKgZq/GUseNHESj0vCjdJsciS6UbxDOhvYQVJupVwdXp1xq1Ug7bj/aQcLvk20
+mXR4oFekLEi0u5/lwXSF7WUATOAREqeO1bWSa4zUmLV0D7AsEafy9ICUth9wicY/7DCGTgrPF37
SpHJLma8LQFXoEbNCuBxMlZvPEaH3jpvI2DjcZtcZgWubrWvUw0/Z1VFGYYXJ1hMZoTvuQTF/Nv1
0TwhUPjg0l5NCpFXdaiR5Oql2I4jq2173fQaC5w87PN1t5j3OGtTZE1Ykv0dHAlVZ8WQ+joQcafA
FmNlBtr91JS2mci7qyJtYwEtEU5s0MzDdPr81hDxhHGumjEjXYHwDlu5FUE4DAxDOhuIgU3PmoYB
xNAqB7xFgygV/BuKowJLQvADhtMNIBJtYoZOoPaM1o7a5Xjeypi4JFkrNp1aAIl7dwUfuV7sG7Zc
RGvaknBWb06fH/3TQduZjK6z2u1FDa98/GUOgZwFF2lEit3KtbefMcHyd6YFhzMULwnSATfCVv2x
e6P1hkCqBHyy3Gi32wX2Ki15D2cQ4Br49wE/b8QSFuL13yPpj7iUMTA1XydRTwNUTdmye4TZNUVF
8y5ji3SMrm9p7FwiVdT35E+FL9fbNAMN+Xejv4+6aRyaqHBBfEwyQP9vv1e9aIHl4KT0wdPBbfqn
bZfT4xYOMoWiH1gRr5Dj+j4Hchkx+D0BO/DRNKhBtFeQegzJlIKW8veDvyk4H1A5UQJODCBOYSQd
57LAP0LFh3Fe5w7/yVS31HhiuB0oheD1Xy7p86VwuyeA2mGmYz14KsoRtXHyZ8gjgDII8iCV4C//
GEKH6DyQfb33CoWiXQEopBjUOWKwX/GLotbyW3dp8riya6V9BdW3o/3zP/acOlZBE2adhb4Y0FRt
E+B/ZZwJtZsfkXlCKysbZspxgt6fgtV79LhgVwSeVHbNyC5XzZitK/4Rdtx4PX4f44YuGW5YJMmf
RSBLEoeBMHFZEKS3XaXX4V6kI4aapJy/jvAxnLVIhPk7cUvbLCcXsh6L6QI3TUbnuKF50QJNyTBW
UQ4MUrJv4xdXpAgF7cp+PLihyk9+2bgzjIe9p6L4VvqRKmt2POfNYgXAMqtKJAiSbY+bBr5dDQLh
uQsdolxSZM4ht/cPKH1tDksOzK8r5FLaWrfaH+IH8td/mcmydoKFdG7JnfnZD1QNcsaJbrLIWAcb
qRkaY63wNek+eMBhFMZunAYNTtNTDVLRJXPBR5P8JGkNCR7hcJIYozAELWC3j/1YGUUrRwB9eOBZ
hDGj6B0Ez7U/4sjuzJ9/ZWW3mrY7VookaCjjvncId2UMZGXE7F5LeRgiJkAqputnVGPtD1GRq5xs
1C6rfwUKO+/EBac0jOvTZT/LbEFAFcO0WIA47vmxQnGATMbBVcbftwViImJZwZqYsWWS7Xt9zock
fpmltGex8reM44p6/HhusF0YsrracnLyq/H4E/XW+jr548nA6sPDTZfpRBRCYc4Hv+aABSHpBhhj
Pu/2Utxbnjvc4toetrorSMlmXOCMMu0NQ0cQpkU3DzIfRdRPaRXMdD6BMbzi+WzCfGsL3ER1NdUT
tJtHqto5n3FpqAjuob74StL9RD3FX5v7StNG3TxJ4ChxnQaiSakmap+k8mvdEcd7409DtJcFw5JX
pDLkwEe5pUgNFSfC+kl4QuFXqXMhKP/wxqEw+Ae41ozDHbjyFobBPInziowDumMptMjAeQ70H7+i
OQO3nlkyGBurP0MkfbzmHYE0bQo/pWcFKB46ocoja1sb9i2/akh7UpqnHVLHPwETK30BekCG3kSF
Cy1K8B/XvoEK7gshOZh42jVFQbGge/6KCumPHch+m9g1XWU8j7M+08yzvgXmE1LX6pcAVcQIeDh9
YAzM9ZNRTfKaXLWRzir8jyJh6zWVP+qv4mhfqklY/ZIwZ7XtqMOhQ2bDTAy9f/LobrO/5udRZH0Y
zda+MOCigm+/w4QaeH7KXMvNgLP1YGpvwbSfpXO/iHwkw/RltPk//qrUmsoBG9lI0ONL/7gUpW9W
uxZEJuFlfV47eknggPkWnCK6xGeiRgbf7I/WqmHvf3FaK+AkfmJ24qwkRg2svvvtH1PyxIS6aorD
dAcYLAv5dgCC6+dD6PECPPMIVz+FHK2hSJ4TadTEJBBmLvdHoGp7eW3JxUS4t3wVcZUVaWBxwxRh
tfc80Z5YbsVyYSCGEW8x2aC6TfyKiEOURC4V1NvEnwT0n1QveNsvZBnSAIFRPjJpCw92FUksfzEy
dnJLFUcwd6uhdiKtE1bK68H2FDj06aobQFQwIbzHzAI20XPXNWxMf9sUytR7Z/+6Pqjy26VBI4Qj
KP/Ezp98svDOKbPq5j90Wn53DEySlSk3X6gREeTqvgY/bbzFZbevJykbMfKS15LbaDYZYdxPMXs1
bkLyRoVzEHdLmbf6stXE18zehVZJSOAJKa9O2iAqZ9V3pmbDuzClES/NWRiWBTPwJ/uBArEQdBue
h40EQrP3XTeFB0Rd9vScuzQwxHfdJPR+81yGerLQjMxVe4AnST/JvYq+alef56FnszZpmYOSwFgN
4NxX3V02VO2DoUI/vTwUh+o9jDr0e+9OB5FLWS7PQceXajtW/dJRO3PIR2BjtqQZz1s5Q6Sa72ox
92zfVxQTn36pkNePstmb6pob7sbCtEKUzrDywpTj/5q+WgsgizQhPb+E5p+AwrDs2YpROes/2bvK
DaovldmobjZHgjK52i/8urXTaE17kmHDB8NP2eI9Kq3F2zSUx6KynFntbJB9DeJQ6OzprS8kfcCL
imY6lo2t7p6oVh9x8AraoJAYaIBpQn+vv6SZBmxyx/RfafSIjCfS2LF7kKC61+yhiA46oiA4llPh
WuiGz8aytmXjdFo6q8eCdgSL/W99chrYZXhLB2LGysH8DJlYdE+J6S/QwUbRgchkErDAYnauwkon
amR5+yM2E7KnRGeAxLlf9juYQbrL7oNOl14A7s9ILAjmXZfyYydu+ppJAbaSG/NGH87EqGvrDbz+
G5MFUT1XoPUYKsTTwOMevvhofGoS+Li7h3pS9zi54Ox2IoSoCABe1duTiLux9So9qNfbD5SdHmEO
deqY96V3EQqzPAF7vfZeyQxSkFn0Jkk8oZFsXnNSOa5RprDHvW7K/grCjck/APHowySmifhJubx1
lKuM2JP5ltxBVI81wT3HwvB0JhzegmCzbfO/m494UCYqi2rK9URvv+lK1ObhGQPHzMpMkzIp9EN2
s/nqBNiErS49Bf8gS1CR9d0NmxkiGHuTLnnJ0LKJhKeXPcFsj6JJRPGRhgB/q7MiJTVjv+NP9tgl
XjKyYpdq1BvF30ZLD+53m3CxTZQQIRevhQrgj7beBtZ5jXmnVXjUqSs/8L9uAkZ2BXn/Ag9leeFR
iBS7+dxtOBoVmtmB16ApV1K0AzcSMLfV4CeFeB/5JCVuVYaN6F6nK5lC/9Y5MY1J0h7vh4LVdD/f
3tFueAoz2jcWD01qTb6IMVxc4DGw8vxFbR/uyztLUBDRnckQbTcZxSls3zLkYmfebmMXaMnZhP9Z
2EfCSDj+F0lLPC4bOWzHnFBos9yMyaDPXMqogcIXTs320L9MaJPh/L1oqIqBv0QtOiNu4dUwqreb
1J09SonfKmimV14SUcf2eXmgudnfpcx+D9SUMLB/UHa2o8Sm+07gAX/2LrjkBSUcZL/L0dAFmlsn
+9O/CuxjwG7f9ulUBVcKGipmVQkkOs0MWKjHuMBU2N+itKCT4I6R62Z5XERD6mwNW5owOFt6k1Je
EfWfTSjGaU8GFy+I+3S331VWbAe61X7vASBESB1eYzpx9ZMfgRD6Gryv4gy7YEvrdZy0oDtbhL5a
GaYQNBEdjZGmBa0QW8PH6E4LNuSG2hhtudJe9cOetJDgnIUmJR+9CJJtnPlLa8SzcXdw+zqiefP+
DntfAyO5f/t5eaFVdRQmJYtq1cvXe2QQque+UG49bBoW1zRS/31eqXP458ABKvU/PK2D9OB+0Eds
tRx67n4TyEdzT0jRN/L7p8thHmRKvrkeK14G/qFzPY9zwkiHds34mZauZ0/QvZBG/lbsFCSjqWwu
b6hh8yV1Wfbux3MXJ1VLFK0+57OISGETOwhfRuKBntqx2mPkfpao1V/B7AP3PJikmYvzMN0B5lmO
5zNV27jzl032tfkhHhOqPtt5hixVYgekum9yeZu8gpCEyANmJs9+RtmVGo8/dCabDqLtLVtnwpIA
uiCaFczfeRJC5ouk+YViUNMx4UkP06X3hcjHTrhvbAW0K3w9v3W6hEgCeqmfleyqrkv99W1utJEi
3ALEx4ZACL16wJR/jHcB1fg0LC2tuQz5kC1Q+xxnp/kko0Mfpm86VOGPYPv7rE8zdH08sHt75OKg
EhJULJ/86zm4kBIq7OW+rvepPJsTRAIwIxAK+aDlLkZ3VXmN+7aw2TEmo0iGF6liEsh4J83hsMzX
Ld1503SAdGn9R+8o7bOsr5I/g9K9yERbV1abbxIvxBaorlOgNPxNaj+o8GyJvLNqBjhBW3IiG1XE
MwSYjauTmr1Mw/ibgGESelJVqzwDAzLyG2rGKICW7AeQU+vKAAX6LqT6kxZwebRfrBX/3cwA2/4k
0KtdAjGPjyYo+E+tQ46k21GP7t+2AsXMZSJvENvf4ugG7bKUFAYXoumhSZPDcSyI5sVHNGhWZoLP
GXHNTdVLGPPZlq0FnHr/YcdgTLZdX3VxUxbimeOv36WuTqg5I82dr9vZDhXCCEW9525p0HyqUpuw
srmnRSd+H3GLyBWWeRej7uHjdfPMMXWc7yyZickhtaXeyeN9ALxSPbedHHWu1w/Kc8+BTxlQyJzi
r8FOfY9KQJmKWcOc0PEQkE+O6wPjZhiPFINWDGgp6YEcPy/DdNKuUGeqbCpyOa6JJ5YAkIRAfMqa
trFnY/9cz+yYM4FhIASm+ZuxvgAcbOOOgWRP6GiLPRTrDwV7nrlEMUUc9JujnvBU90Lf2HObzmg8
Ghlkj6WN55IBzQZvESorONT2SkvWLXCEh01Zjl3A+hsph6CMDNpuqWfX3BwXfdLTHNGydGtKr8s6
IAq64vOUFRek9WvzcXXt0yjQnRSkWWRyUXL2KtOCvgpXG4FG1rQdeT9ycevIkNdZA40Sa0F0zonl
417eekUzf722X24dJtNMIdF6/ZqJJdpd2qPkmBWd4rnbhwu8RJaAJhhAH3KIC07evVknWw+s69c1
4OS+9reCEAH1AZldhi+hGB2oHCcdl0xcEvoJ5u5dymMGiS12BGfF6yUTz+rq95y5aR2Om/PRTBOh
ENpHU7bbjLPu8nrS2Je+QlAvGvv3kZG27HnTeLyhOuiBYjwSWVL3oEgbtHUP1OWnuCTB8ZhX2Sjf
d3ohbNqVZyQKbx8ptzzCVP3dBdHdOgz7Hv3jwOy0NkN9ec+DAXtmPc2QrHvlRtPilyQzmANo9kpu
OWUU1j1yqzdIfU3801HdwlOPHUhk+wtJAYF6PnrfoDHTTC0lNA2e9B2PczvjGPSWcFs3IZ2v4Jf9
L4evzq2+xEDQlwpX/KI+Xd0X+Tgv7pV+WU77hGY+4dLPNUMepkAaVU4Ty2YNRIEFj83VxoDjD8YM
Xb0mBC5qdOcfUAdx9NtAHAdhXaTqGCZFLKVOngX1Np7B7quzd6n9rPe7LomrZ4IQsoFh8SjIdvS4
pMf/qHysPzEBUlFXSgp5CBd0JjJcPPzXehINnMcGZzRe7capHlAJwxUsPFy2dwUp3F1OG7kRj5+b
gYy6z/SrCKDIuvAYexdnPxk/Eh1q+Ja89PPTOIr5u6xGwpZdz676T6ex06oVZFbHJUqcbWI7PUfX
rAfCWiS+qTfJ/Ui0xzqmjfYUeLhDWOgEPdLZgG9Uv84YXRyshq8VG3zTIZa+nZLIcZ0crV5jE8Ic
575xWL4ESg/iFK5VIw6qcDXZg8sFcldHWxvU7PslCzD4aOFHBTn5Dhk9vG7ohkYABce6bZNb0JP3
TiFUdGnCmGia8KP+JabzwJaFPTtgmS7XpCFY3eZsP96mIpVb24zMEABJaLk3NNjcD8+v0OsDWZ/+
TUkpomXFtpolJhMvsNrGMr1FZcwyMJnLGkJz5giZsi+5JAbvDutejcnE1OXyt+soC7RRjQ7trdqu
5nAjauUliOQSrslnENGsncpvKed6vnRQ91reVh9QSNI5WgD3HiAKV23ndxgWnNjs1zL6O1g/B1Ja
jMOT5EdEnAA5l2TCR1kz+b+o4yFI95zxCbH7dg+bCbyjNWEtEyKuPJX4z74dJYY1GnSJUOYzN/t2
eQAR6CygT2T4L5JIg8z1jkbxxvaNZSZMlwEhAGCrupYS9HnBuRcWdEUC6rvr+DB5UWajVqY2Q9dQ
MRWAY6znykm6YCQ1fxTaA1ZS9vYwGBmgUbZRSravmkK/2eFM2SJLVgucjH8Gp5TQPOSjZc2SvzNA
0Ox2Y0AEGtJXzfB13L16a1ZIexZTxn/PvZw4w+M2EC37q/7QI3Lg5prTiW9eMalz3qyH1SqVXsat
4aJZWJN1Yb0xTjMIQcSdnAxAZaiVhdNmcVWd/f0pwxpdawoFHcMmHVOF+OtK/+XvoFhMiqwAPye2
khVMIc46uWxEW7YnX9t8MPT2wXLN9N5WgWWkZiLZdo/AeEAdzzup2WVoDOsvP9L+WBCl+O9FQ/I2
GQwT2hfyKZ9aGqz8KlbKI41OGU2AkMhAqFtA/0JnBqkg5UheobAJkUM7g4AIp2ex2bJagAidCMAI
8+MLTuBSlYefQExdvLsU1ZL7bEKvZhMERiudYOcb5xSQf55SIK/fPSaF3+ovJpS6tQEYjgOz/pi7
7s+6OeucouMU54+bR4gAJyMvkzXHjewqoHoYBUC2QnOTgvoDIjN865cYaPxEChXnMksMcYZvx2R5
uHDkBO0THh6gG6eiXwMY7sxY339NQwH2X7V66/552moDrK7pVMRJliX43BxRBIiBo7Qo041SX4sN
KbHYayVcRxsqXYRIsLBH79UUZ1G/uUVPOF5Radwp5JLp5s55fRn/bUxqtzMFBbrPbSzdj2Cfy2ld
DTaozQs/t3MlLZrd6Rn8a283OqXXopkhRrY2wG8smEMq9/CKYF2Oi3F8yRMsec2ZK5eslEjTIkxO
cJHI7Vwxno4v2KDJiqPiLWVNJJiLD8L8GqoOr5EW43y+PcSbAYW1rfxvdtCAtJq0t5Glu/75ZBde
IhkzXG0IJ7HvUEwgJhd9MucQhmf7ltpWPY4Lrmo0JksZgDMK0wwPGRfqaD6zd9K6E5ID/44sZUxL
QbNMCk6WEd0s87sqjzc+QzxHlpPQB/anVlCdyj8NDW/jpW8029CXf/e7PEqS/ZsSxzxOqO0EFXSo
uKfzqZR60tLedVNNe/STc0u3Qut57Tvvif+Ug5XvsqnplfoWgfTZyuVPcP7GEe2MymSZmrUGY/Mm
nlXX/nzYlbPaBSQk/m2kmIkKJwC7nlF0iKTEUktw2uJ8wEAc6cHT46KPVP7JqT5TsuNqJgL/DQaU
nBwS+ECTCgYnoWnCtsQoQZG/L88ihK4RCvIbxPZ47mA4HLH8EYddOrWEQ5G36qGdTRudpBMYk6Df
EkN0UVzDqiQytlGRSd52RPL4C/kxUxFEyMEMKOkGA4bJ+LvewtI6Zb75QjGt39e5GwME29BboDdb
Ov938sZrWi1CLU0Ciy94Ax6uGTy5zB9rpbCHoLRPk8Y4TzjGfwkZDlxse+T7t5PkfSL9i2Ipg201
RVzxLishVo2uAwLVRcwBOPw8rXfb4dpS4m9qLlm3MEAVD2rRpCqL72Mo7XUN9NegP6wLJJrhIxCS
cEr8EKgrMpY+3AqHigXLghACiXWYuEpjnve4tcayGPaUtgj3Fb7Bpv2l5dYy/mEDmxNcp1WwyuPg
5d7fgxFjqnUp8nPOIzmbWK/yJ8N+AoWk6e95zHByZvciXaC5zARd/uHEF3CpSC2g2U9aFi5eAJKm
o46Ci8jGHZU4EQLbt+VyF0YB3j57FM5QNk8zhrNt+xmzTCSjI5G7cwVGokzIjQS8Y8s/W0S6rDB0
E+7CcCSlq7W3D8up1TG5FVMTXHMIZUkT3h5+EldmLpHGNmdrBCiOnpudYAopaLaWGDOe8AAtaglm
rvUG7k8Q70gizaf4ziJ+Kj0Et5+drxSQ6uiwwJtCD0R1EQA1gP5t9skEXLKAlWbOQeGry/gPqGnp
SCBnCjv2jwyrU1HuZAdDHRk2dtV7F+xviTbVGwfmEJtk7Ajwj0qSEg4DqlwMkk60XgEgDzOh+nzB
I7bntYwiDpJkCPpKHlM6O4boscR9X+cfAaVaN43GdWDnjMQsckr5bJGibfUgr8ZTlkL6EqKCX6Nd
FGOj+3ZBXZJnNEflPzRBaMqjkeKLokJqrHYn6DkgR5w2nppezoRNFO4pTvgIYlBsuajH+z3SepIe
Cs3JhyzOWThgBVRj5pnaP6MM/nvXG6YY7NsT4tytTeZqRX3bmCwMfCY1XFlWGgvFS5/Kk4KL6CiH
qzhvfrSkYfxXn0Qp922bS/Fk1U/PXzfqsW5aDUG2/rsdHTV8fubd9rmtkOZ0yoZTAHHRCw7ZfLVB
s88xfiMsK93bfSb5eJs691ngGoJeUxL+06MFWmnsG7CcpTjaG565qTxCfYahNz/JaII5OJiGSJPc
grVlJcT7Xy0oDQ187LsMHLPvwLn8ecEdY1ltDKtPHCOefnCWzkJokWOOnsoasOBZA3CEUj9chzBh
Nti8onn8vlYDB+k8cudbj51dnPka0qJ8/Un/hcaRa8HFGbXwOLgscrlB4lTCXmbvQHXE317GdnAV
nmFljUITdjWxA9q4bmk1Xrb2bjRE5kfLraswncmQkTdeDcGyCQOqE4NUUhsmNKb9KEvhHMWCuIsO
EUe8+L3+0JVPJd13wRl10PIjgIbkoK3XlYfVADgs4CCG0IbhTDjGLzPe9G7PmyFUGO/A2KIgdjQk
SCPOEtNeIbnIXcrAp2ioGfxSdRaY1R1yeywzRbKXKCGqh3mX/3QdY4DNjBPvSRbPuGCGHRXENpSI
SBiWH9wW2Z7aHf4tvuIJryV+ug+dFWv5woT3FhDkTnGw4JNfHyzgh25LdGWc6KTtVKwwWcL/dtot
4UNJMcAq+BAVzDreW0vuI7HfCKx28uKy0USdDx5Dcl420Z/IqCQ92TiKK18sZ8X2+i2pO43Kgn3m
WqtGvgSzZZYoYytHQfh4XBL+Ewc69DCdc8Jd7uWRnFodH7TdJVpgquBZSspHfmuKnFmK1D/8aOVt
aap+UPmplIw7PbJ+WFIZhlp9dL7ykDywrcvNkeqt6sF1m/X33dL1wAdsUvCtWIxWfTv9x49h3I7J
U0upwOQ7uYqe+PFsNxn0wpX6dk4c6g6k3ZLmTgwn+xMte4i1fpCM3oB9Y4xxoozPR/CiKUO1sxcJ
AeQj4RzkiBaC6AG3uX5J1Pexqrl2puhegyIPYsc1B9aqELwzzYT2Fx3X/mulaGJ/jfBDXn4QjRjg
t3ZiSinAaMt1lCjDlMRy9NgZo/xXM2de9vOde+0u25u18OMdweE0M+OmFLYAYA22Yg8tT7WtVaxn
7WJcjzUwqCX1J6Cv6jHnZWkBu+HH60bRx4V7HzaJ9gCTp//IVzXe2/ToLs64/2eQ67Irx0gWZB6l
uKlYFwBS6FrXYkrkjK7SVgJ2+E01TLrnw3DEMFT4j6o7Jf/aHY+Ut2xfCdlYrqOkJe92fJp0Y9mT
feDz/Hjr+j7u1nUHCKW9/kNdNcLO/BDc3voc1/SjpanKMSuQ59DaMxZb5yvggskccH3FXPkKFf0B
24aOna9+AkbxAj3Hkzx+01khDcZQKnZ38rEguijqHWmeWdgFLBHNn4ufFCB+/tm4pyUEYbxPC2ZR
ZaWV+L9MDxjkbPvNA7ljkCdifS3JKeIy3GjroSlgJyaIMdyOu2O3YHV0YwYcQ9MLPskEA0lsmosB
nZWUVJnLjDD+eWEK1tl/YPlZV/Pb2KTTFN1TmTqjEOBAz/b9NSntvzTIKjt8xqjtdxRUF5PAcyzI
NltjxyS7FvWR0ziDHPfEwFEJU3Yn0FrLjC+aUlMcjhbFfEnidNTMPfr6TnCBqxmRdWvQm5hn5R98
6I4Pww6ILKI9PabPqzocBIsLhUn7UPmhfKoROYDmiHLIGFaSK9rF7w5B5tICQ0tRGwoflDruXQds
pt+vgA1fmruaKji0f3+JtxxGgnwtXMtmhat/xwV0fxw2LLGT5bOb39GAquoIJ1YhfVMPFic6rr9T
UQVwnocjI9iHCgCONimPLrhSaUxgEHqCsbs7nucNFYA7nB7mGm+s0njMcIh8H+mRkKr2EH4WuZhk
GfZGOvUh/TcJYeFQvY7v14WhcVylr2bmS/Bf2gQV5yKXTZjspk8DAYGB9TkA4LW/qbFo5rpLwcz0
/ylMwkcyvM4ftEo+sf8W2dLy7xATj1CsbiR3/PEzKf9rcdtZ0n2tsAiwLFbjSUPEZYs5DFprUB5q
78LVoBNOpTheC7luqCbukhWV66U192TI45RtEO2bbDVLehdAdW8FfkSxXj4WMfp6sDY26moGsFyo
9Vw8CUSNqgqRqibpGyZ2dF+O8hXPzIrIW6xxhWBOmQO27I6B65tFRIY2WpmavdrUWMU0GuxVkgvn
X3kDNyhpjYCDZ/W1XVNMr5iMwZzy5/VQGNPyIVBDpXpL9RG9C1t73UnqWICYpRV+LTCofSKHj+as
sBPtJWqowxUkaV3KR8TKACcfuu2T1sinURaUGEU+ysF2m3tQrPWt9yLPr0/Vk5xnizdsbxDNlGbV
IumgPIk0SH2YPOlLoTsgyyTYBCAPcK2s5vw/uDnyiioeDZqNP4czIc3N7kWa8BjZMAM81X71PXLp
HcoPwtwIYqbXCeQktVPHWRvky6Zzv9VG8M2Q/KHoXF/FJQhzdAE3MsDmTolt2U73x5ePP2ySMJb2
qy+z0Ug1NuDkjfBGauHE2obOUHdFeMElIZ+Xjiy53iRLxBzfL1oJJj1qyXOtVDl8ohPWzowR82Yq
XqFbqbfnemo4RFvkz6YVXVpIwiDZK9vhz1rxxN2sBDhuimJ2nRgNMi+efbX1B8tghN6vs48grqLb
HtV11OzSU+m70EuTcWzF+v/DFkbq+yLXoNOHGoUHvN7WAXwcygyBX5hPy7vuZZWwlsUCRwSgqnTN
E7ndD7282EYWUcz7IKtbYEofsI353eONa9e5CnFh8sc3d8F2/QTQmhhw8hxV2R/7rNONFUotGa8K
hEtaqWBXD0q/g/6wK5VSnpiG9pgj7buj7Ck+by3qrw9Hz8Pbmd0JOscH0+VtUedc/R052rqhVP/r
piSbziwVBeyIVJ7OZDjfyBlIflpdomqb6d+x13fq3wpeHTq1d1DSQx0HvcESFVOUhQa17VmGwXam
4OSlXnr+y++vKBwnIjwv29N6gucA8X1CUNOgjISI0l5tB5Vvyxfb+SGb34cxDKd3tq0eDh1u3pzd
m/iNMXXis1jqyqbumRDsxRHDfR+O/EiH/ylUyGu48m/GFZesjFjZbg0at9JdenHjClSkcQLgGN6n
ioIe0uBHr9UeHgte6bQl6/1SIXJFWNueApYzZLl+97oIhZvG6/QdhjtJhHzRAezI7mMuMf5DicFq
pkB3xUzTXFoB39W6MokBLVVe+ktljMWoAbmzBbV+rk4fq7yRzNZ3BDW73jaac1U0c5IZ1IIMlSrv
8z8h6HzaLgz+oo+HDVqUzUZb00y5w9LMbI8f+mzrRcMFmzjNaQNO2pIvB5fyLc95UN60LyuKl4a7
ASEScJsbdhtRHy+GHS/qzZgIEFMEqYERhpUO9PozwM0USI5+1HnqGmfUWjKLWLDXkiRhCasR8WnZ
hUsA2P7OaTLMOLyM6BBSeyJTTNlD7N9wQeGWhYrPwDJPB9CzaoXnFGk4yBsKIoGDJoEJ3ulCF6NP
NsTn0YaZr8SAduEByjFM5q98GHaYHCOx0az+Lqa4IfaQK5KyzZtMeEmnLal9xW5td9vjI072mla+
W16GQM4Ax1YYR4GdhDoShG50zI5/xq4eNROhlnD2Cn8wo1MfbAPFmBokviZB8+m5Sjf1UAsPpokO
2HpbewoL+Nts/FWQSlronzxfQ1H+zzRGyk8baxMdv2wkOTOUiEeajU7WXo4RLzpfEacNSw7tZECo
R9uyMkvNBBZj30zVEQhuxoEtKwu94lQDLGj4Jpr2jSbkhN50uXJi823MV+eUHqIP4co/koTBQDeP
NLdgZ5GcIUNqw/XibaAZWmgsFJXkul5K1OAYRK274nRhs+qxhuLcPzI022sI1aljWVQZW0fSQDA0
7cfFtSn2Lne0FKT8o04DvvXqFGbe2j7wKgcGZj2GktKXL1Uz7L2oBwh4kNtnAmefYRXeLRfkGqx6
IYZLPdHYXAX9gQCc3xQju5Y6jJaRP4RfIQkO1Tm3eBX6cNdCKsg6wXhiLFG7244H4s5mLvmp0UNu
cl+aL2PjaHye45wLed/YIocNHi4Q4RrtqsXpLBhik8frBL8yI7RQwwRhywe+ecEafAs4sufxp2ct
1X0G3eDEOFrc42Jrdvpx3N25VqoNjXrGMS97G4BmUOSQgpCyOyQxN38XY2mSRnMrBkoib+f1iaw9
AkHeLs7plX00hS8mUpHD+6ABnNIetL1tzeY3BYGPTXz8yb/leZS5q25W5GSGaBQjP9onXmRrVStG
WcK7OY7BfFLo3SPeRIBjYQhE5u9/+Bfa9bkpOG8bwfJ/ATeQOHLwjbQ4Ln0Fui0Q4rf/c4RRPtbu
PbhP+tHp3+l1lubYiACywfo9JHUK63nOA2a4pOEy8APm0LSGWtqPTDBwIlbdTGCrjWd+euWDOMFr
W0iChS0RzV2kdLAABFVAGGTWdXyryqekir14hAHgbj5ZJuIkWVusVrOYLBHJ0srR/wvMGWaRpodh
CUvRs40CWGEe9H/FNNoQg0oAC8JXcxZMtJkfWVY1iw2g1sU5Lk8CageOAN0vycEPfJRHGYYxAU1w
nr/yQjpkfcrUlFSfeXCGEqq2XBbbg6AyjDWFuSIN48waBQ4HPvKLLIdWvYX3Dy+Ermrs0XXiETId
GKWyaPlBJc+3KL+UDDBNZ45P4IurUeU/ER4eszgqhlDcDAdlfjCKYxDYgijLkWLmbUztp0/OxDjV
uMNsnFUCkHHNQXowvtBig+MTekudJsZHSIgUJ0gyM16HIQsrtisSDsSpoemjUpBOK3WBC3IU/kw9
Fk+esZkcd3Sj0JPvTyP4fBkCfHJ4csIjPrPqaagUpSarE1Hai3cG6BWhyovZsCQP81zDC0FWg6pc
tsEIfQN7DglRqEmZ0sGK6zUx34cSNToqHZfWcFBeMccKyBgnsoERPNdeXuff4QzONRfLuEk+E7k6
+sbRtShhh8GhqHDAZp5Pd6e54Jp1cKZw3v8RT3catG+1LHW/KuJhN/dlJIV1dPirEC5vMLDxF4ua
ZzszK0JLs79xoT8nMAVsLNu8yhDdq6ymrAv1lueLAi/VdtCkYP8Q0T+PL717cJuj4g2KjyiXK7r8
mbrykpkaE060IU6bklaktFf0hS9aFGB05fb8Z8p14t10d233il2BvWd38HQ2uaMyOCuBreayE8aH
RpubcRjeVBvaxBjKqWTJjUjvDgbhQvZxasbhpZCniMGWIFIR06LDflIfjSVEFTgvLSVr+1OJ5TtL
Ltk0eSQoT9uyZZMrwAUgKuhqaxitZWL6C6JY/0vj7ACg2jW9aXJLGqekxDNm2ZoKos9cAQPvKTc9
Cg6SuYwF5Ygt4yeJrhPzAtiebMiPtZ+0n6mxk5PKEKVeRB8RQ+Fb//nKnKTKMsXW68yWn0h8NHh2
aR0+VKp1uExcWJelpSekBZGah4sGzvuAQD4R0skVtrzaRD40YieMUZH/76/QTvRfbBfdcxQQRNM7
XkuOcOjG9boWunGqfjBNqNqHbMdFRNFtPkHHlzApCi6aPMDa8o5C2gOrD3Y54mg6uXXvz0q7Ogsg
7JWZFLRTeSmsB+5PBSmEiZ9sG9sesLsqllvRZ/jIiFFtiO259jWQjZ/2GL1Ud7oubk6E8kh+3p2R
dVTD/9tz9LnJw1mWOH3ixEBU2y8HZafVOaRd5mgSRKSGLfP7ESTot0S8rKgz/v5fQY5T6fFLnAQT
Tqf6PpxLoc/Rd6coUHQWSWcMuT5tAbABxxzWYAxmQTMEdcvFPyF24iGE1vzECYb1Oh//1Ia2n9Y0
//36MC+U0gmGLWAzGsizABibTx+1BkWxhnJl7yQpYveTSq9ziaMdAS65fwbyb5QBJ0zrGLwWakr2
RTfesZaqTmk/G5ycRvbh7ebrg4y+ByPwVVUC2FW9qWtlw9ebS+y82MRfSXM0AXuOLbecbMe+MUTk
g1gHxqlp41TiQKyYq+LZAzKhnqKLBrCZwNvg55pZD8OSHHXcmjO9txa5vVPUyJb/a72KbM8PZDxB
Tgd/DGrTxx26plzcf8WIgmweIGQeoH7G+Rxk74K4gyCe2WDCpbbnmdxG2zkHVq8qouoWIeef40/a
CVjJ5pnrv7unM63SxZCYCtquL+PcABgQEQDhnZ/bhgWaXIH04+Rn4Tse6LkAfEsg1mIe4s2aatia
MURYhjHjxJn/+hkg1vF1fcuPTR6HOzLwKqiLjMgydN9/tsqqTAhI7vKlupAZsR2OdMx8xMzSsDJu
+eGK+1iUJ247MT0+hEyzy2DgcsbYAmd1UO3gq6TfBpitLBbzfCRQ6Ll5PA4R9/ZltpLHlnfKvtHf
6Yi4q16Ldk/FejLCv15Biw097e800UsNpC2y7oYA5f1/jSiglslccqdqq6kNZqBWTzZ6SYIcAGyn
Oqd0RdPHGOkHXbpYZY9EjcZwTnMPmT+SuJeQPM4PolJ9r1K4dtfMm69ydjgcEE3veA5lu7dq7qSx
RjjgLXecODE81+CKKeR3b7ubMdzrdKdw+/4f6o/v5p5jBCVQKg3dZ5sSvjAqjIzmyQ2U4T3uuYsH
tlFJWpzO5/SvPNu7Up+PALmHvfKU3jmE0Mer8kKfE3kYkBOky85XfYI+/1xxaiiIxWteCDd+CyrY
LSZPA0KxecOSMfGF3MihwijJqbJQr6Ny6iKwcmoiCiNPdqiWkxRIeTg63bwFF+kfikXnnBQOsLX1
O3TSFWeX5F6iuaEGKNIxEry0y2imM8ff4ttbDROFy0gB1J8A3g5A/LcR2upzZ3CFHoIqlUGcnFlo
iGZKwEPY1KizyiygWCWkF1995uMPBTdNW1O96oqtRszXAGV79bRsmkGJ0+4h3nhdzKpOHb6TxLRe
0cyJKSH8/trLvcIG96DjQsJChLNxnYw98/XSvNiX37OY/zUhlC0VPfIk3LGEV+ORhcPei/1x2wMY
kh/F5HXSi6eUX9VCTelCRKxehPNriDeLy3XfEurifCbdBbF6J6ucexvwPmzof87f22q3jg1e9ohQ
OK02ha5sW15Qyi7DGwoxzeaRyS8dyTNKfTnYXb2F9i0CQ/bUF/pJxyTVhP+Ru+zhT9pvqKSUP6Qy
2Nr2VsLiz7A+/McStX5pmNwnRf8PfJCi5S0LcMOK3NHs3zoJKL4zsWWCj+QUU7g9PhAUwN9maaBO
mtTzGzvKvCulhH9GRH5l2/lbH30YDCw5rkV1wcGKvYjZ5HgSyRRnsHz8bvOuTmwAHe7uqSCg3TQW
GCCJ0DE4ISWOQ2HkSqJ2A0XOSRs5lWkvw+Cn52OAJJrlqKWEIFntD5l3bOULGp7N+bX5UNY6Vpwx
M/+34Qgxs0k9UFVaEqyqAcXS2dM+c98Ttslnzks8qsGyWSEfUKd2NQbgLbr8fkoeinK8YUZgv8Ac
LRcSe1wBxsJUOOIdsXYoLfuT+MUNCk38ZM7hers7s5K1ZYjD0667E/XDpzcYT/PHYPVUUEm9cfP7
Bw0ES74A4FkMLOWOjF9CYflB9CBbDgGshSTAE9i+viob61tYgaEM4YDs+ZqemRMSD1/B9BoAEqa5
LOZPNRcygJ5xJVty/+AwrDkf2bO3Tr4mg1tiK1oo1si/V9/V99/s15QEX4xxnuO+tABgU7iXBLL0
KzSow55jdFFo8sExoGnb91phc58Etc/45qr79QdGbXPvKzqfki0kO05Pl/pHOfClGp54wRFX0rdP
VJGjT7/zbSsqJoplsnGWn50n8HGDqDYP8c3Bff1nXcApnKmqMn199dHA7mG71YHoFIeGpB+mKWBX
4Zli8DnRH+a1Wy5wEZFApENLCUiE7w7dao5da57inswIVpyppUkaxcm+MqWFHykXLhO9ifOndoZg
LIraZwF7bRnoF1BtcKqarsQUzwBT6teV+pM5aDQxjkR9UxTQXVGlgV8dob7X1ZMGgn/qt0ke7sQ6
DKw5xLlMIo78N4sAtOgIxAfOnDhmG7P77H/Z1CEXLqGi65vZEEpjhrkqSRXnBTxTwc31yqRn73mA
Gpf50u4cqb7Y3QDB6pf3BFXJTRE/gfLaQACn0v8pRE4f28iafc3UP7V8/SY7nCduFrR4D0YWBDAk
4AoOIKB8nJMXxSAXeMhI1nziEkT48Uo6+7xdUgGGHuU7Z8xMmg/IhDgxW6S3kv2x1PIlvNwf4TI9
tAoObQVJCOjl3S+KwcrFZ+jRXl340fi+ZZsa++1kDtJqRLP/Z0P3OucoP+R+f9dgD38KdKk55xXR
SGenirymEQ4uzPqQ9f9b6SR/Dcv13Viwpfgo9K+DstKmBT/2XIoXgtYXoJnAP2ijtOQlHdE42s14
JdEN5lPqrn7Xhnk/lAzaZQmxYe2CXuzcVgJIBZUJQcX9Q30A1BFrrPaFd5LlTrjdLvBwwvbdDfTG
AbjYNJuw7gp3R2AdNlK+Vs7rRvotmqE/Qtl1sRugSNTHfVAFHaq8kVmCJKydNaECPPS5sJYpz9W5
dxy4/mGibtGNMvrcbHQJPWPNK9rVIzjKPgKTFFR8t4bECR9Hvo0EQNL7XgJg5bkGNqTQnhzQoOYm
YycFgcimT/8lfdqaSMlNFRTm0+G8WPXU5G4n//evGsjXvzgTo2NGgrJ3aHR+OkcosFrML7C4/SQT
vI5M2OFg3cwrAW/C27GADgtW0SYoSEiq2nKgq7fDtbypF5MHN0jelM8BF/VgBnVkV+hvJoKkDtTe
TtRLgWphaU3xAxr2puqbDqC/CBAQ0lwAupZmMomGzkOZyN2rrDJ17+gQ5ibpjYRPwi6bPCYNNdCg
jVsS6a5tdRrw4Wj+HOPQeXdLni+HgDXL9D+2gMGQw6CPlcDu+VGToJgnNTJKrE8zuolnKAuRhADH
rHfxLxTTdkNSID/GZjzvw2N3di+4mbbL32QK2tuUU+MnN2r4ZnV7sYZ4uHa9oBsryDBPBBP5v2HC
INmfr++1LvoB0q163HeKYfmjUByu2ujxr6TzSp/uIBywJfeequgRJUuc8i41JxVtI7BizI9YShZW
r48qv07MK191NG2UJzfcMR3yjtVD7n+9XzVg8vIT2+3RSpCO8hz7uOMMd+QOidlweeE+vVvEpf/m
gSYZGz9uqZ3Z9SdlDMOGnT9hFxbqtLDOOqwkOvXPhmui0ez/Lq1KsWojDtFhS+PTtZGSuVr9eVpx
uv+s63H5B90S6W0HuBxTNU7+HXJ7wkRy+3rvP7icBRAJd1U4lcHsyEHqxjcQOprwge4bZzzLpnps
2JbpLV4l/0ODquuRlVu+/2cjyMm8s085ISM7Htqfax+7AzUYvhehyID56TOz5d1P93SaQNk+yOSU
dpI+k5HXhqR9OzblW3TLG9jD4OdJKXEtJB3LScn56+M6DauAj1e0zDPyD9zXLM0odZEDzQNNbw6y
VACiU/IYM53kp7UbGNlgRUCbsyedB7pPjzGUj2tYYu+Lq8rkWefO4VoN5XHObTEm+NyYSAwN8Swf
YTVFn7rm15IkGJx8QgKhH5dnScNh7hWwg3eVaJ3/lqn4vTpahek+xh8XQIFS0fJousz3VCjANAjf
PsSXSFt8uS5fWirogFCCsG2lIqlPRPpHbtecd5h35Y+ldb+M/Nh8QJA0k+uogKj7Tsi/HiU0bj7o
DtR9OE2SK9mlggoIYgV+GrK1utB4kuL5BKS7Js6NjLuWSd+LqytXvVGRVfExaUtg2yoLufjzH0UI
brbIFhi2a2cQTq1hg4iiC5cboHkvNh0w6cM+YkR8hGfvdPjJmHeyUmaXWAoG4JY4/IdKFNPaiRDm
YPs9iKTM7ltOltd04lFZFv3QC7jg8mVqTEY2o1/ahH67a/8W0EcgFeWQm/E/v/BeCsuTbPh0BbTd
u7nZ82cJJ0vwycEFNjFUYZaUNF9ToVd8tJ9x98QXXROcIlNU9jJqLq1S5xZUPyN/I92PmTm2NE9+
oQIY98JaTsL4zC26T8CdXk1abTgISJ/YM7j6IY4zWNEV78AnMCiR51Nv2pqLmM5dhYg0428drrnv
H0o52LX6cIyTi9SN2Szf9rke1b/ZQXI/HQuIixtuoJQQvTCHZaKkfKRRoKiyLFb+Mampsew+t5CX
u4Y8r5TXRrmr3Gw70+o7em/ZlTuqlMFbAgRYV/8TUH49diWIrJ6m1iK56juBm3P7qczIzmBIaiUQ
GSdbEbekWq7YZSAclg6s9xQn1Cp7MEP9dvzjmtFaXoRtbhX4IkirKlZ0nMqhUBLHotRpYTyUg9ka
Ib7BRHm4ltGofLsnVRPSMgVkQ4NmikiI+6/uCnnvXtJkc1PE5YcRbGeEtS3vfILddTlIZv9kPf2V
IKN1YopoSnX391vKjcdg1sF8ZfgPJNmsLiqcFxC0Ir6Aqe2qiywBtPEPDWCJh6Rh2ceyE5R6CsG+
CU/GoidGAtuU1xY3y70d98UvXqGfnVNnXchhLXuTrIg6lUM7s32uDNRGppmriAhAOHa8Nes3fPkr
+OcnUFWIlndPJoeyguW9ZEfh7hgw3Lj5v699ptSaNJt0W+RcQ/od7LAtCOmfyHpRlKTbQcexto3l
cpgNIR70sfhyDi/qgOt8UJZ5FV7c6kDNxml2pfbtk/Fx+swG3PjemUi4mGrbeiYWeuA+pAMwK9AJ
eiZDsorXogjvzWUxE2KfOCERukS8XLlzCFIadxIvZTGeP7rwSj9n6Fh8DiWaKBA9VKnx3HYCvHxD
/kZOgcIcMrRcFIDg+QxU/g4ReRMaUg6FEsXc3l6E720qklyOk4nULuoU0ThUvlZ7KD/A/2Zgua3K
7/gjheasizy6WZ+/5IWuBYalW91XrsBkk/wZnRQJefSEjwTfCNqs19p/AZjjAZWm4OFJdt3EEmsH
BGS1pnOTgLn/6i9rh9TC+w9g1FUq0IZVCBfDBLRHtr9k9jlWjidJyLG/PTnFC7bwUW19LxLY1+S0
JrtBfCJUvwKam4rv5L0EquDYS+HrBDVrXpeAtvmNINRacq9OdEB1UcoQXDfabyAMXbWLRz/1gpoe
YNpq7yMHA2gNU3r3rqQrGDnMkSMnzUTx07k89/e/ktEIsg428NGGRFwxfRavNHt6HYKUd0M6UV+s
nfZ/bdeYe8AVG22T/ePJ8+I8F1fj2oWZREcBke3hkJYQ+tejz6Knnf7o9DwdBsUeRRXyq1YTBh0m
2nr2TA7kQqtCDkb5iU5vRJVYJU9TKGQ4hs1AWtSJO0uQTRsg5Oadkzs7lJlKTLHu6QQ6H/QeHgWn
uEhPwara0v4udYS/QEzIt4Vvj6DfL3uxH6zzsEu1V1aI6yoLPq/g+6OWR1dx0KV04lQ8Ii9oK334
izwVxOWHfaLxQR6uDhn9e0nt4QrLLG5v1gQiKa3ohkjEVH78yhSg/iCkYwfJdUXT/qDQGsdVYA3h
2499VsU/ZFI87GaxNgg1JT5L5qXrQ5/O2KGMW4bEpE61lrD8CYvkMHE2uIZsvLdCItXL2JfQmeke
ynYjBGFvCuT8svyvLCTfRoF/F3FGZ1EWsvWtDtlWTxsRvLqeeAdGKFmfBPv0T+mHfAbLLUkaax6Q
+MKQ3xNgmqIJwinaoTJ0ur2mbQgc8mZ8TFYOwX22vlnDOpEA6pCbC6xX/iYGjFzBX2pRxKkKLjYy
qhQKj7br2GnIk5PSBkzkkB7bUfPLWFTM3aPNvZl/5yZt0AFgIGcNJeQzNkMIGFLJwKBslTHicEf8
v81y+cPZU8TYwxbRqPXE8kxnwdBcuAwIbWaZDXBA/OGc0W+Y30FX0B2Mv0x3J4b/PEzfvcNaXaT8
E+pP4YiG81Bu1AHInzOWqwOZxPBe1jKGNKVhvTKida95LquQP84JM5rVuSBOltcE6oMazCTYVH/S
K0C/hiZiojQgtC6jcthaWSNP0C2yTWVswffC+gtSxLaLy34Qh/NAeWPjFVpo6hNLqHo9Zi/UB/DC
9fxP4vGx/PwetjrR4wegbk9EBK8LCrBKuWYlPzUaUph7Dw03FGT1awtMLURwDFX1FSEqVEB832HF
cS0RgyuViIgtUVR1asZfjd1oQOt+KX9BTSRqqynOGoe29YiyBaZudxw8vbhQGRGOIiRk2DztafJc
dmA/p2Ey+3BzsZc/9dfTzKwE4CFKIvoYCceAJHP22R7kE8G5VJ/VgWEQPRmXomlMmOKU4aGgTbE9
OdgS6LPN3wQ7DqoRaOudg6PnVM/TPKGOQvfRHW+ze3L87OxyVTZfVD/5KCA+xWVlNDPwdDrwi9/u
mm05IX2loTKgmPKp7aIcNrB0QuCzobsAbVK5zRN87vhxK+O/zeCN71nqOnCDNp+ZDHn69MK7KyfB
Xoz+BNHvw8FC5QNYDjBOmUNzbBOWXwvLjrKKUEgyTSQjuNjRmaOPC/V/x+wOID6dG5OJyynh7KC+
j8R9B8pSyAisbQGV+P+ncrcCydIC75f8VZQd0BTJx8Dekp11vFqizFQXLrxEdg5Y/y9pNP284D8K
MOE1QWBXYryKkdjOK4e4BVCJNyeoYBNdiP8Q9fus7b/BbkY+WaxD87lkxGmHF6mzRxWu+3nYBx3y
3ZKf3ydBaVjc86IL293gQURKhJDBqDftyWF+Q1Kw2rDMUSiFP+lkW9uAZnNXHXBFXYPFgK1ZFle6
Aq8+jUDqni15qr0Ggr/tlVqwmj4Ya4Fxfr274IHA0fMBx9GI2vZ+mo1+Q3R9DNSBzhxDQrgyrTDg
p/F0wNRs6nAWPIxE+ZUuBLxVtWbOuGc8JtLK72LB98vF8i1vnzK7DrGjSeUP/pnxnM/wIq76/owV
C4uWzRQzgJSCmKObSFsu4DEau/6uQqrkBt78tAB5qpSst/vQjc7MRPhYi9UYSM5mCnJXsnB0f8UN
0JFKVy4AH7JRVQ3thYwRPV8dW1JfjcDAYNCCvXoBPWiT092EchkLMORZ0GpSZ4vuFnvTpdnDR4XD
f0Cx1YgnwIXnGFPIjdptsYznuCf0ewAJto3V4hFb6zP2YMyzciCnf4o6/eemKiMRvO7ioKTBow5w
pnrEzuKcfBQ6DBi/Zath3d2UZ3BYwZXe/sDZ9BneR+sojNaxwijgtFMBqfNfvz30u5TZ90gAr1Iq
IuJQ4zWGZpdia5f3C39Kh62jxR+XHQAPICMT8WbaOp2lHLlx2KBLJym1ENSZhcTsRAeztD+7WxCI
YSlnNeLBo82IhBtmBzHxE7Kik5+ul/V2GS2XzazOdQZXg5LtnIl5GTnpf/QV+tYEU1yRi2QW9qMy
M9xkkaOSTjdxs9Ko7UZ344tr/FIdJr573lC6dD+mYFzA2rfX+8vGadaXK1KRMr8QbymB156Z/eoQ
pO3LxgXkzxH4EVdT09Ri8guwJrt5ZtypxCrrtljCRob/OG8Mkiw6wkD048iNm9riB/DSNVDxcW9P
JddA/K1kDSUu+mvINcX4gHVnpNq0xnRXrH/dVt0a5pM04tX6pLPHqX+cqkLWKjKMImA82j5huFUG
bqDH8wxhSMAyi06wSLapx3tVq6elBT6FTrgFAZfUQ0VdKSRd4OSJmFDKEoCD0dEzGftiQlXq1DWy
Hvh4lO1KcauQUHRaINmkiqgstMqCzltdjr0xRqB3RHJMp8IbhQYXnn/qPDoto1WuFCWIHsxMXixm
xnKcE0WeMftxk51QDJJrceU2bThXev1McrRfm3kMTj/MRGCVUMmEa5xElVVFAaiHzVVy/6VV0Ery
R47ao0Eba1MCRbu6hAHhJPmZjoTeRSA+NnI+PGM4odNnGJaOsBIbrK4NahZEoLEWzlzlfzNKTUbI
dvaeUt4tK6UUVGFVKTTnUbglOQx8okdTvqrJTaEgoBY3kdLjqeyYLF7MIwkSyV5X37DHM26jyna6
OsU3v29+Rx5DO+okfYE8ZevjASzveOtHSIs/xng7qQqwYiHS0M9AKM4WZWnKg2lidiVFzUN6WexK
EeMOC98M1uNMOWw19c4ty8a4yhKBr2wAMTSdEszy0EBqze835Ddb5qehjpHxLifCkgPsOx6V2g3i
S6hU/YRm8vBJj/ZKbdeO/12ZTUbW/rgqKSywZHiyrB62f9CEdFPyWZNqKE2bytzI81G0rb7kz/2j
FXI//QM9MZLCtqtfwJ4/2rVZYtmC8Z9TQMXJkSas9AjaV8814hX5cFoQOQ8F+I72BZU8/oD5dyMs
wAx7jyK8Vj+88ZEJ2yZcpC+yC16HHkEvE3fILJIto+t2VRu0C4kzBlGXifBrsWilwfaj9Op5849A
Fa9eRg55nWSsCNUuaBcLxCNWx4HKl83LnSODRdJsdRPuc39ASYMBUcG2tPfA/Iz8yuufPFmlB+a1
tWfF8T1kzH5HfcpCCrEA314sFChOr3oJl9Mw85FQlRn50SHnepLI3u1MviTl1qT3kMujxlamE7Sm
+91xteG6i3v0x6Pb1mQDzWwgoJvubC4z23kyXDNmUqddK4U+xAUSb3BqjwkTLzuMFBML3lP/wyTl
7UkBb2Z73LHFdUKnwVPe5jwvWInFbnTGxKMr7cAKQBQ1LobUZj500kfElTcu63kWeQJujaMulx3v
MPo/E55lO5xzlX6tV/S3VFe5ejJnn/Pe8VvJsu0pMvz7hAewY/i8xt4fxffgDDqt+7x28k8OapN/
h5cw2eTTtZ4RCcXJtI15bn4uP8p4QWw7voMn1uAJOs+kWDizBEa7kfGm1WV1cfTorYlSDV8nGiqp
IEi1Orsh/dQLzraqR7HPIgsTBLpel42NtJ79taKX29AR8NX3eYJDa2WCI9D/oHWqIQq1PcgbU0F8
K9enNiP2wBOaM7N+2ZRmobAa0XGH5xazwKpHc8IU4cV/DgW4FskRniTQamhPNI97+ZVmhRon9xSs
UDdaN0S4mlpnGCcXOKTghSHbzxgvL99m6DwOlQF0j8VeiWQTJwzBLlJVg77PnSZGCI4QdNLkfMtA
6yvTHz8QEJZBfxw5/ur08Fkpzr3vcoehiWtqcaVSp650kvHN7mwqKZwagad6w7hgRJ5gfl2c3a23
qfv7tmS75uyGzMrOvms2QJPZ4rZCMD5v50yo5ZJTvHEt8lSl+6jrFxWriJtIl4mscMJOTcBeVSu7
IvQzFSkRCPXn7X2nGj2ZHO+wpaIFaGH3TsQ+T35Vc6Q0TmTVDRNJl0LFokdWSc2rc9COgrFDkBN/
kIz3A+83B2Id6HattAd1Bvvni6hMWgPJwe/JM6SF2+OWzGAbeZCOuExRiLD7Qwmx1RwKH0Eln9Ur
H963QyHf+WY4/nUCOFLrP2xS5XJSNBOBlqQ/1kcF5b2lqqfzP/DKYVTN6vp0MN19cQxsCGB/9euu
TpWBtUl3dqs7hhL6aXR0+lZc1bg/nLDoq3RN8R3WHJmPZ52zgtvV8XfefP+94lIWZ2UBD8c97g25
3aPhVsdLNG7z2EvcBTiRlodCKsQUPWezNerLfEDTagt8RiBRCt+X0eKmqcy/G6/8kp/bBKh0BAQ/
/XTLaEzaNKl3Wtf9TJcEFKh23AIpduWnRQsIAO3vmPIENe4tT9TWmc4hc2la3CBKCf/Nm5RiUBbm
iW/tQzP0b494Bp5kY+QjycRI/kWpur6m0y+Noa8tVsrro2WMfWQb1DpCJj5OO4GWYHOFQ3nuaYnx
xsf9B/+xJegYj31J8UB0K2cOw4YuE1g/El8PYMJUq7adxyiLRy5c08uCjWhJ7JIZptjgSpkyXeNq
NSC65qg3jb/6rgrRMMH4N1nBDwaTkmweTKkbboRKdu02dgAhW0vb5Zoq60IBxYOoCh+YooTGS6cG
+hsPbGG8Wcd7cwdiFOVZxU5NWtEeROKPR8M7jL+DrAIUmnlO0kt1LMUk+erF/w/0TDVGDXywXtgh
wFLNlpuuc84xYQ1p3JORPrWil4ZixZTIw3X14Qos+BP1/VaoYSQdUM3f6O6SCb4gTJHm1TzuJWwE
rEKAqwvu/9ZyEEABGw7SHObdxaJLsXfy57ezNTULamzEMrxSZHdCRIKLP6Q5rypqJCfaDg3Kn0Sz
Hd423HuJ37MEO9f7svFZQ8Gaka7aoE1VPZyZUuSf2sq6aFmzNbLJVmid8LAgkOBl6PKSS/23bm34
WkIs2SJwDxm01gqf///0YFlWz0AfuWlYkQyG3xWF94eSlJfvG0PY5C/oW0RMALQkhxg7F9ebs85J
D4rQw8yWllTjvIo18YKF3r18vlUDIK1KKtyvvh4els6sVPynPDpbeygVfsxeNmMrp9zTRHbnjLbi
oGa55m2GBTBjYOb1zHIsCO99Ze0fhMsaENWi9cfW1RlUtZh2NeJkjR7NoSJIxIZ7CCt80ZR2ogLn
0pA6lKKc7Q3iDfs0dlJTxJw8ZWI2q2ZXR30QcKmZ8uVbR5nNmvkPRb4OkK3q86S2s1fQBUOEn7ej
JGXvfP+uNGA4PCFBRQishqHyZQ9w3jrYzulXTpMAeNMceuC9waTdtEE4o1qD7sNeprf8A13wqKYm
75SOXtzkiXlAiGRf8O5m9RavUayyEeg0/vSXFjw6EEct/SDKtS3IezdcGbTnuCcKZn5fXKIAk+LO
2bv260jpjjEupVPGEBYwF+sPEtUu+WAgNAaK0zTjrhzfNzIAtaEkcRAc6toc7e3JwFscvIMjpRFp
Vg8XxvOoz7N6XZfoRE6cW2GephFHGYwiV1z7Pif0kJ6T12AMNNtUOtQg75KdsySaKrqJuE8ApcqN
oO0/V3k5DKf4SgQsDbfoBlNmhnJu+/MYZVSEKssaqj4A+trPVnalnSyJlPeRB0Z2Aa/a9xpFbRZc
9l0p96IlBeqatBMh9PU+BMkchd9oLntJLgxVltP2YSVFAhWvmxOWQW4omrxcgwqVtW2Rc4qh+g40
o4LiYHfKBUE6f0cBXE55C09BstkVzM647Sd74hfxAjNXxpGROnoBiKqfxcUfFYmou/EONevVIFM/
OuwaDJPLkvIQkpl/t3OnFOSZ6T3mtXIG770+XfBFCHIYj1QLemUPs4MQOUDuGZBWkUkVup/xQY6z
HHBWo4nQj9CfhfWpo7x95gnvxElF4M30pmMGy4EPNoE9Q2opVqeKFzuZLrdeS9J8wtKcnLhvzGQO
7dkMCNtnYZDyTjR8OoXLBPL8TQdoM07QjqQTYfl4iQL+f6h9hvk93HGnnDdYnb2qJuyCbNIcOnUb
s1Gzf4L+cdfBktpzj9xTAY4n5IGuudT3p9h673jvLSaUwSTFtZGNw/oqCwaPcNCU/KSOo6RO/O8e
XS3u0V+7oMcns16YZ7ZAWn8ZHp9h2dZhGJIs0mfzGO32olpa0Dm6lFqXdlQOjST87em2L9Fd5g+d
1CZXwLSwOo9OjmG2kZFpvwcPpDUnnPsld8I8557m1VW/NaJ5sJGoodOvxARLe8Mhbf2e2vO+hi+i
12baZSF8Ewb6PU9PoRQvCy//5X3Gi91p+dARhm4MVWHluEB5JxK4Ht2SAI1c2w40t+qCbJogZ3ua
C4Ep/LyJ4VIZwMaMQ9sn0vGDUF7bdySO+jR3n1826q15I+5CR9fId31Pnied5qW7K08KLkJ7Eb4m
Ldrcq8bvxnJey6xLts8dw1M3xbCUQTkxNdZafhmxrRN33Ebe4oeaGHV/GFESIEaSXmAv0clLBJJm
IY4+2qPJLdZ2D8SHQZh4SDAImd4IMlI3RjGry/M6uJt/V4nLp8euyi2iTBt4iorhD+bPWwg7zPV8
LajzmLiNT3Lyo6ljiYN2/ljMVf0Rq32rKno/Math4luHvbXCgZpnnN3ZvYkjZc9C7c+zQed702H+
7tohLhrIwJGnh3zr0GdcNigwoJBw17upzAYKNviZcoNiIcHxUeNYvFsDeyl9OPKLQ+AhXsYFivVj
mpC7xV4nZeX8FRn7iX5mKcKG6nOSWytdbbzsKWcyecW0hXx3pzA36lWnfkK4Ar4u+ZmZoMumLlb7
ZysCOkRqybZdktqKGFRIAjz+nIbd49Rug0MQVYurN1Mtf1DrCjFDqsqGhXBCjkLUUpOkWTZRvMqe
+dPKX40NmISFa7JLak9Pf3lUW1HSWZF3vpyi2d/3vRzMhkQFUK7cjeuAQGQBFgJ8Q+ooF2cHSX5n
jWLAi9YrdgIYChs2omfEqVnRIqMVrYCwHCeAJ4bqL1WoXee/deTWH/HY8gsiJ2skvDrfSHhcKE0D
KW0z6eD28cOoSkl0EfITPcZdYdOs8IYNm7CQgRl0a9WcghVPWBT3WXUDsYQXkKJyfDP6Rp4RBu7Q
Qdd2dsyc5YdenO+Ipy6p/d3+2N/piB6s7OhYas7voLvuwbi8o3C4b1zDo95FtIdBjL2Y/9Gmkma+
J8gp1HG7pM+mpwxqyQrxDZ+dYOsbl3b+/RhFuUpTvTjHNGl6KLd+6UCwt9Kmjzo6hLIWMnaHJvKI
NfOlU9pntWP8NLdNdo8HS9LeEoWpXxI0QFZKQ1yW8xBRScfjag+4Z7MIUtB+A/mXwUGuKGsS2Kzt
EsMu3L7wvvl9mCKu66mi9XzMDgA6pG289qGCr1b03ccrl+p5JX9FB7xVD3NRDFs0GrYmPcFmNtd8
BNbqinJM/OkbYNubQPfXZ+C/QyiJRc5ok1YPXbdqumVFAXtPKeZbKVUwyyAio024PVFPIOzG93ud
l04D1pxqkLOCuNd42hdtOhcIqLtcRw29ZLE0NLRMoof9PALt3BFemmyLCrko1Z/plLDqITmgZSqZ
IBLDm5KlX7IwNDFnjTtGAAIJhvkiV0jTUxcrUR2glgGiHL0FqipIgY8ZXLoV+ENA5/L6ko1AXseA
HerNOjACk0WEK6VkKrQTCR604lx7jxfG+ey8FQrpmglLO9esEaSxPLY59SOXgfRrHXl//sbkJkM3
WoGE/1/YaQdXJL/sNxH/G8VCAZL76HZPZL8d1ybuYHEHKlm0VQFnkQ3Rx95fkU73gyH84aeKRnKY
j4iHq4sgqmyTLQH/mMK19QKSZ9XX8dzfndjk3sgYAWdFw5PcNChnF6REyGeyjSsCWdZEhmATqxDn
pVXJkoGD69t9t/EOrcpfzfh+7nzBSK6BvO0zbu8VNAAlvtXOxl4jI5fG2ywLUNjoJvvbbd6HgXu8
dPWfW4Gr15xRPrIeJ0xlrNrhcD+fViL9IKwn2ju9tg8L/Xe7oCHbsNGPQCJmKX2JBW/qY6bpTxub
IVjVTAHFg6kMBwytyOrLC/bzue1TwgACrlCPfpLXhpJJxLj+v6rsfDTYugLQVRVP7a1FA8cmkxaM
7yK1U5T9pZNxPOKXE+4HZWX9hIjKJVbaQYi576uCKIM9kUMV90JYTSm5M7RVtL9T/K9I15SbBadI
g1Zep+hyh1JSbeVWrRQfFSg6Hd0UZ9vwTJ7Y6UtmSpIGPaxy1TcMAAw2Rcrn7Pbi+hFcFm+OGYHR
jFTChXs81Ly7ZO8dHm4maPKLUFqBl9JLISf7Agr7ilLOUu4D9ckhOGvIrkgzsCW2UdYek6uQvRPU
OH6SRPoS3qkkuQQz675rulVdk2otKv52AyC3rfFy/FB1tI5uqNFnGK459Iyf+DIhzWn5DoRgMXti
fwEBLnGAg0smDgrNPpHJFUU4ExJNIQ4uvvFpRcvUHgZSpRhnQ5aMT5igg14KCtZ42rWXF4zQMJq1
mCiK2KZBRz1+sJdnfbITFNlNaNwINCykg2FVoMBQU9qshOjyHSUmD27Uv4gxSAc6WMniRB5gkxEu
A9JT/t/oCc1814a5pJS5Ynhremz6dO29gKiin9I0fyJ+vEt7fTq3LChUq3FAYgDlZmXE//6oPn7M
NfuWWqDmbUHkYjg257xRAK9GCgpy6/f6PcN4BC/u0zkkKz3OB3Db5hZnpQsS+4mqzQGPn9nTA7Rn
sFjbDoL5bgcGNG3+nwBUP09lHPAvl757tI166KbpLr8hJ2l852vSUZAALy8uTSfIWRIxHepfUrsf
asnSXJq/K0H4TjWPM1WMrGWhPQ+kU7PNCHr+YMnv7ejTcOxGlQr9m9dbkNI44sH7FGUkLwcch3jJ
eOdmSE2m30yf9L9iAFnK40oxBtxNZygg9sTfGa5fIcXUqb6DE3jQzh+FpLzhNgapFS6TRmdBElhk
k9x1LxXd0p796++8uNwiaeVEJxm9TweDVLhqXLuckajMcjErmGrU6DRuAkErxamDzQsp0ZfJAT15
eX/nfAF/865nVqftUYPUhcg1J7AFM/8rCiIhOHMZWRrI148ZCWissaPEtN3OwI9ezMCmVb1oFg6l
DE6+jk247ui7J04oi0kAX/JrDMowyJ3PAYuGFiZccFi1OZzMy2FSnhXAUKlvWtyUxuoOgiVSOi05
pI6aMYKIqwSI1hnyL1zLdz+6dlHyyU6Z0B5ZsG+bo0NJnMcJMhAVd8ApRjIXodqZaTRxwb5i3Iu+
h4uhSyD4U4coYeZ3TvWcgKbC/Ug0JumUIXfQi1NRro4E4/SX/xZwb5FyI4feZFDTWkbil7tt/1oW
RDRbob6WPClRsGh1Nqie4Ks+vgDZhyYdKcyBbb15m849sLSWs+BqK0nRSFWcwiCAe2YyBcS/NaYc
xJZxE0QdByOC4fTywz80jrOkdrqsHpKeeiu5iPJpsycbP0LaCv7GuOTv0+nug1iUj5JmeZW5KL8P
Lwr9p44d/Vj36u5NTWgYgEyDjC0LFEVag14QhhvapCIPapoi8VsmMlF90SVLIFDK3z+uJ5N635lY
yfUzPzvRqdFxokISvb97Wam53MvdKzM1LV1GA5hnQzAZo6/SmHTvlC/qsb9LCeyuAQ3lYwkYgt4F
xu4q58p/UGpcO3w7mfmZhshYoxowvrUxrBTOormDfgqHeB+sBMkQ2uYswDVOGVYVTppNXa3mAtQX
34blfsJy9f4XQRtQF78Qt+XUxwsqouMZBniPDLFQrgg5N7qE1feY9eOIP3SEqoa5XCeaAvVXiWpX
jkIKDT5jPij4J+/RFTFX0AAOq3cVD1G5wW4UWKfddvQRR96Q6BT1FLF4JjaS+2oZbofqMFAoTQXq
fCY+IoczpV2m0NCcdyuMeA/nbpOF2DNUDlEIrEWozMOAnOJ8dKu+fDLOMQF5b+3AthF8t3zZtm+M
wvbuJRBbRscjbD/C+8vFfduhF6aDXoUdlJkXXBk6Q/x8zuREnxH538qZVJtO/a9CgqxajUiL83ad
6eU9r17VDY4y/rM9P0dVIBk0cMx2gVsglx23dhJKmqyaryPxIu2zWdLsYIKYNx49YZQrazInyTtt
onUxDLa98STv+Kkgv/4gzbHiiip7AtUR7ecNs539chA+CCPM4b2lD6arWJzTgbgs5RTDAlT4VEW+
P92nvNUGWVoXZ0Lfo3ao8uzOv9Q/uVknRVBrfju71JYZ+i2UZxGxaEDFL0FxuixqRDqzWLYjvXeH
iECetBMAcQE6ucUPSyreJ4xfcCozIaPIT4Hrc4rjneFz86aUayO+JeoESSIraZFtGO1OP18FnKAW
J4jdd2QAhIuUpyn3NDkg7C9TM3xD5vkVmhhKnxIfXmtscFRP5t1m14ywvyrovUWtlkgcG426CIrZ
HTJcZxbGcCAFqzE3nVXlBqvl7vdriHYHriZ6xbsjhHfE1yt+DALZJ+gMAB48autO4PFyXehkhHmP
DhACIqqXcXX3oJESKOvSVfSMXFh6/Dzbh8BHL+vvzoOnLCTmSCTBmwB+YgRTsOUGWmXzzjYxgOhF
Img1L3TZg3QKqZhDJItSpE3MLciDg0FNU+pIn3ygzMWEabvaTkqeQhZOl16/fJGdPWe7NboFVbGP
PoUXkHwJm8ajiSvbxpBiivtwYgJLus8PPcNWQWhkwIskaY3oB9cO6z2NF+Zg3ir4lGVZjLLz6NB4
/TUHtphua6M0m2DHzVJUlGkUyvZcuq4fZ1S3vpzP/VvN6+/ESAu/b2lrAOEsz1eYYFIurbjVgdGV
r7MxRa34K+TMwwkXCaQF200cC9O6yOiUiKnT6CMhydzrIEeeBoDk2HW1ZMfk9dltx6c3Chl4FKoT
eLuVlKnjb5tXkvARs/0v0q/1xyYXLmyS6XFU7Oh6swZROBYQob1X97HNYTZdwVOnWtr6liZN79+N
nbQointpMa43wKfVxmbNbCAVRky3LmmiXQ5FJu71w3z8nscGwzykRabCzXMTz7km8iajN4IB+Rwh
H26k3uGagsp1BPJxPoi5fZbGt+xQvCwow5y4oh5u01Rb3PRvL2+eQCWfpWvjU1Mj5r8FXm7wkBx8
bpVXEh+ZSreBa90e/tvYhQGi17CVHBkbzyKHLyxM3K0+7inflZHdEM3cPRsAyzpLTdF1Ygq12lv4
jU8hGCequy03kzvlIo8t7i4YCd8S9ZGfqeGb63gTpxeSIaEDstohTLI1bnBVt/SuPYGPcFT1Up8r
Gr2Psgko7i+CpO6bQKlCAx0WYNhC/u2Wc7TgDrCq7A4fOBoKO6EILx6Kp4u4+Xf+Zan+OV25SJeI
NZBqdzOsGQebwArfaD/I8QoImvrS9t32w6lURok4Z7FvZftb+0aApFAtvZ4UKAO4oH5dQSIpbh46
DVQTmLtEu842unyrnrhMmk4hUIZSBnsduzBhLlNOBhon35hcyT8NuYDYygLtQagR+Lmx9JPKH76C
8Vf0PGPKOzzXlKl3KRerpcCwgB8t+rw529tINuk5eCwvPOFXl2FNkSJQNaQ5EKa/2ifNC7rLrS4t
kZKgTNNxixFG8qFoQb8TjDvW4pZQt2d6XZgR5C/I5Jx3T8fJgteu/wM3iGzsvnrcpYiQdq4BcP1u
LUvwTlkXZp0/AvcCegQW5QTtW8y9qHzjBgIweEBb4nShkfu15CtE5mxtfVeMafJqhImO+3AxW8bY
8Exuw9JS6p1fX+FXU8xhecbCu5cCOUlk7yPN0BSBh1ezeAptinEc8BJEkpwvxKmPBN8XeRVvEA9H
sjWFAAuBH3bdn5jptZ9DFUBVa4OwR8KXGqJCicQE+tghjBuK4j3GaD4cANzBRyzUJRI0Cwfmmqm3
MYdZpU6wXnE7TVQ7a1yMAbPAXgWs4VTbyyJR/vSTup2rhLr07wA5RrRQFfCRJ1kBfAv2tE5/SH6/
r0GfEpHWkODYkdnd3otdMphD1u0vycKkhlUjKtstIqzlvfrJkNOUxiWV4DZJOs4X5qf//IU7d9J5
JlJvAr7UE9YK37hB6KrSWe6siCbn7V/NrsotVM20oSvtjKwaBpu1OLDMBnJqMG/26HHPeuHwXosY
bFhuwFO2+8QtAqpwyQDekSpHWflfAmxEQtEF5L81jelruupdGnBsNVbJFZyy2DEqazbeibJRMqh/
wSg0HvGipRft/suiLcSU14WJTVcXEH76d9D6PzuGYEVNmF7ZhEbVI8F8dkEfUzbtzz1vUN+kbVJV
rKyHAQnEgPEpuXVtaw8ySJluAi7aqxf+lLByWd6flFcfTaFGmXLVsA0nOtus+9V/YCzrLhVOnx55
iW73cLgFbuv3bG7ezjIFPxjzEBnXfwLNnSBTh6OVQQI9gE1zkQrAGmh0F72NfPWiiPpFvV3RiB8P
lGbjpBbf8d6qsxjo2FEv/+qnKIhRVd3aBf6Zrc7r/jhDRHmT/0bnI+cHXtOWfIBCZMtRvO34CW/T
LkIVbPWRv7loq0SzqajV9NYZmNAQ6QoJemso8OkG/kus9HxW7y4XlHGgHR8cgztf4yzbQGMFpqo5
kpB5zguENctt6lHJbUfP0hOcO8CkL/+cWzV2B5qtGaxSpVgv1/dw6uk86TGHbCt4jJSve88nemre
McOptiiiPWzZCbGI//lSCKI+4K6jSA5shd9A33meUBEf7jGevw41E4qbRqLSeIWMBo0v/A0pHD4o
6gMhIfopjgmlZjC+nInl+Y+GxalygowSNr6iUc72gsdCDbuWOhGH+cwkH0DUz9S4r5+QE6baGJ8p
0uh3gZb8OueTLLr897e0sKvR7ZOPyXBHqJgnu6V1SqRdemg6tt+XRZENwMNioCkENN6iCWFE7OQf
USxI6XHM1HDwUE5/eLyhW8tQpay1Dk+97RvE/HUCM0w91R4okyA0wcW1vWTpPL0qM5xpEwcsTbP3
32rp4OzVDxSEtTmBxm59JdF9X4s5DDndsG6sbJ8iUPTxdAu7JBotkGI0r2C4T8QClj3gzCSZJiP1
IEMTYUubpVMloweDsWTRTAkpKbdzASpGOlR9TvT6i7d/7vF7InGg3fvB2ey0ludimVwRSO27Vn44
y2YvRGpurV7UeGMKH8MqjcprKMBgu6DtHft7ZMcnW8dpsNXYcuw54rdFTvP/VKoc7kU79Tb5hBqM
CDqLhrjKh04eY8WN/OXNm5ygNvAK9gG/XX1tl3bXEayCIDb8QQyBhxDpaqUGWymfwOdTTCKmi4At
iAo5cgmoywW0wTQm66NvHFKonJO9bLIKtmLqVRnTEmmccHyHHu2Yr/q5PPKMij1yrsWPILFeF1/O
V5WJ5aChEgRz+uto6vLV9EDrdBaXGuWGdU3sevPlIYL/4yMDAS0hp45DrelZ1I+00VPEp+plpI+e
r0FLkKJeQuIvo2MVBIn1QkdZgHI+9qDeH1f1kwlLNS8IT9osQ6hgc2rhL1k6LjcxlriWp7xRqbht
LVRgWkN7RFt+AYb80kqe74zAZobPG9mWTNg9/DdhtDOMN8/5oq795h05VpNfr0x+UzGuhB4ynyvJ
4QprzsEIEGFGXFS3gT9cqvPVBVGmw5WFRhOZztNbufgrzzbP72JFUCSmWR+5+wezaJZDR8U795na
i6CAPk8NgPAU+WVB8cTKJ5VlCH/q+NX95ePKtOsBUYsMFCEGbBfH8ZYJuQ1bxFCNCI9+zbEdSz0E
z0SrpMH5E7+f2peXK0Wnuo3yrTyWinuLikyQDGVBpKwymNwktmQfctDSC2CiClEtk2Qqsx86DpTY
TmUhLzVvXQ6OuTCOovJbb56D2+wwFDZ34jnj1ZR4NfGDAYZPRHmpXjszgwC6/3b2wGtqjgA8a7dQ
/NLMgiDkhkmnoM1/WuhtpmqNfXOD5TzMNVjLljY+ZGI+D6UTDukxzMFDT87ZVyNNoMYEzwTSwcZy
/ecy+m14QS1mA7y+CvaxFQ5ch/ycgYLEqLWdZnmaUKs/i9dXv562Z4spfh8MdzYmLobXBYhq3Y5X
OJYS08sumHP4PX//KsEwiT2UIh3jVcLqzkUHi5IGIPQHnwThra+L/D4pAOQUaRVmivHjEDf0IImz
xXDTUEe0/vgquUyfc4usqIT+GLx5/iEjtQZ8rVGQdIzO3NNo8A887OouKRrhezjcCbGTYgaSHSbY
sPR+TOcPgoYaDVyANPl69YF2RDZZ+xKsfqntyUaPeyqEjDk1knvyIj74Q02PXWaGV6roIpKdfto7
x54zI8tAy+I1md7DNnN+zpVk14rtB2C/T1ZBZpxHJEhPGclOWA53qsdgzG/9y8/RHFgoRbzFAySr
9TytcDQq6mLPx5C1BpcfRBFxiz/g8IY/HzBNDZ0BNnIRbvg8GBrcPYNFhZsk4pnNv5pstIZnHE50
F9DOiR2oHo0PFL448UVHplL3YhCh2RhgClLvRWglBM6WrNREcoD/v5T1GvTr6pltFAQebVH1UiTT
lpIdh3p5z85lPrsmoVv7KRp48lkVsAMe/F+3n8If7B25tmZ5T1WgIBBLTJglG/En1AsJtwo28BUa
tPDEo2baZBQA9WzUGDhzNQ2dMUD/A82F5JFQKW/F6CePJeNJQcseyraDQRvZM+aCbytWlwACNeqk
v82pXHslDKGjIKtyf41q2V9RNqkQB163xeElXvcIKA6RLknLJFBMIlWe5t0SNcFgthOiF7ndl0/o
+a9gwd3hyFkKNNr18jvyyHm3CEFbSd6SxQoDUf3+cm9Sc0UW4gcy4cu+sXTWxFtA/91cntnNMip5
fgWykrlO4brlmuLUbiHLUTMWly5MDVdX94atBfYuIGBEcszVLMJbCASWpOCjRt1slzl9r5EPP+JW
RQAOKyrC0GkebMCE+McQOD5HX78+kHJw7SJknJHnOioJ1IB6FeYefK+O77jzqM8+7SfvqOJcnSW6
tAreReFq+LbOFzx/THXmzgE5zIT9bEZbK259NbODVQ1d1f3uIELV7mzUZzTa31ffoKWzOB98mW1n
oEhsQAoXVOMEorIJUM9jk2oHn3LGpxYUkmBlGfhPVMhRla66fF1kYpEMEYPWnj1kukwoaNwHGxB8
VmKCn7DBEjTfS2dOz9VcWEnmccBjFqwIJO8VbD9Xp2DwLUyUWtwBARjrIYq4fxUuAapPwfwslrrU
U9ywgI6iGPPXqIXwh1wjUK8gu3JLzI+19h1eU/40vwqKTVXtbqUm+wSNffB9rbHSReoqNsuuDgE9
VPGrRP2SIK0dg7rtjpwqwzq1AXrLXvx0VtYxFkvTEZXvYgpFi0REk/MfF2LxMPRoWV7GFXarGZWZ
VDxJOqBsidqTrwY/j3XEBY11yuhdvgXXP5U/zENfthu4PyyWquJFryPvlEh+Oi+1mrXmJEKDshy4
WM4H4wWViIxuSjoYbAJEasOBeZvojdjYshErm4VlpDn0nKMIA6KvJUcN2uWTIto5HKvHTMaEjsY7
v5QzStpeZhoEbHGQ28xt2Jo7NxjCFoN3MuF7YLQXShCoOGn7X3QoBo2PSiMNKhHbTmG2CXyw6kl/
p+NOLRZ3FulRQpEw3KV5tJ/QsBKtbIwJKCId9wTt2pkSbf4MnPfxTstq8NjdA48oxNfdDjJkWTBC
GW7bLRclh8U8ELLEelqD6dgGa5sZAgaVfSgoJJbc7nPHthiNGFTA/cjOrElOSn/KECCdyXyZhaCx
3WMVc8QlgGIt6dxCj8sJmz+rP9Upp8IeNAYlT1vdh7oeEpPlh5ZzjEEFZUlue+j84hXuDkT5r5b9
AUGATCQ3nJD3vfiFc6v6dP+vaVpf1EKvHQfyx269LbOdzI+3jYmxMDeF+6bcIr2GdAvPr3Y/uucr
vHF/pC7VQyZQS14qVn3FSV1vzlh0S3lbcjMq8tgnJgAqK7E166NJ1a6MzP+D5WNYOnXDXT+S1iwT
lQJxy2ReyWvpgDxdNWN9EqjoH5tol0Ag63ncACXZUKDIlPZYrLH8azVaRYu5rkLNJLqQYw+oVinv
YyWs9O8xGU5hpHWTTQMbnDlEd3BE9RirkA0kgdIpqzJX8+tcNL/h4kNr54QF1uQmS+SGor2e4GrI
y/qaXC1zdc/gShYVN5xZo+SSJ9Y+8+I4jeQ4HcSEqZx2MR4dy3jFhZtHrzq91/CwKYHZIpqUZ47H
ityVKALm0+CUTrvGjwaYGhZ6nh8VlxVccqs1XTEc4WhTVrLwGgfcGWo6rQnmjluFWzOXpKyoDdsj
bxr+/Ck2Tobb5ZuH1/XioRU2567nCjyZ0eu0N857edJb6ZhOeAtkPGMCoqmK9TzPfGtjUz8DrQRS
QLNW/mo/ulc/xA3ajh8a9KaLCnT+Fmxxst6jLzYj/7ZqI4d69EMAs6GV945YRfv/8HjrfxV12uwH
vI4lc8IoxqfF9h3NW+G11WK/K4064o5pBs7EGrt8U47+AykkpGjHda5HLhlk8UJo94cTR2CzgAzD
hzKhIYlnGOV3PFcsRCzJxjfAmeOB+J2Qw2jnpN5ObhZLFTlNvw4Vm+5im3ZtnZ+0sDsw30iWzqjO
NFOAfH2mvDDAAwnbT2+RB/++s5G+FQ+CnXeacOYAzcB1AO7WH4Mv/2bchHTaVngv3D4Y3j6vjSgy
XGlKH6HYiybwI1MZlrzXK74cuQVLJcpBIHPDzdfEeSL9cZ7TnEEpEsZCu9lT9Fj0Z3fjz1pzpbfF
1du8+piLMSMUijt9lsaAstyrpDufdQ6v+wU5VoQyoDclBljJjamer3vcJf5F+GHcWWBw7UemjY+Z
ZdsCEYRgsXwQTRR+KCPmFmY73iWUm65/pz0/eIzXZ7bx3VUu0Z/ZojK2Jk1N9xTRytETkRutflsq
kYF0XW/8tcjrza6M8yPqw+eVVg/FhGHpbGIG9eJZhNeDGFgfOf9aGN+UXsNYt4JsEyJxCRnttTxL
UFS1zWB/A2a8etx05hJoECVqZKQhhLYNwthJ4xv/M/O19+qP4VNz6QSoHH4Q1c77j2fhUIzTE1HU
dt5x0/GGH9oA9aA1ipB2/EQpS9i8HDUADW7KW91TlyqPxO3T3/M90csWL2BljcNG2haP1udjpzMP
53bRuELBPqxFIM35Q4sv6j+aoe82e8epw9cpop9V5+lCEVXtXCUka9ncbio72tOLdsBNoVv/64YR
/nVyhGZVrwlrmXQv7s4Sk9YE6KOswe4+KNAMs4tZb5TD+ylqokDgjVGr7uoveR0VwGKvf06EH+kd
ypxdWZ00O/a8abN1P+BfK3R8smr3C4RKYZBFlKE/xgyQGapc3vuw1sCMxVd6Z/ZZH4YR6BvOgLXB
b32kRV666S4PpMqLVq17RTNpJzRuo/yYMxqnd5QdyuLHDU1I4KZ1TlMD1bNTCVH0PTCK/u9nuYFz
2UAF80+6gauZ+cVLLfDAdG+Ei33j+JYb57rga/q0HcGwNwu8G7S+MIk6as3P8cU+kK8dNtduoszs
g1vXzWEyj5t05AscX/OI5gTNo8Kv6V7B+bk8pbZKfJEiLTe0ChHUOBN7bGOC/cE8o1lxez+9ba29
PlYdPKWEUSLzl7MHWQYdi6CxwWiTV0OXY2sHd6OWCGCp6tmWqw1vZDAkezam6IZxDuc8fnPL7tJu
/vxelIOcjrb3hatHWx6I+UOMSujk2BHeaiv8TMaWVh7BJGcPaOQsYE5wA+NoSYR7pDBwx+5lux8G
uWwYcTnQH0REukowpRKZ4KLb79Buqn4dkNHRKGkUlJDXb+yPR26yaY5Zjmct09iib1tWQ5VGda7E
L4evWDudX2O7qrhEncMTNn9vKVHXeNu4UoSSO56PYQ0BOYczdh8gNbnxWGBfWqjpmwvxS/Amrotm
+7w/95eSe4vaJzaCpbCv/tEL0BqaXO5PsKPs9CB+VEmKoYZ7KhsJ5LnF+VYCxLthMuWI9BRhSIyT
pgWLQedHLC68W/ImzgIvo2Xm64j0m4wBbQvn++6RJ3i1GO+dXTmWVDkyeIrlyuIHLdDToxPVUIy6
xko2A+fQ7xbhACpqaylKKkXTgvIllW54zWXkJ61HoecKxlejknNCRfkQV5Xff2Ternf15nRLjwC2
1FUUplKBpdr8BSniiavDdU9qGBICmZNbqO1Nn/bUJjhtYzenKvllpqytXeIZydF4t/alVMJfVsEM
XS8NASLpxOKOHHXy6mCXxTbgqXIU7Vp93r9ILY8WoT7kKlXJHHGVjHTGi2jXQ9VnEgBxeLb4/tLz
/8fSeBorCTYJr0e1xdDnnzPOmomuwsBQMWdntwl4yomb7jmL+CzlF4B4b4W01+0BbID6duqF3WXA
/urf0NHoFOszd4LmcposglI0ul6RLA4ARicKi1PO0qf+PqsYZBUO95zOtFw0VjNiiqAFb5Nz74mk
gpp6UJZ92I1XD1KR2Alw6A6SKgyuq/tdfD0Wjy7E8FBlzFjV+xJN3/WEdUjkNXAyWLTm2wYnrNmA
ANegLgw2f0gtgoOtcMAnw24KOFJl4pFz8S3iSvR7oZUAIzBK48WpOZTCweOJ5eNCYSSmikIz56LN
vUxvepdbFbAZZILH9zPq2ymClafFvG2XLoknK1cYgGeCqNp4lsUp6gFUwQYl4qzaDYhbGdLhAoCf
KI53QEidgpy5PeTX0h+82ofef0MOie44Fb9pLGQGJBbYszle2aibuOOFAT6EzsJ+RGeHEmuJtNaM
t7SI8iuwTfvT7qsTdM7qweM/16rCgUeZerhLQ01ZF2zxlm3pdpRO8RbGFqms4UiV/psTPfX330CW
pTCfztm63Dv4cr+RXO+OE5wTaiZf3OHvl57XjD2E6EPyxtU/LB6FH3stIIvTzPayCyH4cVE5s1Ci
TUPK9d15H2mnDg3KZEG4tXOEg9NkGq7+Teqi/oeT3uIMlEy1OzX2xnf3qnd/SuBEALBQOrHX7Ycr
R/f4Zg75vHhWC31lof2nc/y98tsT75W3HC75g2guscvlPHHY3bKTD5LI/wj5gNOSOK8nmTCkN3Zb
xsirxTUfeU5JepV6gyFOZpUDT9kSnhQ7rcQmLQto1kilSRKQCHuFCejw+fTXQAK0cwa3vBISOots
zLQz5VeOx0NC+Pek7RkWwTwT+tM7JGdvAR84r881QYHXVUVPW8p34WgxvPz9kiP+fZsfuI+eJ1gR
jJdoYDNJNBx2/wnVZh2mkazUXGf8Hol0vhj0lRAK4yF/pSjAu8b8w6qFHy/xr3P9OIl6Gyjebozx
CSmTrzKJOxeWT7ifygkV8kEVx+DYarNo81lRSiQgYl+YH3UVtlhiQNoZHJrQFgTwcwJ6qRPlTT2b
C9CpsthpHn4gsEFCigdRNNJw/ZhxbAGWlOasgYA1GAM2qAtjX4pUd6gbvuODTX+H9L05fGJJvUfp
Jcm47KDj7OghBMWNl6kh4+mfnP6Dfx9QsiNZpahMga5mer11omRtX/LC9akxMp4aIZaul+dZ4bJN
8B9KlIpA4cllg6qeAavkDvCd7U8zJdMTsBaFtVBv0ic23EafUuWp3NLjNoEa06lh3LXZVy9dlDAb
vdnu/hJClEnaSqiGnPuBNTgvnRwuzR4i+ff+kywtlOy4CeZYuJVgwtlg4wbGp7LIzBe4DdZBd2iR
fxNWurOaItuGteaOEDofYhmvLIxcgmOwwX1EHFea+EWaejcTirqcCfhEKZu+aP8f6C9gcYDrgIHb
8ESDSr9hngXazlJ0rBSYo8Laua+XN9EPW4Yps90Q38Y69RkU1T99F5s5M9vDXKRoimdqO+Pt/BxX
q0j0G3wTmFLJtbaaFq+O5g+DSUYpGbWxz0DwUUvKzpLGGXFWi3kYSTUlm4g7bHtSckYWLBiiBWu5
5Su1iqfJ6jIbphvE8Pw9dcknTYRFcdU67bsxXMRA6RnJkxMZjMgMnz2MrZSmMOB/s1DPLwrvqr93
2VJDI/dOz/8Ed3NmOVx/TFnCIz0LNTint3PY1Zeg0SRyeGtl5U03JCf9/U1TLTulQZrrWy6EarWb
HqF6YgS84BPFno6wvk0Q86sc9Elw9dSj4TLcWKHAE40v2RdFFOU3WRt2ysoSnahN1o1wuMefhfzG
WDTeV7jIwXKx1TyxIOwM0luvewb6Vl43mkGPj7V1snCDl36jn2pgHPHTzHvunMkhYkrCGGm3RKOw
kyWmGjmzOl3n+4gsW8/wt1A+d9Ic3/zYsiojRErfswncdyJbt5aLRV5B8mL8tJM2PluDv0Z2Q1ws
qXeyDklZXZ4sWjluEHixqp9AWMA+AZPFR2Pf7qMZGapaFI2P1Fc7wGhvZ0kSHL3IjHYAYIibUKbm
wX7GtFY/XEP83yd4uKk1SptqkAPTLXEXW7o9CB5pKy1ttuE682Y2evCQ+eSHW+X8GlCzKiuCxmBI
NUUvHAhH+eydUmqeQ0k822cdh2pj3r5lhdToAlEadDUX0/loftqftiMp/uEdLuH+g39EN6Pvp4F6
E98aCRcNNnV5f9mwuMcDUylx30k1UohV+FBYE/+ZCucokt0/pRpb5ocL5OFeWlht6e6xNEnvxqx6
WsDA0gVTVum7hhxFIJEotr18kvaSxF6x6zjMTyHklrrbpvOI8b8t0qsiCdKuw67acqmpSeKIRxAX
BdOA+f34cpW1nfkXF1Q5S60KM69ZLTiwfg4cSljqW5cIjl4gBOaxZfcn+NN0K4p2MVY56HNDAh3B
b6WD8v8S6w17/KjX2Ph8zstHuGL0qncfdDeUr24XB6MJ1ukfrMwyu+RtVSGobPXp2C26wOXOS+2h
yAhNP5I05tdQ6Vae/DcCQO1t298md9S2EtIz+H9T6+EWzMTDP7FGb2Q61HfXwxTqxwDEL8bYNaIf
wbLKX6jyKrTrYcG1F7fAd80lpAiYXIsjMi+XNHuF+I+qeYw7jE8AmRzhZEj9R7ZypoPBAL1PiGfc
21sC8AVp1xVqK6ZMqtGE9VPNc7AvaBiVdBKpP8b1nb6JU+2xgpgV9kJeAUzzXpAvtfEYvn7dnNpM
SD9uxi+iPjmWZ0P0uZ4J7CRuwQ7/NIyRnLRMHqBmrD9dwsEh24Vm63z7zzZk4jTvQBqmIHdBLxkr
PC+/KOIC9N2LqKg/uAM4+Fl1CXLBIkOE0hKYPgxRsDdFROIQgje5lfMHSzLiBTIT0MeCHECcortg
DCjocFRvbIp7O7Osqblrmt5dOJoAu/hCWfZvL5GqWxTRpUDaMQAhi9T1pt1fjcSgEZupoJGQIN+n
MEESgAdf085yroMLP+ov6iJLRaK1yyfrog1c2vaESbAEc3kZvXNYy5kH8ThkFM5rMvcKZ2Tqfzdp
Tue2dKPK8HG0zLxhqJnbXoBzK0LrMPmtkGPXBbSyIApfy1SWWF2eyBoTqRxbxgA+2tEEt525GsuG
UUAECdid2RJKVYnWdFxaARcdNmoO3uXSVaKfd2DMnFWScWjGdqZnFIztP1BglTsOjJn82gvapcKF
WB4RYjR8FY1kzzgpVy+0jmZd2huMNTjen6r5dlKtYumWh4gI1usGIVVDvdZ9pwdBAU/aE+OIuejl
o00o/t49SUS2oBCudQ0N8Hc7+T2JZtM/bGibphkTwq7sAhXIYpztaIvdyVOnF1rBvNvNE25DJjRs
H+DiF6CtNd2TO7nqibx2cpJkglLzAJjPFruVwOwS2OVBy9ml19tzohGNVg5eaJ2TWHzGOnynONYN
D+8OBlPwE9WduvJW+ifkNMPsImrLioYx6QA8RifXOXhU5+p0E0eS7gN7Jb7kB5rFtVpobe3a3Phf
k0bLxmDDpE92khZbGKM/XxM7vAicFFc4R1EASH+V5Gd5hwBx1lo2F/TuAu2xujzSIAkRwtN4HhA3
ebrjdbKsZaDBX+5bnq61bP/0nIU1jRkaaSChG3nipsA5DgdsC1z22rCHJKZtKghW4VpLOP+e0ke3
2GJcWstpNfp0b4u1wtkU8QCWI2DkqHtCj4o6iRKbvdGbmEMx/EWQ4mxfK2J9yJ/D9ozGBr8sNlmK
pYgj8GFYgyRIj7jY2XNwkCzlYNZiu0TNqSO1dp3hOjeJfzhOLcohnzlkQ1+rE+aBWTITl3RrjB8T
IgyzaFSAwIYFuE8FAGcVhBCdnBg40kuR9VS15ps8n6pjx3Osz4rciw9r9r6PCrUxM22cSzBjEj5d
OBAoVpTczRVFpEtIergotZsNatQ/iRMj7Lm3vtul43izjlWy0gwcvacmkd49JorWAxoLD8Yq9V1W
LYFDX0qc+3p/42fsS+OCnmqNu3U7VMq0Y1I53qYnzlI2YEOt6BdfAiGOdnYwz0JHZErwtAFJWUj6
MdRKpJVV7o8jrZcLHjNyGnU3N/OsF14CEmrbhaF/wIyyw4S/KwhxrqyBpQjODKFu6DfxUGvcLsDm
JLQzUBGVUR3mKqlgc4zYq5ov/0UV7yAwdUdw4q7gzYfTTSPj6R860KncS7OdJouvTdBUlECk+/3p
PZwlcLF+RUUJh/ttvxKM7uQRZ3etlLySzCdQ/IuI5IaPrR3KqrsI6PoOzeNJS99ToPjsDqYpHzX9
sv9ukox4ttXcNglERnnRxsYSFBVjglher/DDdQ5QgS/c1Vwyn9Rd/bdRbBRUJUrtCltHPWLGFyHc
sb5kJT6UmIiCQeJ5F4XG/NAOek/5RrbNR73zfva9ZD2fppIoxA/bDK0LIL87pH1hAA772v2HqEV7
ta8blhbcjguMWatZqmy2NU2VaaI2A3zUjjczEJQ95ZG1bejpNKzoM9NcbGvFUlFN1sqq6e8SFsrb
+QHHt7bkMx+3yKig1agS2fMO8ZPKTSsDYYAFweneaf/MF/lQtwnfrWHxiW9cO5DB4XzZS5A4V1M2
nU7sQoj9AQE6RhBsW7R/xL9028Y4nKn9cfqcWSP38aUgkuKdOnfFQCiA1V/DSFUCcwJpGInDtv0o
N3RejkRn9PhQpKtIqiiRhrElif2tcFt2p3ChTD3okwLyvbX9yPDBZ+bK+iRaOljQ3XNBRFatVIjF
eHctryHIa6RC09QpzSR+RiBDSNITeqNIxpKIanEuVdtL/fzrYCjOrLI0blZGiMk4cRHAKAzGZPCk
8pJcId8NU4Ieg9kaHQ9R41qvyJ+12PJZA5cRVOpikfoUFSwZMjsAWtuOcp6TEPUdgCCT47jWKNgO
UAkilZ/8PfGEIZbbURrGIvwQEDhg968R+x/QDUIUR8o+oGUIbI5P+GhLH6Pno6FJBGoGwkmjaF83
jbkbhbga77dgBL0FEey1AaiG3NU/FKXLCzHkbLL6M/V+qBuzngwP2IVafc8ZOqEQ/+ULG8mlGZCN
1g/xu3Zs+gJE1G6zkEzBCHTxAn93YFRhNvBd2STFY+m/qzXSP9LYM660tjubWhSoXEl6a7qHjk02
fyjuo12sseJuiv3DyYYxinAvhM64eL6qFg8eeJwvi0QuHO1BFJLcsXtT9Y8P++36WK71PyysKj3j
duRb0fsZMb6EXG34nU6/h3erSpBAAvgV4oxJB4dhU6shVl3JMv7xB3AL8p+QZqkZK3vEQHwkHSrI
VL2A2JpDX3rFATUgJbpu81a9ftJSIXbyAj2mPPC0DroqqH23usRmbk3/mC3c38sv5Wm+UCpj0jnB
GGlg+Nkk/Rp084Fcmbo7A+vFFDforXwSjGd93hTHMcrdgrIrFvpUgu2Dck3GDOKjGPncnidXSvYs
3we7dsA+AEIbC4D4RjP2jnasvblUDBhX5aH4h5ZbD17zPRbnP+qfxZSYRufKtidBGzL50aoS7wpU
WBqqAiDAhO1blf5tbKA0SfmT8geqOGXMGr8hPvpr8oToXtLhn/LaROMWlGe3WEDlKiZsxtFoO86R
4zVKnDB3EEPifEMviKn6/vgKZCgHSdViBaWgNRPZpDW6g73TFYyzKKS1MHxDuhM/W4iJOg02rUom
0sjU3OU8RS6TsjypVZ1KijympK3B50gOdSFqzpt5csQlGrtRKC8mc4nt9tT9qs2n7p+/wo5bEVKT
JHPK6cakatqGyomwg+MutwBnwAcgAbAFE9Zmddf20NQuM6rEF5CG1mtTUyBON6vniM79538dEDUA
JyGL2ohSpKjaZj5Yjossz+osVsjuOey4v6Kb+qAJw5tnLHZjOMolKjjYi9FMDq3Fpz4fKj+RjXQp
n6khIm9K3jKAWP3Wc0LGuVL8PvdKLvaiP7IOawxeuQXUEzlkefKBJIey0OrTx7H7qc5E3hB31zm7
OrMku/VbEELAWCz7RsCnjyIYr7DpoR/ysXYPp7URxwj9U7qZ7bMKoJCBui5DHqvyOz7EY5FrdQOr
hfKww7F7vk4EGVjYRrDg6iU5Qb3nLmtxRz9m65qBatEZJCYZwHWbWV8VrswkUoV2G2LHwg1C0NBM
t1AqqrH7AxJE6VnnQucDQW5O/VTjKMylBwgxnbCZJH9rOmQOIO60RLmRP1YjnW+y8ydH9iP5+Wcq
XicS57XjMF7PTDHAFxQ9RpMAZvoOkIXmiajLx8bO3VD2olC5AKHqiNvWeS+XBwDYpbcN4lqE2a1P
7wWENh/WjN3xragmp/vWILn/Gy6OFtbFP10eHw6EhbQLfF3q+XJksKNSHWBrnztbQB4O5I0OOYi5
eAsfnm8gp8zaedJxuRiZw2D+vZKMdPHKEvpoOzg07hqP3Uttivek0dfF3LF6JppNWxs9ZOptfKug
Pb0gmEtGSTF1BLHw0II20/vVZPHjzbganhYsS93hmFo9pz/0lcikdZqKv73If84D1gmbuwVsEAyp
09OqYARRnpURwkhD6Ka/be3v+TNsiDRsIIkTqYu1rti1lK+vv2LGYontQqK1XTQJ4Ajo7ew3fYAL
vHWYKyVu0f9YisoxeMg4vdyJzzGDzB0Dn8z/y0+Ys680oMR0bb0lm/eUQ+KZT9K083t4Uhl+Rjv9
TmwT+yF6sc4SH7zARKpt1UbTAoxd9bcZonzE3jv51aXBX1wN0WiPrELA61yC9K9yvec6LyR0V4wG
rJP1/MjhXyB96LHUPpG786ehkA1Rnn1VdBYzL7f844v5LmiN7SUWrzsNzdYwQr8L2pSbvGKjO3sh
63bbDcZVI9o0w8IU2SKZI3od1ucnvCJZlID9HF7aG34ROeyW/lvVGsM8f11lklzv7tn2wlDq7DzT
5ts8qtHtyv83HXrWjKT7wl7xAtrgUxaac1BcP190GA41+rNYuik75hzYICNr+2ME4EcXOKt/wzhc
kLfHKKbA+uZyASlgXW355iYFjEysyRbyfCQT3JabfJqcWYdy9ZD0y4Q5njhtyq1ql8WheRNC4OJZ
aCYQ+p1cQ8Ez2jujOSHtTIF1J8yH9fqxJPIako/3E2hN/RsGJtSrHDOPWN3mLF18aZ9uXu1v3nDJ
ivv8jkOtv6sKXjrQwV0bBNjk7xF6GNrG3Ma0zF7xi20LxO67afdiskNpVam/8mFmsL6jkFEe2UPH
dtEt2y8xIMS6H6FaYRyNLsE8so6kQFny3qiujnFCYRStgYFEOFx1O89aKwCTuLgnmRxU9km0Aqqi
UIfBSf3hPB7Zy5ZELrp9PbSVvZj/t3BiasNey2adPsG5Qejpg5+DfmDwFTn9g/U8JreZTDs65IzD
Z23CoLY+HbV+JUovhqhxqzmnqtlwFkI70VXtBtpdoq+rD2WATXLexIRlPMrBVdY/U5nTF7Q7zUXK
mwhO206+H1W6ZeB4bODfvbqdwdSeQEELX3JOnU0WTNv7IUDcByAwfA9FDwwxlISj7yWBtsXx/GFs
N4uYyxwCaDjE19yv5avZCDk/wZWSufx9pqEyPbDXV0QUZQtPgKMNHysey+lRiGBcsBCmRY7joz4e
FGkY8lfJhLufYEDqCr1DpfuGMa9C1g5ZVxMT6fK/OC0pC1ojl5CX3OhOhY8WbuntNTq67tETX+2y
dpQUdhQjfuvppD4rFMb7VVjC0yKNQKmLmrEgH4SBJcDRSXbiELM8RS9eyck8dAvQY1nONVjFV5Lg
S/iHmuBv3Lj9M/DYFtohs4BliDflGiPNf/InVo3TpnFoINb+kez+SAbyDLW3dcfLpTbgKPix2qYI
ox2aGrBP0psRSGZAF1TSjzuEqq7P+owBnp0Kt5FGQgxBwl2ocKtULem6VmTPF5EiEJfRNIwUU+3m
LdlujNInnYlGvU+aiviM3GC04qsJtlE6940f8add4Q02r8oCK/4nYW8utzLguK0P+yw0Lt5g9DRP
KZ/sKx9i16z1VfpkxvIET2Y6My2kZLw/4SpWnpOMvcJbKbPz+HoaQaAu1kORQm0ov1G+ChOwb+R8
N3WddlU8UVXhAF2avRvAmv0+SPove8x3MjW07OApnH4FwKVPsCW2BjuACU/JZVY7ULiTOqsc/Ol9
4k3IzodwX0qqxCxj7rFpUFDnu3ln+v1tTSRwenSDAzhRhqH3b+lJamLluVjUnlAagBrBSEPYymuD
W319c3BZxUOOZldAEEEi0y4AoDEZZRIaFuCobAfsxkn5CCIjZIuooFFOSJdMcy4uEYSXQiAdm7LV
XjOBJjPb7/6vt1jcNwj2EtQvx0cbp270RvpJyKUH/wEWxR6aNW4sNREujRr41tdZplJIRPbI9FLt
hDDHxyjZAK+c/pwiAK4XJb98Zx/k7zs4dMU2gacXhrGrTamnnYj6AY4IPCskzPf/GE7OfdhVs/Ft
fLLbwONtd368R26UNAolJDX4YnQ1BSABhgC5VAdOIvsnLb89oJpoXlBqh2WNz74bk0gw50VElKDm
e3x/b9msCULFNH+8voPG0eZY2R2iKx49hnEYNXngqSHeKbOzNxuydGJlscpCPWynrIjDxeUEQCxZ
1YUYKCz7Ep9smXd7doqVyLCuu08NqjtL8w2jguWOJjFcA2xZZRKDvmQ1y1pdbpfL0lHmABOhu4iH
E9KHO56Rx9IUW83r0/SmFFaGWsFdlhCjsAMpHaIpqQJU0IUg4XahuX9/jg3qrM5dmib/wOAFpJdq
AEeugPUCnKYzjvmLe86opYe/ulUGWnl/Kk+yuCcqT5/tus26udhOjAllXxj1i4XdUkgYq/XCfSqT
R1V5WK8RVzi5t+r1sie5+LXYGYVj/BZIHFQPKwG+3MT7xMuHiirWYogQa4yGhkcgFiUHd+7XBmBM
95UZQpCP3BuHMwfourlAHfzG7sPo+cAqAW3ZvJB3KrvQ1KqOvdbgKdAwwT5R5s3ebVRkAnFDbTrs
DC6nfAq1jMXxrfe5XJm3p6UQDWxpFXfsMFWWA88BjvYdsoMSKVrA3muuHBoXTs6iC/pcvXmbSsF9
28VWGF8mlYIyLvjUBL7I7MFXPNhHO98G6H0cQ9OOFVIbq1L+v/ZqzgdPnGswUx2C/uSxy19RGLvG
BAeBA7lpyctga6QOF4W/XDDuI9gDq19p7ppEyN74hxomPLpeacaEbPfrsG0ZsLfxSW313Fgibn9O
ZfyfW1aVDisRFWAVB4MHzdIBVFSMhuoyWHQiG3FVUt2Cm2pXAKVRvHj1A7J0V2z/TN2dmuotZuXL
f4eCOWtAvVXtFXCkan0Pis0GjyqxVn/h6vyt02H61WYpVfTr1nTQmGHuEo2+BEDybgyUiTZbpkPw
sFff/YB1P0dRM6d8m/buT0i8ckqvHdbUkc7nHwFcKmlRUrBdQMOm4r4JIw53f22ej/6UPJDPmTtc
CFlGJlRAvypGEBzjBX05MRFN7rQjJBMTntGkcAGr7oqwgO2/dLPHzEg6zFGg7JT8aoT/CNG5XVsH
GfA/iAptfXyALk2dINidGkNG5fwjS79IGt+sJ2RyUpridHJTqIA35ui0nwiYGTlCwixqTASvQAUe
x4IWOVRVAIIiPhFL5oYVGmwhroXh6YAqk0XXZakCLXMGnEEgU86E4xdoSDTz8MxVKjqArC2xrK1j
ekzv/D+cUwY8jfp0rTjflq8ZWjrQev3OTKnwwMNmmor3GcSOTgQ4BuHRdAmnuspx/nZlSbcgHWMn
eoQe1y/AwnxrtN4S/vBezEYeHz5mUi4hDnWLc0ZY7D9LLNgts+fjcD5cBz2r/PkAQBvXwzPL2YmG
Z4IJvgMERwPARI54BBqag9oUTR7lPUo4IOVK2RjlQP3dSjYYaxnuMq1qN+qHVzqZcjBSTA8mZdem
x6V5lNBL7SgkWY0a86Et8Z5H+7Iru72MN0GW+9ejUXCSBy+64MnlAR87M5+MeIpI8tAMO9nJToYf
MA0erWUMYqbuGEdKdTWUmfIECGqYgVeX+jf8PQlb/esRt/jIWBnjcexorhl8rROYxQruN0MkZMr1
jr2czVNdFVAK+6s28J1XF+pyvVJH8Xrt6jircNAT681c0TEk+Mai5lxCEshG6DmZeYBNgoeF4SkS
AqSjLcibd027G0DJohDWlSEPMUhfoG7jAjqVH5zrZqsiNu1dZaWOaiKGmV5MuNGohcDViKnth4Af
GF2EnYK9IzLIVH25nDZGpMVEoP0XBqW+DTUkfhRGszgxa7slrVzMwnx3Z+8E+Egd16a4jc2nUhe2
wx6tvtBHQK5G7rbxSpCrS0IQoQpvaPL7ncG/MaSOL4p26nqRHX/OE33tXt6Vt6wipN4BC7qRxOKb
0XK18k3j163TCofgYTXchye0IcFg/i7qf0/ENXF0ONKqLEaW/Okl30vzu7xoWJcY1Dl6Km4Xusa1
ubc11eoNMP1mM1KJLsuY2CKkR1WfMlgcQn6lPXkgJn2GJwpGtAwZU7QkmlpE/lkPsuqihiDL/5Jz
sDtDnCPGJBXh5UKbHiYkjfK2Ulpgek6FvSzjdM6WdoVRU+RIygW9VGZ5gVABnx1oqikdC1WFRpwo
3fSSM9cyGXbWyV5pv2QGeHf+GAINmg3oAyxApnd7g6pIxAsXnFa1jXQQOJaHdwXI5gUjIki8nUSA
pQ8MrYSxgR9e98P5Hb/6P8/c0vP5G5eJDPA5vD/S2xEAQogCeeT/TSngYljUq3NDypVArutoSic7
r/B8xCkE/FPTOeEOvLgrkvEB9dTBfgPOL1mXpIpIAuCeyK9j5mLiUzloqclqrOp23ZzpvhlxJHni
K+KIWZ6CR3lAgvUFMmJk7eERXMYAL3JXKZJF28sdMIH1akVgLP7VhJ4uLz6i2hlGhRYfmSzbCPVh
C34/sIGOdQznPi/F3IrsF7PW1ye8J6NgAJ3crR+Y6EHAZzj8yHZJOkqcXKB0YvmzUcmT86g9xQLt
iSWPi4xV5DmNuFlC6QkxhbXrvssncuUUYAO8t4wqAY0RjfiR+yTmqATr7ztvi8QsQ64mpkgAGhFP
ScJ8iu2Fu35LR6e4/3Yobn2MvhdK8MG08z7WoN/CpH22S9+GDIh5/5xNH/bK25bbUWuv+WLNSzO3
z+h1m8ZYWQESfFXAzZMsXHBUfOf5ErboSt4fwAO5zPwdyQFCtppu98srFwh46Qg7dNwv33yc+BPo
eqxZ/xXseycOSG81N8+FR7ByYirTk/UkhPZjTzBjNHZk7gKYBHdX2mboWDp0iKqiNtU2ZhbkkoVz
EnhwHJfmWJ8VSCXSLeuvLTrGX5Hg7JttG4X2UTTQ2LV367TZflXfdlKIc7RHkY7kYtOkiylbhEbU
BoPmtojnaGs79I7ZCENp8hNDKuYOWn6dFLYxh2MKUDXwFzU+kvp/NRQLHoqFSOxPe1++2IXofkc0
b9XXc3tiuCuHVGuxFA6pKf0Wlc8W8sM7oHTDYiUPdMuJP4vA+IQKxyrrWbnhq4kzXBJUwzjOOQXr
TDGHdz2fM4dG9Fdnqg/V0XYa6pLDvmxhNMaw2Iif6ck1pDwuR7cKnX8bSG74TCwwUZ9nzP8/0l48
YDBHu8GjL5TkVzx4wQdcBCucfZKV/1n9nG7SKZ6reeuZ6A+Ts8YhRbosZEFhFp39Hkp8P802qF1Z
hU+ZEgWMxg+wfIuriONZsk1bVWOlMN4gHCUK+odi1s8Bclvd9o2F5ZsIYwkO5IPaUBapLunc/tPy
JSPIVDwYpMvyHnLixQlehIzf+42Ih79A6AQSypxkTlkl3jCL71Os1y51m+/RU01QGCCWVpqxaoZL
mHR4h2W08sJ4qc0Ks9gYp12WrYVWpn0WfoRLsXk6m2mXA+ZGL6B5s81rYshBdRBlzwmJKKMHoec6
+W+sI4Qg/RQezroYZRJ4gFqDGrnvnKqr1MibRL4dsLdbpyeg1Mxb8EbNHsmXPAh1di1C1PIXKZlc
NZoAuj9Am9eWqMSlvmhH4l1UHBMm3NFFm8zqNJDB8eXLoDLe36mD6CKp5ZHCqZNLYuf+qr2OtMny
PwppjScK/193ys6sbeWvxSa4Henqi99Bdv6LSTAshvs2356bn6JBUiEAkQjUeFtGFRBfihBHCdT1
XPzg0Ey3v3t6Yd8cuTbIhpcdwg6R1pM+LnAbokH8poABX/y8kpEHx0NSY3cCQoPqYZyJ2kevCswu
Vo+mF6quzsZkMOtOdDNdCCfL8aR3g5lKKFVh/1q65rq8rU3LAScyHeXnXn6XyKTo/sag/liekFqs
xu3svsu44LTfV1DW5n+BGY03CGpOoR3lw7LFq8fr6y7dySN5LkyL8Eq6EEM1I2q26CoGlCQJduWG
npQ3LhR8i7s/OYUXBVvmQfILcfjOwSU0KIt6E71vVbRerChtIN8EyzFXv1qasaq+EGPAuCLpTsdB
9aVOng/OwG8LK46Oy/V/ZE4zlxpB8247N92Ac1isEduKwpMuM9aSvT+rmCDF8Jx3jZJLuWpG2xbO
Cbjep+P3MOj/YYclNyP14lTD9JaiuwrrhI5aLRCBVuk6Fkoxd1qP/CpPy4QF/j3IGU9PWN7XXoDi
Ln3H0LbzHFy3pgM+3aVPFuFgk7VdHCsOs9WrVbB5Dm2Rm5WfMD4VcYXWcsCup1EFpVQGS6U9AQgq
S7FSSZLLO9XZhbaUkf0yrFlX0idgEP5giGwJnIoUXywEeT7nnMFcGUkgrh90sRLoTIzMsdgdw8yj
oDV1HmYGAaS34rZ7nFz151Oem4povDD6mVkIIfkTDGXtKQ/xlQmnk2AuD5ZEKxn3DEADHYdItdZP
yN548KoR4Uz7Mz0zZb1SPvsadR5VHxree3UiKXc9WcZOIgFmmpkmFG66ndppI2Sfr5iQy84u+YGP
dvEU7pp1LiTKwUhMwDDeICKE8BIyscEKg7xNE/IO3jNOQNHT2RHGFiu9k6qFk8c0lqgmgZNm/z63
dJiMK7ux8659pBWCaG700dcQlChm1x1ccSKlGcytbVP4oaDJWjaIEe4kuNiPvB9qVQmSYSvRtKc4
u2KJSZSKogzlobow9paD7lt28wSv564fHdA+x0ePx1VrfH/6spdCzkDsMFtloyikOYUTOmeBRFBR
vIGVPAiFfx4QXLWH9Xl0nVxGM6oU7e8TpR5PYP9QRB5rptvX3DrU2GyH5hgXXLMq88q38ix7Tw6v
u7HkdTQnsOArTGXzGmAKmmR0a76/nDGZWxVkmMkC56ML/RJAOgLX7WiTS6bKsioWhWtSe6pYKtfn
1rjmkmyQtGAsadGTRAJbrhLGMQju1cq6PgOX5zsrpH9KzDY4aYVzEtDIo11JUfRcTU4uxKZc2oQg
sb5/+ZWtqt0yJR+QnE6lPT466gfz+R34LXCKf/HLmDrrheJKyVRjGaEsSGlXIkJtEew9XQqHdXQf
chLh+vI6ezjwccdNwOoTVr9FYk7iM1B1oxN6mA3z+t+8ZBNPrNQ/C7WcOqU6FLtlzedBKvsjAWKT
57MPHWfigOCGiMDI8E2rOjO45nx9AEMSjnsH6Cdjlakj1CGJ8JXFDR7NB6BAdKDOHjLu+e8+f+Ex
e9VWH00U7pIn1YHqy6p1EapzXiHOsruEyHWpOG2qpXX2KuHFe/J5aChkLxH56b3c+WJ09vp3JSuz
mJ2fqakiMLMWzNMD7YtWR+Mv0G9ZrQtjMP1b/n/LyMEH7N9rJ0byv7Q1uHWffT65CqCMWr5cNDKs
WM8WK/V6SZLI1RX7szrdTYxDkRQRm0AUwkQywxHQB51r9vhpzVMj6jDVPpNrJJRMwzmOaDaajKAn
XEpxLemHhMfRlUDdt4XxqcKHHnPHJR3OFhxppcwnBWzRwtP8vVv0dcEczAPtg70Ya3lsqFuQS0GF
gcNnP3mAhE29pFpsqRKWd9PSqz89LG6XR/HV3HcwueHq0pcpNFwW7uS24Qm94fSLIljVWFwTGklQ
Wh8KhZpOyD0v78XwR4KD401MFu47wtEEG4lPNytZvyCKudq4BjQh7AWf64NV67m47wYPNkZJUJ5y
wbP5rthGJ5iiIZYDkIKGtPQzgxZkUDR9TiOpCUYy7QY+JSf+IlcV8cJc2lNoZfPNQNj+2iVexKPI
z3uc2m1D9fahFzWXNoHnutDapZLJmG+Y7y0lJV5t6/H1lhF8mFUMzcAG4+261AWx1pzVrFC8suP9
rPBjxm8zw2a58DE8D1P5QmNNSNOL2n8RF8SofCB9u2MZ5XVou3AB0UQ7EDFAZZFeNrp9hbPrfypa
dUvEFL2AjsLvaFK5q0jyTKFAHRYRunLtEIGIIhALTHejm9rNTL0TIkyoEPXPmQcnBs3H+ASCyHJM
x9aq5JMTqJjs4YFB9Q+Z5MKGhcz0UJUHPB3VAGNE8cgYFmSoE271Bd9aUjHUo+UV6UboVXIWXjxa
RCdd2ozpB+SSKOF3+TjfURQWXEDsXxJesZdNBlpmyOB2/kW690YFj6v+BDQkWqxTIC6vjvTbvfNx
GKi01UFlIX5ZRCNExq6KOdKRG9NaBcuzCR/LC2ADRKeFPjHFZ1V2vXPBIX1WBYnmug/7DAm7EvI6
iushrE6hgb+rmkmdZJTQ7nMcz718xs2dCg4FsDozNZa2/PGmClTG7DpecCZGTfWu5Z/IcZ+XbryO
+/p+ATkGmrxxeCqKFhbTWKuuqSuS3B390dFk9up8tL7LcuanET2/DdUrgca0dswawALM11HBnVvW
g0cwvUn2+0DBUKeAuKKA1CWEjhbRC+5s9lNg8oOK6dZAHRYy6IR8MN7QkamHU+zPeu7pcmk0EQ9X
splsT+/cgYF9iVQUReKwANo+4UHONxPjkOGPl0+TDuRhxRv10mpnNHVIHiPe661joDN01zS3DDDc
ldSBugg9tHXGj8FG8Qlo4f0qwK+jY+mgdibbZpn1nz7VPTBVyrb2Hnnrke4DtwK8tRufYmADOYPf
m2zPsyVLdToQ+E77Nhi0hi7eRLbZK9UZ1RhX1Oa89yzxzOYDYKIaqcfd3oNO6yYtsTeBJozL3UAL
bHJ9ct+dDMhtVITToPgeJwVHzIaiTA2CUOvUN01lMR/rFbbkARiENyFzeJwNGre5q64DiFghGOBW
69edRA0Fbwh/xkwrxDh0tHGnuG+O0Hk4uDCrh8PMHD4Q1SDqwxF41G5gaM2ypxF+Us+Ho/9H3D2K
yV+YZvadN1SpU3g2gdAVTS0HCBhkanSV5Ek7xQgr0y9UBDjBLhBWei/ngQMDQoZNswdLDaBd9AHB
djVAIMWGAMDVEvaRzsx9ovmkKsc3ypKauN4liPF8ciYGPNin478bhsDgL+D3W5dXQ5L/VgYACPo5
YlDES2sj5vC7AcLqyl0glr49SzbZ4Kbh16BRjN4pj9hYbVEhC9s82yoTu9vf5hD3YmVTvWbD8Jt9
VgMr5PfAE37ibUNrkeP2t2gtX4Uz1ER2NwvmW5lzfcTN+O65PZETnW/4hX2AXYyZa2hj0eGE460e
8nHMjyZXgU2vXNTgGN1IBFPEfillf75+Ew9Zr8EPTGM6I3zYueOy70U5W7bCmh693U+x2qR2DbXI
pNIS1fcQ0UTK4JVzcdqcEOlgsF8R9j1NO1rH9vFYneb0Eu25RO7Ucpn0LGOqSZFo3HjE+RRC2wOb
qTIWjS/YQXRrAS/tucTM8rRV2jxe7ZjAMYfa0XGPS3aQyUgruaGdinskFTrL0lf4mXAlZjU0Pg73
UqqN8t8HMnRyOSWL3i/QIGecWZZXCs/1MkmA+DCq+JaplicDqJR0q1qg5O473K33bvr/HiWKwEvR
qYzUxpnPGJmHhlLWDWtbbtrCLPQM2fp2i/a5FPE5DjBWqtREA62v7UCiu7UjJZg+fFz6xkfoh5TE
imoRoGl4dZRBSrbo+RvpsVovCTS3/jImRY8yfvrdNMJsvO2Ko4tOhdU7GxWtCE0FYFysW3gdultx
DlIhY4PP30vwNALlP/FwdL9SAmV+0QToGFoL5Hs1b6wtTSPhtK70fFgViLqa87qIgyRHR2bBYpYF
LatGUyNuNMoJ40YPwDtBtVA+0nSWrL5eb/acLylHSzetWvk+CTEUkdTl8acJFgvsMbFLZRt0GnOf
qdq7kWYemO2zF9KK1T8iyur6Oc9OGtQLx68Pgt7zBaQT5FCLM8pDEw+KDVuicqD8nhj30fTADZd2
077JcmjvNs8oNbUeOcjsGCcFkqItLQz5J7oMTQa91dvCX09rDDQI2IYbc6LVAMEZeBY0p43+djRv
0xJiDrVwfVClKlEL27LNH0o8k1/x5OYl4KP36Ivo8WBMQFVBlIKBveN22bkf+9g50U5O/KdmewfG
r5QueHoqPpshNac9AniyQ4JiFwyTcXM+3pJjkrBdBVXEf8/eoIDwYjFtToW8qvH/Iv2aJG2whNWY
2bhme7QZjzDIKmZ7j0Y71KKFw2V+iu1sUjMdYQZzk64z1nKEnFMvfvuumw4l6THQ09qkFcM6byW6
Nji4BNqq0oJFxxGaxTP7ng1nDmYgH6zRaKh+sMnuS9wsh/lUy9i7osmGqNAa0lk9sqMLU0Wq4gpC
Gb4LnB1yhGeXqpTc9kZ7qpdwRLNYMjE1DWzrpFZamPmz6e1SQ6V4SmTsZBfIwsF4AulPq2XOiaO7
Fv4iYrnvdZNQ6/KXQyOMoHkASs8A2czXpc2Dk5pU/92W9MCSy8dMu0X2VByvBYqnpa2V9UGthPg8
4pQQCLJUvhvdkuJvuku9i1KdjGyqO0+hldi1mHGdPB1dWwyS22PpI2Z55ymu/TpbPcyIW3HUb0Gu
zC7KPXpHqQCMgaFrzkVlwc7WRQdtqvbLiPbsjXlUbyEbLYiFvpywKbfVgkl96O7tgXgPFqXU/GLY
UubK2JRSQsMTJyO8MIAKglFF7wRwnm0Tw1dy88DAlB/64EG1WJFifpaOMdZsJQg38aBAa0NoHmAA
7nrEGJoPLP995bVH6rL4uU39EUw5bykFUFilqRI2vw0+lq+t6FzF8gstiGBVnft5dIUSMzEIGqcy
CkaEdbuminAtb9QQJKD+fhJCK3Tv7M0ZYiVwBi6ii3ks1aKJmum9v6mju7z37nTSRehCJwpnYcNL
Ch/Ai+GfnO8BylgHYoS7Xv4UsKJK4cmk9Nqb+X5fNPq8ZkSLvtdAO2KF7BfLmxh3KqWzkOhwWn9y
CRAV4rgT2U5/IjK67l2IBS3MsIrnHldxRa9sw24dY1JB+umJ/M2abK4soCKrBkk2bYrVvh+YTtkb
wcYci3jioLhKYNSQwzodchZUk5x+w9nv0NBBnTo5c8Q9pgTvCefVapXKjDqjmRU2i799j8k4ExlJ
2yeWKId19xdHuYvgBrQqGWQ1xekkROUWG+2FL9UF9FBne+D3FyQRkV/C767NQwkoRU4cpFqrHGCE
NOOb1HHKdpMXLXaPk/hC48nOB04RPOUJT7LHHz6KhwY8h6j0+BNLPu3doxOszyU04QNNZKWczTNs
rhL0Xbcy2ZUpbnk7gI87dtec83LKumV0v8FSajZsEfVbXzqEZbQFIRrX/AziCjeJuIUPMCAnGYVV
RvVtNuus/yB9pfiu0+FTqWJzaBOLp+u+4MLpCpZXMVQsAH7W31iZg24gG1gmJVnsS6Dr2VuKqAYl
gdX0ZAxEAkv1ILTqvSmpxMIbXd7GPGJeRWiQgZkj5xatM80Bu4EgfNwSF4V7bxvfVWDQvQXTBz0J
Oo7Vk4Dwl6wvHJNE/pq4H206uNDaLJMyzowRdS/Lb31uH/sJ5moPSVNcvkvlJRpNz87jIfrDNEvs
7bXETPWpzPcE+uzQLSEGIZ+4ANT7DFH9tZ2F/B+2S6NHIO1gKSnbvIjVczT/PdG4lGxqqal+KBij
3kVQuwO3dzfkP5ySg+kLdjGjzd4abi76ebBsE0WWNLrawtMRSWQmWVi7wvtEG7CsRVHSrAcdeNzw
aDUSYAzD2JIf0TfVf+9ijlEVDOiSYwTUJP/X2w1DWP7RbX0BKIjIXYkOxos+20BuRPce4F69usvk
rqwO/1hl7ydJzBY3Q+QwPwLyoL96pFM859WgtC+7VC3VVbE0ZpYRhULQCnbRvim3bJyTNc9djwoO
m+9cCZT2Ulu4Pvv0aWkb8gd9z90TsqTs8IzBgFwYuFfc3iby41BCF8zZTjbFX15yt7gMxDJke6mH
YD0Xsj2apauxjEaqv0BmYRwf2TiVOASsz1+PnttDO67vT/K2mJDzmoYlCTEozFFjS8Jv24D5MTIV
PVaXf7iMyy3YuYSZoViaQJtQ1d6KEuW3X4j7/+Ri8jvGzB36mQlWfUyZzoU0erVxXbXYLolZ8Oyo
mY8EmyYy3FN/834FZ4PQNceSI6Zj33F1sC+msdwBF7AxooVeEwSDG4IBnpvU6ZT/SWJ+wr77IiH+
KF+0XSSmcPYi9aPCSEx4evPKpha3X5qn5LSwVP8XMWG+xUMXZbKdwu/x5Q7SIaPJRrKcglqoXpqM
2lPiZRpFr1ECDNNH4tWal2SsVy/VI2o9qg3VWyTPQULI6goE/mkuPu19XE43IYTwUvu1hEyVwlMX
lN41GjwqEV+WzGH8C7IPy2K1rFStsBmLoY19xbzGVTvIWkd6RZwFzYi45+OyugUPPzRvJftz6yRc
7ElrkLtPpXwiyUKnOzidOwWsgzJC9LK6nZqfbrOahAEfEuc/bc+Im4ULk1Psj4MTfmGeGGI1aghR
mZ4Kd6DifLkHTasW1Kj8oToIwEoGXndW485QCOo7zdtKbv2XTe4N1E5kqwzGMovmZbhd7WvNB8KB
/1WQzkh9rGMpLC5ySp/7wE29cggyZquNDjge5R1GDNHGU4vClcP2BRUQcmbn4aoxpsXzfAjO1By6
8/yH1/J+Yc/nOCW6qbBPzI1MNKr42JbrE0ywGLfJ8wAA1CuSIzr/l6Zgs8COkoeyTaFq2DL3C50r
aaQvqfFVjXZxRKTVdFE2z5JczkNOon4NrnDbd7i33yYVX+i3dctbStTcODmnkDfH4efRB9FvcDeK
c7/C6IStchoHUWvkO+PKTA2XhSLcBmKZ5DWy98yQjngUtqFNSwzf9Y2dmzabwJdDH05lznDWsCSx
mvgt3IyaUpcSVaFvsXROGTe7d73t2BisyC1iivJd8oy2o2BdC0Dp5PGeSk8Y/GUEPqE6u6+wz6Dg
4/N1w/FbZTyCdEEkS7mbcoSGk5Cz2w8Lpnb2PDFhBBYt/rFdoPmxwuwnRVlrDcqgmOH879KG/R+F
anhM6F8nPmN/6tMFZXZxnU6T5tKbu3XqvWPOp2qb/1g3VRLltdJBAAkAx6LNvN0T61ijnrdl0Tqc
0Ikv8N+BZpYg4/M/8nSfSy+YqM5I9k5tUUGXXwCR6E2ftmavwCz2XnkUT+gzqwvE8mC2c5MQ9VNn
PmNhgLd/7lKOfISjLBHvguF2iPSM3/Ntiu/UMsneKNqSJZvKIQvdH4nWc+cAY/Cpw9vGI0pgrYju
wZPSg01eADnq3V3qUvlx6pIs8bFOYqz679ahXgVjVorm5LyzAO8qGQkpqNibH675vmuMEmtktBRH
f6rNu2O469LGOZddFyFHZs7lPqojPkxeBpZRkYAvY0+NpxHjWtSkexSk7pzVrAzNRToLfZf6yQvm
4J/t/9H3dtp3Q35OuM8Awa1OdA/rtf3BiYBpeaTPQ07d3ibusHXrKX0YR1RkYHkdgxp9ee5WV+vK
on92VLQJGRVi2eSSOGSYSHOCvixPNGbZzIoAfiK6g8G3wZ/LLgFzFBl03DurpckDNDpNdNLTFIRw
p287ScxCiD/ubgaaQy/64iAtoP9YCq5qlq+mDy80qhrTZCTpDNsep6p5mv+yChWN59C/gnRFoj2g
LbqB0fSOAcN3mrlJFcsGdDspDDBuFiI2CitIzo3eRzorAuuxtFHDFlXyO81tH3m3fOELklW8upxR
qLq5HKfKp165LUoNJrq3BZ6IG4coTuNZOXsGsB6X1DI1vR58qsBvv26qI6EgPRFbq6YFUa7UkHOd
SC+p2j+0QKWIRzvM3RtFK3svTKzr7/hov0GBG7Vo1oU5g4lnDrMbc7GialN4WLYx8bFFWIJqpUxe
fGxx1x/3ZX+yAEfgOFKMdD697hGZFjapB1nc4IKd61SF2tjb5Drky2x5UktidZEDXiRyeD8Q3gol
akhZQb7eGZ5CDmSN/8sxNVGoo/rhZA7AfiHo1v+KUYWSAMIoy+NZvgUg2wzkTfQPFC+okX5HauDE
bVuu90dsCOyE/EfUJ1TizxOkHd+B+4iu63oJ+a369nbdEGbLK3opEd+PePGRzCzSqcJuSpR5aRRi
wJuLaR3AR4/bucCzFyWq0uCJOIMnM0R7uvLjfuS3QHwEhK6AnCAL/uFLkTYDkqu5jYkifgWUp5pi
FOMeg3rV6WlzFQxnNQpPUj4dUcOLqH5Yb5r5e4S4kQZ16VTvQVWAL6R1z8UPl4dqhM6W0o2h6iFj
z16apKZodvy9UpgDPRIebu+yiN5nB+Bc+xYoSMJ4JFasIGL8N7ihevmcPG3Aw2VU4SI0cCeyqAGb
tThZbNZA+wI7zb6rAWoUNF1GTe/Pg1++1J569Yv+xZvzXY6po1VpZfgnr3dKkpjQoRzORndw2Zxq
pzNQVWVIv/Wae3N/GoGGRNq00zbR+mw48aebsWcpbIC5T/EMMxvLOoT3zBVwRIkFeVzwKubXxCAX
SDt0MAs+ECveQ1XdPsSXq4OF5HEY6XzHqLwRlTQuRq8VX/strLumyU2g0U2VzSf3n/R1MXs0DaRp
3UM6zgkD0VI0F0eSuPwMioia7GvQ8Zl6bkjGQ74lUP5ZVZLAzh3LYRwMmxIqh1sIa5ErPP2ObeRV
dzevNcO0qt3T0Av8MsMtVeRJx9qGRfM9OApnGxrZkoQLk18AxbFpW7bGC3abkFgswg7E5gTgfgXW
lRiy6204hMe2gtdpv1aL3vKJ8NDRkqC8jb3ixUoQmIALtvTB25SMz6BBzrDwo+/c8vrbjcRzpdb+
iq1SQrBAUp6+R6BpMUjQMtjDsSiTN+DrAyRg4zkZWhbVAv99LUgjaWZ/KfTV9oUgi2rsycn9hRuA
Nfd6/oal68p6vS1bwBbX6EJCmDIOa8+evcKJ9QxhxCTHOiBIBAS3xe50mbiK2GO0DziJ+ZSU+tK0
hvmxCVJlPd3KEnWGaKNAJw6x/QJ+PuR0s9C4Bd0Nf626yJJ5+wKSjZ/TTznChjefchTcXcS80t4i
jcIWGNXBUvoyop5/gw9Zzd9qmf9BUXazRUlffrmGqkkrvQHV/5+rk7c5dMV1Gv72nI/clMGw1qn2
26w9x72w7EQgtji4ADQUJ6Yge+RU/770zhD+uwmeXG6Sn7rxjksoHmw64bVxdAJcvMySf2OOsgx2
6HFpoSTniekSIDEBCfzGUdcP9o/F5DLYlmXkfErTgIMVf3Riy8NpGvy66P550y5Th95j+ORxFur8
TlVAAHuXVOjxHT1+gvcokP6gqOV3KtyyOFk0JUfDGqBURM1LvgWDvk//DVdeo1wM1FUdv28+310V
9B0DT5z8MaN89+fEraYONE35d4xkcpVmj6rrFdAhoyj1o6u/Cg02RvSK8Ge8+SvFydiLZeqxtFP3
1hkzFcNYtnvCUNaJlf5H2FGHGaQPVWetosam/OTsO+q7khrkXsBE0Kym1HqFB4iW4sR1pe0OSi63
VUHhBkyVO1dneQxSdEVLaAd6bnJlItMbgNngHw5uVo05zZV7c6fIvBu86kSjTddBTKr1NhMWi/kD
JUpe+uVvfk9F59VxHhZ5uSL4neRIohIMxfewSiN00nFIBPCcQ220EiHpZqmP6aUGD9CI5D28VFb1
InEAXEGOSaY/jKEOkCysw0GAhzmWmyUqCQdVcQ8F0UXWQmzRmDaUNkSo3ON08hjiWZiOW8Krki3b
0lRQK90zGVwBgWBLkeg1ZhwaQ+wt+FoZUx1T4fzRmj3Oa5ceplg9UhKdcSBGHqv+j9+3SSlFVZw5
SMTf9YxoRBgkxdWpv5vfWDQQvXlWBeYlIKx8PZ+t+JPvvJ4OVtWIKp53qVvESoiEiOPrWIv53Gp8
j2hO+ilO1q+uxakZquKLCClIw/9VT7XH56r9Pqj6jMrz/lKdaSXJ30QO4uJWH7llPCoByr9rpc2G
qzNnTEBcJ/1sXjHLM5m99bB1iUoLRu1KzZgqjt0/FIpMe5W/+BXl3XSGtbIhpnjWSX+I/6L6EN96
vicethuLvlBp56HhxlxV9wxnx9PpMBJNrCAKHMRzRYvbhP41pd2TAhw6wv2B9WMNGaWe7Ux46S9z
7jyo+t197bgRAVbkyyt3kUa55VBCHchUTiQ/YKHdwJ+8PQLu8iYtrg73mNV73++xV/0B2mMmVMvh
Wsu0cY/2wzK9PefwnY6YbBls3GiR6fH2I3nEknXfHNFMu2mNyDJCDjSV4GbyoW883fy9RAJUIahC
iO2440rMjx/810gLYE3bfjUIza8m9I4tnIAtM+Dd+fzMG2pVyQDPfs9eAU2z6kLqRFy1fdnZj+pi
ww3nQm+TEl5RSudB75bM6IT+4z6hvkuLnK4iqmj6KaCoUdizAU5U4UNuqCbyDwt+2Mr27JTDYzwE
xPIhcOAdAGZlA4VitM3yx7c3H3eD7ySfGEABQn3B93nv4f4thQx+PFFZHwYmtJO7zs3b6mufByQe
SLnYB8Mwap6uR97AjPJTEUL7rdUgENBcPubRlZKtckBr0pSm5sNrhcTanpBoWwV0tV/Ibtgf6R2p
PCi+PBxwnSVTc+PBLc7S6MYwfvtPqWzwnxK8IhybL8vgwbatkffTakl9yYEpO3le2U7KQI3PFjED
tIwFpiP1g29lNZJU81ekMzDo4uDdOTPgUIQMMy1q6p/Snsl3Z9jf/LcEFxwTp3kPoXmX2bWJeJPQ
rLtW+FlFZBE9YJJ0wueexJn5jyOsNgpNWXYvoukThEva55G0+1xNqFolz8RgCm78lXVrCQkc+TmE
OKe7JEAp47TwF6nMRcVPrXnfGL2m3c2LCCtZLHjPXDmXdvZv0oJM3mRExpaUjWfAMvKCi+bj3xST
5nokknUs7UwMkKU6zGCyWuHybw+TeB9mhFH0JuBKMrwGwXY5MgKQQ2K1o3KSlIXzI2nurWoKj925
n4ah8C9ttvLFwDyGW9UFClq11x61hk9fUcfSfJmEL308fwidDUA+GXdiE0ieEUMW5ZAtW6LX8PFd
YqC931BEy3ZiyIG6gYSCD7HFPfonZYC0G82TXpRC2r4fO87wPLAqEA0uG+6ohOfEnO7oyXhhIXe4
2pQ4boCf0DnISOwEl3lcqx0qMg0SYfmVXGLmJD1v7wF/QWYYL2KhntWn+kcglE6dUqVAcGnK+vBD
mBU6sHLWbKZ1OVzkRDChQDnuHfo1lVr6xqEJZbQcAS4M9Yux9egRK5Xi6/i1l4OdpOcTOkAAjU2W
Dcwhqf+nLvYkAXPzNq/NfQs2u/ozf1hCodX/4LzVy2xtjz5MIKdKW6yht9TaLm9/Mutot3Pq2oyM
nOMKUSml4DD35tcf9W3/BcRIlSK0xIUuVuuu9iaRgSctheDmJu058b369/qfVtjSRpZ4SCrplmKz
9XbxFqsIh9nbiAndcGnbqyIgC0+ZNJX43hfFIwMNirtId/tqQu8iJS4mRcgI75DH3GWV0MJE4rtU
4k7C/skPRFyEnbceGUEinHV7d+Veq7qffIBEXuPViWVLTCVixiJntRkxDFx7cQna0PW17vPzgqk2
9ZNqvJ+hQA89Slks7Ud5PgUhGFhPiqLUL3PudKyiUimVZtYc4ZJ315vXGXe+s8tbVyiYPWE5ThFY
dp/2WMsea9OVWldbldyN2tKWv08kxzXus0yvsa5ak9BWpxXZbq4wSfaPLnu5zq914e6LLAkbGnvR
lQr81UsuPT4y63HK3QNMtNazQSAyUlTsPvCiTkjaB+ytJPd4MyBvJVwQbF9U505zJoeArCu41yt/
Tlfff4oPUIWx64wmSnhPVItgrAgP5iKeqrPe+vN32YMedNwOOHmjgnv6F8hzzmA6Mr9KQwiM+KhX
HKF/EYxRK4fftG/TQfWRXIEMX/dEObjFqDWJ9KZYKQNZuBddhAetU5rbVba2MArSDusQgpqMzz19
4fJOjo5OThGlaKl/3ZqMIZRlagGMmAe0BpiTWNYJK8uaYdKdN0AtAcib1UzQau7riGTEP9Sf3PTj
1wMBcS5lwb2IN1SeWecddcdJO/niwcJrb/WWeSuCK1h3vXHG+2OnlJRYjIu3rSucYMXeltyUANf3
gWHg445V1EnsBXPtRrQOoI2Mg2iLfHbc2aF+8f+vGEnq3Fi42+wPsFSeayDLjGLr/b+EqXkomGfD
FmCufCW1ScmlyUEhg9aRu1bALJJMBscgfgdoU0jfvcKXsKDggk8TPdxi8I0JiJ1Wed1bEfjWvEO9
a01U82I04GdjT+fh+208THgkmSLzKSMHB5uCc8CcZJl2bx6naUKrY5AdniYQmXHYM2MzUNvoU44g
tGBG48+5xtTlkUvK+VfvwLkgGqBTKWGp5lhpZFfxfhOjtKmM42ZP+miBGwQGM7uOUQj/njWVhCzg
5bhvuvwA9fYAJwo7n4TX28BRmbOQhlBwj6hYyQ1VQNCCyaTz2BiutnlM7u6niOWORJvTVTQmgaXR
eGNzn+jJxTAPD1FoQKj+dCP6xFmS/Gx5YrOMVz9BdleRzIc095AmFuCZQSaNY8AVF5ERsGjt9dq6
KLaSfUC4sAUZmf5jpGP/J0dHPnBMQwIyDAZzTeoAkfzRNosX4cDItKiVCSawDS4o0kFPyNWfH+Sq
wVW/KO6zjpn9SqQWKVlEASFo3YiNLNPFRC81w6e/MAPUoKDjf94AOiemUXNtpkyTNwE7W26nxigA
ddh9wErjdbT1Foptah8lJZ1rzu2UXb1JEZAacqdWWxNLrFfPgDYHTTgE0rzsallJ0f+dy8KatFJ2
26Ut7m05OBnA11wjGcJw4+ENI3L9LCKlXGF/u+SR1hX7lslmbA0JWgpJMEpj2UYHdw+CLVP/tFqr
wFs8g/3xfWh/Tc/nudFSoc641KHmkMyvVnOeSz1KYE55Hz5+1C1NUHsAfGZO+DRUPoCKc1TJ+k0L
dKfsZUHhbBDiDhLKf/1ANDauoX8YQ380RPoUTiwUZj+ySnF16c3acqW+Rmpw2xP4/RuWHQKPx0SP
QwOKRJs54DzbNcEvxYPijlfW50r9QMVwYqeV/IYVyGBI8dp3yp4ZxSSQau4dcEIbyJr2BDyHq8yJ
G7rmorwN2MK9ICB0TcgZ7qEMxZZfBQeTAp1sAhjFWSqpSlLjC46f/naayuJHNR71E5Nst8eoNXTY
9OdT7P8afLqCcDIN0r9FPn1n9jtMtp7iCOLNzMtOkPw1vLMKbjevngQF18ZezpU8xxhsAo/aAq+W
XRVGKL2s8ScdoQ1PcD/8CNXjHf1vjCa/jo2nROSgsPGfvC3zD5L4Iy6Sfus5BQDHGSgVCuDKMOMh
Sj6+XtnGyPNIEw4787SB8V73+9582iuJE24Hgc0HVzMS2vJ8neC+6gsA7OIz3sUuUxFDVN3bQVY7
QxI7B1Z2WYG6aKC5hGdRT0y8PCStc3cpN6RyG2+Zy2NAufSb/XSpDyAGHa3ZhsZwfUw4soMfIBdh
u3xdkZZxJ3OLHX4O2XQFMapJqKBfiVXwe/Odj9sIFYWpghgVTqbZaB4MadxtXAGfkBFG7V5vluJh
0v60+/+O8ciPxyA0r0YQBd3vo8CKpGUnTzZbWqvhLIKJ3PnywZKjjZXp4og9wpjJsBswvSnZPPyi
DjfQjTdeBmLJUaKsg5mTSNJVeNw5nDeqI1ajGPlXDdyDdnWofIhvIKNxCuvB0aQLkP2tEgy+1ktH
+HWGJsPMGaVaDrqcLb+nItkstOdy9cO56pPOOhefR/9f7GGu/m2+0ZLYV9kbhrwgaJuBpGSdzLLs
17cjIL0KaV5CVomN5UitkXPSJgudwNJff+IAgtezllQ5X3zbsyQJjsWgQQo/mbyRbnhQ6jro1AgE
3xgsq7syPtpPMK59AQnna2Uuto2jMYvc7GnCigY6IUi4y23su7vwwDxJo8PLFjH/O9fZ7T/54bHK
QYP3gGFvGu5RQfoaxMLbkL8cOSPVO8x+c62UYJRYxDtL1Sl8MMn/YYAFujUeDJ/vbZx4L+wcWKav
adeheoffPXnPQxZO0Rql9d1bozMzzNaTwxl9chIoxCaHxX4gSh6iQ4nStRrviyGQ+rWIIEAtSuI9
vdFKrgev6sAVnltqoHZEt4lVZgGa/irnw8d4EsQ/kkRM/2SbjSFgeT+m9BD9Xl79urWpfiG9keoR
RfldtJBoDTowH0BmxB4UVXULe4QRf014XTuZH54JIvvEItHHrXH6xkMoldiLjdhuFWjPuKOqpJtF
UbZgQ/3kliaLjxcaS2G0jGlYhSVWgWMFkQukPu4JFf1ndZLZppB208oaJkiIOWLiVZQDtG3xCLbq
lG39Da/cXW+dx+kwCKmqfrq0LgJ3x+4e111zkDA4V898V7JVIAOjgfHdjRgSBdDI+3cMtBDvt0eW
mdgP/SGUjtcpb95oGcIUZiStoauQtPCdfHovsH2MVEr5OvQr1rQzt7OYJ5tkG/8ajT7kakb5iZpy
5eRQ9BrkQRE66bdX4kad5jOqAIKDv0/7iopMql5cn18XRlK7CnXNo6pGXZmEipbKNiYt2B3qic9c
XX7T3g2QaC8ZzRG0fWT0QaPHjkTwD0G72KI1oyJqxxEvIoAultw4mEPUPkB5rTKSIWDMtWJz5JyW
+j7AW63jY9GvztbbW+nlj13MB2mpi9HL/cVwn1OXQWMWr6CD+XbCWwUZzDe06cdHs2wbBKimmf1T
1nzopjRMk+wJy+DLMOFopzmEUCSGPHSf8JGvoaJFFKG4hKuKCDz/bRT3M05K46xT3ck/r6vDEAiI
7HNbNf2WUSEok2zxl4y3EqegVWOKOPI9g1tG3M2Clm/E8nyChaUMhL3JtYsrpUiP2zfMTNL9jrWl
GZep5ZoJV/XKbPxWD0+xqQK8H5Oun91FKYZ2wL3fEwStfM4/+J7eJ7v+N1k52zm47/VKe3t9btFS
bQ1zQ9RooLeXN4OvtD0aSxvScoBW+MYyn7pLoG2f5dT6GzvmJWvBVJLCRLeDgJTAjdT2etiaBtXu
ZcrKYf6K34SnRuyh4ecqeKGSKhSdneA64cxI0xuB1ONixDXBxGdXApff6bLiKmEm6O8uhLV5VpKN
UK+288N5Nj+a11U1Vh9/dwplNMZjfb1UITlDYp89bUWutX8EzKaEkRKszK3q5tkU/6KZcl24daPY
xyeYXsqIw3yai2oP5ZySGGANo+AXeHzxteWebakVEbkiqur32ZvWcT3atM6mHrSfuETJ4D3xbOpr
5QPQ7LTrAw1kGZz4pDJE1mqpJT+ljBbixnOmJ+RFEHxQFGh+QVLsyPm39hHKk/zFyU9jSQhd5JJt
/gHQOVmz5MEhDnhgLpnVxGWIiO5Bf+sSUyJ5NmljzV9jj654w+o4jgsYxDAQOCyMK55GZYGxkdGt
U+lrd7JqwS4/1cgmzsWI3tpA+tDp8/cAGXGPtf28aOw/iygAImM63hvVcT9A5orChHzNkjsc48pR
an5fZTYpnuyKerLnmuNP9nKaxf2h/PvJzRc3Lf0qAnT6o9ds0z+fRusXh9wPxQaZ3KES+5rEeQs3
+rlfv9itKn81ebH1aPuBJh+lexPhfFbgdCkyd7CEAERGcxG3b2UrAXPY8ons3dd2GSe6and33+QG
/TaLFfwKK+xkkm4loyFkA1hP9cVhS30HeK56KmnTEUxK351f/uYkgHieWYPDBY75nSWlhYVItn5S
SHBK41xSJM4SzIE3nglypITwd1v0SgRU9wRKHRNXwNxtzr3FIArLQcSK8FkFbD4Orq4SmEHotzmh
Z1OCV8vRRm3cEDCUg1SBEg+nFFxhVqwjmz2O7UoYn1a2nc2yIox0EEgvDKctoc5mTVggNCNvnied
fTo4TEm+i6tg79IMcHD/gdkz12PBIna0ybquIZDYaSwl+O1BaSge8P8xzUT4f3T+q865rC4GoNQX
42Y5JS9jQoYB4uQ9lp36OB0P7DTiuomkAVxe31PBEJa3gOihtwf2zqjAsQKzq7ydB5mO6DXU/huq
RVIqSddRfZl8nm4tFipl0E67f2Hz2T25jomEjcZujA5kNOJZEGWegsW8vHXZ9FN3Qvu2jtvmoE9Y
qZw80iKBYSiouFeFfnzESGGCZ4hDdbwkrTgo058OzouIxcoxDKtuZ/fbg2yhuN1A05NWKrKuJQ+W
jEeP8casTftOJzYDm8JfXRLs5SGMzWweHxlAQIivhX2uexGAYCTq2Rcd+fCuBO/SSx4wgH+CjFv7
g2Fy0+YKDHO2tH+JI5pjVrz99VdBoIetbDrPJ95vhJy/iDzwm7lr5c3WA2zvzPVyqsXncgDVRwbK
VVLEbPns6JUtgdZAHnSSIAMClp5GAMSa32FvWRHGzOcivrMYjPkxK+a6YaeLd9x/gKnJ2/AYDNbh
w9OsR7bBDi5l8jRH+YelyLmGIVGLgzSvqz/GbMecK8wK6sRmJmQw4qqLooBW7wkXoAtoXL3tmZlb
JHMCVx5aOIxOlNqzcSHz1XXDnSKZoLmC/228bGSvY0bg174EfVKcsCsite0mrnm7HwGgZQ5aZmED
hYSBRxCw5Ypi7IWw4ppDT4AVmKyjzS7PmsR++w2RrkQvsMoFujM12WyLHfOcrfylY7ZeyZeDCH8t
kUWPRiWbHkv7Ra0UEe0va02JqMD+Ut1BbF2TkwbvzNJXQAab4iome7DwOrhImaacjRIlWhay8G3j
DrvxPPWPxOdekK7YXX2is2S8Uc9yztbe8SJD1sZVoqVhYcL0K+AtsBL4ogm/PAN+fmwFkNxHj4g3
FUBrviXgAmD6TtLP2OhBO6DqElz9c193K+8H9+DGvPapvqw85cLjsKlGOrnn51Br/PfBWZfBj8CH
8CCzZ651a4Kg3os/cPIOGRWZPepxNJHdxhd6LKmumiTkcS7ZWbqI+JDo9qqypQ1Li9A1rmiW1vxW
Ltz4RLwVA3jmCqAx5vRkx+V4N0nszW5nig8w/sdr4XR7xLe3yVWLqDHRIJgvBSuCMBxVngzNlYQo
vlpZYDqh7HV+f2clrLVeZ+jRAVih0m9ualWOdpt9MGmQJNhkh0Wv+zccBs4s1emYXxbjsXKpAZVd
u2WHYBjAS2pFsmiapcQN3bY8QmiaKXfCyu9NWdUD2zNaqv/Nxd3E+S0r2GESQ/x9fuOd8vFpKAzs
yArZ2QzvWt82wlxZPhzxW7uwCcy8hDWNJOBLK0zDD62ratvAnVoVmAOf5JOZoxZCplbUFF0yRJkH
649INwAxAaLRegh8Z7Iye6py6bEsZyU7aBynPFgLCZH3H9e6uHxhu4BT8L3nf/AlIlh0JKhg9SlK
KLR+S8aKboVLKcGNYOh3qI2c7q4Nx1AVXFaHd0yn1uQUkUecZeZ204ueY5n4oHd6VLxJgYA7nhBe
n4UMzVJQ+ZFOD/y4aZdfbIwlRJZtfZaSwP3lSmXNIirj2t0oz/SZQPM8ZqCRIBOXtRpuwpUr4zar
WT4RbM6JkEiPuntG/HdGwTbWM6o+vgXAjDDEb/fIyFQwPvM8hzYRD6rAVun3uHBHnS73AbDG/0OQ
3pqdxOnwtqhZFLfk1x/CUJ95a8/S4SJ3/ex8EtK3xXv9PJgBroEXQ+FKjVATcV6XwlMmfxLbqsth
UDWP5Dp90Wk4etoOZgHQUu9g7LL/bMhx+1BibT1DyNs6NIjc89DUFGAH1O/rtVa+1fjFNVd+2z31
89hyqlG9+zeAuxc+k1KNsLNIZNYtPSWfl/XFSQMgrmq21+yEFn619+cp5Cw6pGOeB7K3HT04p+Er
+5Cc+qFyIs/hWs2+qUqv9YYJBTtTFX1rUZUwZq0P8PyQZPMXcNXm19EmYKE40n+EGrlBOOTj/3nB
VAOxpSpo00JNDCoszDlzgHtdFkiFwsjNAAHFCs6yxlrfvtAMYZwg0/5GM2e2m2LVOSIFZDKTMmp+
4nIchJmOTXsZUb7ZsBQy6gE3dyTIETjrKvrAfAb/XYMSFSKkEP2BSsr2T+CO/NWAjUfjaMhh/ZYZ
8wjeNmNLjy2DqRuKdWUNyCya0Wt9NwhzLSprT0FRk5hOAVB88YdrLsDbt5W7+erpPAYUghwDo1eI
1IlYhV2gjibFX6Mvmm0BL4tpDmVthJcWANYtTdSKcr+WxgVPh81+1S3TFpuCcaeZqoDVvgavAwBt
Iwhgva639xsen1+/bJ7/oPye8yZrbP9CzxKSRICodjfgon10lVFrxKI2R3wnsOedwwhZjX611f8b
0klqntOIFhtDbT9gozYQE122GBGnxoAJYoVYIkgsbyoSd9qQKFwD+XLoRnqr9shtU3BPYOgkaynO
BYaCqCscmcsDULLH/iy4k/x6o6Z/IRsXKMXU9xWuipHbl52tUMR4tchZjVcH2oW8hVOnD3WhIeaw
iZrOTsqHSgGWr3QhpJqT12z2+8eUw+nr0AES0133ytAgyaIq83XlEOrRpcq22MplHe+IvQKHrk/0
b0ckF7avO9nd4fyz3iESiQKeyN2EES9yaluTjYOROyNQ2Y8cu4dA6/T23jm1IrzZWRYwHAGXwHrL
+S1+1d50tCkTCETzh/wx49ZlPr+euhikUEEZCSBpyBMimmP/rA4yNF+EVCh5lu8qySgyZQFVO0bP
ffD9BRTE4SmbK3zdtLuHgOoYoG6uHNuVEGbmT2dsINN7tDDW6/Pbodu4Atcn4KnZK8pELhwXMbXy
BvOj29oolKqoIaRtf9gzh+Fp+fsN9iBZhBqNAydeXe+R4vqgwrpGHUhTO/rQ9jumlvHbKhKfkyNQ
JdnVgUXOGTsf0AVQZY20D/3A4MgFSslCbDOgFQ48GYI7sSEtru8Iw3d6bhkR0S/LeTv3T8Z04XXp
8jJxniw9fkfHDX2Dgu/GkMADa+cjKPEVLap/beJYluJB40mGz7Uvp+hDX2h1Jv6rXD9J/WyyjlX7
Q/BFeTjwo9HdyGxFI2fOHp/+HGmPvzZiP3GEBqsbXPINGDyGY5N6CtTDJ3lHRAV7zuCrRqTB8fp0
BGoVVs0cjGcxy+z6BNAo0AYTzaP5wxlXfA3UbGlbuSv1rFQWYkMjBbOqFCIvHQdrZB/f3xn9uf2G
3JoUJn7o3wS4Gibe9o9zBab0V3UJu9WTPF/141RkOmY0NGD3Rna1NHMJkTdzU7rU1D+jVjinNv5A
8bvNLiDDLO+vJ/MRvYmZlZr5U0aqUgoBUPJTXmJmLbZ7uVLmp5H9b0oTbH8z2A2xRwmxaXaVxk9j
xrS0BeTd98Le0f6ZmW5k51CVPmORPj/1rgpSgzvpBVFL9FSkIZO3Qhdy1F82cEgddBj+M+t0G2SO
6ClwGzuQKl9jGyKrxUM9+N2Wa9htpTVyNzVagLAYkQQHdUdOan/o5wo4+U9Rf/xAVoV3G4faqR/M
Yg8wLSIfuviUUBE20IfDuZoPDt/XjtiSrWcuSPNdrq4LFIlaswv0o5nJbA5EfHGwfEuXy8e+zpKC
U5LNSVzajnY+JLXzcvvh8O6QrWjd3JUNEFoouQ6jlLGkRkWdCTAA/b+Hjgk9ugOcz7pitGnVnv3O
dmzeTKDZB9BOkBffrjYVnggpVgFA18efPzIHk2oOC48r1S+M+3oZOgF59kNDnDCTRBuPGwjbeOvk
8Y/deqi6/dqQlES055O4XMwvkTjM+zHY1BahEzm59xftY+BSAtFjAQnm3TyCM7puWoyj3i77mciN
JnPr/YN4rleIQciP+Ou2BdZZLyxTn01eCNrpiMB+yratc5uqkxN2f3u3ZTDN1MQ2nlzVaXDuqrMq
fjdMSijavAz653eJfKWi360YFZtkomUWBUFRAYtdqS5guum9VsGtZOnQ7vYyyg9rITTG1b/Rf+IQ
RIxTpv0fJE8Knd6rIszWkRk+nKgPGeFVWfgSv/6rdJIqJAIx/fXkhDum2DWDQEE/eMz3o2Eya1/I
LZBn8TSAw6raXOoJCBVVwUo7haDBfPU5InjAu/4yRzk+iRWgETaghwbGtSKnOlPLOSkMpPn+qwVh
9U/poL3ZU9UZ7aBAmYkToCI1tEAG/jQMz0CHy1JNSn0SvmqB9O/BdOUUdzXaIVJmXH1RyBFZjIl6
9wdAewEIYBYr3XuRqOC6S4b4BdgcBcjPSBYXuWPm1rcegjr+Qwh8E5Whw493DK0FI9KEqsrUsiEO
jfZ2abiAzuaPcEwp+EFPo6BGRk5zFt4BUsAO/PfryXJRbJXUxZ+ftTCi/oDxhd1o6mOTI3KjBoDf
zBzqHhpGprXDeZN0pvChd7443kJV/ntgca1i29epnhUJndioK6jwzsBFxbqT4fL9b5qK20f1Fvs0
Uai+DU8Je6h/vh7/jmif3pdIZz58J1MpC7TnMoeJrRDm1gR5ZP+CKdKYiCCyz+5FXpOt6z/9ZUvG
+AXsyb4yB+GXaoxseolQIZEfujME2bFb0wcZoHTIfKYvbNUKzvYYP+yrIRTS5ol3Twe+VENEN47z
vPvxd171nWJFyV9a5fYl0i50aGOtTf3wHLxBrMCZufbnPZSTYCbv2PQ4Fum+wcaxcOiCEvpiczO9
9cSVR6sXlHndCWrKaO+iT8As9lUiUmJPhvjyIssl/1WM4dsCXB2ymvoydRK7Utqig0D8Glh/2+CC
hjAZD3D1qtv32Y2G4Que9dRs4kc8yOhb9NjmudFEuGFKpzLj4Hnyh6Aj+H4P9s0HEwmfHM5H1HJa
+HnAHxxhkFzbm+zSDllQzQKgtcP2wR8+ZzSttmwW9pFrWKfeAeZDpLtGZsLAgLDQ0sBMbV44lwcB
H2yuU0/hz4bjMc9RAycOyfSYVrwrh7hqeV0xY4iHxMF4WNlZ8RnvqiSaBBkJp25TwRYKOkuf/Axp
iEIaoVwC17niLKL/CFVhfr6gRtOEUojwkmSgDDfm8YoEO98SQPPvDcLTsVe36RC+E/oElrqMdSbT
qwEfUOrMVnXP2yDtZy9rW8KfEj9lSLEre6ExEOHN22korCjUW7fE2Uruqb93kM/d6MfzJmBsriIv
QvrqdvPZ3BG8IpjPxzFZJsb1Y6BiAxiFmceaj58K3Wbr5Lzb2mh20ew3cynTA9CaZFszHZW8FHfQ
PGUGNgFhhHhRZWfFr5nRs8MdcHgZDEl0rGkAnJ5jwCSWN2iC8qWenH8+DhrrjVVEks85uZoCdF/l
pmXTL4A/k37jl8GQZAofhkOjzZTy04kSFjVNPaREW2iHXcId0CZysLPAZlFSipa+tF1f8bR8aEf4
20/kEi7A+caDYNe46bDfyqs4HratQfK0u2dJ9A/TtamTBCB5li5n5gxVhYDyLnOyTY2kI4NEzM44
vTV6rDOW2NKaenNSSt9nukI2QhAtXn19VKKl3SWMGqliKYbyo7unSCjLSPQ6fMqTgs0GXmV7HygH
pKAK+0C1ycCh4kx4lxSSyySGAL31SPTIv3CqbSy9wkyL+2WazFftUqfczYYv8na8WvXDQ/sc8gkU
1W6+f2QP7N8C+bboDWjEnU6BbBUp2OTiGXJKvoLb0o2vHZFMEDGQe9m2//p+TFqBV4O7aeL0M77y
zR/eas+u0xRO3Rbz0IPc6Im+8rU7aKwxNkZZj0o2t9VuNXwdEy3p5IRVosyAbmyAUT6+3Or1FG/T
f4qXsuLFfGRKr2rIEq6c5Fv7e45n8M/Wh3aUuw1ZNHOyId0/aadIA+feRkIicpMNaOqjlLBsKjzH
G7+g0NZvSrQjz4VbtwZz/7vl1kAPn6jIUHAg/oCywiX3Bwe9S8YnTxYfndJ1ZgS7xRVjEfq75tIA
zMWJQVlEk/xXZtbmsIrGXbH3/2PjM9pxpbraNYXcbzyWH9Ojf1jhmdXl0nIZKCfQSRwo/GQ5DaQJ
5QJCSM0g43Dn2Pkdvu2X13FXvueHpEZEK+KyxYJtZu7i0AIf9NLbEyY5YxfsGgQhBgv+eLpvNNFx
RyA0Xk5h8eLcTm1cQHqiYwggS2N1+SnjwjBvlZt6BQlmnuDvfbjlmTLbGzHCoO9JMFjgbQdyfYWv
B9Zw27XHLQsQzpOapk7KhORRvLSvjH8JqNhQ8J/6tiQfmzUkrbL/OtPeS2A9FdOQFkPkwrbJE+oi
22e9H/jlPzkXbPPWTMpHE5FOABFRdqW7DOTHi0TXPIZJjarj7HDSltpcp/FDukQ9f2HI3vfYHITV
wsa2JqVT8WH2WqbuHK/kuX+dG2aG5yYzw3anXQcvVjDAJLBJukUf828aAG9hi5LOrkX/gjTlxZkn
oM7vb3kxriJsinPKcXvdbL5mfrtLYroTYuMXT0yzSic3GWnqxqXMay0e6yhHn+unyMz0EoKvoLfA
JWi3+c/0c5WVUSUMR4FbmwixomgVkzySHhR/1j4QkgDlt/JDuQfDhRxZ/jKr5Aven8Tnh0D8JDsc
BbxrBBBA7TDCrf/NILLU1IpM2OdRuS3baZ+WWCjhIKNhp0WInNcXE5TpSpxzl0X5ms7MdnSQAp51
B4AVEFlmjKPiW/I7QJ6XDn2w3tRWowXInRV5OxpTZFUfxvobrg9LifhhHaO2MxJzAfmZN/yeN19p
bOqP1eteU011MOclanCDpVBjVk5xNL0D62o8CttkhA4L/3RcP8tIejwe6Eh9wnRCdhJ4bobZScDs
y53fSWpsLClklXqDVznU/YOGVYfZ0jceXd8EEvXa2Hunlxw2OB8euwaByGK4abV40g/Z/LNDHkfz
0XqyuEYQKm2vT12gAqx2TkmqWDRKJpNP/xLtt1mlsYl8mB9gl7WPFw6cmH0N11mtE9x8ZjICtenv
buVT21XpwblWpCdjMt4eUcYORoeuUvguOVjRG7jf/witGACyTAYrpTHE2efLC8jIwOFdU05JqYLf
cHfJBYmw0P9pHel2cBTo0SfF2uJqeNso5E7OrcR2y7Yvf7HH3J8bfYFpE8Zrs+JQtnqsAWWPgLiF
qjVoItjHBtaz9PC466+KT47M9O/iEplkBn3Zh3GQs5shMdK0dU7zKIxc1Phv6et0+1QinsbEyVAe
+p6tpC8FkiDa/gmLq0DBJ/jsyJ3KkCRwAu4oPQh79xij4fUBD166RprN17zRE6CNgUE3i0R7QOVx
VCSKyemQMGv7l8lVzM09t3YUfgmuSW5063OqvdfdtCOEoZ7eQogoVEgIDdVxNJfDZXxvJRc54dS5
hgUww/gPAf5bV52MkG3X9lwgjlAUdFpDz3KUpGOsogasJBKgIWsYMRbLACZcezjlvwx608yamD3p
xDt4gwjluoPcwDDuGxPTGgi0thGhlqvBf8T6gyMjSvDC2S56wSHKX/ZN2rDCg+KycmgcOjSlHMkx
cJzmRMqm7W0LfGj2vXgLqdkYd/fYoJ685XGFs4aFdzZP9Hja2oOswYrkkIbFc/bNcbkZktBfRkXx
erF5Gfmf+ycbjJunxwiwc36jrvboZfkmWuVKcu9VfuuCRoRiexi8X8LX68KAPQmcOpHZLII/3Bl/
BbKx94MA+UMvx2mefyPtwsLcrgwniV0qZkekcUhj6qiAQWtdwtB2p0tlBy4PgkO0uCihUmjK4ygA
piB0tCInapBBrCQjBJY/Ilb4PiYxI6wKM5cIm3bzYkQxwOwr3DPFv8Gzj8fskhCQE9xek/uVHnUF
CePMzeFtK7rmLWxDluWCmNu0Qfed0Nx7B7S0sb4LXdMTzmLaLK9dkNfd1wDWhoFxNqHCbQwp7Dns
hu1rxUq+Ng0tlreQ54z61gOhfW8+bPf33s8C0cHLXx2K+pfmwhp0JJIRY5Dw8Xa17D4fH5vfQU2A
CIi9c+BUTjGxxSKOhrczkkaJdmxrMRJqP7TQpSjXLSl1pPnU5hj3grFPuXyVjEqjo+Vj66jK8qvd
ap2WX0g1aEQPa7OgyLRagYlclIPfBgVqozrdmH+WDUlorMBA2/HCXzsHaIc5CH6UbxXT8/gGchrt
1P55TR9Nx3sSPLJa7oCPrhKA1c0BZWE98WDxRQWTO1Jf8kCCiYO+dS4gnw+cI8AnO55pGiqdgTSY
DZLh0CZYyA8it4BYqzsGkd1/qEBzMyiLVy7l1MLD1iHAFilQNm2oLSgsDgZtLb+xXQkq9TpweOrI
sCOmTS9zpUdGjTA/1YMyBxT/TJQVWI4E7DdcAqPcxbxVkAjhI+a0piAai1y0Bs1g3QW76u/KczaP
K8FRnNqLNKND2WqHmfo5OzwI0rPoPpvxObG9xg8iFhGWvr2eF6gSzWjeDJXQUtd4FxHAZ5wrG6md
rYJJ0f8A4cGTS/TD2I1nzra6JHFuEuVRIkrKim+ADuy311q39sBoi9Dfmhk+BjxzXT8SLlyb4cR2
LbScozoMu03ClaUKE7DGpILpLSn8URPEbiSEmwf+GsLk41QIdhm10jG/jHX4MgTWxUqaOecLY+oE
8Abc6Ov2trkK1tnrsYxY90U8MPzLVG1+hYiZ3O6MY1rSagesI6b0/DbYKBJ6QGdO7Uq73dOj+Rwm
QCj87BecEvO0YPjHNl1BxMogjYIZzGlLvlmeXfVcyUOPArvVUg9OKyIMBuSahgY7x7abltKi6hS5
90LrGs9yq189Jrjhh8dI+r5Am7TyY+6mm/T9+ZCW7MhoD5idSE4lzFKcPVtKBSLsy1LY2zifDdEL
j7YV8bmUzPJyYGok0OGPtbDBY8yBRU8uIp/jWSKu6AJ2kDpY7Lq6rpYhr6y4y8mNv1fRELsP7LSb
Qm2/QdVtR68VjybDB+p1qtlLQ1OosvXLfcddrBq4IEGzPZVt0Kxhd3N8bg5Z3qxL/qfabDfAi+tY
S9sjjKUb//7C8BZzoIdBpXuXSMEE0CPBcoF20MvZl3p34AusrKY1V6F+MchXlhWfK9zLvJQS4seE
4V9DCHUGPaS8Oz23qTkUCEFqbN//BdizcbXYkdOrM/DV9XBFKB7lie1+k++0EitINGijD5XQwm8U
aERebzvO1BRsBQ5+J56V0/kSyuTFJFOz1xRiPhJCNF2SQdHdwYygkWvlsiHw6h5ZaPQTuOMJxO1K
Q050XwcWiEI3ycllEJ8vBKbT/IdCge4/PBfS57tLd6SYyZR3vDXdDhBE1RRAGB6aZ9jVb7v7s/Ty
6f3DyipNWnJ6G/2+wsOjFKGbM1EawxgvZqtYAAGmNQj8ZOlhnHoCSrDC6f4aIllcQq3dhA8vBEYQ
6F72DTt6IrNulmVrbhd2Oa00VqEXotN5grKc12AoUbY2aZz79wSr5N2G87ptiiEru0i1N2lvW/G2
2CbK+JOsz0Jx/knqnIiaX57ONLq9bi+v2LBS3U4QgjgB+zRDV+WHhzqO/rXjyGAOTfVLDlKgl1Fj
A6QlOjKyfZokiA14g0Xiz8EuqfL/ZkYp0wqYrb86buepJUFg9Htm4HwsMT3/hVKGuASZxAsAtMwO
d/GbYdJyxNiDCjHCIwAWR4gbiMM/zaK4tJTJmfiW7FPOYQCHSOTuDO1xqnyifT0Dd/so97e1EfyM
U9BKIwnQdRcIA5+ZvbWJXXiYn0Vb7Fhst/HL/gmy+bDjlMKDsnbMXwvtDNNxNejpzyO8/fRt4xR5
k9jY82oj8MxzWUOYyfHq99WjT/A+X8jPneKZ9h/XMexFP3rWnUdr4BxK03CjnkhPj3uAumlZ0JEa
78l+c4NzRLFKgefILhapeLaR4MjEsRLP8OxhYUtdgcfP63QttSe8JFcfKKFhi3F6sBSm8+o2rSG/
aNw/XC22ZbrhUCI7VLEMwOv1ucBVn/OHxsImJeptqUWNg+mywDfCq+Kf3LEXSjRnF4dgc9RiMUFo
pubM321bhwU05yHs+RG41X7M05sh7Ih/m3MpBNtH5sWG6+8sgp5pRf8T5g3e+t6ZHktThv0WiR3r
qACo0dD8ZFEYiU7PllwzJnp+7Sys9D+KB9UbkZ7/dlkwo3bTw1KQ8Hm+tOONzzpP9sPn46l118Ae
qM2wiUJOc7BW0dwqAW2cfLQY9/uaamRv9EVM3bF+2aDnUVdEgA3uIwoxTxRwf7I5XegcsvpfNGPg
4aPfc3CB1urdbBOVFpuCUHVeLkOjoRu6WB05hDPjxC3fOJ0L/7tzy7erZ7u5WpAjGopRDSVncwcC
f5dSfP72T3dYZQhiugKRO7IUfFAy+MdVBknuAbPE+MQ1dzrDvP3tJE378U9QeqSwqXYq2P1lHOqG
A4wG143rptfapuMzS8Kckvvdw/PCeQqAgj5PjAax5+r+/BLLHfGwBidv6VM+HbupsANBYWJKzFA1
55W2QLwjiDFTu3Ii4wuqxm8Sjkp3GAHRGVlIDOInVAwiOnXJFyoT/26buMtiEBRwpWer4Pxx1bd5
JV9/qqsVj0UiAm47Vd/upyPyPoTpGegNeXIxpbwyUljGzUoo48h75rVhkRRhecrbLI/nTkjPbmIs
NrwuSblBhCPFE+p86Er0d/lpCvMVLaeQUQzI+mtQulSvEjgvFNP6f1Pqd7cL5+HiWRlLwf2qiqrd
2VActodt79JxB0pNs56QAeVcxlCj+7XkcCPnBd0SlhA+nRw7nI9gUhVI3mIeUbuKgjiOymevwJVe
8sb3W7YAMvzOQJdAhhhCKVNZWC6NYTLQRJxC1Q7gVViZOmK1IwkY7vxaCsnWTzVgDbcKu7+5ZWXd
eDHr6rX5jQ6xo2Npu+YXs43i13JXYMijMCpue1A5UGsfcWb4vcY3MzS5D4ivU672Y3OPmZYB8Lbq
XKrVXlG2rzXlhzv55jtHB5LScs2J6BZh0zMJ3o+ymo1EpLesJL87yArp+2JLMFMu33eeJYzDZeo0
Cml4d81Kc7wlHt7TMMAKLxdFgPGUpjgObB5i3T14eSCiJrJ7if60SRAVDPevrjX98wz9ArFQ322V
RS4PynSTggIe3aZBYA3avF7F8Eqhj4iIq4GrdgyTE0G+Lrovu7xDmwlIPH9gQTUdF4mAnyk5Glgp
ZkiC0yJgNqveUydpRvlLV7jrq9pLbIjKviH2gVxayi2w+jVrSF3KxMw7Wd3s4K74axt3/sD0Hb69
moxmSphDbsQZUu0/oMlR2+lAE5bNY9WdGulm9iuwOMZS3zaDRW4y73QxBfFR+c9/3EN0iDD5mMdF
U+dbNnXf5ad4IEbLiAIrMsONhYIyF5yK93hy3m2L0HNoI4A3M6cpsxFYUetN2nnZM/d35RocNcWC
AbiMrrdDi6smgOkJOpw06Hu8JewYT5EIoiDcgKOcZc1U0P2E4B3DWRg1DgpQ4GZ0imMSztj3QeA8
4689INGGXZz/g4y3Wa8rPw1kZnDfqh35oA/ALl2tfmOsoJvyZjh3WQAaeuJA+1JzCkaE7KvNDrUc
5pSTHrfZXAiJvjut9iHvjTLHg8JeQEGIpFpdDNiq0XxO7ZxJUo4MW3X0GY0rw93EdqB0RampPHnm
WAFEiDsBFbDT0PXVVVGxSvmfnb3V+0tI5z8JmoUuarwkce8Jg7PRbUrbQeB5zLw6BcadD2JT2tEH
3IyqLADi3uTTEubVerUFXtRs3PBSnIczwwAy7xVTE4mvdFOPjJxZf1wbTf3AToX/sXTpkLcerGao
Ssj0dQ+6auTfXWeOZaL7RoPkpcN/NhJOCuyig7ryGpDqkNhgxbnl+jLZEkIsGj4NqRxnXM2Kmtx+
PIanlz7YAKMlr19vr4helPgjF3zwpRiqHo6BcGtGpv38NGTiTP/Oj5xdt9+Qajj6hBY3Pf6w6bFc
6E8IzDtLteayfLtp1aWlrY7evbXheBJFi/YcKlMw/uJVvS7QxIZzNWSUfweuB6kZhwsYZ4lMtIIx
x4+IHJ56YBaWxmmEJn9cNkHgH913a3H3nSa/zdpWBZw0f132t1/stZQabJT0Y9mQLh3d+nBvrKPA
ubyEdlrnsy/jwEy7vVooD/bQlDsMYZbJLbdR+7pb1bvgcz8uA5YjX3zvB5FovoMJLcYYkdBsBhJn
EFv2F8Dr+/9bbY+yCYh2xmwjBoj8CfDIOxX2cji0iw24pYCaPZFgmkxQXHFFCsSX1GRp9o9QF+oj
OwStQvjhHH7B7oaLJcifrrXceVlBsuhYrbKN0YlmAoCO4s+RrsnxSeM2703XccyiPbEQc7RgdaP2
3xOrtLtMu+DyqezHkMU73C+oJ0A7rl8Lg8zUy2zeIj+eWi9NLPT7YHLJbAz94LM9m1bUD4/3WXcJ
WU3J+s+UmYHZ82mfDFtwppU0xLiRT6izTJfHfboe4MnFSVA4h9D35E9ZZYpDwVScgU8pB3nMmwz9
We7ecnKyeYsXS585hQunhC8eVaIsrckL3pNfd/kjXp6A/YY7CEDGKrnc1iDw1rtx/3vtgfW5yXTK
uMw2uGJVm2ZJPvGnlv5N0DWdans+I/LwXJwWezWkg7fK9om7pmt/qfEUponFAFsVGE4boYOew59W
xNBvLIrUoZwymZWqrEsy/p0ZhzOzMm17IzzGw/x/bmNOvP9REgYcIhZtfh6b7+XZMyV3MNbXnwJm
Tb3GQtS+06NZi2+XzCPlElWhP/coXSl2OgR7pDzz+yPiXsdVnEdUQ2fPfhWtXrNMx3C+XdUdItqs
USha/n9ptW+3xKYLRiV+/gbn8ohxRQw2gZVE+kJgSHhOG7nEZKK0p3SOTUDsXVxGMbKPmCeCgs0d
9Az8XvqZh2ECota/Iq8SJUsyDnnh71PmPqB06GqD13Fyd6VNi/PAyWrc/H0pVu6Lfd2s7QLHGRws
cds5qVLFbpHrZVIo9FRHyUmP3RSfWrU0gwW879dcShswUIoq4zLCUqxyGrQSTV5bFP3tThB3Utv1
sXit55GQjl/LIPDck/8K/EPr9M3HF+LzN6naHf3SDWfFL6bj2HjfwqpPz9WZi+V0WnqDnQCwVoRt
Q0K3m4CNMOY26jOU9LtCUCPq4o6UpYf1S2g/C0M0rIlAZIUsGYw3oYF5GmJz13hHXpjjavY0FGbG
nch0IaRa9pLLcqya33/1RDkOc9XV+DbvpFS0GCjQvuv0atGj/YRgEWbtUlLba7uoOu2+zzoA04T5
cJ9ZGMSKAsdc3ZayAP/BzHrX2rZ1/hgwvvNUyf+2DjIlFVDWKkavnPv5hQrwM5dOVowGskKj4RZ1
/WQlKgXqJLHAbPHo7+CQZwyKmAEVgOZuK/4ch8nJRDJ3DClFWuqwmg5n9Dhx48vcoVF3/frpW4PX
PlpNCMaPUGWk+27No2d+AWQ2C9cpiD2mi5jzMj2H65/+vCtdC3kzyvYtUAm3ohXxpBVgqcs7UBF8
qSQbfCYiMjSNp9LAQ2xmTrYlAv0RjgqE/RAylFYCvyB57B6Y/AcUvDvkVCrw0qgchVLjFt+jEZVP
ODloqE6znxnNRSVHgUvOyemTxBz2BBSeIXAc7soJrenFcUo5Pmnx/LD1VJNuLobvPDQl9Qf6e/zy
RHdgUSUAGGfSdA9wjTjCxdBEctmuVKsnKTSRUkB5SBiKh0GyoNWHRC1wVLaFdoVuUrfSq9I96/xt
L4NyclrcmWvMMBV0jgmH1vMVTtNMiZberr4DNCiTcaYvF8S5crrqmSSAuuDbRIk6MDNXYqU8jVBk
pTr6KyTZruCstdlR3nKjbvTH6JObYv5ATVNq5Xf69w3d8PHmpbaaC0G5A70vgFaYVR5yR2Wc3iyN
CE7CgG6sFDWn7In1EnfwZzhDnr3PkLPqa18E12k6nwDQx5pwB9J2Tozm3Q15CcXxuLb8oKVI2nKm
GOVTMoemGAVm4kmr/wdSiytDv88kdxOSa6jChcTudYzTduUWbJeCqr94MhsbU7c5uC1oJRVl2lKU
OT8fAFILygQrbZOvxjKFNIizyB7l+lwXrOg9wSejT3BHRRF8Q3yadcJTlIkZwErt8oghNvSIompt
s1zJTKvM+JFi/hPIz0qOeqmrvyvpfBSgk6pZtnMruXtdlqVQ0vOfOag33JVy9OoKp+mMnL2waYaw
Mv78I368jhOkPBZyTWksVzeGUPsoBaw5+KNp91b+IW3E4BR2XNYRE3DwRPU6vZxjxarf73jAQyQO
Qt2hxyLcyyofASBCzavp1OLab/MJODYpwFr6s6WioYPA0NlR6SFXwHIplwGVsZOfSU3j9dC6C02t
SaAiXxEE2t4Ivd7PszAoK0anP1FPbMFFqNSKwM2w9iaNvU6ZZxUsuWUryl3l70SlSC+7yMtMEaM8
izrW3Nj3q6H6Q2ZEbVoKgoOpZ9HX5gmmah9THl0wGwQI1+rnPKKCwtcgQpAJSFRANakbYoiUY2q3
3SMVbKpWlJrqfoVBZyKXkinji2yYdOWtEF935o8TjRBsoX6xJ3tXuK4DgG8ws0fwqYWZo1d68uiN
b6QSsorPUlVn5kzM/hCAP7mSrDScKhJ/UlEwLoR2N3CtNx7VD4aBqYRJOukYkK9O3Z0G4swViJRP
exWa8+KOL8KZfxXe038a57Hwr0T5SBN/T0aATwjc1huOeeBWIbyw2N9cJBVdzVd8rbRpp47nQGA6
+iLr+RhWUYG/47sNBuhpWNgwbJXMucd7HB2XqREtoGhWS6ZlV9h7273Ge7IRnSH+JEABlXhhCUJ9
9KH94iJ/6IxKbgcVGFadc4WEA60uO8LPJ6n8Np6TIFA7ksZcyuv0X7oPCp6qXbz6yNv9s3pMq46c
JPYRBODUMwgx+ZcFfL3Ad9J1UqV7HW2ORwZ04gPx44ZJjOMMrg0UWHUXP/gLRv40nSEPCcHklEhP
k+FGyKr+8OZoYjwlAXoKxHRVnVvv3bvDSlCwGP/zySPwHUkyl6oOhU14wGq2MUwhImATEq0ucPNP
TxpDKdClAD8QBR/glMSPthR+fqiQkuZzfYjjKWjDeqW8JM2+5LUNUZfe+wReHWe+xmIJ8I6Da7/Q
xdXS7lEwTqjdtnMMVuKWk+ftbAmA0vqOlzucSNkyYmw2oHrqXcHnNOgXdWvjMve2n0mNqzQgINw2
oAHKmMOasam5b2xDHcA8494ZQSUX68i4c1ki8mvnt1WytmM67Cv4m/+9zh8NolJYkO51EqtTvVZT
Ok2whiXYOl5fW7coIxxB6Fj8XUpbZYZAfUExaHTH/DSBX9fW76AIsGUBVbpkQACRlvXdGsKt3Iik
GX0XsOP6cMYyxqNV/JUv60uYrWw/c3zKwVr2VUMkOPhMJQTkJOTW8XYZzD6uHHczPlJTAzFb+rKf
Mdn9Rn5UlgBPJRg2p0TSUnN6nPbvaM25Du+ZfdtznsrOVIke5GdUBsDanECuCoW8rvlhR3Ubvu44
zJuNifp437NY0d3rTL+6mPmcdInsFkbzuatIqWABbzcg5oLGZClODxWZ9ThW9NZBvgMTkQweQk4a
mmiQ7h3NZ7itGZr1uBbVUU72X1UvA9B5Hnjz9kuVFS6navnPfu+zME/gRSLhAAWm0JIAnYWZWKga
OGM4G6/99Jjtaw3JIndX7M1T+Y4Zbo2rU57opaUmZ60h32g182h9TPLMduBDo1puQiUvY3zpkpJw
MpNnH2J52cHCkZ2E4V132i0hZbqF3A4r2UWIZrxAICQPll2NT+fvIgAi57/dZb4syXtJ8tL2xZAk
u49MAcxIk5Mh59u1vIsJ19uv5F8y5i7SKltwmEJ2ISkmle+fbhJD/+IthEj3THPz+WTBDdG1If4e
2vbBfM6eba9cvoVEZ5pLgmx0crDe2a9WMEKjobHb5GpgWF71040o8hhtpyGCQIyV0sTliOqn50lG
fWCkfKdMEqKid5wOvDHmVrNHi8oAPrmOqu70Ym8Pa8g2NzaB+SUYRcNB5SPNoLJ3Ybr0hA8y35SH
6ujFj/bkrxOjoF3CjfoFOXZbHAuYAAPXkIx4/w5cZ2EqmwtOOfIszsAebztomc2JV2M5vWouX+yO
nuHc7cEFUUGEJezNPWmPr6x7Iv3KoVOEAwtxtkNJ5QOOcSDk2kAbzMwXYIPC6QT3dJcbNyfcrgB/
z9RFYS4AnLaHl1wWT47VQLO9/apf4KU1MR3iqv/Q02WrZ1YNfW24l1h8ZbCnEXm+z8mSufDoiwk5
NT+1zGot9EKslHZJZ55v0tVwBfUjJOu56fQqZFsmPyj9UYtxHprmZ3/HIC+QP76sHEQj/R1wAzoY
rsBzJMRc0X6i4EBr8dXBTprtuWbo8xN4Y1z/SpZL7JpInwxdww+dUSKUPXbG0eqjpvDhxC8GP2na
7HolORt/rrzvwoCcViLMxUPwv2xyYoeC5liWSLERPePEPbFZLFyQGHGepddw6rSIfxGy4AhuRNO2
flBsPQ4CsTaKRoJOovawGtjoEhCvJ0xPb0haKofB7UB4LB9flz5ZZ9UiClqLEaoim6hCnI0tuUHy
lQQ1kVIUrE1f9XsNXQFmhDZK22EhDTy6my776X1YWxN+lJuEAxGh5H6Z6Iw2VkzxqKhNky1yf8Ot
Q2w5BYvAKqvQ/9On5A8Gy8xupwTFiSxccRcG7sn9S+VW8Bak9SnXLN/nirekCr7Wqrpq9bsdORx8
/mFumSnn6m5up79IyOGqj2iLSAtsQzWvBXjwdAEyqV9lHi4HQd9h3ddiuXH83mkyC3vJ6Q7d0w+5
zVrfUZK29mIwWpMAiPUA5hlQmYBGGbRPaY7b+IMaegi14VmcrAt+irUKX5r8cJihfdcsWmmXQM4L
3JwBuDrMo/vXd3Vtx92Ufbb5EE9aeUATzaPd6GGTGRd3JcL5Ts41kxM89AK3blzmLGST+FQkQFEA
4QRwmqWKqYarzgB15sj6hdJhz51S2qoyuOdr5O95C77i3nd2GcaLA/1AAMHZ3lJLBdfXMVMJhT3k
+Ain4RDp3PGSgEA7mkZ1vUVE4XPsXMtqmXWiFySnNmWPxwV9EcMCictPxzLCd+iAP0wgEh24taVL
wA1+z5lol9oQPwcQPu7OcrjcJvUCsjnsEdd2MpDBp0bQqGcQ7pSpEKTNzAAXWVdm6Tu9K+TrTGED
RFGgILyMkdZM12J7MfVOCIVdhV/s1VwzSeMxOVWZeZTBQxO7JBW11PWhg5zoLDX1Rd27vIQX0CDS
ySAthOVIooKoIrbOo/yknu5fm9Uj6gGHXVlRnPmiOu029QAGhSPHMD+GSruSyaGPscDTgDfM76pu
WyiRkrQ4Pctcgm9Ujeq+ihP+R3LBCDzQUY+YucMjw3ok0xxPV8VDcsndGPXpfY8wMvQBGJvR605/
58s+ZiBircU3Xf40GqctZVTtku5spo+42u2sI+GvpbI9D6vNtoTeaY4v/GBI2MBZbIcj8fm5Ejif
OtCDoy+JQ2NIsPivdH/YjU3iPBaB51TsWrZjgVjtjuPGj93MUf2ip7j30dIv90EedLrP1fmXV66L
oBb/oUbkgrKdHTmwGiBTMRpBe5d/RYIs+zeLWzbI2sFhxK4zzst8wIuapYK797hEAohOLzIbIGqu
IQJMsP2TCWQ7m72XGQTorbbPC+0kRT4eUHQ6BjmcdNXuI8P/6miPuKPjbVLuOVHjBk9uUuz58UAL
cvitMg+ceRvGWsP45fObtpJEevwsJR3H2LcvJ677n2psmsFTjtQkSwTeufvtfGbLcigOTjtl5Wre
lPviJxMvCmF8YKkwaANFs4oc3HJ3wJbobzG0Xa4+5dD0r8fyr7uIOyHk/fjx4HI1cvV1+vGJGX5+
kJqMH+lX97bs2i4xZ4s3rYilm4VECQzxU5Fzcq+l4u31Jb5QF1dKhJ+RPQykWZgZFrx/yQMJ1QvR
41a3y+gLO5P9aTxanJtt97pSa2aJlSy9+HqiAZygpMgBLhzW5PG35GZ75fHrgga/h8TD5D8qrBu/
tuZQ0BZnwsxaX1xqzALlRuC/7NviL0ZcJwr2az8CGdtuGT+rrQpZN97CsDh4+MZ2stvR7PMIjxgH
M7k63+eP68rsoO3RUcLjVFQpgOIU1gZZ6FiIAbVRPkNG8dh6VwilGUpmJijWmG77Nwj9djW9J7xH
M9erv4lQALVCI3hwoMXDr9Y3aPIC+5ZUx6heUJif/So42sx26QugHM1ahPr0DmLVa7Z6PxlL+D06
0vcywgg3TTO/jaVieSh9zldb5U/klBmWc+XFUUGPvrHxXAfKg6F4Xlg9ww/IcW6NuqRSvJS1atKG
eXni0izOObdYSjvzdRzUN2043f7JLNpFLGHHrDd70YT6xISQ8P7pLuY3cMR/5jAhqgzX41FofYJI
EmiYzEZJH6EsOlU3/qCQlQmz2kVdjsFhRnjsRE0afkRJapYSyohV6EkYBAPvivpuIsZXTtAR9cgR
mmByXj3dvr1VA+IgKgBOmf9sQWhwB4xIVGi+toggxLaRFnL+F0kVEdRDYq7d7F2OjDR8zOnMkgVe
jRCCPpEgr74/O4KZIIt9GR/yiphY+YGPs8Wi6WxYUGuBU+bgby6TJVmch+faq74JVtnwwRv6tOc0
/a5tj+XMDt5Q0GQCP6IwkPRL7dsIpdtDztIADtC8S4B5OEs4ofCuTVfjRknJSe1toWhoHEieS3rj
YYaihZJNtY/z+t8e2DfYPf+KTHNAEcnM22iYJszzJH2ilsVo5zDPP2XCHmdUj2GrM07WDCRmyOex
rWOLo20kU5AFOpoAe02D3mazKYPh8Io+oi0gbcBlToKxKsa3MWBOiS/pJgt5ar5Cb7IZcGKUPFam
RKSIlExjT3mOFD7K8ISIhhBSwR1oZV3vP26ygWHbIhN5yPgJ1BkhaGXCD1Jigr2/9j40o7NMIg79
8J25oRnTF6PNzymmzKI7XPgde0J19n9iM5pjpBG3eEL8QqLhjQbHWAWUniNS7Zx2Z09+3ZCTkm/m
yZKqqOUN8V0UzR9nQLOMTc7pkaNbzCYcNnHcopltxVkTVosgR+AiXK+iZEK6bA5DJgHMuw89vMUf
XHxIaknDBWp/p3u+XuM9qgTj7laCGfYaf75rCgsn11gjTy7Czpbh2LkRzAiZJ0nDd/xeEU4R+tUi
S7xQFpaqbgJ15PCA1Fo/m1c1e8EqWVjPv1rHzTIliE4blhtTlCw89OCkzL5I5OXAXRQaoA+5SkxY
4duPBrDq3r1n3qxByBxx5yY7vxEwYm2ViKjwPo0in/5tD0tZQfbL1b+pa7rU/HYa5/vPG4C7KqoT
jpl0x/66m9eskzIvTqCu0f325pNhHunVqC4kb+xWzfG50YyGrug3py4opN5zhcwzWQNQg+4jql5x
8GAtEHg1pKi34o797s/g0ZgD4NuFojzNYnd13v0RlHjjoutZ9FyMyJs+gFhHQaHWpqC7mbNFnDvd
gE34Ybng2jVboMLhnfOVak14MctdTWZQn9h1GYK3NxL/fkL0qqPnkeBZFBTcMvENJDc9R1GNhRi0
8wi9St/dVbSTgE8N9FjEew611w3bCVE4ElJCE2dj4ROFSN7NK03uTazdXzFjF2Xp5wRpML8LGBcf
ASUr+GgNHXH2Ore3mwJYMpYsoUBcC6lwWf91fcmKUpOe1s0tOXDKAl7LluArCuSpPBhv8ybE3EVZ
2dKuecWQzjVdMLVzt5agCuEr2mA6Ceywn3dG1N9pEM8O00TJ1K6NbBX17zjziC+6tpA0Oho9MB/N
khaqHsayb5TqFk3S5oAZzOaBKLIFJtLipKPWhtFiDCycbmx3oqDGfZItL86c9T8v3rzWejfRl4rk
wUHgoDpQujal5crzm/uS8VISl06OCgPVErFbJZHOhKi7oK/KfTs6x0CbyVnPusop1XNs9OuyNnsC
g4G8PIV6AVGcbe/iYa5HKURapdBNif7ROZQWBKj1T/O4kagDGRxk0N5TKHvWUHZ46T6kEjkyUVJu
3uDYNCF1nNpxpd/hrF2+wF520j+wm10EpB2NJiRzv8YI3CSXkXYwK6yok71MRzGkln5kwCba2YkL
t94xk5LkQKiVc+CuC/0THsuXe/KBO1IImB0PvyZpwH4SEOcgR1mvDSuINtTVSSO54+cXj8wdupU4
PXY2W3iiqumUM7fODb2b6dq2cK8SIW2trwyive9NVkyk32tjXKolEB0pJH2JH3PkXOYKYQysVj5e
Kdwit49UxIcBe9UeWG0ecw94csDsm9ts0dZlqq48YR/3a3x9z42gJfoF4Ht5zDI8qsymIfvaEZ2Y
RCMX12VNMD2uApdEERvNX7u/0bDxnOD9+ovKUcq+Nm6s45HKbsWiLEkhawqh+EBhoQL/Kpbj9ioz
9glTXXBoxelTcxjw5LWoPkJ8A6RNBzlu0+UpN2wYJ2SStNeuTjFMw0X8LImJqP5g9+PS9HmfhFcJ
OplEK7KkW3VzfwXTXxjmERibuW8jIj7XKg5Q5fuwz0PrQeTlPB3t7CCvDNZz4NKG4jz2/tRB3zze
BIBwyFMFJlevbIN+gARaaEmm/0op5nnhrpjNoJEo+ktb2lHQCkmf/6mqNlwr58zEcDsiDabhzZps
YGZu+WtZW9BmBpbqFSyvH5TzvoRU/tO3gmawbVneYxxjME3lpqZ13jWwZpsJFmFPjyAu3B7S61BY
BiaEF6MWhj+UW2e66ViO5T0TB+xDDeRGIlQ2u26FMbGr6nRZ/Nd+7BQ80KYJX8In1sZ8F8Zp24hA
p4HXliCylqUw1FPD0rjaI9Yj/NwxUDMtvl9NnIFb1akqt+Qr56XJpvNmg6sE0PXIQN5zJ1AskbXI
0Wcs9qYTlLGReVekWj+Wyr+JAEr+Md+8szoFmhZPLpGiK/1y60PFsMDoZEru7H2gCZeJmnP8gkXc
wlzwjLwykVGLOa7x23yR3aR15FwSEz7Nhu6liVO0ISaBql0Kj9MFsPHxJNJ1vgFzod0NJausLwm/
BviYUxQfjN2v68EUMydoYNR7lI7PqjK97GeK2pHUCCNNmAHLiHc60mmrHyjIBCdthEUtDYYKPy2u
k88VMQrSeEmqfl8sHA/mPt8SPi2yGttdN0kZOUYUSM0Fglok1aCxlGXHytEBJn4VeMdUjqOY1Skc
VAm+o0eNaPEUJgJSTG2tKySWDPYdjHiqir4gfDA3FAr2wGF7asMX5n241wGJTfRWt7rON7cDp00g
z7UUUrIvLJwYK7lp+FM86y4KMPqJIRGjEJpqXHmaibdSxLyqgwn62x4+eVXlxIBi22uJrHnjal4R
3vUNxUswWXz+0ieWal9XpaDGilzyjVp7d35UAxcAqhcDVBUrwRiQbATR4g13A2tLLDlYFIArXo3M
Tlcv0TiA1PXtGQWQA5djOUdbPgZCgmYx1l9cY00FBtjhhXew3M5KTyHCMPO1X6i7T/lkF7MPGpM1
Hk539eTOeu7CNcjBlwZUQ7pXvYFt+3NYfwRMQJ++9hyja8jyq7HfbI+hjMEK4C7BoUg6OTd11o8D
hJVBetl+rSlxizCh9tFBH2ZxPHKxdMQ+dxa4NxmyXIZWLX5tcvS29ouzwFwIXMkPudRwrzBrZJNu
2lYIS2RGA0A+5XzUOm+yOq2i1/TcRVP4S+tmR7ORz3hawqShOQPmyX6Yi3/lnTXgFM18YC8AqqfB
nzoFDcSCqP2WKhV5BVDLDxdJZ6zfN3kMafy26ssCo6owHvoOrZYcQY0kzcWw7LSeXDo3ECS8KWXa
Vv48JTNeNm0w/o8iHG6nmciN9Anqur4r4FifX44hpwMki2QN/ZtMwoXC53jujUY0XeObYv+v1v/q
Bc/ZLSuAD3hk4/ZY6PAJCKowCVy2f6dhvMWBxvGJtq7cnxZ3oq5pxooPfoBXWxbwDwT81NKwzVOI
WaM6/gy4+oc0dkWWwjETuOEg/TRgB172aesUCKSQ+/2DIt59ozbiAYDRmGWJxWZEMQ5wrQLlhqBv
L2Ipo1nwt30XCeQxBjdVfpwYeCw6iS431iKofIxNnQ0YO320Kg/tY3RzNPrICSRh28qnqjDQMxbF
lYkaQYftUw1i/8ENJMZ89Jnv0JK87R722g03tDqIYARQhhNxO2vTK11jeLV+1E7zV+XAdpKY9kuH
xknk/MAwyFHofPyif0cp+O0LoHozbU5QLtKeOgfBp+/PknMPbk8VZ6tua607UcLu3YFO50X2WpZ5
TvpLRvuK+JS890Zpj4I798nNzjilZaztC10GX4oRAT7Bdw/5S51qNuAuuh4I+J1pgwQeUUfpYs/4
JKnZ+oNMonk5ZQ8Syoq9WsRQOaVL9jL/HXbmIwlw2/7kduWu64JI9KuOVuCi6b0Hjc0ewkLeNzN3
9fUuqw4Wb/K17PzFX2jw6V8JntNGoJXUZtMQxrkbTnwD28vUcley3RgeCt+ZIc1h8W6YTKeRSo8g
03vJ5ty/EQXUjeus9uVvqwFzPpjWdnO+3cFLGaN0hW80VxNNb8r6HWcfpy58fgRUTA8jW/HiccNg
piD6xr2wAICpLhgiQVFmo9NVuU20pWPi+rAad9FWNQJsMPMZjBvSWd7yUn2EHjAPDcehAihHCVSo
TrGaXaEC9Sl9bkdkvIINawfkyUCpl6errXneGIvx+rPKyOQY1qhGRnQjLtKE38TnSelkpxZtVmtM
oHpl4ZlJGhjZZkpid5Da0nZ9HqhfIfbDLJG/EfjnpiTq7rQznQ1NVZ/2T+8UNlIKxShWe7nnudGy
z+zAMh5bi4pOuNH32rvJAzFyYAtOgVQDzso+sspEM9BnUCsqFI/Eel6PtzYIO81wzChNKLvoQp2P
TNHKsOgoxGlPAO2zJ/SgbWA87Bj7e9LJ8lj03TZ8upnvfTKtNX8hz0LXcSgbRy+ASmKL52cfOwg3
zqEsfL97lD18bQj9KFw4K7oNncAvcEfwJjH53fn+kNMuNEb8/BXNZtTITbpF4KPNVRNe+4MCpaHN
jAu3UNy4ni6UDzFYaFrs9Tj/p0It82QjH6SuGt5VHwhJzPBnt4Gd0vI/4KT9jA7jxClVDVfwOXDw
kB8LkHkbN4OclAHFyOT5icpLgVxnBsykBL0qlbVTAWm+2r7VyQizPW+w1hdKXvkyaasgiKDumJrY
D4mX1B+tk78JRRW9+eLvYRHi0cqWcG23YOXYFEtELnxS+fxkVtSMcWy+X+krPMAjGn6x8M3J1K5u
QgJi7J2tlg0wlzFNbfQoUuN7uLxiBwwarlKcA5F+BwdYCyeet9GY++ypHRepOTcxA/CZqj1z6Utb
bG2sFRofoW4JavkI/Tx0pYH1ayRsFQMzn4dCs2u6k7LNlRTM6s+2pL1bbW32li2bx2xUqmmLHyUC
8pNWQ+ibAj/23zKiw3k0DOdzh4gM8OvTyB7dvmQnB6o9TIhp0qVYlXD/HgAn95C1pfc1NO8OnRfS
MK/h/6ieu16ZHzxO2hrX6rL7ZVJ0EfaFoNgnZQe6XbJJiAdhJnM5Kt2VOKAR3B5QzdxNZXSY9XhB
MXpbym5b57Xb/cbfIvxn0Lssh22WWjtlcrFWkkIU553UvGQpogtZV08x0Por3mj2Rcu+BZgsCAxV
WIUbP2OdbHSffHkNVPKQ+xlrDMEDa4EawCTCbzHxKBaglzxRFk/xX3R9TpeTHB4UuK9RsBVWdCBT
PcZCceNIDTuzSnbZLaf5kXKQSHChV+TVdDM85vR9RBO6wf985P4cLurMGpMFH1x0eG9p5UP2aqtq
b7NZToVbSTb0YHhazdZQIgrM3rjRBbovgnO1hYfWc6/LAZq6VaU5kdDYa/3Ojhm6nmmeO0IBMjpE
X13yGCXCOrSIGsnpF9qUvgtwgQETscOSTpaOyl+bUJGSyY7ek/fPje/+lxxXL+Z876a6BnN1Ytt5
Zl2dOPNYeLOThXVZXsiIfbCzW8IdxkxWLtglck4UnDLfchIp1R4lFVxL8Jt6U8v6iQ5EoZGnb5pn
6d8E0jBKq5CAeUP0FOAOpyYpRCLpG4lh1nUV2gXQVs+9vNXO5k1+kTgSoC0/MYf4ZNjiyGrLlE0j
WcOldAXAK20sd++8PW7L7OI1XkgS6KpZFa/AzaCdag91baCp/3Vo9oXfkzmncuU1V8CejGT5wbfJ
inb9WKGFNNz/3q9n34qWOQvvbTqm3c8IWE7h/3kJWi5Aqv+WuwiiE57tkRwJcejqU8MFp0FWmk9M
vfjNEmWXXt5tS8kHUse0OspmodYgsQ2sW7PhqyQeoXxzhmKY55VqN+n7LRrFvkGpTXqyzY+GIK4D
to4ouUvB84JtLNE4VEWJtCwlCSVatobg2jnJpgnZOgXdK/EIW8f+/hi4IYMJbDAnhK2EE1+fwL3B
AA4o+nlbQuHyypC9ESNC60AIC8TJ0s4F4vWS2CcGNgtMQ1KP3nJLPL4UItCWLPHt+UhmGD8PxTy+
MsXM3kvc3amptErnPlz4PvYXWhLEaiFZNqGaKa3Na/Bt+K5DLag6jj99nZqyg5GcMVyE0HxJyKM3
zZt/Pg+L6ZoFjEphdsh3KjCDbDemOi3WvwshGcuka7WuJquVcBgqeoN9fNKy1tTe2X+NCoPiECDC
Jw6V+5NLBZok8Djq68ApCQzzTYexqikvzoZWr4sKalutkFxaEVNxGdSDkKBhMXxmojD/7JxAMaG2
WNPWwXZclq9i5Rhjlt+SYDP4J9D5G2XHtXTV0kp2NI7c7d3av0Jo3M1ZHGUbW68EoUg8AmcCaaqr
sV/wOua7s8QtSHIZsCsci8oyXpmNdINfSDfox5fCWTF3yRY192RIYtRm9vQdz5HVpjoWHUWoxtIv
+QQv+ru6attOAQK/QYkhxGARGHgxjZUO3+Lu7QAex7bVs0zkoKjWO9d6FBzOCnrc58bs44fwUaBK
VhHJA/NGjnPwCHl6LHURBcWGpLxOg7i4ReXzSWDSFTb4fCe4kIr4Bdfm3mXbbapqVwnZ7Vs5bkPq
ITx1m1+tzW7n4cpdvYzmMxjebJnaEZDuHQITV6JonoSO/b8DbemW82RnFfAow1kz0A7Q33HsDcoF
u9oTMcCmOvmoFHfabxHJK5ZSEDCgf3szde1wuh16HzguBAxQNG0mNnVQzXsNfJxqff2xTOAcJHru
1OOkgN4dp+Ewv5rKK2sd8cePP58C/m2f3iLVIMmtTlypDyW+078abea+l69dtC2CLn94sKOI/38E
Y4Q45AqYtOzwtRUNCCHoKFoRhfUondKUTJ2CUdx1+eIZbRsDZBhfLFmg8fo0c6kcigUVsZPbkjQl
btk1GnKc7ZLnLcCvQzyoNBOsvjzggI9+kHD5LnSL7va08q5TOkA4xLmlvWyA43AJZ+GUhB1GokDO
/+FTgWwVyIUAD5FGkvCtlA+Qw3GVVvda99thcbHRGSAapLOdOmlOlyndcfFYNNlHshRHd/6zJ3go
WWcZC6zjz0L00yswv7nEZ/JUxaYMpj4MwLa2vCFx73o9COyQ9x0phPvxQuMAPY0Z57GNflcAnPsE
ktWo6zcg+AHzwHLqHlAWfywILEKFl2u98GuBUHVWTM2/RIU5EeU0I1VJ+AZtO+CUCaNQdnXMCEdp
ztrBA2G/eoxvTS0G0yyb/bJ4of2y3i838OD/h6MDE8Iv6g82lIKiAgi/vVS8vI6fwrS1pLR/e/dK
eY38qPaT8MSxhofuv1KEZqt/NIMDbszKqHkgv+84Kf4+3jEB6F8untSDdGqU+TMt4xT33dQE+ZIR
uHUUKKYwF+sDqukwVY7Bp7KTYRSOkfaws6qcCTD7yRtVEaRN+pOReeF1Ys/N5Fa8K1bz2q/z+5+G
HIcwbiFh+Sf94wUmK4FPaFABGSrrLEPi9RfhU8OBdOS1mYwpKPgQ1JbmQzQWMNkxokAhczyfPgJC
4+2jLj/tbxZG8CoqFExm7pG9oI4k6X6tbe4JQ3fWwprPguBtOdrgNdye87HqZsOaakQhplVFs0SL
+9bdnMOo2vh91LFsN5cUsN/pv4pEVZgA/i+ZbZ4HZkEbYkleBn8neP1f2O+AAMdWR8AfswKM8o/X
ZtkXUuaZPdLFwI5ZCzqPX8shcNig4EgmiHC8q59JppCsDC1IN6ndQcCgAVnNdaJNgJxnKNZybFI6
xmPOfhCt13eQkBW+TiwBSr6o0Qeuq3dwVIxfWMck2FQ7NqZn8+WWX0BGeS5gMaSlgHaElJ8KvPex
ATFOBb708V93DWXe3XBd3LyW94YXCjUR5wewzwbl/Sbjm/xLPfjlRgdngt9dG5cfb4tYCadO1H0w
8HyHyXpwIK4VdmyR3IQ+lRyrvEYntmuJPbiGza8gQYl6bKVaEg1Xc2hF96AqFNBZSpOEPSLRxUZ+
jdsfGV5iiVkVTzr036YsCKlSf5HG6erJLYdelqcIHvjG+H6KeQQVGmMzl1Lk62B+HKHKT2iklYur
i7HHlu/039a9vh7FbfMgfRlxzUApFyXBHgNjRN+bKSCHNOQORPkbs8nEq5tEWvgfmhj03wjePM1M
zrJF4Z8bpgx8ZLmNOwfhBf0gLTSe3b95fJX/UIxez8JlY7RNPUrVN5kIw1xooR+Qtl3qpKeVfXBg
oA78GMKsieMBwYgg/th5HZ/rRchF7+VN6cYeYzKL9fPZaJkPKz0+8y7fM1MsvqgOK0e/8nfmMRzQ
MjaWuUMGKKbTXTKSjTDWrO9VGs4/a0V2Adjtkk17Ff8K92dKcDiK2PcInF53XRUlBrM99QA20p2C
GyQRxoPmKJrz8gS9fTni5vOIF3TcUWMWHPRMOmXvxGIcbzt+4Znxq757sIHKZG3JjssC7cxSNABx
38y/Zl8zO8sBBiArRSN0gB6ZL2B3vyWoVx5DnCe4zoJUZeQ4URS3Tn8ArWpXtrMtvG8ZPPbYNIuQ
piQtJ5bbVDw0IkSc4kWuDMD0GyVWiUgZ++qVJY9ppjUh3ofi3/t2CEMvZdRv7slW9mwDR+6Ztb3U
+wy5JC/2fEWL+WAmhs91JAzvUpcUWYsli/TM0Tr++BWcTr56V/iQK/+gKJXcXEtq+wcJkYTWotQG
cpWbd/haK24OhcXPkvcKcW1idtYNYkuYbd4d2rGgIFV8nFZIXolu8LXRNAguTzqIE3N2e1xstA6K
xOv96fOVi9z8sRh8IgM3byB/wyBCn0lJC6uJsivoAcZVBpHqM0ljXzYENnt8kPAEic6iCbmjyB+p
Ej5S5NWCkW/VdVSPMfF8I+F727L0WNGtBwgoAXNznIeH2456FlhA9Oc51Ym8RS0mmqpn7ItMKjOV
+IfY+RH6oZT88m88XmJwFc7Xa97CfY8cv346MPyS2tOhOy/4+vPA9bnpJKo3gnKBp64Q0UQVSbT1
ZXaBbbuUVxwfOSw/1QPlWSABT21rE9Eew7KJ3kt6Crzv9ECwZD5BAd/oyprjqTcxRxW7FhWMBT4a
XSqcHzFsgSVVzzuAuKdyIOwdW9H0I6G9Ue2cYCs+z+Wx68JpcHuqxNSW293ibv1TDzKSgULalSD1
RsYF92SHwCH+UTHVj5yiUWw/DFlrMgaVELg6JpCVbPpQpGOiWsACwzIwUT55NVHpiXufyLCAkHZB
8uzr4jj1u9gPciPEyrUQVQ+bggiBf+wPKqaUDBzVrIX/X9QqsMQoN5iW9eJi0q0Zz/T9cpDHjoAr
Kkp/DgMpgUFIQDfY//OLEXGnNHgN++wnt8o+GSdjRN2XcGEMf4DAqd0TVdqqRh90sBqXM5U9dccU
Wn6RT8cX3b7Bjgp6IS4HRAq1XkI7jUYMf5omcLzJyEyZi2qAA+OFhAXHDYU+aCtiVRgYM5VrTquj
QL1gxJ82trCVC/Rk3y76Y8nfUoYAjCXdzyzgfz5TeBWThsWIYjnA/XVHY8kacj+whszfe4gdkdht
c+mvFMcYNi/Er9r6e0NOoV5Zf7rZxMJCWfAiUyik4yP/itWhB023zk5OosN/DsaTRTrb9N6MLsN8
P5a07RKJgkJ0abYiscdLOonL8jb96xkv+6DFk4B+JwsQ3r7DAwOfzUGJxavQiPpq/wmyWn2YYdEB
42i1q5CuESQCDt5L8hWknKbZxGjuUWYoPtHagDX6mYR3yGM48PyeqZI7A/IzcBbRsHFGlPzWxLLz
GkMz2sJLfLORoh/sWlW6wqGFqACJea/PLaoS6iPUH1VwI6c/+LBh6Tnjw9OuC1SzZHd83EXCnYL5
GORs6NjlB6wGOAwNhN29OtW2z7NPZappC3FdT+DOCSFL+Ngv2uJQAUz+dRX3VpYWjCGJA70kzhdM
JALJ6whHAGx0MCyx2M739DW9RBoYwoMyPjosni3+K4DfUm05ICC931iTK94U8ZU+YLaT+gb31E1G
p6EL/m7CQuewhGM85xCc1FtcE5I70RAI8QU+tz2iTCJ1X7kzjLgodfbLyUbWMxEUVtI+Co8HY9Sa
UVS8O3K7IMIbPYqzv279ehhntsrEGcKSahOjNInr2EflYXeg3vC8u4K0Wynnts3Eoxy7YJrQNTCT
JXDSNCl4Ui/4RaRNDjwMAJN6PbSv4wnUp1S/3/2hwAn/cZ0/K/zr9P9e+OXmxvFCy09uxMCiSMyj
7Rj4IHbN2SknYlsd/0+ORsNMVvE0dWgLZ7oBlNYlltk0X3FPcsYHldi6xSLXyxJazlejXOjcA/17
tsVZlh8uKAvNqQPbqKauOV2Zr5dosmlaga6qs4Km/wuuT0hKZrbkmRkqLK7YgSalbLHDlsIj2MYY
fQpQ1DlOre5Wn+Z0X2EzesH/hcaGPWb1yudncvOQ9nRCLbMfpTEVAzhhb7QUvznE1WyT8W4/K6zL
dUJcZrFlapNJhQu72fQylI9sACp0b/T8x+0MiyBEvjARJRn0Df4IODPYAEZl+eAOWg6Lsow/7ZXZ
rrhlVxEZt+WtqaKi1LIJ9Yi17SO+dNcU6DSiltGOmwn44I1JT7aN4uzXHJdrs71y0OXxPHZ3dW6H
DNgr+JjTzeTrNzyA+8QRHjpRHC301RpOmKq/tWAAs9UX6TxOg3xlJA6idiEBawvgcxYl56LkdtOo
txNkjBY/aiJCa7p+EmoTqII6XkmjjojIt06SpEuvdaVVW05s4CqbMlqQ0og4c7oNS5N9AIHHFxsR
U/l2XjCJQpj/d5Mmb+6RCBpjeeY10fi00z6JUKZ124HLgFeNYmrJcVGw2cagUxqdN4XITy8LwlGG
u0ItwAOHdsIZjwdlA04IMNxuxetwjFqQ+T+RjrC8xdpSpnX8fTauz4CMQ96enIeuNKNhVjKsCB+E
lY6b52W2BGnMYLnLmC9JUhf5Js7BSbHQ9R4bUsJ6mYcJ2hGURCI3S/gj/jZHOQBmXRNGVfH1nYHV
mzp85XE7yG1nWIxpBKoCO3iKavVECuq+2Qv3Cb0n9zlp/LW5N0/WlX5Q87LUTuwgyV6bk+rdIn6n
YF3DxRA8m5deAbkp+3uS17N32qOZQOKoF1FDIHeTfEOKNrJljFH19MTlQsIIiLMdZGkPQ9IY8EZi
wszGVEh+P0sEECzE8krPZS/3EvKqM/RwraSKPbfLt08CS+OM6ENS+q1NGo4dXoziWc2ccNLNgFR0
WMy0uE/NnYZsYYNIx5SpMYxvjSH9iLxqOwF9u4NDta4v3HH0RNur+JYTk/sy0fcbjP7uqMEzQyvy
zeLW4aZDtPGaosYQsiAaz7VBpdcEy4SqMBA56PqZkDUbi4icpxkndqTPmEzyAGgq2bTPFu7e6AQq
9gEIoGpDVqZllP08mvVxpXQ+ATVZ5K2DZI/WyiiruEyxUTVzFYtXg8YlY85X9tGoKz4LV29iCx9/
g8VcJQ/R0Xd8WPd9oxllWr+2QK1UMcp4ZWTjcOi4LC2fLs88UTKVLJYGhFCe1vKN6TLraOusxSxX
boYhKyAmiVPtWuTTrj+iEvnZv8iraLkEQ7ZlPsU9FDPqtVfuaCUfM5YwfZHrl8/xj5VZIRuW4jtz
/bVL1y00o+LbxLAflyrvu6xYyztOGrPo95ijRIDejd0J1QvpVTMkqio9+OnJcUDyQcKlGcRIP2bA
DZLsQqVJyGiT3f6/oIcQ8bcn4W99rs+9Wvjt5QR4nmmWMU5oRwgDcJJt0MBe+xA+ZZSB9G8xjdgG
wdafi0lFYwSHinr83DLMVGIpSdjFtNFmAP1cGR3fd+3YQ6+UBEsn7Erv7v00E/tia88PTOBjF/fO
wprCTZc390eTcJ8odf0bLrzi61IrWkiAA9h1tVj8qt54ER5U0xWc2ZeeG0u8riNZKH7yeGcT/lu8
mKbqObVe84pUITzHF0IC6HTG5Ymd3tbjz5IvlMVpkhPWz8no6KMcT1n2RW/BPqSHXLyOC3UC3kLH
B+3Ar43FDRDiAaSTPsFlLI/7HIFG/T/oFEhIIrbeblO4N/u2nXPz93eOFUCjqWBt6GlpRJ/Z0DmU
LDjMyZwSIzAfKC+VzDWEnQaJvmdvXy/JX1YQ+Lkj64Fv0TjvCw3Jc5pyngNabqZ60dJPQz5Vg+Wr
OVm9wBknG9WfXKaoPm5vsUcCIwnVmZuKeovOiYk++bilUtWuGGaX+2dA/1fBPKo09ftLvu3P9SDl
AtGiVjTrDQivYc0xFiBAV3eHEpewTKeAfLhf+jnaTvCbUEZNDKInkIPcAuOLGyxNv6IuxjaMctrW
n20Ppf997admmcgMbREf0L/nsdKRhWVcazPyYSL3I1npm0r9ROe0SH0DAtaPwoE2rcpErLSn1m4P
rD/k7TLERG0C2WSbeE3Red7VWJoEBPb6RdH0AIObWCND6Ba8iFswlI50z2ypRdyLz1XqQnyyGpWA
EK3+BpuH1dpf0JpFRCZKeFcbEBmDnEy+6jNbH080HgIeYK1NzjalPAQwtCbEF+vbH6Pub2typEo0
EIEEBiOLWjBV72XJnGHm/pdxDY4eVfRD8DoQCrN6M1g3agLDlIvOmaOYJnYTxpI67d2z0rhV5hCG
L1MkhiqmnSdqB0/UP8JLWFnAVyw4xg3+uk1dzuMLuwjpwTuBjzmGTSj1ZaGp63h6apOXsnklSmqi
JPhysgCEnAd2oUvhssPR31RX4AukKSReIvYXK23hhzRnW9l+GPIjYZ6abnMMM5negIg8N+HfDuqf
PiK5bXK2l7+RdtPMW7wBdz0Iu0yMFf3FBU1bbvW6ufUo79C89clgvjwk5r5B2nJRxc2ZCODfzm4k
6MvWSGrJSfn7cyyMWzrEhyBy35+F5uJn1POGRhEi2+YlMK5O6g+uGVT+R/guwINi45qbwhz6q+kR
Hu66syui7B5jKKlRTnP+Lee4gcyOzq+8xeT33s51fKUOHSCC+mBrQzljHA5eOptqOq7E3uWdg/7Z
UPnoCbE9vCwbfinzUG8Ip3jiIKzRxWkJDOspMhGT37AdFM95Hb1IhxxxrSZGS5gxTgjVDRq3bInD
8oTuatZko7zpdr1gPq18v1ke4GmR8AwMHBtiF6HxQ71jrUSkdWM5vh9wfhgDrrPCNMag7I8x6OLT
qT+4Snc2tHwfp2pQ2J+NbP+JL1PPOuUQKgm8sptn3FIBtES8MSSPRwpvwUD7ZBMqxhap+OJs7FDX
Dn8cpFhQ2ZfoU2iLyEo3dlML4E3+fLlt8O9CQBjG7Mx5/aGM0oUA7u+UfPsjsNpaOTltOLn0BPXV
u+5RaayGSnzpAT5u5nN40hOHDsA+e0l7JgW03efWkpnD+fqw6IvOlDcDwd9V8kqYICNgCp/jF+6b
6ghT/gy2ZOrqxEKbt8E/Bbufj9AUOXmOk6c3fvF0WaYvL1nS1EvF+0wcg6yEZ8A6jRaHyFRSjXNM
8pK2PqBLSZZPi8k0pKhSVk8580u/6GCDNH2BUPoGsU+Z56IlVT4Pme91V3L57s/8CJFbgM8Ke4Di
/e/9KjmXwVqGuEJjv8I1HSedzwFH7zIqbBhhCpaXcneURjlBpKlgth9Y5b+PI2IM4D3cv0WX8rZp
gxPcXFyrjFqdaATqkZ1SNjkkhm5AqHZQxRE8whuIjZ6eVdzIP3HW/aNcH83eejdzD8K4QsU/UgAR
5oOi09/fZKzUrpMVhUAaEXNs4WnFBGR5qQZxTiFPN0onKlplHwPb+GvumbGp6ieE+aQG5GUY+KEc
AADUAdqZEILZ/E5SDdSfOsSq5qCqXWVBqV1DHwiSXo3dkSrM2B1RvHyjk2PsJcwSXdJ8sLTh/7Jd
iVHyQUOqiZ1efoAWwkUHzClUEYAWUfZ0AMENG/Bdt8S6izhTl6V/3/M7ZUj+GcqQrsrU513SnUVP
bNthrb4TXQrb4XT8pgJhv9zZqNkmfz2Ny9qVWJ/EJ9dgsvOtL2EGMrhZ5cvw1wuXAyo6NPeDH8cV
Df2twihJlTg32kLmtGjWdxYY3k5Pxw9akyIaJXw/G4HAyTr692s0az/bM+31KZbpJcGopOkKT+L+
BxGKHn843QofO7h9z8xmmvTd81/qTdXKhWEE10i35587N9RFLx8eETfLrCgrmjKRK8Zst9vjzlJm
66qzeOS8wQYodBwnllr58MDuW4Nrr9DkgwLnFcpndaJjSwunFsIqflGr0jO+yUZwpvP1mZOtd6Qq
+qK4SsV+PMiQ0SyOa3LkOOUFDPEBDpBI9lKwuOtoql+ganC0Y0IxgTfPL/iIq8BcdjiIJmdVvNh0
irjjfgZcZhSA21yvVVGWBi8MO5xDhvn/frPlRvxfAQaUgZwqDQtb/iM+jvu+uV3S8Blo4wnei70e
p+e7JEEcKmZnVtTJIHpG9ZA3hPPu6ztzYy9KTZ4A5W5USQg3O6uFfVh1HtrxB22JCffnTAPe0cw6
3EjQmaPSxZ99sxa0ZGDRHaHyyUq6A/XozBD0fihcB6eSgLgpb73VQZIK1tqjsk/3xvSoX/kZGGmE
qtDDSZ8qgul8w4ru2gmi2wR+JlQMz9CKChnt/RLK/u6B3qYeXSu0r3MfeCmqy42bfF6E11y0wlJP
8r4NIEuHmEo20Yy9V3+6bkZqCqPbmSYsmJ3IgmMgCRcd4cd9vSu55fmuUvQFZHgS8A7sAO0z0Gtk
DlbJPrTiBE5jWOa/I+jIk377yDdNemY1aZS3/s63J5JnJDJZ3y5R3u8RPn4U3qtU/diJ1X87gWHM
a6mC76AHt1OPmJrkKVnn5oCFU4GO4Rd/4+u5qBXB9YdxARKpIQS/g39Dlz7a2PKS4OGPV/vRSncB
O1Abz9DY56ZvlZFEqTqqXLFPO5hsfzZNNvlCvQ/wRau+B9QY/YNI/Fiy6zmls8OvXWehuRMdTIty
mN+6qa/UN9EQgSRJU5vTjszvZRiUtmBEaqsc/yHnr2dK2Bh+KsiTw9CWcC0tLBXynV1jppg2GuCI
u3fYH3bJHsZ9PJsMVZ6/ugIdi/cmPBsTuChZufw4cAL4TUKrj+wHxKfNMZabNp6PMmoSKQcDXuKK
Mdw37KYRAzM9IVpbLkVtDcSvLfohuXrp+EWbjr9iAHQRCiZEmN9CS9oEtIdpfRSfNOAHm7QBHaXi
pjtFOK70nMnnH6PtllYd1m5L0RIHI521/7i2UXfU/Bg4X09bP+JdgK1rQrseBsjBCf68u88bUHET
HQ9q5dOmSTslAbvcUzPrHdRbu1NJPCd45UxIheajUOogqZan7g+J4TU2U+V8yLdMIpcSJyuhVdIM
flSJP8m0QlXl9W8kaBtTmuoR4G7wns5SIorSP2EGFThaw/8dhDQyYLHn+m5ghC5E2OF92PQJ2bsI
RuDyc8i11BBq9w7SuVN5/aT/hF27MDua1YatRxQBU5gNv42ADoZztOxh919H4ColSGIsTcA7WzT2
eJwqp/jdwO/pcX/YTyALSMG9w9yVWCmvlGlElZtlrSqOn0WSxTTlL0ukCX44VaUIe96uLRj/bGSu
TXJLVyhKSGJae87duHpM+expMb4XQT/Rh8vl92RxseMsrHqbb51AGkskSGHoIU6QGM+sdTHTiCRq
pERpGXvFtx1HuR227zw09WpqpeUpu890/KfFX7NeUHEXALJzUgfBmpdW8Vppbt2fK/xlCq3IFbmj
bh6phi99kGvoQLGUMF/FmckkV4oxPsinzGYTf96rLqvm9g3kf1H3R5F67ixecsDvYK4lYtOW/9rs
lQfk/qVBto8UNYBUbvNAec6NiLteKI3+QGCxi++yABMXV+xWmblp2lJYf6VHkeMuaClaGJ3Fwrrp
DCi/2RhN13aZCR++vgiPmVijpRFk4Xygn5jy8HhawFwrCfvb0WGkegYmJCHHTy5GN7O5yU6wii1l
H+U1MIrM4JWYSCAc8Pkz2CEfhOy0KHyXNuc3zZLZIcPLm+sZZX+sdBQBCEt8xy68EpSMcGRX+30P
fZdd44lrkCZoeIrgLqe3woCy9k2bfa54/M23z8DRy2Sz1C8AslTB9d1bm5sTxjZRj+9Bxd3f24qV
b9FOzIAsmNG78tN3Ng53eWMO+pbbrjFpgjksFG3a3nmjhOrSJRFd0PYgwVwdZt3gQ6fvzLmm7UeG
vw84BGmYyHvHy11N+Z31etTLsvML1M1qPvCPJspzOiICtrDZBRamrzhbZi/gRvbzFw+CQUjlfpjh
cl1dEKL9UY76K1RKsnPvZt/VMM+0YOuO6rlcOp0whUsDSGtE+EkJlk/jiC2L3C1xcqNDapZIQIvB
j8NEBbXEkQ7JLf3OVDcVQcnwtOF8ccAL00BiLls/XO+1V8V0fm5Qfw9gc0mYj5McFEmD7w1uuo4U
k5yUQiplASFOmbe6IhOUjUPVaeGTEhLd7P+IBO3muK0ZDaXT0fn+Tkz4CclWFKMqjUvNyPYGk117
GSlmXHUwJGF4wwE+XsVk5IYquE1gia8rjObm3xNAIG87dr3p71tyVt+TuVOHpXNj7N+9KfFLvUCJ
+IHgW8r7GHZDiUa8TWliYQL7RX/SbAspqZfu+RDtkwMHzGmODfO3TvDyPs1rh0+DaALtl/7bup+u
PzFqDx6OPasV0zSSJogrlhQVn9qa3tQqT96pjHL2rJ/E723fzUeulEjAyKViZLgUDUAFOGbyp5if
N6haYs/LzaNDndMQKX3lapSuKYWrYYajevAT2UWNPAq/N7pMDnW3NX5oDoAkell0tMDUEjSHbOl6
bwvskEUkoNaUFyNJ4C74OmL+3PPFHHoGCnuhuSClJO7sD1Z+GAuHhmZQq2SDOaA0Umeh4Ao9LUOZ
rUbUjsH1g0SLOhLWIeYYbmWq8OpQf40l89qx7wjx6lt5rlhoOxub6Ylik73WyRfuZNehtfCKJUAk
kExC10WNraK4XI3EXcdSQqMs6rqh7flHFbmD//RkiTd/azIrABCLGs3VAADsnheW2SFZ+epal13Y
KAIgNbMoeVioid7Ecn7Rq3EqTg8WVsWF2CYZwBqmyD3wx2ic7U9PgkeRb4ifim6YzGGIMf6zVf7Q
iu9RvM7iEI0jsGX0eSxKdrb1eFfhEdbYh5FeAIrAwlv1EZyrTx8IcHWwauDhvsug67MBwn9zVEGR
ktmeFjVLUNMI8w4Jnd1po1jMEtxnujWkirsk3GziwE7KeIVJLHLTFbLhIEYbQM59LlCzImlLhxYi
2gwGgD/UA2lFqjFC+335yG6cGLzJK59N2FU0ZdEy4vOeESxywjbzK0mFha8446gLf1NC/tANGl4k
pKUXWcDSZPFB/BFVtS/U6lG0ezsWnRQL1wLtYDUNDxFB6n20fRjfu6K25V9uaSilikx2LHmi+r5b
mQt2qIRU4HGato9PMQC+MpEqkdT++dNJuwM056Eg9Y7DrUwLRT4oELPJT/lAgyhRpvGjmMQmotdG
TyliSlHer76hnGBXiWq2gUKiFxZlQjVlnK5SCIpo2Mf21KTB74lZnSh056n4doKDv20C33nQYMHO
hvd15Uz6VjtMzVOcYlOoDlO/I1OBv96K6jH5BzHQJ4tvM596bCnZPOpfUP+zWce2qMEKJwNvJ3BI
/5Gc2gk8vNzuYOB0EM1HdAx1RROpTtgOXUs+LhfjCeQDnhTC0nCwSLB8UfvsrJXq44ZGlIbel0zP
9eiz+DzpxeVMb8ftG2ICOEVoQpHbuK/iDPBZ0GX3iPFEeXJF67QSMkPWxHjcz3qwOmQy89D4lVnL
B57LvLkNmo3xqpasm3JHHppfs1CAnnk/7M4tAwFBImuu3LVlsojKICR0itAExqS6m8BUp3xnlEam
oP3+tJZwCUvEM77uyg22TviMcUdJhxr4VHghfnFRdCtvCtbSjIquO8EOJF2Y1jJPJVbcy2GW00yN
6CJDResHTHJWZt9UCU/Co7csAYhJ6ulNrBIyqGQsQD3e+/ot8i/aq/NE15ycPvOqtQgYsWXx61+E
0QV2oeq4jzHrur29LqWQpQI2H0c4XWRTnti72RhhpyMRlkJHrx+KibuMqaMHojBViNrgAqn12/aH
oFDJJL6KEhDj7cz3ZIi5emQ+A+vGNgrs8v2FctdV/leDU47/WbnrmutSmTjohGjzNmvrpKJt3XJS
o8ISS0dW+AH+G9j5ohCICTpLix4w6J7suLapi+YCcRmalg5PmIZA1KTJcx8XLn+pwytf+2suyfGn
k22VzulrThLK+KPf0X8WRjZ5P6S5Ua/sDaFCiC8/CBRXZd5DcaqIFkNTy8FcRZwdRynt8lV8Cpa/
y7PYC9geK8BD/YgEZ0SyCWs6dusP+4sZLgYJfXtod1nAuyT7mdHEyp1R4usBZtULjtYgiB6pCSh4
jm5tUKezYn50vYZ1amRMBMHdwDW+Lv+htPjw5qSZvyAQ91DzgHlIQN7V44hpTdLkUxW8y/nfwHJW
08gLh3GOkejMkDnEPzBF7lloMabjZbeesndzW0x1l5dLgIeyy0bCc8Wyuj6c+OoYhlfR6bCCyhvA
QC3Cl7FZ1HJQGgJEFe4Beb+GNFDLhDVYdBDGqZwjJL+gkheAwHvC1Pjq+8Q7GqnS45TncIu89QcO
RtEg3ruSdYvY8qoojqc0+jEo08XESL6ZupDUnGdsD+sG+JKsiRUgbbEAKuKNU5eY3xNjNhK8SbVn
/2l3qyMH1CT/hR/xlDucYXbAJT+syiLXYjskBhUnL3GzgfyT+8KljKMR96+AjAaV6JDzrpaBWfa+
6yT2at09arZMlFH/AoiYrIASGnykfaX1T5wo7UdjCZKIxBRjFy8hWcnVMngYOV9q6YT21I5qC26P
WfvljypcJCUkVOhHc2ZJQaBSaF+NXpB5304O/lJ3kos4Q9QI7Yd1i5edM4cxCGX6DjM/0wb4n6kB
s8UrT8AQtW/cLpRy4V9rrI7WYOgb9zjBJimAhqCsaN/VYBtkNSO1OBzRvWIJJaLo2fKfJCCkd9ow
jxcMrlLm+Fg8ll2OOeE6Zc6ZUwhsDRXyaT0aR3BdJT/z1Aia0N58svBk2ywMoZh4KGwui3hPKFP9
ezHLHQtQXNhNJbfvNGSGohwSrKlD2fUXJF/t89l/wF23o+52dx9ZoRySv+AUEbqAgIK17rooLbrb
fClZmVUinM4mc+Vm4ffTtG96BRU9QTLWpXpf4gsqNcpBeP0e+SQq+fPx9iCLGGufnWoDAvh1qTb3
FQPlNcUdADu23sM/hmdTKog86jQ/1n21lKuiLMWG6qZ6rOcKOS2IHoBFOzhsSGXg3B7I/azMQM1B
2eKvEQS8wpKon0cLzIyEDMQSObFUAo8jQvK40jjbrhzG3YUuXGnffz3FXuolDhD9dgFOMEfI3P+g
iKcvB0AagJ3s9GFMr1hdpwwBZo5DabzCwsv294JfDQZDKjaVb+MxcwOTcOOVZsqyzsV9NuS6pKdU
ykhqAMFQnlgbplnBLW/NxPuDYPNhkObCMEn+ncYeG+9Dl4TxUmlHNx8NiTsQFLQ0NHSSog9upk7S
0kGDNGGIleGdORuOQckCsJklSfOcMuqJKlSAfDhw2FqR9AsTH7hRFeo9Y/7akWGbZxYNuQzOse1p
DIfClAsFwJtx8v0R/th9zsF9A8K1j6jsYoTnJY5wXTdkcdUI2DqEvkxrS+nY5Bh0boZnxHQVIuHz
269C/m7vcm79nddHNll6tBIKoJMM9l8ZLc+7OsaKmTTaw8Z4GvkF1BLn5id94AmfXHSTKCGRPfqV
2kS4XuxzUI+S00XHbNkeqrcnbcEq9f2m0GUn+CW9cV2sIR7cS0V0FafQqvcJL4Iyee/2dng7r+8T
hbnEalH1tANsyS6YsRjhvZh/jKQqC5ZbPPgkvcvbHz6PqxCnU0/G4Qu7XNW8UgWxcu8Vk98wPCih
3b5CSj6mB6kacg2uMyVdAzkYhsbn83hKw4yNEixel+q7YeYyuBjwEhFRKA2e4PpwLZtoMuardrRa
ww1IHi0O7yJ4Td45J3yOnG7ey9NFsEu7FHJoM4I/vkLLCgR8hkpq6WZrVB6nZ1hDVyZttQr6fdXp
REQpB6ewSbQmk5lKl3ex2sPfRDHwTQUOE0flkqGaAnVTQk6Fcenvhn+E4+Blg9XMJPI7o7JaKKgG
zefhzwGOn+eVajE+8Fi5tg9W4x3ckJuSURi4jKHpLi6Ee3ivEGnpUCvEAMGDHL4mN73iP6+qkBpT
blaphjEGgcNEQy2P3/WaxvWLxHYupWeOANCcYbE7Ar9nv5NzGZvd1lbpCKOqPWsUD0Thj/G6We99
qUQ0iT0BhLS4WsSGX7/8I/1jKFOfotwIxWGVJ2vWPUkI8x/Rr8IkqKkkgjraMBTOh3GflsRpmjOo
iSqv5F2ttRmasmg7ID59M2JPgdPhEZ3EsZAVRnfzsmK9hZ4PK9JMAvtqCIh5DXxaJQB2/A+pWQmy
VMWwYsYp5+me62Vpjp7oJa549S0lg93pwOn43V1JnEGwx6xwjN9dbi0nADwf0Ob1ipqU/isUt968
AT1fewbV/GEBgU1Yhv9cGbjNDvtJ0pN59ygn5T6NAPHSjx8/ww5rT3CNUGxiGo8JE3MSj9hGYxij
V8sySjxcN+TDRbA7ex9xUnGC5H/D7YiSWlWYdJp76inKd84Onu5qDntJAytvEGz+3GsmDKNh5yhV
eaepQnLsIMu76XzjbTFqr6sH6UxOkZVsv0GXXq1RIr3KPG8rOuZCBdQ3h0YXsLwjxYVsZk8YjUQ7
aFiFImH2oPz4XD08i55iOYzIWXgPQ8doCO3RAYk/UjCHRRHZV9Efbah47ukFJbW5ORJTAC1pYWTi
38d/oxp2qCWdVpzLXct74FJa/k842e5I6khXgwF/75i+CYFw82ikQnBSM8I9eRdBwdW23N5Nj3m+
7TDS7xv1237KwtnjIxpNTjl1S2Y/YIO+RtCnMruZh2zYGLKCgI+QS+GcuE0PHIfPtV1N/kYj1e0s
u2Y4Z39MWvx+x3Kzb5hksBmGngHV+riJhm8Yfj3o28dfeGu0loEyU2yXRLL/vCjKNGBNzD2o+yfk
YE5yQxZc8lr1vC1mFpYW/Mo/0lWjLqvWbnaJOB9QvOv96igZgUrnlKSAJY8s+p9aE0yHAnUa0Knz
wdv4EEAy+/QLePOaJZreGPJL41FoK8BVl4g/RUc+bdJGZUw6Y66G9685mPKeEaE5QSnrCYdFzCpS
rZ+AcdHsvv6qXj1CkiSzj7K4dVt1sjX75Y/88UyDNkRgCVgBqWtm+vfl9grreXgXZa8Jk99ZrXMg
TQaJQYYDIfccnI0sEu4kc/1thKxbLGfCY5Xs53EuPk2ljQ+OuuRPMjdfg56D36/GN30LLH+INmyV
Pj7iJFv3a6eLFT228UTY94jUt/Q1dhhMJnPKu7HdsyTqOY+6e1aVOmbWSAAViTiMFW2Qmq/F/PFU
19aXHWS8ky7FJY1TqFklDxKSqjxUXEumSuBcvyk+fagn4XX6AhKAhZDP5u/Eh/miQxR1YwEv9s16
pANTXuCgDwQz2wFLqBUR2snoG2OioVu6Gzuk7i6OQPw1zykIkIO3Oro3ZanTD17smB9kPEPw+A8z
EDL5ZPy+8768re1fiQzB4j1J3G9CkthSRy3ZvCugj4D5Qfr6kUb2sqIobSZ1ufvUhpvKq8gl7Tj4
eUBy9/tOSvEhsMECeC/+nqPGqImNXDdi5MJgSDDEAE2UqMuR4EKk5LF/ynQHEEORIsQJCp2GmPEw
zZa6mR8sPwJA7kQWjmYSKOtwR280Is45Rbxx3xwfhOUxLl01KxSRwA5rQ0unAlOP53TiNS8J7Hgr
M68GlmAEi7WSMU8QLMUATYsrvH7u0IRhe/1oGUDq4E2k4DKnQsbUAFAHTLzUHeLg2VUPwACh3PWI
OT9XRAY8K+9Z/MVjG9QbOJ0yD2jgMEmrn+KswGUOrgkMLKUy15dlZjmqVQnc6TPvEkJTlxKdUE6R
YhozNphC13xrCCA9fF2+RjGlbucr9nv9vm5BSRIyIKjgvQdW7pt31j6VFcERZe/8xAfm1n3z01kq
UUeQJwDtj5Q4xZ5VKrN/eg4nSZLdVrnEslkd0qBelY+aeJ21z2AfEkXGTu4WbXYFPwSDbVBCmRmO
jo2zviRkvtEPKHh4xm1+SmR9pfkzjpSeSo9R5J4w/FA/SE4g/GF3En5tRESR8yOIgUk0x8O36IXP
8oKRJJ4E/j9jhTcYSFlkCxJWsORA/Awjxo4jWvEkq3yTYd/8z8RD5Jn83TyAQKioxdDcf+nb9P66
DTPsAnDY9Vx7FZzuTiKSHhYlGc1meVMTa0F8ahJ19pSbmuQ4WTGil/BE5Haq7VDwRqa/m3B6cUwC
+kv61050Y1T7oF4wC4lMZjF7NwVPBMnDe9wMveEOvQFXpXOgpZDYJG79v1RaeFfYnHTptoUMS2iB
2SfbRSVDG/wbQpddW4Ov3ConaOmknaDP1JLgQ4p7he8pzf9/W/U2age7TQj/2rA/QuRAlaWQ4Esh
GE2eOrYEIg1f0KfV0S52Bs4Y77vxOvlz1KQrJFceCk5zKejyRWHDppyrQ6qF1g+gGXklqxEkCMpi
kwrnoW2U9gYz2rC+DJgQjxRLnFZ84OM4UwZgVdw2Yk2DRKApT7k43PmQT/n0NcyiqniPUmwDfU5g
Z2yavxORyTkSQtA0VsCaGOK5a+hH9uj6F7PuG4Jm4wek4Bqe00RcYncFLTN1YUmhfJ39ZYc0UxsN
KGT9Sk1+donYWxb9bjz11VfXV3TULd1pzj+AKuZBqeCubyyTYd1TmliLceQWD6bVVz9RJqR1WT5g
rnwMrX1uJDWE2CGDuWWHV86XWo301m46+5LmuAbELi49ksG+VB+nd4II0EdQ+Ih+BvUGXwDCtDCw
aCVWvuobM4x8DQb3R5fa7OVL0HTIiSlNPNFn6MoqXMudvkS4RGMZ3WpDIOF8JDUMBCxJC3VUXxJP
5/tieue9T39WsNRjVr4iYgmVXbXentkdktze1+Ys42CpKvDNc00LAP2X0kXtrgo3eDe5v7dzwTCH
pCReLlJRFoheqlQbJQY1NZDTdLv7vVO7ZN2gQFodKrj2/ytOj8zk4uIgijQYNtmQ/McFDDj8V2Bw
ZoGn93nqV1WbyFfW1Fjv+AVjCcfYaW/+8kOr5aG3pzoEtwVstfajtuQ/LglOgMoql/AKroYDqjho
/jnqkXiTx89h7bYCeDRV2L9/+pnhODfXY+n6jUZsqD6Q3/JMoT852XbxA4Ir1U+Kwla4aycyjDEg
y5l/4hF2stha3A3sTrmwPYJq/CuvHdXVQCl8DeqwR2mTZgzC0p89tfAILS5b4GJ/oxVBDu1LCXLS
J6muur2ejtBFjQBdrRuHYAHi+jAYFq5WSPCmMStw2p6v2MGOR9wJYToQKJmpm7PTPLFDsnm2/8rf
eJQ8WZ463G90LdTcNzfpaS5TiqX/U+uWc1G0InkDe52e+34kZZjCGALYLTbM/W/eEwxbuJyuf9vx
ziU4+cIjnse6BTi87hF8FzaN2ezyOJwo7MB2Zb2OBeQEM2T/QTf5EbEw/gF2o3xIRyKe4tqmlsGn
mfwRDvZqI2pyMR3uyW2DGOwQgS8OcGEqQi8QFcKC0BO1LEqQOGs6SjhtPqoJU7oebTPAGYM+OmPq
zrxRCShphXCmpM5M1TVgMZHiQLlqmwn0H5nep78JGU7oN37X+KpGhQdE/gf3QCEic+ClCzAs5v4W
itaEHfZw0PVpLbPpgTC7f/qFh1Al77gDd7YsbRHxu0qTcM7RI1SCdlZLx68tRDlwuXmIGsX1/GIg
EiezRKQ8cfe37VK5Qv2/FUtPif4uhPejNvRLDO27hjg9/3EBRwyuoaeyq1wzSBWGIHnqcqRn1TKe
wK/lBNvXw9dhdfqrRiwvmJV+L3c5aPHKRqJ7yTrscsT9iVm5yymOmUHlQxDc3VJyBpT3cjY/Y48I
mrtb9Aii1bvDtJfdV/g8WKAT7dT5GXFb+e8QACwOHz1idAd4lkED3dirwvjp9ElfpPwVEiPDN40E
0IZtYPlCZzONu8fzroJ2hBYKc2BbukJwXCO9Tui0wXKPTOJRtXCrfzOZr29uCgWy6a5g6E4ZsQdu
cVBULoTzHyTlNwqXpvc+3ackSpWdY6baEDs4Oh+tjlqd9Rs7ZP9DDmXaY0ySIxEVpcUu+558rWbp
rVr62gSgdi3Exv0HCvkIU/ZOaDsGPIXtq4PNlbDxAn/25iVv74zaoakJ5x+qILh372GXxhJuN2F6
ISRVf/jSlj4nLIYEJZtDRIGF+gBnqohH4yl+jjQi39/htNtuHJaQ2N9b2aS+qkekr3ADgdLIleW0
9ho97YLRxU7FkmkF9wzA7l2shhd630fBgxyAE37kSgbjCRkSA9f30HVYhwl/g2JOLSFDXuK0BLFY
DJl8cECl9q0pJ3/lTmzkWiNOMoLvjkkzUfil4gM45PowsdlHRPrfe/vmx9h5e1as8/eTSVKsTEZy
yMwAOIXvW6DuVvMQDoJc+CUXR0BWbeyq3uYrx6bQf7+CiQ7uzyXrMlKoqhLGuUCdIi5Wyq61jpqs
AUSOPwBQN8MV2qKidHU2RPXrgkO2uDRYRTlpzQ2n7VJ66Vcp+NAc2mJEuiH82z3AiVoMtW+3dnv1
uttPHNF/F8Wg+68cDRg52NF8Z9VM2k2Jw2rODSbXzuiPJ3JSmd5rZrNKGACEFp4+ch3433q4qfgU
OqqspQlFe+1FVzzus/L+jvoH4O/JxQuEiKCuXIAqzIUbv5GrfeyW54jqKHzimnqkDAKRfQsJ83+y
yJHReTOJz8eFy8iwDF5XQvoXT7u6AvQEs7ZonXH4Jaal85XHn500quiqeewdoqgOPRE6VWyBhRGS
Jz/T+7aI7JX2peK8wTYt7ccQAtdOsC3BIvl8aGOIQr2nImO1Nae+5l+g0Hlj1+/U7WWYk7q64s1i
ShOxMLK39Sw2AzOvJ+4Y+jhtp0V6PIVdySj6s3OY/Mkxi9JypMUTzF2lDbzci7qHCsoEMHGC3w6G
CZcSYEuF5RqxS0eG53nOYvpYxkmbdmTYr99uKnrVE/sbwh8FrAGPgL8udFVObi1/+W1DJJhzUq+C
SfQah0NnzzNDgio7bJmS52lnF6pGpLlMFHMdDGOuqjREmk0pMsvaBlgrnUnzX+F+wuVB8g92usfN
YW2MfExh8rJXsikENqlgcoalR2HKLms2OCY/M272fpxXEBtElui+4i6cj6nWhEcQMzW+bf8bqHzD
rzTCgQ92cTEVTFIFgS5EXVORbWUIeMfeE/9g9MsOJyHv3AeDCJ2U/9xxFWlCG7At5irD+VAht6uI
dFldAcuEx5xwjFIZ5Y4PgfjaWMA3UsWV3oWh+C89u+4S+3ra8fSDvqEZ4eGVj1EDWURPDlyuc5mN
fl8KlZHJabyptIswdYfobsNJy3SYBNd0cWOp+Ux3V1afU+OPtbZxx0yWl/0baiDCcvFj95bs4HM6
qQsL6uF4mNSZGhVZZpVuY90RfgTPOl8t+1QwF/TULs4zoLBjC0DkYkrQtAQclW6TMm9UIrFwdHif
s0UZNtZvFisk/GlqFkJ6kTsGGcaesk8+eaYDUErfDgVJQGoGPIHddnX0/uDWCQqAVWXXa90fyaTm
+ciBgszrosx/Eha8uutp3cTJNMEmoxgABJ83Hn6G5eAPi2EAg5xnD6unoBlp89GUB8BWGoJF/ZHD
mgJuEZL4U8W9ti0wTM4Mz+4Cs/KsZ8IDBvuFoBMarR5oe0WDq7XoPmZbPg40SJpYwD67cy08sjxp
htY/ZZRRR47hwD89sDsSyIJK6lwy18r5xUEOaz49Mlyn/HAkGV5ZNLhpjcQ4+HfBshjqtZaDNOJR
lfDjwWW5rsec4q235nNmS+gAe2ZXsrH/HiLqcu3elabDTgGkoFE7st4nMKPDJ8koR1r3evwjWzcL
33unBR64Du9xgmz3rx1AAM12g1/8yeqLM0IsWa7SY32WoWZxTnCPLMNP4DNj2TNE5GPO7Egzt+kp
7dd3dx7FsVg+MjqwBqdgG25W0FtxJe3hYwkcFU+uS9ljTesAPAafJMH3WC79IKIuNKEWEvxGP2W4
vBghL4ddg7/1VXCpXle3KuLTOlPf8exE31HxsqBI4Xl5vGsFhsEDI/xCkRARCbWI79+tjcU6+sH7
7JqXpwTZF77oGZyXd0fuuaqwNiAX9IP56xwmIfLYgYwcXxHqXqXvr+Zd63oOX077OhwKRpee3UKB
WNljovKXBkQdCW4MCHgb4vm0ZBA/z8FrT/g4ThMGdIc0XXV7dN+Gb+VqDjn/PSMfU7PyIprgN3+Q
JSAMISbGd4KeJpL+HTwhFlS46IQR1AEZ53AgVjq0gNszNXLZqyqpaaL0kssVeHvfjYRVB4B2jziT
9kBghnM/91yjZKUaJZD9W2rToQQy4+GQZADvFEe8RDxyAItB/ZdzHDlut7QGyqnq+25+mSGF1RsU
ldX2QDekoRUYwR9qnZfE5ZMod0ePhStfAhDpVwGoa3KAEDBw9O+zTVsOoy20Yjn8OG4sNO/VYsKJ
Of0qzB0K7TMoPzgQxErHJSyHkTqDQse96lwaS3nquD2Su5oeSgkk2j0PHAW2kmJhjFvj7VjGdZEr
MzY27S5jn19LNuqLS+nE1qQ4n60LOA1D9Zq1UZSVLrd65h2/rv3l641zHdptjYLAz5ztMl9yKyjc
Byh1fA0JG4vCF1YxSo+aBN5sfVvDUEOmNS7PMDfWebb2CU9AGWOT+ZUm201QsR8ShtK3cixb0ojh
EmL09dfEA9U/+lIK6/5l4q73pRCcE6h6w2cDhiYaQWPqW/SSOt6TZOsMNHRNvPbGX6OWx2oR1ElN
QuOiDcVzxpiCbUsmaptN3U3dqh4od2f3y+dk+m6g1cFIe+3qo0sZpu671fMSlvoMxbn5Hb1w4X+/
K1uqUaJCz1xL8H9gB0MtL5XjEosh3+pDxT3XuApNQwwkKQrA/cn2EJyBW6oGq83ACxiGoAQqCN8O
1/MamW+I2hwWgUfkJ+RCnZNt5F3DYFlmmSyimfAnJ2LZ6Ib7s5nqns0qqJy0i05eWO07V01j+x0R
zxy3oAv/RwurjY+9gTM9eExfogkxkdfb38yTD0Zrb9J2HgoZtctOvjIp1j6H+GCcsJgW7LEEfgXS
x/5YzKIwitRyMWubMKANJneU8FU7MMlCEgL1qBFUgmLjWKLzrT1NH8Obs1EI+3/+PrQ6qD/JOFmk
R0VpJUtjJjUX/KJpTR9xiHNaeVOAf1gAKya1MyLidpUIxN33ICDAZBFmOdS7c7829pbPuMxoY1Jw
h07DiSa/D0to+swsIZsjdReF6SAe+2bs37CNtbfItnLfoyuLkuXRPPb/nnRvMHb/xwERPBRrXYPr
cQNrRAbINYgW5DliTamuNClM3pFak8IDxsGs72DjeagxxSK2gLbfOspLgQbIQ5J8+mm7hwxlIi0a
layeprgECa3AdE6eQcV4cVfKRWelJora8rdDd2VnvYzwownV8E6B7fWMutkvbBOHEHSDc1luj+y4
0Fpmd1JBwBAkNsEc1fpTHuthgs7V/y++7Cw5zFxjk9ATc5k0y/53SIbf0ZbpzlmXTqImKsTiCyeZ
JALm8V7wn1iHhuy4J3msEweB13lnkjJLVLtTCDL4kKsDRhXFJMgWcl0CKoUgpC3oeFZJ+hR016z/
5BnwrSxtY1iqXkCoSlI3GrZ7aAZfG2zZTMX6EwCgQT/zGpZucRgf3ZhhQW0DbtVIDBvcjdyrJJJv
5NTpgsPN+3XGQ44G/XwiNqdixFdfg94JwO+U011ntOVlGNTr0u1sfOjrM2899dnKnssACbtrbl38
w3sxMKg3Lm5CFp4IdtZN0FHKn2KCeSbK2KeBaT1WXdlLMKCQAWethQ+8x6FT8aI+hoKvLKHsJw7e
P4NaCemFo7nt1g9UL+EDED1h6gqIjHdtwDaRovlkLUgclDTZNNfX9wapG2CPeCn8PTJyfg9xJFPy
kKVL2qGfsm7BAtELgCp9StjlAw/SFimUngY8SpzAI/W6Xiinzdt4xhrDVBpFzZ/mKLErAQmtmYwx
+0rC3Hll4FQTG1XKlBGlhOYAip6hWINP9atzZotkHEfuPW601R4I0kqMTvOBo4yIESPdOQlHV2nL
r6zKfir0j6+nOFtBsoPhav3COQVvOwHuE8+jtDHPKdI75dFJ6PftysECObJqI5bKKNqXehb9FQam
H+8RaCdqj8EADHVKeAzSIRSsdIurIDv/ySx7bs4sLDdm5BiwDKXhppwXmfGWOCugv3Xh7z5mf60a
Euaeqlp5cZ02Fm3wH5iRBNPKb0uYkwJV/J9PHQz8fGsHTLuwCF4/sbY1jmUgQ977Qdcy1fYvLX3H
2W/jvP0/wmcQfwjNfl6eMTVS2fUthDaN/ljhgqlSO1DaVfPSazz5Esl8HhH2WEVspApCYxgOi6GR
GY0MHY2CxERJKswiHPgWIKXoRd400imBTvCKZ6wZMXuC36Ki6MoO9TA1VEbDOmR3ms2PiYWGvqJR
P6mYRjvaoaFa2xBRT/ErgK3B1VVDHRzmpTpiXPQ0H8uXafjmpXtDUyGenvQ37Sftd2QeIj9EG9oO
U2Eq6yZ63WGgn+HJn8+MBSRFG0OganuqC3xVF0ht3zaU5++c6Phv3ajOuoycPPeCGYpiKtTNa6rQ
ZblItILTDEtY9XUtVkvrl+YqApIftCBbt0V/47w7y35ZRAEg8sHxaYjkChZHBV+HBES36bcUzzGS
YUJ46DeQKS/pPui7piK/0Ph3zNKou1KgjxZHxWbGEuOjIQ/E2R4LLfcYyYA+KZTMlo4qrAFM1pDR
e5dDgNDu33c4S60YAdEtNz3ZXafafgtDDSxCpAKJrXRIsIZo33TuAZOK9webd0uMT7YZY9LUPkLT
SW+wwj+/oJ3oM925pspq0yobV7RBSa3WuQcgVLNJvWjfoHQVWTBN3MZpPdKbwrM9DIDyuP/hwoxp
zf41VvKzYX4NtF8vtZwjlZ6IDE83+bPDvoJSTV8H4xohuzcSP8v0hFW0h1NAR0CTjX1qW9K0PC28
0hzfmg0Xd33HWLQYxa1r5CqGXom5vqDlhSraI9CnjCHOVUyX/Aw+bdaM0n3qyQesNqmrVsIng2OF
n0ahEBzzDbDidIlOFA0FREQCZkboV9lT1AtCVBvbKE3BtopXfdIaGPWmKJBcDkIxCKcH5n12kv5V
hWCs4LNe5/FYO8F1exOBckQ+OyKUvU6Nc478v5gY1YMBVMgPIPFXP6tYQe3qozbBwBChG+srdaYU
YOmj747rKZDGvw+nWCA7lp6yHrbI0ZtuWkritofYexx4yCV+dFn6bb5GDPkKTinKN+SuX9fVGeaZ
+Av+eabVxipvaEBCyGM787OAYG1ldbE9273mqxyz+rqq/YB8GdUpKKMJk3VUFYpKtVLl2xYEsXLd
WPyqwn6yCY09kGBkqd4MfPHp+QL1hbaiFG6RDmHA6hlZNxG77XrdE/Le1j1LCKSw3K/mQRY7MVg1
4DWfqbAPxtVwFgyXMgCHqiqS24AJHdpDgakcGAvTsRd+5Y6LL78nSsfQ85MPHYglrXqbJgOgz2X5
bCSRNYLCEN2HrtthkWn0mMZf5qm5ckXPa2pCJapqboajpW4lAnKlEytI9L2esyudBJviGAnrg7e+
L1rd8bxAvuXyrDDJz4XdJ7HUTAkIej8VqCtvLu6ELkfv3TqwgyuIBv5DXP/H+CEyfdYb/2m5Tx1L
7t2BEaJJAjFoW0ECxy4EXuh1OR4qMV6ToE681y0zawNAb5N+cxgS9PGbSy4nWtGUX3gR0enkELM8
1qUNM7I/8cEOICcuY2WQXWogTVHDEu+N+wrPv0J6J8BZ7zcf/1KxrT3j2hJpjGr4+RmxGQMD3MMH
X5WfpASDif2fbacFn6fy/M7mBCeYlzNM/clo9zC19BGlNPQH/Luu+HgEPh7GO8mavkSsZMJ9/shW
rbiPgt7tCzZ4aCKJA5TVpAC0PBbBbMOkP/GjMYo9w4JM7kLWa8EMJEEMRqJvVAgbV9eBRnZES0s8
+cII3pUXddOlwWcElYzF74R+o5ie/8ytpL6wPdEgjtPRc1AsaQea1HNCUJCiGMz4TvOgkRVcvTZM
hHKoIz733TAU4OVOW/ZQMHnzEvEeHq1KZekmubq1lrEnECtqz9nQoaCfsNCdm7/KEVyo+xsb6lLU
5+ZC8ePhP2slazWMu8CT11RhTifCvY2AgWtOVbHvuhlQFbApt/Aj5X60R33bozZaL+16gAFTPB1D
myDpdwExSxYWTwHNJFqQYfZ5YmWnTQpWQYi9R2/bgjrXDYuqPADGJ4WKLU796y2OwX9I+rK04wKv
d0WKv/6PgXCSV15PhLgqwDPGHfSfnN/735t8shzlIIoWmSMLShExzTBGaSVDTNAOAdpSxslJajnz
m3Zp2fCJQDr1HGK5s+WVNBo9QJOGaLWJkw7rmfQmgxmPxdZp5IZlDZasSAIp3u0xUI9MWNZbNiX0
KiI+t4PsHCVt7h8eFCkhy45J9cn0qFeecQOl7XzHZNAjDXIHkpGlNJvSAONZjlJWyj1jU0pyuztb
EmVjaRscL6K39kyi37NNQ1g6R9f0HjowM3zE0ggM5Gnf4rAKR9Ww7/y2yErY+EQmtyIX/GK5k8kT
nHTslvKwVMgj4mbfuUzIuz8Oimadj66Ntx6mnuIgthHM1vsXK/jJNQjMefS4GYUDaHdRlILFyNTg
Pw5S3XtDv7iOq+7TyBiykjeFZ8JxIsAR/F8aDacIiO8By9PX8a3rsxfFgU7l73EGLGxaprx9KBOg
mZhr0QG6eMz5drNcXgcNFAvWd+LZwWYcWqOUJNSB9OJa1yUN1W9z/BqKC68wwSljMu7XAAW/OA7/
ipOsWQpTbLyhNpsVR3qHWHfAOY1vEgxZjkhet5Vv4n88VyY8MtpE3d6vj1aXSX7dFU5euVamKwrz
VkEeqbw+EEoCBeeRjZlmxlpDHh3JfMeA6MDcOIMCmYDgHMnpKVv5d/EA0S8uA++b7ltpa19PJZ79
jqxFG2/iKKlmqg3KjS76ajWQNnCuNx3wN6ATH/K8SAfjkpbrQxkq/Uzdfq63B+REo1iHYQyEXENW
Py9e9AztCiibR0ZZ5eD9OgN/r+hdjHfMKPVJZWrBytn92EPRL2C+fWhVfA8YZNKaRbeNCl5N06Dc
qcXOA+tgBesgkfnnOIjIc9TUQOw1FoqfPqX7Rp9hJuuWaRQCT5ImV3UaflCCyYaC3VG56hLYD/Pb
WC7BKSJqbQ/S0B80fDfukcKV62W7QY+9MFDI49ZysWwPktEIG2aQN8FzgNNjSA03mffVEcDu/XdW
1hFgLTg8IChUgOEwEfCQgpZFY2GShTWx9+QDQu/ygtw33PBmc8XIoAqr+jExcxbgG8nic3n5MOnb
QTKmNGpMTU83b0Z0dRHwjQDKyKjtZ0WuTHtriji7XQDh02yDwu2XCDY29Y2un6UGV7aMREcVd722
+vwURm5DwlDIUW4dnAKQ3B0m5bkXTBp9WK9GEDfutiphLvz3Z2Z4RvuLxAgk57ONG96KmP7+Jjc6
6TcQkw98mcAk7X+qbt5Bx++gp5nqhr8ARyVbL5yJK8IhqNKAAFHq3KPlSWqGOeeHl8zWmqQlv8wf
/H9i014ydlqO1ZCK+vFEPNCdYa17EA6RLTFXTPpb3NjzBKNH3eBLpvyDezTVnfiYEaXr4rIrLm1E
53Mmf2eIU6f0XNWPaMgPc8mXfDSgJRjFyuV+2kkwCd+6cUDjDuH7ZNt5WPOQZTwdq+VapTagoyGt
A1duIOorjSpNo6a5fxiYci1SRh984Xu3qGOPUikeLoV0FfX+VoqcLF97PtW9oHHbf4MwMhn3AvvR
yJo0kttRbKqwdcr+VrmysfOxsYOHn1jR470c0P3ZN80EnlvTgmd8lQ+VM+MrIK+s6oZEqZ7omPpv
s0R0K3n3dTfJIRsqkAIGi8xhuXOF2j4chtYVaBCwiNljKYJkwJ8KMwMiutGDrZ5uoPhIrhPCVHfr
AgoP+n7tjGb2qZMdUo1C6ppwHZkW+F1ekRvi4LQwma9R+6Ef/qvFqQFk0DN47zuZwTyb++7TbrAM
gRxJdog5clQmHpzNPSTvodnASm8tHIijxJGQKJH8w6x0RIg1h3YSHwi0oqW6/Iyz3tH6JmB3IMft
uteXKlmAY1OMRTqXpnbk6a/vMgcJIXzIgMs3Fl3lmVT0dNW7Eo1+9MwFZ9oenLYpOSgJyDh9R0j+
MLC41F7ql98xASNbvuNbBjZuiQkTztbT9/0+iI0FEXPhRLkAomgNLdamOSGEz5kR6AL6ih9myYpS
sKIfW12+h8qWA0ekbw1TxTW54U7ubgW9VUE9M4Bf4s2y8Frwy6k8oA+FJAziU0Elsw95DobgLQ+3
R4UZlQQ4z/vcEw1HKW+Bc1Xu4STA+2RKgGYZoMR9Enx3Ntb0n984pZkwGeHhdtt7RoaewIg/aae0
MtQhQVkekXMPd5cdjLNVdyr33zHkCTp2ZK12eEp26kI5tsOUpLhWJ060WmHPUrhPVRyxKMCtOjSZ
Gd+YvqbXq3xTM5N8MX2NFMqMH/t7UlrHApwYdEBhqAdSZ6JGQMhO52D8ZAhCdx97qbNbm9xa1SAc
KWJMmzoeEJM+3Pjs7hbn3GfofdvTQDpEQjo8wc/1pFAo/NWZMHlDF8N4dC6CnFe5GVxHqKY/dJaQ
sQLRB5ee5D0nLIXiVXPWjG/dmmXBYs1kHLclVGKzATEUCF7tuwjiGD8KMJrYUN5ej6nLld58DQHl
wZnxByedw1od0/mTSUxvVKfEOx4ODWn7+bisZzlNjHa5IZnBskCJOBE1xJyfLVaiERofHE/gQsZo
+ecudeRZRjGZzqQ/+hdoxWOG8wPePFLtFj/7iVM+hQ3CPLYZ+2bDMxfLL0iwYyvwA464JnvNc5n/
AUi1d2iQvhXvK4e4Jx6p4vulUuUns8eFSwO1o6+EM64DUR1/DPbLuEuFEdf/N4e+ARgaLLs4T88x
TpxS1TMz0sob3VKOa/LeqFfi3WuZo5NA8uaMjT7iG9SzGUgZ8xHM72S5SziHIC+QWgAdnOOi5Xgs
nyRRYKigpBghZRPaWkfOEmfk9Du7Kox34FNa6/6gutkgHZUpUnAx7uCscfgIbyrO0FlVoRLoFfZB
/01fFtJ/K15qJhAVlC2WrTUh7PCTs4jxUBrAM7UVJG6hedybqlErw2tzSYQFocXVsmTuroV3Lz/s
lflSRwagbNjuSxQaJ9DFcHJY9tiLPYhz1Q0j2NCGj/V+5KXp/ZRIOAsGykkmj1jA7IhLbJT1G1U4
6IoLbKgTajuBuU7Tc8hLLj9Xtcyr4ZohGkXi9of99oLjpUJLB4wNUbKFG/K0tvpJZ9qYkwKHRavO
ABn7dSTR2yKz4H6Bcj2mAIpISXbbRL8JHlt1nZqgPxdR8HqHQfiCieQCwT8/5Ho3s5bmYbiRdLDK
JEkX+iwLct/H7msoWywq6RRHemQm3nAK8i/Ztaah1lCUkbAVjZJEfpE1RNJ1easK1Twg0xuo9uPP
t54RRAgvXr4YMcqZ/WrxeRRi7mMxlDVX3q3PAtJMNsSv/+lqMhjkOcSCUEQOiefkOePeORPA+fDv
CGVWgeQ9wl2bQ4K1S/nTn0jnaJpFKwqXGnNv2uM0Emdv8qNun/btBcWjpYpQ6ddPdwZZxO0mF73b
P53hNMcggRi1ImGwov9GrSjXc8e15art1tMaHHy2xL6MiQvwJcmsz/vITPGvV8ywRFwFF7XXoVOi
QUxF49YXAZ3Fr56eBHToDbZmDJnmB7IiE3imWoFzBuGN4sDqH9/sXJNgCmJhr+u7NljkSwRQ4dMD
uYrKWU/eqHrSzk0C6iN1foF6rAS9mqeKL5OfsYZ9KcGIiUjldcDV3GCs/Nr2LNvk1l7jZfiYpS5d
bJmUoWLQPgYSTYhzhKxySG8NoSY57Sw40IefE1YW88w0rjudffIUFjL6yabqXOJJpeamSQwbc/hO
digl2u41C93trbruUGr/6skSJeX5yNVJ5quLAtvkRQXCCqzwx1e77kMJ8cijcQG+t8ZGfAbEeH11
yNv9PG9XesBNoy/ffV70jCB5XfexQBnx4/sbzX5GSuVawb9Wm+COWIRNHBn5r7sCmj92HTIvUzOt
yOgKbWv8UWb89r5Jq+RxUyCl6DK9SPAxWXqqbJ64hPGkHsRLW3DHVjkAfZKIqM/B01Zq5RLA952N
UvJMVMQg74Spr7kwJvnwrCkIk49rLU48VUo8N2YYVAf/MeZMg3IqoOZ8KOz6e4n+KDg7r6iNph6m
q1/mxJ0fdiS8tilJv04MNkOADJPxIHpUOzUgHJ0Umy8G60mMonXm0cER5ACLKojtnEO659pA6BT0
KY1U2Wix5zukljz/1DDsbShSSfybSPqWypNcrc1xAuoBpphUF99zNML9zihv7dccEoito2O+Wl5/
eeCv3HYzZJUMldPObqGh4DOgfkSrfxbIz/bwJvtDGi+oLiiEkz3sY8bHHY2SBa7nme9XCwVYJyic
HVTxI1J4p50wV8QF413r8wxNqdLr0/s153fy1tljVoAh1dtRMXaFT9w07sh9NGN9cf9R/Mxt1jLX
avTa4tSBDkTx8bi3vBWKqg3k0Z4cS+bavZ0Lrj3uvR2Rgkhk5uFa4EQu4Ipr5hR9dShR43G8Y6Uz
gcOizSxFzfi3C9zJUGc259vTkHqPy6uCNt9XXKDJo0tGNVzEqLJ4FP3UdyXKLQGJgvkDcCZpJyul
t5yu8uaIlpeGNIr1lrpAMmEGAVWFlVJk4fTY7eNAK4P/CX7yY5SuEiz2PvjS945RIoKsmZ6IagFz
fTcYOoU+uV3Qm0nZ7oKDGrjidLe01UO+GLF1ApEXRdcBoOxtZw7zrhlNPeyQzxtveakzKWresUs6
chk9ehKL/Mqb1UZmvQvQDo9VF5Ypsa3pV1AzTtr9PoT93l7xzLUJ8R5uwNZ2Nzm5jguhUdMvrujY
4tA56W6mZw4+8FfP7otFWel2sLz7lbJ6wd+XlpxMsvV/2IhP/mN4rNMR6Rf1m3RV3beEKNznGE0S
lB+hE1OP1S9RD8FP0o/1VsI18g8nr+fzH70S51V/NwdYTPODVDFq/92t20BRwEUXcO5QRLTdjaDB
b1Lqzaq+hRbhBS6DzvYji9OrGA8oMEYqb8QVjb40JJ4Lmee+wR2AnoUR5HZVB2yaTRwaMfl2QFYv
1mvOBl/hysu/20dYM+TpbZdHF+TYATrFD7GW+DNqi5tu1zlvxKSAVWJIYc80c+JvnEM+4HUGPTMG
/DSN2XhwB7aAlHFPfh2IEV9DX0QzqmuoCNRkzKWgCqu7watGhxdpXY04C524g5lGvTXpy/wfb/Y+
I/RzjjgQLF0PtNStkDQY3pEcpRk9NlY5AtBD0hZnF5Z27u2VPhqroNNabguRsOULJm150AcxE0r+
/W/xZ1y/aFJHsIlp9LIiT8hHJ9pZ0HawoIuWUt8kRLQOLq6Wv7rf0uV0/LnCVr51dKJGcMChdtRt
iZO75LLbey4sJNCpL7xwB/OprQtObIrKRYk4troR9C2vQqzBxSbBUvwfyXpsc00I8+mKeL4KW+zN
w3ege+d0EGhI8ZZqJjLnWsh/soQGpIyDp1bgOmee5U8gaufJW3x+AsLJg60qnp8D7jgOqXSS7+b6
Dfir0j43RZbDA1XvMdPCbBsMVrny80euPg1BDquoXH71SwI+t5Xaq2xRBmEJVvdV+kSLOqTjTHBE
LZBNAL76zWWqBBXm9PSJo8txaZfC2lvNtk0y53NjpC2ahHtd1XeJhUtmtruNNZ2FBIOBbE0svwzO
mzk+QWfS6QM0f4JdM2g4xgrBAhDKnenGuzM6YPS/9dkKPv3NYUB7FqIwLnG5HyrnjrhzDdJUynPf
3ODznSeHF+/Jt5NWFQMKo3i6CExr/TechziFcAWk8bZgQKQkUl4JOwCiC+0zcJpgaOHWQLEZik0a
9kje3dh6aLKGJG/zHp+J6jJQCc/ZaFsFfgxWJ8Cki9nJbYEO3o0au9i6b+tAF5UcH7mKg9Kbgt0k
BrBARV5KaOMtpPNZ+aBX9GBtlYj68kjhj9gFomcf6VeLzQYjW2DHYRzKG9b4uoI4oxVpHNCLbiGX
iXVXRXNAZUn6o0/5u2uoxpy/eSnn+GXpAspV/CX3II+OxdSbSGEoCKHy+iyTADw0hdPJeevSZy1H
sIM3RpJOqRZWzOQ3NU2Is44TGTb3NObTRSFCc+IxmE6L+3EOhzlJnYftFylLwEdRWpJUce9LsANF
tQSXa+1SQarapGTseKin8HPw7gOvO3f59KRH2UuKA/8rqriCwtqdU2LXhBx6kwhanjZOPhUMBBlR
poXEjS/hA2CAVXfj8K9r4JP449b1g9BpbwePCzPwwvAEPBtPQN5EgnqykSdTuXvZoqF5QItdvQRi
7UaOBFB72EorvyUHUxQIJs/56JxNz3pSdbm7m50BMfTcEdWg9yElPloSWUJYj1qxGbOGfxRDqE7N
fA4BZVd/GRbfMgq9FhhD4kPaAFZXuzfN7kkFBRV/vGBusdiisa37uYVtAcMFyoGtn/UXqaV2Re65
w4iSYo85mz1OQapeQmZ7vvjGtzP7UCEpPInoS71FZ4igT1YJ4qoskzb3KIF0tvLJ1sqfpC7HKLAU
V0Io9yp1+Dfdme2NjZ4FqPaNJ5qnIIOm3Jvm3r4/n70bP6zbqvt6tOx4ecN3/owv1lcqFW8zDwem
/T2Ptf7EfgIDU8cYk3lySeXTYFqKqDhKwF4RkrAp1DxGd8PUfjcXJqnMwMKoE+GoL42ami9qj3Cg
X0o+uSvCsnkWC/qVNNKyCMSGWrXV1okvA6VlWpMwWtsCrnCp1UyEXXSAX7u9i2iwVlYzae6YE9xX
GeQ6mBl8oaK7HsqnO9XNaI4K2oJ1qta/gCgRyzm+9rsB2MrcCmGiwTpZ52wDPkKAPfi8jp7qbtrf
T2QdN4FjVqpbifywQiYqweSTZGdyF79Cb+bXgJr81k8QmgoP2KEaYw/9NcVnx0BaKOmtPVmcaqrb
7XKiS8xZ2FnXXSGwnJhGMUt9qGiQnIgMDK2OPoAq9XazJiCeB+X/a6BHAKcajs+bbQODI923WdEV
FwfpQmvAhXBNPTXB4qqX+eIES9AZF1S31nM2GgTKxZbilzcozeQlUUf61bx1Z3S+KUlYU0nGixFh
uKhM7+zsjsh5jWbBXzgSz9AYcfh1YlWYNgmEm/1fNV2FC+v4SHRKJoCKsrX/DpqXTtUlHCPigGsL
5uRBU6xqh7xLjLU4mfBQwdDi2gQvOIjO26AMRrV7Bpj2nh8tCQSX8nzNtg5M3qoyeOOdOiNukx8j
6OZrFwev7H877xgarJtg20ei9CVZmr/vNUoBYd/nrhu6WZyKFPbh1rtmgclXyJUE0wJDEaT2JU9r
P1lyCyZLiVnfbWQ4kRTRNqvVurdN57bbBEAUhM3Xl6hWIOS/byTe7dYvU4J+xqWMmVWi36tgq6al
JFrsFjdMleAiSUKZCUbWnA0zwvXoyhbqBHXpTeHo7LpnAQzS5lx3sJcfvfu/PXSh2noYhcvLQH5h
EeZOoejLzHqlw8NecdPvJ9buIeSpcSrh7F9UZgWzIz9DkUGKwsllCnnuaKu49ppBo+JbZ/frpbpK
Pavn7JOTyHAZy7Kh/PKrvc5TlUSIcnWXLh0Xy0236VoCYFAAlGCzTGUeKHKeZBtNBBnKCZFFa9CA
PXVeNwA7gM7+7Jsxd2j02OUXeFvmns2sKEr5LF/8KMAtCYWhNcz1Z0zL32tMzfd3A2uMnEOpYqv5
Mp13c51ZzHcboGbrCYn3IVB97da089KRcMAac43nUEGYyN3bk6SdcZt3QvzyMWmjgpr6+5O2sES0
BFno+zzzrM5swHMHq7xK1b444kesZU258BIHvp/9IpOq4H0wJRfCP86f1GI6QNxuO9ocsn3En5tp
iV42HBr11v56dV1N1FBpSK8tLF6/dObPqkrB6VNVKGyFPmSUiM+qLMScDTXT0WqGttW5TwGuO1js
/7AHpg+Cldo91v/aIDYGNxYeK27IIJ1ZTl1RqmeED+ehc/Jy0k6DonqX7qHTqqPegtq8BB/3vNkf
sredVO5MoP3XNlejWgD7rJ3DFwArzn1ssbLVUFQPivZc5Q+SLWWIk1pRpVlRUVHPqilQoJjo88Ri
42/Td9jUjv+0VbhwrdtCeFgDpP0G4J7GXTQiabNr0tTC3TLh0Dl61qyQy8U7PX/cb8T/GTnDJcWH
jc5i/24L5F6cepijGAMQ6EY3yKhw5xVh6qp2iUimK92EvTphHuvynC2OO+24+LLCkVxgqrwDw+ur
deWVsz2/zHSqku8s9oNzulFRHuP0OKMKibDatJb7TGsQgKkBo6ZBxlH6tN6Iuk5soAU1/H+pL1Bg
lt3MbT90DUKAk0Zvve6t0SVDPvVik/4vLq+nUU0pcrpU4L1IEj4ixkEdkXtIqT05F3sLWuF7OG5P
Qie94b7vYZdXw5CKyxhTZPRRqDb9uSvUUd0ZXFzQBgEiXn88hh7Ve8tGjGScJgWhs17vkVV6Delx
ivkrA+l3hDOo4I3NQhvVHo+k7sZRdKTgAbb2vPMXbMXXvSmfJwfpFuR4vpApagEzIQp6k3WlKm2e
dIgLx/LOSOE4ZtYuzILCvurLEBYDg6rjj5BjoDk1XD1kX9hCo1h+SNyD6smDHpqaWA1JZIAR0Eh9
ZfBh9TTwAkLO6bBEleO1XH4H//uWasD9y+/wVJfGtr2936nVYV+vlpBEYkSFSGBuoFa+STZ9VFKE
d3NwU+ftC6ZiUiXoWDi4nDGeX7HpfF2gzCAsjgp7c835pLUJm8/qK6VjPdSRqDICXNMnZju/YqJW
go/HNe/2ZGpQweXsOyQE1GIbz4LB59n1T0FrFt0V35pjJFDK5E1Dx586+x75wmLHP6MM79RCWK5W
kpcDcN5dFvwHoisWJpJKsDEdHSfXU70p8B0z/JGxzRGQ4wYB3dDw+FLP4xvLjPsduDxWO1zUX3tn
J2GRPMMJqHceUrhkBTAhTwmr+V7yIOnyrNhnJrMVNxrGB5vcHIKQklqueCpMVWgPi6t8jzijTYRX
/RbDU7DTX4jNubI0I/yc6GpzLxmKRpRwjuUXTQuqdECRW7fJAkjmM09VYeYx0J2HDAhumAIGlGDo
6HuWjIAIH5fgiAZeE9K+IaQoqVEt38xEkAQ4LCJKro/j6evtBxqJZPHKCRFo9Hi1HJ2KHbFkC5Fz
t67RW2kT4l3yyj0AlTyEZ0542wa+L6ttGnNotUEXdeGcl7YLm7SNlp9uvFkOA8/N265TcYgQ8A++
FS0P8hTdEB6+8Tx2LDugSETGSgxc6vFc7RGqpr0kLogc5G0awilV4pmhq5kWbbNXwGyDoF5fJRBE
5k+HVoYl7SIpODwaJaCNP+7IqUMQ06fAncDcDmt+RCj2xwne+ju5S90DA1n0tHD5M5t92WWqeM6b
u0ktrFA8Nq0DP9IUioj0AvecPIXJQIGNfcNQSbmHzshMQytRov//hTZquSEZmzo5upPfucWZQQQW
GAJtqHNWyRGqkmSrcATI95UL+bde3p84zTk965oE8Y3368TwhLj9QnpfT5yKAI0VgtFVAQ18jv/R
yORLHId2QpORf6Vqqd+V70eDSqqlDGPa5SwYExBjE0DO3KPynfhzZIm19O3QS4MU6iVlzuHmBSsw
ufPaDKWoF0wiLJoJ7/5A3TpG7+lHYEaQTGNXWD8aexDYSwHbqjyBrQtR+8Ez3lhw2tS3QUkUf4EL
2xaG1Wui2tivf4MTumSqnktUjJpkb2dOkfGjxpqXpxHiHWXcmzINL76kBM1wJGqpG42UeZxyDblX
2zuTjWDCOBm4BudvF8nlUzRE3JMPV4C9+uC1anJL6REXKtQB2gt641gx8muWrIsfv0QW22jdj++R
7KIx1cXe0Ph82TrzB+1WGOnNOQOrShgbVvazPv94muby5WYqJorAF6nZ1EUSSwXK+TAW8AxUSyiU
N7m7eyHvk2wTaUJF6MGGecTLnlJAodLqVk4MHelOV3GXmG5NHyWUY7PD7sW9oceHQu9CsBadDCc3
+qYJ/IOltOBttloQfKWIzHMWBCzAD/yPP8j79s4lCJomr1Zs0K4XB5LC89JCp/sIsLTBUrfvDdsj
wwkbsEXr2Uh8jtUdZJfBPIpbLH9kaeEdk7+o8nLxsKGLoyxeFefHD1XNP8sNmLdM2zE7WORqdOst
30bbNytRuMkkVaMmOWEzQJtagzXPTzmIaojn8wFLZ8RADnr/iuhHDQ2czh93lop5TW4ULX/6oBks
iSZu9dYD+fYJj+dc8aw4GaCPz9TIOA6WQmnYEmTAoR2lXpOhqDGwQTUq2vHfVdR6vCTP1n+9SHgV
UlYFI9GD7vTU3egKZ7VnA+VMELFzU8COgGCirwlNoFeg+bj94aRlfESJIsRykwJFjB3EDgt4hsD7
YRpy8yls5d5oikTvQX+p0TALV6Ga1ef+GnlZb36sBAw554cVX2g6gV8YHLleId+8wxXuUfyW8I/d
suN8m/N0cpTTWbsvx8Es8eAllS5lNlZzK/ZUFWd3py2SmLKvbGfa+jpRuplr1AK9y84dImRHLKDP
vCTB6aB1qo4ah/rpQs4tVZ0LzkXw13hkw4gG9KpxCp5EdUmNUozukE8uva43TGgjb+akRN6dGa4c
AnBVgX1V59g2VzErxmAQswV3xUqzKijNI/gvzQx7aue9EExvjDFDyU7W6OnoJDOFAehOLrzHrhm9
FN17ZzW0n+9zjNjQpYpYAqexmDwfhTeBU0wLWKI/T4tWZN5g12KatRdL4BfaAqZL38jE31iafjgo
i8bGGstFj4orQSExomCPMJVSLBbo2YAZw3oxo1UT4M7u3excQtrxJPOI769PH+exaM0qt4+s+QdT
f1G5ZuvXSXD3gBo/G8XgfF3OXCObHXAepkXz1o03Lpl7xkAVoilzqWj+xdb3u2fyR1B3hyN1vwHx
x0d5SXTPC88SOc2+PStnFsrvHlGrpKvH54kOh0bf4WWKcyb4807LM+Bnz3tfl4QYm7OrboJcgWII
UzPCQh5C2MI7QsaASIoAc1LM/urWoAY6uD6Htk67WfEYCC5K1mVRjZvX/iXCwx6aO8GOuqS5UK5J
3u3576o7jAH1yoR0ZILdui2a+LcuGz/U2SAKDZbJ5x2NjZFnRXP7eyCsPZ5D0mddBnaRRcQVMiJ4
ebt6l3w9Qi3+PMmKidGDLzR1QpYAwmrR/Rmpoa8rV1RHO1OKbY3fhF2SBu/tu3EcBRLVDCObjwJC
mOUtypNRT57EiuE1g28VbZfX2XNmmTUtMbWP5XHpafIMipnfzK7yvpTzoQfp7VWqV9YPcogERt+n
k8VmhD9F+xKvUBpP4vjWdf2H8XdrVVJaSExT/9AHI2XPFYEHWjViDs2VhAOQKoZSMmGfEke30+Eo
XoUKyjDZmQfF0hBqetj12n6oHqLk+67BxzcMhYWRRy4fp5+DbVKXAnxgKSQdLgyw/t1UBl53RNrU
e5lWZoyHhOew3waEO1ynh43qZ63b27/f6RgN8+DumggJaG/KH5PdUQxXf5c0nNR3QdnyctXccudr
fsGFeyMayT3papoHTGqexlqrsOYZ2V1jZC0CAYvabFpUpuRC0ENS9byTRJoiFmCboGzFRKRWBXBS
0fa2n79VzMgKOD1JcBXnqb/QxaOuI97M0gPfyMERN10cdHqZILGDGYRaP3UkvfBRvxS5z8sr60PB
Tt7vd2fpsPiQo3e5V4c9rv4cDmK7OQ8Gd9Iqp1K60wNrx1le60w8CsmM6Gi5MdVEvV18QRA/z66c
lsZyeGD46U40E0hiy5kgHc0JdLlmHNIkFyRAKruQLIVEaXYTRplAK6QntHqAOsFiLwUnrWe7EsJa
gh1lJntJR9nurZx+GE/IcK3TDE+fxRbmeoVmqzco8O3LiEZ5qZrqd3WVy7HhciNZHQ4Ic1JwePpC
xitFEstRpw2i72sCS/eXdJEjepFSMLRvmZHj//AoOmWQKFiw0FZPpNXjlxlAhVUgQWMcdfY0/1mS
gBN49aOrzrMNq9c7voNkF/GtrMnNTtcr5TjCP/C63oPZGBfkZ2krgNh34QqB5pwZLE1vlFpZeI8l
/lGOh3/rRupOll11Q0w0T5+h181csadzsK1eUI/+nHcdGH9m/y4iawS3MRcYnPtU2IWH8yRe974X
P3valFO0HQTqkBLBC8SzhgtbAXmq9gPOOGnxDVReS7VDKN+Kaxs5EHY3wiPtVZQA9lOehWIcFPpI
lqukoQhj7drZVINDp11Pi1WNhijP2+8UiWAepRS6dpi14C71xdZjQhePDJg7Bw+s5sJk/AayNsO/
IIs/eNWYCsSyHRZ84rFLU7sGP7Ayi+Qidruoymq3O+MQ/aGhxczgYizyA9fuHkf3NRNSdgTL7gy9
tmyBcxhA2J9/b1qVUsj5eUDTTMtrJeaBaTr2MgjJIrVCUJh9DHZhQUCjgVMl6w23rCw4MvIywBsJ
6UU/E2Ku3/rm17YaE6TPF4U2r1sTd8iHa5vhGtpjcv8jvokdLIrX+zyj+Q9bmVTOJT7JctVBamqN
Ic3BH61dWImzOlwfrc1ISvH97Y9n/swCPFxueF+Qbfko5qQY+qLLwpz0IJaabCGJfCwFIr5IENSv
YKBVFI/zKFARGtwe3M0pJzCTNXR9HlMEbS5ZVG2Drw44BAP8h6tkAGkrc9QH+7oj6XPXnyW0vJVr
hyJThXb3GquGX5h/JOtqtYCBfAf8lOHJ+bwm7/iNw+yp2DRzPU2QtQY+8DwgOzDYwiZFkzRL7swl
JDLhR5aVqhLjVVqPzgeEGaAEcIq5I6DWYV4ihWGHoATiWNznyvYmKkjcDKU3Mv2/Bc7WRImrAgXg
2M3ixc756wRp1Wk9bzM24iAHLCZmTyouJJ2uohjUghoqq+S/5TKDORlaWOtnryWeNMC4x+jrNNk1
aNVr96QCzZidqSMyz+wA0LozSXqky4gTAkAZacFfFMM2K0F4esWxlKxQigXn9vNk8qqFwqQi9jY6
MYShAqEy3HYUTnKBpXUXgZBrySuoA+KC0XP2yS2MK/oBQQK/QMTKgI0coD62YsfRslBNq54jemLE
k800351ZiiJsfPMaH5btUloiGf9prq3ug/EvhmWlwoG2xNmUU2ABbMq5Lpc9z8akp481V4ca7hQk
g6XlZ7XNnbt3df7EGaeFqSIcY97f8byoKEfQTAc4um8v8DsDz3kTVlG1mgmBjkZe2vYxRoum1Eca
RQSGCU5b5aFgdW8ObwZd3a+yBi/MdhaUinrSBHOyq0Jtm0LN9ma/HuU1DfcY0OsUei3RQRgMSAbi
8zYdAZESXRGXyCkIcb7vwjh1JNhgjEDPDDdnXy6TRVSQhQ+AqqdFk+nZSWR0ZP/gkLpOkXtbMPNl
Nj//OPWqlyir5Ar+19kFAAQaUYOjzoucBLN93A6t+zOaVg4iJYSeFgNXedfpDWUx7Mm4dFAN4piL
iRDUv39RhQs4m87gTpu9BQ+XFHwOSfuZDGAbkQo1Gghd88AztJfDMXkPaiPI6viE+aJ/VKZPXh0F
a7TebGQREW8Eo8FPZvBFFQA/56vGfutz76ks1circh+u6pTJysUwIMktMkFvSpnxQlapsD1XUJbl
ashAPAYTorRgjHuJ59wZV2ezUt5Jyj0rmGzewsipXGg2zbSltk31BcZcu+/evEFKUJmHOFNiIjeX
JioaY88EAid0f9sG+lW1cfqAFJ/uO/JWL40xrISh/2OCxp7VcdnV/Ck78PtxGljbuWIRXw6TGAXU
Wo3BM9GP3GD3PHfJxGC4uBBRB+VCrkqnI0TNIfUJMqn5KAAaehVibRrTFxsLuesHL+c+TdYafp3k
rj10idUI1c29zceRg5xK4/ThnaI5CNBOTbw/WR1i27ax8XjDDLUAd9JohU36T9zn0DnPhxj4FHtB
fnwG/zikz2pP+sIdojLz+aKcrNMNJZS1ZMN852YXUSCHenworv0mOHbYOWcg96wzpXNC3uAyfLnh
stUv0dUtjc4UDgFx0QusYT4gwox//AF+x4e/49y62gVkuvpbMLzR6lDzRE1GxFgIQ90fegqlEu23
PL5auQ1VHLWx8hb2+B1Sn+UCSxjskq9ddd88OnTlOuz1aE/fK7irNlRvGYy4Cfea8psaX03Da9sC
qL9uHTIY0GbSdx8ceynQl1mWVB/jXujSLE6fgn1sfDmUD+tPEpenXNAaIIYoUMQ7gCMXM6nW80xq
FnAPh+dUkDeZQP2twXmEOW1GlwZSZOd7SfKOSv0VsC3K9IVZUUv/xSWu8cx8vtJrURagzkVPQ9cG
gtx2YUag4Pj1PAQR+5agx9KNZgQZBa9b2lxMrYifSEV+DYL6j9Oyu3R+5ZYaUrI2rjtruRbkqnPy
4alY3W1MiymdwDm+tUgyAUohRAN6DkPeMISfONNxk+v5yRMYa5Y/tctCCC+4RHB8G52oNYrkLg9f
fd0KqcAUnCXdLVvPAmiZQEJgm86yll5qFLRtcJsfjwOHSN/FLGqqh/RwhD5ELgzi3vAf5qu3wD2E
82AgVCwJZ5vLYn0xEt4TrkFWNUhhFQ4vkpVJW2wcdkRKDoHEGSDq4hw8LGceWywyRYAmZodZP7o7
Sryy8I+26O0/4zy6niiYpUNQeqayTUyO6g5e3/mcmWknYVUB75bpFcONdrfKMsK7+T5sDuCYNap0
po3EeLGLejc2PX8AHY5saOINef4M3gYRvo2uHCkFLhr5oeFs5QuC6BK0Pn4Xi1UZjyJLUKlalEko
RTRHrNaL0yU4YE4pnG4cDZbiHRB2gr1u7bohZd2qYAyhLpzD+ZGW4HNWLlEbgEn+Fwm4Q/yuSBTW
UHHjGsV87HWnI78BUHK/Gv1WAupb+SFYN9FMv0ki8KFd05tpf6ce25YLiOopXdgJZ4VuHCuBLPJz
Ih+vTUM4grn2dNZAX4DcLTQ4MD20kmxihCuiYOm2iUrBT2NK/zaZshg1c42xmCrhpoUYy/huz7Xa
IXLohVp5pxiviUdaLUi26CUC5DhtD2k8vM9fCrirpJbBSFiE6QJBK5HmaYzA6Sv5Sm6gWVkupIZg
cbIA3K6xKXRK+OIOoThEmHtOw405DS+Rb9erdU55OZg7jQ1WN89u652fxR4hVMFpBV/hj9In4HK+
DCssk6eLv70jiG4WnOm7bCtbMi/lyuIZ6jzO+mLosaJu3PcNV/pO2ZaUq6zlkeIzq1pvgisc34ko
Y+Ia1DQ3Hd7alXyBtXGTpsMiAyZ9h7R24I8a1q3dxivLYqK9hj2A6/fbLLErvMOOf/3TWZIxdjZe
42b7p99RD301vGKQ0O7KteC+a42QrZefcKGgOxEXlBiuTPMM+8tigR6nEi22OZe2kV3Ctw9BNONt
gj4YUyYOPSWAPm06Hf2lbpyOawQIivggfW79BbvTXkml7s83aFdU7ILVFVBfl4NKhhIQgsGXP88s
GiCJmpxKkXB6+u+M+sfqqHKQI3Pf0XOBNgI9H1dJyH7xtEx9kCVN0cmySx2fJxIllA2JZkj9gn2S
aGebXZecczqJp5nk3qpAGJ7ZZSELFLpGFnLMZ0YJXolP7dPcUN6s/Zt8bHxF8YEdxcnPPjevd+y0
RIO4ig9fAZLmp8NdeGKItnU3W0CSjGJwwRjDKOutG3SOlULIYtV/YO4FjPKqeA0/3rQdHDW7kNZQ
dUN2iPvTtj7vXIP9RttjKX6nzBZI7E2djWJYvBP4YkeOafpruxNO0GhvIozDqs27CAJE6rhUjGjZ
25G1HNseUXzC/AMsB3Y8ezii7Xt8BIH+giugOkc4lpcfh8f+bGyw0cym9J0bVV3cxlZCdIoDLjQN
ErAFmd33OafDRqXJSiKQLeKO6IUYty4EH86N7m+xBtHoA9MfZHNis56KLZV4p5l1OqIzuymOwCix
eQuyHCi9QOfKnyxm6/ncWyscD6AWC2Xx238KBFcAMVcQ1Yib23iKMdPj61VcTNhUuENXX8wED28/
e7gKwgNccNZF8jaKF7gQfl/y1/fbCSu8OJmx56fhoPwYKhF2396ZZA5bHdASq1zJWmdv1HEJlEMn
6obUoM6wXjggDwUINkaeXkj4dPy6TMam4QvTLrIPVHj8kFfGv+gMxoUR8a5tquULgsickK93mK4Q
9TZZMRbtizAvT4rte59YQ/6P0URldDkcfGj2Q4IaLjqTVPtzeE8g96HWBGQjAnjcxCC6ZeW60Npd
ME+7CHy8TcgDI9X3syfDUY3bzWfYSTezI9QS2Ax1NGX2O2Fq6lITJzMgObt4gF8EapOBo8iRfYdC
edc1sWXGSRZnScmX8hFCVVstZWNVhBeZAd5h5WlEZrh/Ha0T4/Wjcg05jS1xKie2KU5ByhH+GGWx
ODTwEh+zkERYchx4q5lAoNqFxrGpvpJe7L6vP+BrYSZ7mIv7KkAlV+MNCo3FE0LqDA7qNOnADX+3
FqFDzMkn/JBdUmBHILHA2jevvLwJfwTUW9TSV5jAy9qAw+nZ9snjZ7cMoRbtePR2L9nrjMUetLey
pTyfd2qtjVZMbmoDWI4Vm7Jlo6nDl5V7QOpSl6Juf/by2b8mI/q2O7bVTsm+dsBiPFnS9s6Da1ht
/AKm5sF1oQomVQFq+6U2qgZwxPY9MuSB69yWHDOuqbWhv6JCVTow5L8x257jbPapDC6CIGyrjfwN
ZhEUwPOfspc88JV9gltF87+98JyjQHru6m0r0vVzblmmc8jxqtUnbNwoYkp6j4uriRMKGI93lugv
SwCGsY4OT7fRKMbFke0XrLg4hqKsyNckOy/mqhvn+phabVZznLTKZxlNhe+lB3l+nA7uKC/FnGaD
Q/GAt8a31B3RJ7AODDLIvcZmXBKAmsdMu7n6OU2Dh1+ivMsL+FsCUmmCGRrG5Q8xV5k7H5xAYN1f
Dcc5EfnIyeqzp7pd0jrtk6yeyZYZXQ66p/sWltQVh4vTUZ53UXu4GfZGBjWjoWqIrHkkA7OKoaiK
/1HrpqiI03hrXC9XGR3DvwIgoRilQjm24RWzOEHCRmQwWO3KDwa9OqBrld3XmEhYpdXPzwfo7OVV
kxQHLdkRoXatb5W41aSRuMHULAkrlj3sIscYrrN5HV59QsPGz1hh2MWdlCiPfwuE4KrNLHo03NFC
8SVCvFUtHht4wuWARa3rE8o7USX18RCHWM0yoS6Ac/RZEvgLczusb8JkgwVVjMz3KW/Nt+ak6jKx
L/Kr5aMYi0l40gAL0sPY8YFVDOs83I8Y7BCxzSmzxtNt2m9fh4ydSciJEFdCeg8khho87LgnNUA3
Dbj2P3lG8G91tlxAmD0X2QUn8m4lBr1GtBf9WV6cXFXiJCU7xDBN7gXurU0/7iina+WFNOZMUiG5
z93fa6Y3Af6XUMyielhd7dDK8dgqKAXciWjGcm9Ih1eH46a3o0+XRuX/v6Ej8ykAURiPn7eRoLsy
RG1taAwLkAorejCndlRCU4t4x+f1Dj2zUiT9GGU+ITcWzGUI5jzAKOn7KpqFFDpxHU/PZZZ9ERw4
P/P6RYZhv2dqQ0EMyzGC2Iz8UAJclkKVZ9vdA8/3orLTiKmKAgLhS/6nVK1uzRsjqmoej8iPoDqq
iWQWoKSfGOp+i7mi4zAyvEjS+EDH+HedY3ahaHhKwb6m/rNhdEjjUpxvbNjKmLjjty7LCPmIYq4V
ikTV4fOPQRyzh4pb7tPVgq2o21H9FDO1djwzudS5y8ijlNA2w04zG1V8biLd+MonJSXTUkKTQWXC
knD9isxhFrier9jeqyACY3OMnpdH2Da8tfXPjuSIIe1ZfK5yU4SjmweX111qYw0q6QdSj1+voyDU
c58Q0YknjP0dWMyKsNMmEPK9bmFVi+x0hf4E10AZwkmnerr7H6c4uZNEwtjv5W5UFpfY9dR8clFu
rPI6ivw7VuXxChWk6ky8E6pePoT30oxxTmrDt2+A7rdCMYt3sDFruTIf+u5jQFHZlrzSGWFPjJ/4
3VieHSIw1RW1YEPIWBC9i8ODFHTdASM38xacBHLXB5gT6OcbWFYtS8zk2+qUB/JUQPBq1TnJlhaI
O2qg5LRHnXJMmTZQ82fQ6hJOtxx1zYGHbL8Q8BvWas28pQxmfDXmo+1GjBkTFFobRbXjM0NTYzUm
bYNPhLilQgqHpWAstjlea5IdLccnJA22Zrca6SkKe+X3fk/OlIKpzVhHl0D3cFW9TEt8HwaNaJ5K
C4azTG5uIay5QX14La+nffBi6OLEqotjkugQMI+bn2DT4Ims+UkqAmgdOjbiGnfIQFPiHsAHR8YN
Wps8Q0ygaKy6+9Xho9iZ2826U88HX++Dfh/m9vYdFnh4QRHrM8P+T3pLBWyT2wviDSzx7YRyODsN
JrD+8lhEbEHiyP+Hu5oRyDjgkx3qZ1bEaB608nlqk3SvQMf1xrta4w+l0X0kwVOErU0lVqJNn6gI
USqc8F8dfwqNoQq5dk5lslkcjCLxDZDdS1BZHCX4Fe6ss7keSCiUEbIgK705aD7rPELqm0E/6CGz
XM6MAT1vl+7SwlTM6YzVhFGILS09fX8wbvHDG0KSSRz2cOoJnu2dWIMGXSpMRhxCgt4VYhmDq3JM
EE5Vl2oOTVpwakaUgmMXHtFmZUuBwxajLRZV8Fo1NDKXoHS6NgFpSkEr4mPaUtluS9Intb4nEieS
s/9c0GsgrjuX86P9cxIKfB6K05/hG2Nj8jZnDGI4THBzsSLwP35lay24cM/MoQuMo8HnxlUInwtS
S7X8Ng+frrL+rbZL1VtWLmUhYGE1ev+vjUGbTIcU/eSEybA+Ktc3QPOdrWGIS4x1lx+SirhoFw0g
hv/0he8iaCxGbD3xO2JqPZC5g6EGTe48ATccUTWIbjhvZXcBEEq5QIR97Gb0FNmt6mSkKICQqqZP
aDhetzQnLI3tldz+drXOBCMaL3La8O9PHA5n3Wlgf0fAtAOEAL9I3S2KWm2Q5qJ4apyv8PBmeADN
xo+ah5UKoe70AvZTkfgXUISeD3Rkr8TRr7u8KHISlUNCC8iDwJg0iNhGP80xTDx69ZvlfTy1dKO1
RNQtNdsSe03LCsp4PNejJmtU/P3azAK7Djjiah10MH9rn1rKErdWlmo3AJLehJRzieJBMXSnNpWJ
ysi9QzCCh1w7XmAa9EumvGvZSgzXU5ot7Y1Shw6cVfZe5DP9kZij5ZDh8zl73p93M8oHf4H14tCZ
oyKK0OqquWmRFHzo9CscucGLlzhpsy9y5io/Sh3aCfOtxDQPyUJRFCIZ/asOLuBZvBo32RKMlsgr
cTiWi89vBoOtmdAMh8nuUepIlFaCKpsNJbe9W9nKU6CE5WbwPIrYkBVZCW3TqYSS0DZ64nbzwWaf
j9Ts1fMmgdWduFlivkGo3Ea4k+2qC4etkoqQSgBb/SrpBrqXM28UkiGRQKbQHFH9Zh7MwB7UmNFH
ToFoyDc2LYt2mZBL/DS3lwK2InCDgJi6Mo8XdWGD+NNA6kIH3CppZjR2fTlDirLggSZi95Q4vCR3
Wzq6/JJ4P+ggeB60UjD5lLARJMFc77c+jldBz6hqxprfSHaYJaYb1Uawmj68nKpOR2/CpJWYpNgi
AMQeWoDAKai1y8W0sDR/rUbGAcimFqeTNsLT6m1TVYpI8yKVz49dv3EOXMArgR/S1SSgP6N+AJj0
NG79e5hZDKJ2EW4WsAjb9K/u9tGIU4ETfAyLvO6FdsYrXO7m94934bq2ilUS2IidnwdYqvcmwRfD
bSKC8Tl1F9MplqOZygXLSHxgCWzo8ejCKa8OxaFcy4auXjvjkEF6Vpm4sMB5WY4wve5FstbmghUK
73CFgbCsvPcuCCw8NR/ZIvMiIWr7HCTq5WyLIqrDdDDT4n6o8QbBTsSfqwi543zub0LnNLQFu3BE
6hGYLHWKisgyFN8KqZMz49O5NW3yTf7GMC7n3fh2/Tpe5zuvv8TmmG/6nhiVCOt0miyNQcBFoSXf
swLcUs3HP0xthQABDBUY+jggYh9TbdBRJ9cDnfTx8zwNkzzlc8HQxA7DMMgBkk8MChAxGwdkf7Fx
Zn3dS9TOYipqxglLMHLS1Fg3kpBxS65XRqr6L7e0X5pVI/WrUJwFZN574QSLOFbmMfWYhe/y0BjG
W+daURKi9+4p1gyUW4zsMi/Jvp5N+bDbeHK1drg0bm+L9f7Q0ney3ft9KBleHn8X6o9C7nuiaV5R
Q7D9JtYvXtPBXZ9sgM2nmzDhw7EeFltD7jXdG80iUh1NagZYvrcT2XNxYh1Y0Sy5X146vUuyfjfx
sUc3VoWVoJSX1GJTn1uMpjdSsLE/9DDeC/SRewyW5H34Mj7AyYPWJo5mx91OUpyu3N2KsuSOtDee
wtMwx3Fr8IZF2AK/yLhoMCq4DWFkIIkfswArQqu4wU8Y5ET3CKY3uVFH/BANS+RGQiM7/mrCLyPp
y0c2MrDSA9dHvBwZRpb0sYD+gNiKQd3JRXwM3zQL8GDOPaP07oXmoGtV1k9E9rowdm5qV7V1nS/p
LIp6oio4+ZXRGvn3mXdW4zgyivJ1q6WOGuU3GgTAsHrGMyuv1jgDuhZfQ8QfTd3cv/M4P339ku2f
MF4LaRmAMSa6pKRCmw6gtfSY3QbNCeYUYU4DLpxDpRKzknQsIPOew6nJa1ZlkEeNSNFGU3Ith6dZ
MsKeZ80OEsL/sWKcCgCM6P05iC6KEXhMX5mrXpzCDQlRu2iYi2FZbkws810akGP3BvUEDy0Ku7pB
woMd1gHo8IS+V4nqw8oXJsK4Li2fTkzq7WL1jMn0UMg1qx6h77GqcttyikPQ0L9wQJfG8QwfPT59
Hjl1uLBzwCFCXVDAlIkavbYW++xv6jqZVZTGrsvPHUXLQc6cxFr2ui62c/NX3suFCRzrBH2uWg7h
f1wE/fJ87AJdibGMLgYu4AEt6Xk865jb8172yazyK9AUsLVzgTO8jxSOIaNvVs+/RDDjgRJxU//H
K4rL4P2/C7/8vJxg99ROAoJuYZJ/496mKrpcxLCfGUkFKAdDEoyhYIc6gqgKjySNSgL/bZUh1MPp
mVDlS1lgDZeJod+qhJTN7Rb39DcLp/z5gmt3cDxfIZ6a+hjKS8MA2xwYFQwbHK7sdIn11l4nRcCs
D4YwGkZ9Pl+Vl6dv2Mjqc47XYQUHLNQ+WJ1kHkaSYR2/47uxgjPoF+2iSbsZHx8/Li/SY8CiO74b
xbDY21P76XxxGbnq+xXJqh8cxkBIMVDYXxRlGtLga2FUaAgyDGiNuUBzbN2XfDoBp1x6mYz1JSZg
vKfLX5UnZV9U9eSwYdF1jU978wdL+AyIoDe7ZVrqBqBBux9Z0/TTg8oUsTO2j1hcmbwKrz0peUQr
QzGZN4RYoUvYIBoaOPdt+/XnCbXKRmceWfZ3/vjf8xTFQ70izNyqnRGgUlPcXUyFS+k8fd8oF1dj
Pr4I5s2XUYuxVS2X3q7kTTmOrIP1+dYtYDyHgajsFH9TbK4BmdynhpteqVsEcNANEWIAL9ljMsJv
p6YpUkxZDa9lct+e6ero0lUaGoXyHhtJ9cSDFcfAmsowjNZuMMAXkKyIyfrEC8eMtdTTOkFc9JoV
lUBdm13/Y/ihckJSLCYnt8zbyAYDANQxqZSYzX4cxv8l8sUJqRGRgGXypbwQO47mA14bwQc1JJaQ
vps80QRU6RWfYnd1gHxY3aa9bLppFvLm1tN1BrLg7ux9dlUeO5NCMTRnYyPiZMcZQBnBrFTGffsf
KIvHyZ5biO/Dg2kqnpEAlNt8rotqXnM/NX/5DxC6SyTFAlHmnh5CgWNNHlNByh6185tKPUCYw3FG
2Fl5VPNti6vqdsCbMIwT6Lp0mrRmpJ6IXGX7+asJhbBSVnS9e6b+2MFkzvTPhvvo6DaDPJoreTU0
1Iuu1vVUapRdOkNSePYj6QAXnou2Lu6rFf2BoD2+DGeRovBwH9Pc5FeNUIh/YDEedXKeYOqB90Y9
hotMx9K//kizLyqe0JCurXAQTDeOL7TjNi0Obj+G9K/1fSZoB/Kug+m2ViAduAkTgT0pSodfcD4Z
gWTueeDOEHpDKKRrl0+b3kjy41gEL8Q+nF98rOMPnVIeAJBr1GLlKFcPuzsSZ8tPsRtPHIh52srC
Dt7QC21Pl4I75EQNwH9F/Q6pb3/eYcM4IyfKno4eZaIleGkPlfqU7K6MEBvrvoGp5E1h0sS8U4z+
N54FYdBPin4zPyBRHcCw7DdZfYqhkD1YfXZJOuolqt7FOdZ5lrQQRzY/EshsmV5pzmL27RJCEn6z
+lk9tpjyxMg+iLR84N/na1M0GjriJhMjt/EBT+QIYCeOWSyn45p4Nznt3plEDZucn/MUS27rzQSK
BISKH5+yWsCgzHD9/mSX4bG1LT2U7BGBmAMdwGI06mL1jXxTqa6G6jHiR2YOwOTOnmFkr7J31vL8
lsVny+cEA/hSSqeVI15FTn2w5/j5YSDA9+CpXE6L2uGcyghP56RbDFSBA0W1wd/n7AKc5r8lRUpM
80zqkiMOugoyv+GF14V8wRfSXmKDqvew+ttU4uOCpmThn2rCWAAlNu2OexDCpeoYtBsjUOxJJtQy
A0sHqMaoLozp801qbz7kJvtuEmKWY5I4Bl2kxJcdZo/KwFkr0zjXSFzWSXrNgT450EzG0HojxbvJ
u1NydJweoa/1Z7uYk8s21Rb21bY7SNnNlzzNBFtI1u1JkUWrNiZzSl60utPMHcx8m29QZuBZujNs
C5sXcH3bA/4yuJ9lJh7PiBZETOS1DHNBHMm8DSf5bcWzoOPR7RbNV0ZaMY8NAVDHp/tAugOXcLpL
vlTQ72ecLBwHBe+yefK1tfGfUUPnyJs+1hDdsqyJM33HaNprTAFbbktgpbav8eGKqt0Ojs6KTKm1
dn1qx5tCgoX04Hjh0ETk4bK79HXoXGc2vU96BUBmqXjDujVI97fkPkLF4uc339UeX4lIiZNXneD6
OHABJESTqoTs/tB76iJv3Mz68PJpa8p0SJRMhIGZzCXepqLsv+PtkBEQqCY4k3HtC4qgVGYiRsaU
ggSCFaCOfekGw8dZ6HMS1eQbEgab3N2wVLVhPHqV/5W96YE0e+LH4fmlov97X5JtHQtzxRY0DzTh
JlJ+AP2zTAcYrA/RPdIGa2ywBt6cYo9t6x0qVpJjCy2gWrO3ixenHKaJxz7sY5JT5lbzhA+Ic9ne
wo97EFWewvmlCsgJTwa6yEcrVecSK/hYnXewyWo9T5YnT1ZSeG0Esb7ZpPcrUsf0oMp5EWLSGSpR
RLd6hqvJL9WxZ/RXJY1ZNVEYyk21ZbC6IMbwpFF/ZDnl/zAL9JeKqnzlX6JwFffjuajh+6DEBvmx
PljJ1aTRmk53q+4IefOW/C2I8cBd/xBxlUnbM3NedR5Zh/VG2O6jANs2joLGvv12+clr4Xfj5CLQ
t66X4odmJbQnjScl2hF9HHkwzQQc6RBE3+3sQsqMRuauECUDfnmzI7Ul9ai8NUHyBR4Zke+NFwtT
Tl83MdKmHUuF56p6Kng3oe7y/upitBTjYezlxxR1I6M8O7c4V/UoZBZmsnGtI/l0zrH6bwVgy30e
0oynDAclD4llqjbWmbs38+PvAXhGLO12zs152W8t+qLTaKE6g7ab5ekI5TmGR+tEEpmXps2R8BW1
0u/eEjSd0Cj9+wrXai39S1xUXM9qjFjE+vw+78GczQIqrOHGgnzXlytWBOM8stYZ7zF5HKGoIdiB
nPvjqpFCSDDX+2RYRKaqtP5X8JBxmyo71Ivn0DvTmW2rUmaZUDbZCp3LSgB3J/x1atGXc3FoSaTH
D8Wj/pFS6UoEIoqV1ePjV6sPjSlt1MVVXjLulKQohDS+JYYe88N38BtWnsVik0KXG4F38kV9G5Az
7aOdvImo9lR5nT0hrhCt0sbZmZxMys2Wzhnm5ge324HoY3cY0wS0788OSEBXAYSVB0nX6HcQV+g5
uVfEoeJcOBwHg1YuL9wHgJR1C2BPGhXFP2G8ve7LPRsOVb5VJiZD1yZyyNGknW3H7J3fLRComknS
zGNlFUmnvNHQIZ/a47FscBSh4eetDzLd71CASnmbtjEA3LoaZT1zzVNXFRRq9Dfi1YAUkieeY4yJ
FW0zihagHDzydALH4j8H5tSvCOUc8Y9seFlZARMa12gQ6E+UODo34ECXbkcCUdpVpz6EWOMhMd51
Iag6eWeId/a5Bd5jptKCK8FYwph9v8ia7KXk2jkuHaFU4Oo5219w1mvI8xc0cnK4Nhwfa7F650tG
wuUnfwOMASe+//wP3C2/OP//g/sWGjrsvhbgrAe9QNMSy+EDGcU2V5eo+D9yJ8sw8vpXJsbE2OT+
cx5YU1BfnPfMTzPuapibYOfMeH2KOboRw6n5bjm/U7WNZiEGHTJ2+IvUp/yXhQu5c4cB8KaBZheo
m+KKkzp6AzYpWj8ZTEckSuumfjcWEnfIrP7Oo3sy3oxkNZZVPLqdOc2tmmo6iJ7WSG2x2UavPqwh
4o86jopij3o4EJjz9ZD1ervFZgDHg+43hBJ3eGnGSOPYUw5s9RWwqoC3LGXg8GgT1RIT47lUGNkG
CmQtOI79STXHp3td5lWQUTeJwZOF1+1/ivzTWFmtXegxQGE+pvnTDpRZNRDoeRG00OGRnBw73D9F
BCWIvWj9Atx8zJewvDCT3+WTPu59Q6pyyZusCXx7I2vq087MwJ0YaFUkf82BnZf0QtviITExdaDp
YhhGusK/cVb8WN401yvtrgwyZwPlmKFOTtoklybk7o7YqFKx33b7GSXgR4JTlep4Xbif5JY+C+kA
l59uDc1drSx9FrogKUb68bfR0KuS7ulvaKt06uPZcYe+p3+h/OLiRfpKlqyfV3osl4xNLcOYplZ6
5wNdRif5qGOOlw8LoKWlvtRJg2biF4xdLT4yKi9Rl1NezSBSRwLWBNHIbyAEMfXzSHJyv9ifW1Qh
fVMH1fIS+5X/2te45Cq6q/yRHZ6p8tOq6VxRA9IsfoVvbwmMcbjscuNBMY/4LHPnptzrJuOSW3Lj
WLnHgENyujds234uEDTYdaXJ1WJohZ24ir5pGnosbLBEnVcBm0xYkoMVFW3EX4f0wbAy3+n01ms0
UOqaTcIsOYPYyhCGEc9YhCf4KgV9uzB5GTolYmNC7CFBPdQcOzlwjukBMUiqURUkfIBVlDRcixii
90AImxsP8zMtaq1VPbElT60CoGuNkg2AzMu0iOALU+VxKC918OgZPNh1pE3dfWvd70NCSlyq7Uni
zlo6IqaM+CepZiRWjT7mBZdbYFx/P+AYCS1PnzaXcUI7QnZnJJwjKfPe2YAJEsi86GYnzK9SnlVu
iV64ThsfhxVXWd6bPbYOAvMTKu1gTHSqeJF6jgOJneFWEFU8IjCzNXytQPJFcOsefHMLI/dy3dRQ
PW1Ty1b0PK2ZOlo7vfNHDtcllaCFyYPyEZBGZc7mTg614gu+7U2m3DJ36ql7oBmTGo+YY9stm4kJ
AesZ7iPDYS9b1X6/QP1SRlJ3c4L6QlQIdkLtwpUbqrHNnJcABhzfwM4tlU1qJUm/0/2IF09VX8KR
D+g2WHTTuJhTFCN+fipL5XBWVxIS18Vh1SIJBFrWvZEINCDWisgJjMNmzh+OCNwwilaOCImG03uP
pjwkSSTTNgvSWGE65SuYVj52SDbGPDtEQScY5WV2RQUyZHIHnCzkr1/8B0X22XppdzVBWl2Pa0nv
TuNTzXbOO/qiy69S5HQ8z3cj3fA2uNOkMb81hA4Nv2dwefD8Qderv5W49C/HVSQB29Xdjmv6Rw6r
lGMIaoKtgOPylw4TvUkwPpkJMNk5lBih9QCnewNYqYYQ6rHtH3fKFjZ9u8QFlIYgpfjLRxDdqGWP
9RPgBEi+5IlgWeKxIx2EdV3Mi126vE7WwTM5fTLeQB5QmTTpnVARfc7ihZUDhP92bo5Iw38t849e
e7uEY21pyY/HSEkTQPpEwap0re8nnYlfViBsr+nsR4RvfAzoNvQ4oeWxmN0qeodRbBq/ICJBzVZx
OM7h9ZsYtczepaIfMv6T4Uvj5ZsmmFICaXhzNpSojbZYJPQrezTZ2yuQGaX2e6WJ0/Y3nLrz4jS/
VvwGbWWIpshvNMz7mwrCVE6yICuMyUghs+TjXFnpwLRUdONj8UuG8pLjnPw++32i87vCt/QY7wpV
DzjS/dxh5g0QYU+chg9Dx0/AF8Oe3tV39I0Y+KywWNj3FImvVuYDnMj9QzSqfQM7t3PAN637L2g0
teFRQfypbnVuTOCncLuslPNpEOzMfvqAVQnxKfc+O6QcGxRvSLWIgTu4f8vLYGhAMp96XVOuKC0z
/p9XByFAxsB+dfPewvSM+0V9KIAfpg3GhuNXAwB4RA2S3qtKW3UR/Ca5jfcoNfN3LjGIh71V/HPl
TF/L6+ARTrqWX2DBeiJpJsEfunNROBrffBkGFDQ1clJpQfpxI1M9Aa8mlohImYtyw4fT5SdpV2s3
SW2ZRCzCIeJNp4b6+OfPgTUZHcnGdufsYZeaoeZGPHhgDtMJXh6H54ykZhK5y8vhMDcsGcytkWXP
BhJBtXg6zgIThR+6Xj9aHdJ2+j0RD7rh6axHZvEgo5I/dMAhbed33VVm72Of0T6QdjzVLLQSk/ZX
AGGwGToDr//8eZ9u6BEs5NOHYJ3w4vbHgYMlx0TiIuWf690rz8qc1YEAB8mYkep5pUtnkGSDa0w7
AZ6vTBtsROwyhjcTSOTtFqsLdX8fyphewCk9v8D9gudetwRbkqYohhFyF0I0GK9jIOJnk1UJIFiO
II0UkCwdNj3pR0UbvDy2yI+ZSrND4ZSc3/ky/WXxHeEVzUPfxMEB1nkL7jl1YkMifBg8Ci3+2LvJ
FlrPVqSzZcLrisTBpqJ9998k8fN7mtKpVAF6amVPrqIZz0lJ945IwY/3B771ZWWdwTLtquu3YRnr
FDyrgV/SfU+hivz761FlGLiXPriQ1IIFdOpqxQa4xYFuEoMX+JtDBYq0mH3VcIGPia9qmCthZt44
CtXzPZ5mhzEfzcu4nyPQ2Rgx+W4+0y1pUUQtEEn95BduNLYnT2AHMPXyg70svtp3ZZiIyWl2FYzs
e2MN/ZQR5YDqk4aHI/AN5FHpZWanxdcKyHBiX2/MpttNHvENx9pJHrG+It4n7Ha0MLuMwZCagNjj
q3r8q3Ra6hsoS9gEAA37Hj0hND/Nogp7Vkvb54OCJoD/R9L+BOzMWqMrY8Dmpj3r62LZd2DAtHT/
fEx7O3CkakQA/R9rqX3zozzepOenDoVU0UcfZkpQyShBFj8ClchqMTZZVoYhCoLTOLeaTo4MIJyp
pkq+TGZRyGKQrMel4+Iu+pJbZ45I3I0SSk350cPp8Bgn3/NuZuwZUzIFVpWCzzQyPKNuZp6Rui4J
9n8HVoPS97EhoChVmtbx35DpAN0Fl/O5pHVWWKaGBB4J9hnDzt5EwpRd2uIAJ0j5hXsY5CxHUJCy
cDlz/FN6m4zGDF8GRAGNMGXYA3sR7CiePOxM4kOpYWm6WcMSOz0rksNIX0O1PiQ6lHLtZJ1g/teV
oe2NeoJdOPgxRiB3MrldzcWhgCgGVTdIzfH0srheFzO6sb1exN2uH3cdRlwQwKkRwfOO47In1Xpt
vK2mfRAmQoxrh9JtoHWswf+BgH04gBIQafkpoOxAFxFWMe40xnYwxDes759Lmg0ElKZPX/hAPm2/
3nlN2HHXz5Dk4PE46xa4Vyi7aGSkoItb8vmTMqZUAbv6dPg5WeplXtHqlu7SgRJZBurrirVz/xh5
xHWVg9LBAfermmiDEbygz842JEKe+Ub4V57ixC6xafdVZmTcr9Zcvu32suUdr9gwdEN7j7EFEB3V
8TrSuVenGfsNiB1keDak3qh7UbpE75vk4tcKbBwcLxkALlZ+uUzRhDbeBZliVHqIJE1p12wpL3O1
uaW7rDhqaTSUqtVGNjBHgAfzdcoRToLeqWN2w6IL5G+ThHKyRUPUW4/KV1E01KRNB/GvgBwFifWx
1Ktq7Z4hoYY+T6eVeEGLo4S+IBk6o4a0C5gC/XfKomSmDSJrBtGil/cpn8Vq1LTW7YIthx7/H59G
Xa6vU0TW2ad/Pdhul79/Xdp/rSmqWmzvIjPQ9lUmEFKaWP3fxcQ3EIp5CWAlsUPenxhtkMKuwxAG
Qibg2sc01szlZeU4GNxJCY23YYIuhIFlit2eny9YASAMtN0reisc92R3vaqfY4OMZQfCvfEM/s+w
7S1euTG1DVbpYjHtCeXpOpLtHQZTX+BXqPVm4LHS0D/TQxI36r+rJKzD6pW6XA+NxtDgF4KU1fcz
FdArsxqYeZw+0Fs2tCHSlb9hD/VSq45daVxbq5AowH0OV0Gnl5plNntYtN7JBvZLDtRj9gtCqkkC
ufe+vg9njGeTMVgejJ9oIfZnhCN7aweSb8AvEABqhXvGt9qxbM6RDJG0XUKev79KUgioBASxPAZz
qdRylGUj9m8YbWSCIHMmRP2+BI/4ViuSc6vd+5j1f+VsA0AX8fdLDLOmX++isSQxGH7fx7W8w1g3
M8++WlClNxzIGQLtbJp9vFL1s4CUkZ3u0D91K8cPBaNyDwMMJDUomW3NCZM2+wsR53Evm9/S9F78
D441QS8ypN0+K11qiHIMUGERVbnfTSENUKUN7OIngo0nqwOX4Jj94Htvo6SQzg22zp+GGP/F2esR
Bf7xz+tBHIP+em2/+zHoKhhyIaxu9lNXWVut5kHzHiSmTK9fHBqy+GXc/UrOxlSpTAZ8x4ZYawbk
OYEi4h8oQJYFOPjfC9FO8+FTG25dAkzNw3IZJ/J2llLmk2x2N+PQ0PsVeAfjQqjtfCrQpxffP9Pt
DU4+1e22UcY3NAfON4tr7IfWot7UK00euN31zH4pFlmp74aaPpfbYUhmPAziDFwzh4fCM86If4l5
AiYQVr9JAO/Y+qxs9OiNtmRWgzkpVmTIkutEH86xU390z1+H33KfdfWTVwUbhNBpQJgN8EW8Rjo/
9XjnT6toqlgltFJt203nO2lIm6NsOkmrtutVyEvN2RQvNP4h/djJyhL2RAx865HP1ooZseogqDWS
uEO7jZsZzND52lLUVPDRBJmbmS47or6lihApzucBty0LMd6axa77k7RuXZF71HnrHxIE1a15gb9P
ssDI+IMsqG/fsxmouR8c4MzOw7vSyNrcl48NTK3LLcEvEt05XuJejZTT+97+RyJg5R67nco9JYbw
POw8TTUvxxMsaG62/qv7NEZ/l6wCHXIFGELsr+NsbTHBPRxoY7wJlA6Uim46+bTOmvWsDlkH9Q26
4e3quYrAcxgWdOoUvOzDQOD4nZp5mQ2RVkTSKipHcwdzS3OunNhdUDVP7PbHNpADqBrAtXR+o6JZ
4FMKG22t6mtBI/481o56U34KFYNMblIdvrbYJpHwkl0U3TJxQO4On51ycEl9try+MdY4qQ+dTcMa
9/gCTZ+THGbpoDVjlyWeQq0TmCqunPHTlX8sNDvdKY7y9ihzaDGYmFQDNu/vhov5xjrqWEkBubYE
Ha9wNrSxwvY/mhrxF1DHZK0FLxfBQfP1TX0ff4hzU7zkRNWRm+WJIiiwQKy+DXaPwKh99vFi2uZz
5bNovX8pZM8lbiQ8q+so5jRKeeG6Oa56BKbGm/WjxsUEPDMZGpqXdLZQNUfEc59076Oj/DBfqPJW
/j/n2aRasBL10B1wfnSU65Ueui+6o4f8ogxCxOerv7ozkdoiBLgec0J08SONV+OgEsFr1inz/w1F
x66SHZNez0BYf83Vw7su4TXnLKOXV6nwQ0DIRSPh2hpDHBUyRMSVo8KCH6kE7WynFAp/b7aT9fw1
bMsrpTDS1RiXEw1UC4KrElQyJBFircHW/3qVBZcxHW9cbq5dCQlbvcPoqGwmW2pCzVQ4OV0xiXpb
yAjnKp4xdEUT3Ci70pCUODbQQAfbatCGdQUzrw9keP7Ud+dERcsuUxNnZhBBoMlXo571jkoAWElS
hMQnEclXrFBPI0AJoI/8yo9pxVtOfniUgpcsNNNjCmyk6p5jQXTs7B1SV79kd8mA+e3RPZCgznlI
U76SJBgY9dxMuscIgi6VPLsuwj+Ov6tcqBI4krqNpnngyUb0zz8UCyL7sEisSdFwCHdd3oo91sNX
oN6wb/M8yD+7jWrjOrzD8yVruAwdMVCjXfjzXIUmM/lWnzt3Bv1w9EKVLCjiX7WvwSN8nQdaHAPG
6A8sC4/ArdTCCL4oO3OxXv3X8Cp3fy62mRBhWxrsFm14+xsqxpq1VZ6Nosj2/AO+KFBBM/QW4Z/m
NHdlZWCuFoFdo56GH/Mo+53DM5PIWUFteag9weOVVRa+KK6JCdZ7cZ7sNVkHgT9tCSdn4YdlXHu2
EraJkjjMR6N9zx1UEAsvrB7ORutKk/6SVXjfAFPRstlh2GzUIL5zapOqkMrF4GVonj+3uCChgnzy
HJGPPyc2QLKh2yLGetclI51EWvg8oVvMyw1doXh0TWTGBb9PVG3biBqVlT1vbBuEOPw9jX6RKBm4
dUyh/TQqI+HJGFdMo03XHB9JW/puNEurtexIF7xTksA4rNGGpA6LWN4hYhjCl/C5oCAUZD39sxD3
uNIMuVKCqYijsV2ZY/QOVOye46OCzq8xI5DLVY69AMcMvOTZJWam13ANW5I0yKX8x2JYTPNSr3s4
vgJwSrkfxekmNIET15nEHry3IvVSfEQcmyAr+7SwgQIlbdDM7i6ImawftwXznrPK2DI/5/6P5cBj
wlrgbr9uah0WA7uehIcEG1lcmIxuKZMK5tEwDjLEDNm0WTbxdhUQkCHRGy9AACFJ4UbfjkOfB736
30fRn9EzdIiYo3pVVW1loPM1R49TjN6jdeOAevvlHdFDMvrBBABtGLnQuK1TAL0YwkrAbYOsn45k
QldjbzUacAsFGG88y2xAiHVx2fkUcyqD/CLBg7rTOepBZJPnft/7szbqwKY0WMXv7szmehJwfUUb
OODDOtNYm5VVSGrVz/Yzpqw9J3LgZDkEd1tB3rWBXn8M8F4YAVj42VjRZXTRRenmJg5B/2bHLM3Y
3FRO5LQGt4+DhGSsZoASE8M4RcOPHgRsicHdYXPrI9aNZJr603WjVBVshWCGSmSp/lST9t4o9dJD
kko0ggakZ38j4k7BfcXDBcc5aEns9oOkMV+adG3UcYP3lx6+OypXxA8/aOSzD13oE6Rj22QxIFTM
o6AaEP6i4o2Bzmo2Ns4BcIGPoFZpwAvPAuAsjwqttpSxPg/MRCbRpwH0hsYetV9WnB4+4A997Yk5
rCKS12c8s0u/hnWVtoX5V5fseKzPOJbj3+4U3kfLcGWOy97FIhlJOPLSUsNc99ivC/oNCL59c7o2
in2KXnKiyNUl1B87XeVqASm/iPNBkAXtCj/osuONMurtkUCHlaekF4crE83lDqdM1i2HtaRzgGQK
nLX2rpjbrLwjg1S94LQ90wtCV+KsVCn5ZvJpp+Rlwu/UEpEWKBkwet+8gJ6vcTkNLoapgJ/BsKRy
Zj8iS/g4AQoVjlVaO58nCNraf+d7AxB4qf8i6ZcpUbIWKHK7JuBpYyYGOwuXhD4nDLkOrpLfmBup
FzYBuO0w3ASILIuYQ/iB10CYEUd6+otG+RkHJT9C43Bmzh5CGTNI+weXA2hcNar0J/KylsAGgT2l
K21n9TLd3gUKY8CPqrNvxGMw0JY3k9VddNr/fR/EjZQIfs8Hx2YR11Ce3PCd48+q1IPTudxxkC2W
WK3gWjYTIVS9szwcalMC6FF4AkIMcEd6ibQNKDchcjg/lNcUeF+Fr05Qq1Ui36gjkwCkcI6ROB1w
ew2sdMm6zldSXBrNpDv8VIWJ/YX6vjnOUCSyX9aMxv/aGfvD+W0FEfgTQnkqKoKy6+WUDvZJTOM1
MxhTaG7p7LsUuwFJx/y71utFLGeZrAsHQrphLo/WFCPDEUTG/PCRg5Dccwi9F0dEsoKcPD4rR4fG
uwPSWPNF7aOXjrFUYQcQbkwdZK8O0lefeAWvtMuWbJCVQN/gXfNmMloy4iktuGOFgKcKzw5ONZIH
T2Hv60/qXVNBHSE3z/frGA2gX+EKDsjuamLBgwQrA4WeWegDuxyieHEPz+cecG27L5xAbQ1sfL1V
zDGPXcQhtoObkXemTxn6SWj4qbWLIhrbpp8LT+PkkMvawdspkcRnzy0zhBGBTQYfF2aZ0qj5GLQf
5CsvFKZMLFX3Uq6rZ54ZRzSFrXhQe68eJS2V5UQZT96bN6JFLsMMVefs2yUpn6XDw9NUVhSI6/Yx
0YwkdoCIiZcmGDZq1HTv+/MPDjVVZdljMfVtGyqTZPAWRFKRK6tjdDGHeTelSZkrBOSPFEjd/MeZ
Q5PLVIbBkQiCGfrNArgFTzq7GM/ybzHQk8DNB8CjIwefbuvQ1+qaWN52fVK0r9qF0qHbHJiIBMla
6jTwoXG3ZR6bSYHI51zKmlUhtuLntIGU9XnuIweJT7SR/tsl1wcUeQcowKx7UW1hN8iQyHxqGMU8
cQ56VuJYEAO6+vtH9jZdmFrOW8/wFT3T95IHUrWgJVgX+U+o9Qg+08kmGQZ43QLO5nnowZpn5oVl
ZS/PYgSu4qW/pFJnraItavkcZ0MyySYJ8qOP0T0O7nX/R4GKXA5LF8wKJWwlrQ5TVekFZZPCeYqN
xACbPVpNXsSRE3V1FT0RFw7DCkCtAEb1CIYVCb7a34b81jJvP2Q9pOU34Xnf4tKCI8XaT3h3BTWs
eKvwMGp5Zxa928vhwbKMICMzUIAMsDKdbGJ5ktfq5O+CWBIiziB/tLCqG6jnzJC0ADyayT5yWgWb
n5kTr9A7zhbKC0IF0c5XaveP4pUA9bkB0Ww8Um4RzGQ7tVo4e//voKDc/1/rq4VABp5NfYrHvkD0
q4WEY5MJLV0mjYdYQyGJKtiK3eHw2K4gDUycKZqgVa8VX1I4JrW3fzcnUUEaIvSkY91S1g3uN8ae
22bYZsdc98YJEQGOA12oD4+dR7Ayud9X/pvkYKkSF22pBuvs2LT9kdKd7qhNsLXHCqXoj8mDsXqj
Aes7bvTvqkCxTeE1ij3mTRrF6Z1pwp6Dj0IJDepb/ZUxn8sbq6YDwYy9WOJJXAABtrJ1HjC+dc0u
WXz/7XoJ6IzD1rLXHRWMCBXxA2EnRfTH4fGfR7zjoAYLh8HEpVgHLbtGcqWdcZ8RgLN9jUszbRpo
D/dywXiGqckf4BJbwejqERuf9zObA3HRU6fezP+3TJ4rGkoH1+cK7fypa0J6D+dF9Nkv1yZbub0t
NQpM6xwEnNS9eJM4n0gLjmbbnKCj4vZWW/cg3qm73+LdYwSYtKhJojYFP0YhWixe4eqwhDNisMfB
ruGMJuY6WfWAv+RYvmnS+jvimnAa89IqbhIDLWH5/InOo3SOSejPKoeEp0pBfZIkbVezKJmvkJOH
dxpCCKk1D4x401p5M1wSL0ZlkL4mIwd/idsKpG9FcPXSOLWTQ2o8K5YZrHWfuNv6ux8fjJ/oSgZx
JoAuYMmgAbDrx8kzezP4WCJJC39/bKZ6PcMJ/57CDkK6hYBSRcVsv/ZzNleb0yp2rXnjtLhmvTwC
YeVFKcwqRN0uL+s2xHw3IzvvNT7ZSq53uyVizHW2TKRN8rGZ6U8ifOA99m+1UAInKkM8TwArLcy2
tZW1NtQGYfFTvozfcE6A3PERcZEdxEdkCByhAAESJPOj8BmaLNwbktD0hG3vKbP+3GrcoW8QUzFY
ENDitFIoJi2scGAjiXInHoTEeGJGg7gDIlZ1aPaLK9080eXUTTE9OGUJ4m6ZF8f9KwwSZ7fzTsVp
8MZnGVSoCtQQu+4Hot/vECmBavFmJTb4cnCBC65nn2dm0JBvFD4hBzdLzxdX7HGLyM7LldB3Amum
BMZIC3Z6QK49bd4bEv6dbhTr210+b5jXZ/PIetQOZvA58b15a0fPlUvxrxxJMV/5SquOBp/aBRX0
2QCxUXvtS0NhhkKLA9vZCHLKaej6RL5VerW3YM4eksTTxjtAHi/M+c2epbdNlrHCFSmZT+EC2uQs
1OmZ7RcR0t2YG8SJpcX5gIK08DLsaGLqeO44lIHsdKXwPNLS6wJn9f5tHV46QSZ3bp371ypHPi4e
J7cCKUc7oFwtY2R3mFvYq7kSFHg4GiVkadOf5fZqNnQZOtKmaSitZFzuoUApBP1rgJ6sdamTIQC2
Y+QG6yLTKf7mU4hqQ6NvZ2F6uJKrO7b5TmccV8fflbHKzoCrRBRCMnXoAYDrsrugrpX1xaFZ14wT
yyp5c0n/x43RCk3tf9gvRDEy1U2Ya2TfekFYveZLfV0qQzqBXCp4S7k6LKkrrfi69+DUBOO/bHry
uAgk2r6jxrGpGF+Tf0T+VPI8MXSFXOUwpmums41dbQJZOWOLrc1dkAjhEQG3fGc4hLy9OEp55SYh
AJiOH34PvFLFCiC4gEcEZbuTjwJ0V418MvgUtSLOdKBURrzYzzcTXVh5gSlI3m9dTbb/lKeYxoQp
c4mTf7Pg3VZ36JqMDt/ogGsVxJkbCW/QfYbLLKb56qgvbtbqK21knaXd/Lg9JzTIQuH2ebfrzj4F
qFUPGCQcB19pK70uxx4zL2xe51j6+VJ/WcqCRY+qQrJtFuntMMpt41EgbaR45W4CJjSd+/DsAitf
q71szOI27jsB9M+zJiVIT2gikFB/tDlqRmnIodT1a7J0Ux0rsfwhtNCA0d0+5jdyqQvYBufkrOyz
CeYvKvrrW+urK+WQNeoYId9ye/thT9+466/N8ngNNqwyxEo04IZxXmshY//3VEOz3iWUy96MNo8d
4mHLojMx+uSkodYvN9WWgOaJKiOZt6bbSYXBohPGCQzGlNmanZY60ezL3xN5qLaL6YclQ29arJdY
NKi3t0GdSVGeDUTrQoX5eGBUMTq/XpMg98disBbYl2N3l+O1Djo8R7QN+d0u5KwAMImOl3eOxI8t
9bVv6D8SHuzyjHy9ZmZrS0rLKlEUHyWhvXoGBUz/N19XGYK452Gx8eluRjoz7EDRiVs9JH7yJccM
TW7o17dL7Fps/SQtGJt5CpTOVSRPVtiEJ7uFowrsErOD5a3l40h8fq199xp4+nv2f7kQpAd140xw
E3UOPc4OnkK2uSlfIG0b9oB8opqUfIPIT3OoDBsAPIp0+qweMjVopOHc8bXhX3YIU4RH336g7zsu
eLt/K7G4BjHnjWJKgEZjM+45hgN0YwDOX/faIelL+VLBzynK6wuL8ghVg1RMzwMO1Cg26PYIObZL
56IDVyH6oUCWcJEpYcPqymvT4hnuuxcPrTGvHKAsAxODGM1RfUALJCwR9InyUIiKEvXC4rZd7jqm
FeX8WqxYuK1rZkQ81/tju+4skXLHeU98ExQEGCcCIxKXdYzp+1xQGLzwKJxKLydR3vhSXxRhh9Kk
tBOQjYKpbdzxIpxis7PRaSDjPM5AJNeTbcikUM02iyBVB1eIO6/64+yFRfdqOVtf4fK81LNo9N00
AR3CgsdStNRgN5CSoCtCDXYesRDIyKJGSod3Yr8GDjdOE3IastrRvVBVwt42xXpfuAGHsqexXAAN
BHpgZw1jPksShB9pFz/7tJf7uR6M1qPovWXW+TkoPB2N1R6U6Yyf1ObhTL0m3coJz5nVCFGZ5jVO
zFe5g9WO5ShMztAap4VzXNbIGIwTVubmO6HasrLOnTJBtCOzxu6UX+7jmHn4Q3Ty/TKgH63cq4I5
eX1HoQEzMQyWDLIFkKMJ8TrZdWE8JpmQEtAC6kHZX/pB6+3me6KHXPm44NcuJ1gR8DieFMEK3ltD
QikJUBWQNMYDL+ppusbYYi2dyIKXeqXqotxfJ9zzlRydEHxo8/NqbrUhecHgAN50m1tkJcBEKpXV
MgDeU/bCzcONkhFJI98v39rRwx8ORBo7gQMzMZ5I/WoDRjxDqzsEY8JRV5TUXARzSf1YxVo1qLUN
Whq57ITulmBln+/sI1XkY+4uqTyFwr/5AH33fdCXjUDnVuv4cyoZrHYX8gX4vyNLYHPUE9lQGD3O
7kyUTF+lt3lFPoyj2OKihNmACjuEzgy/QwQiAoiZoZZ1eGR0BdLcDf/yH9PFxYvtPLSVX+tFK2gl
L1HKOZ3kCURwCQzg8DJHkwLRcRP/oRTxe7UZjTU+wFf9obvM+jJR+xE6xcSjfAuy4B+TAs/EVtPr
DU5kBUp0K/hTGw1SheK9qjhaUA1vucaCJQmHLo45Q9PzspFVvkyiVLXa4CMqzx8cSQbmQ4fgFUJW
HWwyXfZ/mctffdaCkctK2zOJiRpkO9xYvrc4b7oo4PbgUjDw7aguCqOxkVy/wUmOJg4rUhrbtNbz
UnUz9Op54uajMJZHadb8pQb0c1iDbfIgu5bBfxdvtVjvcPTIDFJCvQ1EaCUG71c/oaYi/jP/az8x
n7U9Hg4zC5KW+pkSBJE+JDJftTpy4qlMhN8WidHbRTqf5/5hjpIHqQzAOAMIq2gRvxyRPA+8GY5K
P5Pbcx3gZJM+v1z+APcvrspohNocQn1TvULyfAxdvuxWAQkq7Lnl8CQO0m7+m/JvyXkRJPCcZm+1
a/sp+GWM+jZ5wgPj9uZSbhsP4gIzce4L0c2C08vxwklhkZVAqovafT55tsfizQt1goxt3kL7xZDT
gdZkIAmuzaVZpQCBf5j0nlimQGFRVpQdatStiTo/DdTrqrBeyS06k3j2Z4fMGiDfDWInehgQNRm3
aX90W/3e8Z9tG+n/eBlSPZi475LF0Fu6KUKZ17bvNi2B9wv0Xlc+KQwRK6ducVv1ohPTk8218IIt
uUMN9cGJEUlbj0kCiWalEsj3nQFf42WJXMMBKUE7yYZREIu6oHq0L8jgeUBJRHvbRir7kszpzym7
5GKPZi8SZOHZVAbbH14sCWGtVp+EkAfhl5Cgag6BmzTi3hqJjcg4KMxsM4BiIxpV3WedvVOPmlt9
WuFyJ+AzTe5CLh+RQUiyTrD3rM+gGqtRoPVx+WKtjviLZvlLiKlFI7JTi6IcaMsz524wQjXlduI/
FI0ICZb5YTdbJDBgUOIzGpMOjvmwKk90M4YgaLyeuS4amHdEUBJYzpHEjpEjo4upMFJ0b5807CJh
C3UXoscT8lFO52nuVA6ZnhENZNA41ZM9sqvSBrchAUa6cvzABCBUsG4Ct0YRrq1krkL6sWirWUat
etCpptyl4lSJTzGUPZqtW4ONiVJPmEuBGfYsDAOnVXbgjO6VD3gcs9EvkxuW/h/pYxCxPcUbPuDI
fGxuxzRERPCLeIKcHVu1Ja+w36TKI5Dg+RJqn+PSZWa/qpCJFMJoPJUOBy/O7pzdV9ljB10InY0u
kr5dvzYGLSUyUTdKeENS4VMul7LC1alZP7mJb+4OOxIdZVx0YxPA21F3PsaFT/HYHqE3Uwa461mA
xTh2RCeSRQo++7YXcf4PYHyB11Ka5CMv3tA2VHO9kwIsdRfYVvO3eVRQimQxV9mOkDv5a+Oqp0Lm
ptCzosC9yoi7u0fICk46SB4P1wNqy5QVVWCKiNLIMIG3XM9uaTwhrs2Ujzs26A0fK7O+tDG77FhS
igUB1LsEbIWYAkyayC6LBOxN2O4P2NE3Ihf1ypWao+qtTSHNwiExDm7RjWh8BqIrtqeehn3KkY7F
BBi7C2z0je8CW3NdHHaSkwnsbt8d/YOc2i1h0Yab67dfAhLeGlNkn8AUVKWiJAh2+6fjHON5gBtQ
sHes3aiFLBndh/5ECRESu7hmOQS8ObLyYis7ZV2r/5zlRENkWN0m8TzRI7hDlrybFxMvJuFs2tv6
WpHgYLuFB9xNMv+btNVbl/Rw/FsEgekbqEG4dr/vnXLguc84EZg82M0H8qy0Tgj6OiATPvvIS230
6jk2UX7N2wMfa1XIiaW//OYDl+2NzVRP+w5nD31E4CDeZTJNUGn2Bed2SDSWY6cF3/ZNbZBsHPYN
PPCR53Sq2hBqZUz8jRfX/lpnvEVuFQCcxIBMWeIHzNMNlPQrSSmB1/D8Y8sIw/0sG3mR5PWSYWMJ
TRS8cXZIPPdgNbJnqgbDGUMqcxASjhiZ4XL+Ub0rPpjYtOuixA8mS5exLyNDbdV5QDQkRxZ8hb0T
DYB21JCf4oBuapS3ETGswxJAoB/HXu8J/ikTMdzWPgENRJQg2FbbiWNPOLmGkeedKNr8ZHP81kOh
DKqIvxsAXJSjcZ6X8M6ALIUFXwe7VCrKNWMFw3C6JblZfdN9aQENqTMo2ETsOJSsiq4ICM8U/9Ey
eH7cJMIuEwQJsDgWG5dX6mrl2/Q785QermH0tWcph/lc2nc3tQTHmsAQB3+sm5yGN+kFXeRHflWh
UPUiXOMt/lYi1zWPxDmIxq7Y6UiuwvOZPT22//UYRcdd1gS2ii77T+br7XJZ6MK6lY153ueykzIb
ZJ10wdL6frZwx24i1JRuLinACofPzGU6McogVJ2Xl9HCfxesg78ckAQnRJ9ZlN0O2//vgLQQV0mM
5Ui2jwzOBYOYysKw3CXUgQkTzgmuz2O71AznCXpKut6WO/02laxz/RcgFcM/CPUI6GQxU9QaxW0G
1Jea/Acy6hajpL2g/4rAwrzMFmsMPFAYyMCcf1rwnqnRpZyYBnCzSeG8oyUNJZl5rTqntasU8VM9
ljOTGiklr54A5GdLkKE3RHuNE7hkE3DRBz5cvikcY65nx5e2UfeSSgxk5fGCtFiM+iJ+UGu4hXzq
yvmzML6s4Z6Mfow31Hq9Kj5kON3IRW47UOiPCkcNW79tB5dAUztATTJV8L5M0+gYsSD72JdZ0QEy
ztJp5Tm52fqTe4ff/XEc4PakyaCm3+Ytn0SFq0W11mYY4U2G2EXEB+u6o6b/5WZ+hDAURh1MXj4J
AxsM0VFEUJNaQmTpeKz0586BZ+9O5hp5MIaNgTkBnodnfxZV92VzJEBpQs/tXCJnsNvzFLy4pWRu
frBlY2nIN9wW13LCyweEUDqfNBt6HEJ/LJPUkfLARHDnvwrm9tDF3/I8Oz9wKLN5awLQxqItU2BL
uSKlVbMSBayTdsgG5dS478kwEInHZpaGi37WFh4LvKwhUGzhFXA08mRxsaeYmar2WNShN3AoX6gn
xUVKiX8MuhejxyCLfYN4ZftMoR40tLx/V5bbkEKBzTzIKZAridBtqymFaCrg2uBwO3fuPQ7xaN2P
1KS9W2+6dp5zNPZT+tSVnBvmOg0W1QUkLfruNqDm+iLkbNKq2DSp/8g8RjjPbkb1LF8R/cvJ7OzQ
l2TeUfbHIRrqivjUNaAwBsGk13BmSeXXLkgNPK6ht3XTjFQ/qX+Eo2fIFRzopmIRRiK++UskzKfy
m6jRbfuedcgkVUKouknqw6xGKW+EqC9L/cx7jYI/UVZGb2GZclH4jhxjfWOe9RSb6zLYEy4PKMA7
Tg0gNYuRa48pDAJDUjMidADk43EeBN1lib98poxeZcdmr93eLzOXq2HNtkwTgaJrvKoMhEmdSvcz
mtAkawzk0K0UHsXkdLiHhn9s/zcJzeunmpAnWNmVjGn3dNTZhPAl4L+g/KiWXWAc3kxrMRFeYHeo
AWGScRBCIk2KbBJTC8sbh5Q6wRyOzWXBiPFJq2u5cVZnGTZLz09+FZmnBtTj+t09R12UKflHZG84
VAj7JWcme7Hogf6r6u7kkSct1VAO4L0oo8AeHO9/o7VmsR7aCuPMXq+tBC9O6p7yth+dk0zSCbCR
900UMK2lEyETPpmjrPY5t1JhhrsT/YmbJZqZJ08964tC1vTP9V3UkIkH9/CtXY1uXTZ16E+cLscH
k3F5xLT+6CugL9ECXJS48Vl0zIyHg9aES1POf2F7VcYlXUDFtySnsL6scUbnSjqBM1joMiUc3YoR
dG2z8Khu6aRminvmn0gadmXXQH+bACMU9AkMh/Dy0TXkePAvlSWRYH7M09D/+jALwn4kfHK3O0e2
ooAWsJc6PyICwI0kxvqWDbtq6pjguVadMzWkA7iF2V6B8qQAbAu3FyS8IZ+V2WyN9RjRlZSCW29R
BP44a8U+6R/nHmBCYU2UH+jyVBb6RTMVm7T2HEi70ar7+hdizFsj3+li2LrQmiU7v8bFUxpDvGw0
4X7AtCsAOjQpGSdZgzSohCrG3ePmL19VPGfAvWmzHqMT9aTyeKmKNLJxTXttcoCfatjL1G8R73HY
mqFy8SxNQitXdOQ3IHgjTyLLuV81isG07otrEgaiYmzU1tNZFkvH5NiM49422wf/NNEnZ6SHztyj
X7K/LAFxARAYxE/y383TjgQesATQ1YLLal02oy3KM+mwfJdkgpiXNgKrOfo8+sYnSvGeRQRrHc+5
0wItffuU54e6AQx20LQApjM6jLyWyWZqeu5jFJk3szt91QGaHup6d8X3dA6QMFPKXQru2mjxSweg
ZkersX8GR4K8W5rMW19+Notv8ig8nuRFQ3XKkYc524bdu4SMiXkAfVUEbFHQbJhIQuYfYqukbaCC
OeJk2peRiSmlmOmoaC48OAeQ8cU/cl+QC6fvhL6YE5izIpbTIzY3rTkVYscAV2/n9m31ObKeBjAJ
zhbzLI36/Pv04VnFud+uvv7UDxPfvuGBZkVKTS6YOVQbcSnvMTQPbXDUOoOKNfBK3Pc6TK2CclDb
3B82TSG0KOGpzKpQE4HKBqy+raSLlQyLrdhxz5vdWXmhkwi96PuM/6uia7F2oYfeOqhiQRVb2PJ2
QVMTfoZAogMRMLyFMueKZv4EC+Kcj7C0Ez5FeICSuEuX+JH6m9n6MiDRJZAky6swchdnFIMFtMns
4r0UhXc4zQNRRZuDTTxAYfVfuE/Cz2/Zo/9EyALnu6veJ62vmSmH3oOB7/d+2OsIu9X4U1qgbAZN
abuX1NwAYe+5gVrkXCxSKmE1P4PKRJSzawXG8F9qjrb9t/XOY111IGiGqWsUYU1V84dVGlkhiFPK
kMF4anpGRLtOOQVR2LBwA1UEsZN9I2nqN96vO8ANkB6XBQ9Ww5VaoRHtmU3cqslomnfiQTlLB8Gg
VBf5jUU7ilPjutoYajr9NuG6ALyKRo+2C5zIOPDN1HMQln/ToRupZdaVXMSCmXZv84+555EUmKLi
6OzSyAvsHpDywxBv5q4lbocVBo19ktu+mpP2rqfVd2Dpkc3p4Je+Mr+udm2KoaOVesVXq9d36rKG
z2CDt4qpAuhqb+IcynS4rv91I2UomL0MpYsAFGrvA54dnXjOtaz9juZkhBcJHQVi+tJJokQPdNMd
x7j1bhKa+B18e4yQ9D7PQOWu/tggU9Os6TNmT6m44dhzQgZcl+QlsYmJsRotliEtYH9aKeWoMe/T
twSxIg941LvGAhQr0WG9TYRJf7GtwVtDXurRxXohOzdU0OEOdM2WXs/axBvAwQBPVJ9tpX0FIXY5
tj+EULu9YAdezkrhJuiasAAnCt0BH16g72sQqOPAjA+ddz2ILAhNCMA0sb6X/ZpNbOWtZMrBfIbN
qPk898oMaFwhbpn6X5LjYniFfYLRijd7inJ7meHiJ5/ZydzUabljMjxKT+DcA9aTYmzZtNhFKyk+
1iKGzxbJjbHx48Bk2dILAMmTSiNLw9YUqHrNVad1UJtRAVbu6MzY3/ho5gymSsWPWWeYGOWekq6I
aAfDbQjuDs/ZLlLo/VG5JVpBredapFxK3TesIy84bMVAkbJoKuD0urqrLUk9T5jR4uMWCZwp+hg8
HyBYGEcu7lbB0Xs5xqR/zYSlnGHEVQ4Jt0AiqYduHKrqYdro8S5fDSnYPf0PWnPK/oCQxU2/G1xo
Smy4MlBM7N0HGup4g2PDtrObEACowjps+QG6sl8UGtrmcmS/JZ6fqHoGn/kTsvSdAcVW0JMkIs6V
VCcS87YR3ADCpVfVY4MwjjIQJAVyrVNEA8hFCVVvxtCN3p5egUXhSkleXjjv3Jv0WZeRU+CO6qL7
+1GTzz2OFSbauDk5/MxgJCtCRyD+8gHnTdq5eNxq3rFayBHRHIbWHzdC8xg/MtkFR7sj8ueOP938
RNqwU+vMLgnCvMxHDo4jNj+fAAchcmkqYY448JEz8DT7t/qRhUXj8uMaIWP6GOnhwXZaIDQkFUGD
ciMIMa3lFmOjGoKcHeSIzcRQYvHv+raRamoBzZdC3BxCtmIFRoriq2rWn/b6MKDXLAdUnGI7GcwF
Q7oA0zn6hjZKKYq+xznb7y2nsLJNNgdEtYx/0odqEvqp4c2myRSoKBTrljdjbwvjMuwYjeDRFx3h
iUKSI4YjdolAw6xwge7jKJcFYAszKZ/VboEBabLAun4fn64Dxlu2KGisH6PfdDgmSEP1jz629kMH
kyOah118KrmVKjG2Fq8nL6rtYJDA3azbcTw6O+E5Nn/DE7aWYNxydeAdkEh1OCDhFSnDF9e4hzsU
JmG6YNx7DggsRsCnMA5GPXpzOE77PuOyTOYc8Gr2U+smJ8MpTpKybzB+5o2B50BYrsAehZYHKGTM
ReKPCljTJEre7amV+GALLprB0u0Sq3KTyuZIOCVWNQxi4tF7A8IKZY4Qf+qMIKHsmBcGk5fC+Msv
GadZJELyaOTWV3gY6If9wL4Vxxx4hO386doJ5Clmjdz/7k+FdWZodtvl9jDPGtUAyHd9GCV6pwp6
awC03YcHgqD1GJs+8hsdSm42kiTSrrNNtsEnkWP2gF5iKxAVzv5OzJT0Wj3PQIsjd9w2G3/wjeaR
lY3TSv3AS0qDC/tGqCiLXCuO2Z9vHBl2yPbphr/0tOot6XTMPHLw0deN8SA4oBciuF866Bm88dtm
benKfBhgBGxeHvaQFtFR4vmxE2XOA8zkJ8wRlaJEiRn6jKaHL9dnJ86nxnwrc0S2gEGKX9cmKaVY
r+oHHZULpPka742o2xRx6ZT55vD0P5am1cJBACLLxOUIaJIyIS7+TIayNE3IYGVhcM7Go3xQp7hv
zBEdrey/S2XoXYTcoLsXpmGNJjGddfo7NIfuLzzgeB1kFz3fQXek7y+Bse1VRnvEbPTqGfbW5ol2
b9YrSVcnXcGOowH/maHrOofKINfeZrxGCwAi6JvKp3zkrtZ/6RGLDWRfxeYe2JysBGLI8VIjkSL6
na8CsRjsdQNtgtWw4+vM1i41Ua8IdL9OdXzyNMQX79851wKWRvk9W7tIoPeEvabBccJnNMSCp31r
g9i0F7mof1tNeX8Hr91UD3Sc9jeBIveVhoiOEYCpTc/IXj9nTYdN1lddjPCo8i042dOBJQt6+m3A
q4scpwL0Yrga4yKKDmLVYo6sz/YucE9AoELw4o71ddwQFVNhh+qqJq/haWjx0C4EGfh3IqOsRU06
UX6OhFPC+tjrbvcF0hJwQbqk7B/0L1xAJ7aw2HP6ecPhPZ84RqLfZKdGsVgTze8wIfa8hpjBTPEb
XGWX9yScoaqwbEYZheB8cT9ICbK15UX4eRUthBzviLHe1S0cKUdK25DngvqqqrJWLPSuY/GpyEdx
p3acqo308WFcdXBHyv554EtlgUKJEIfDsO99tUwP7F+X5jYSwIAhZ95sBBdtbf+89WeHbuXaKZMI
NDKkwTMNZvdUzXLgNxzdL2cwJc7Sy5M8OqgYmDmIk81QNpcK/Et6Jj2QqQbf4y/Zu8PdVh0oy2SZ
jJ5a3y0OvPdBwhsif+MczLFWEhFaprmZidzl7s9at0lkz5aYlfvnwAPPKJswjPWMcWbzVpecJgL+
JiE8lbsjkrPUWDYYkq+TyNG8s5t/BGLHO+UVA7+YE2gEY7CbmwEE/Szw38ohXmbMP0GSYT4XXsbU
EQe7qzuyg/pzoYH2OtobYzQh+E+jqtUNsKm+oUI/jJ0ZpmdLmIpZ1pK4puSrfsIho0Bdt+PHAguC
ZTOgtT+vjgAl8xKf3WsomHTF5cfhEMu3lhepZ3lyzOuOCVwFMtBJH4zlkMDjWT9GKenLFWBeHs81
sybzFQHc+xHoNdPGYvWoRHxoJd9Ps5RrHGEWPGbFe7iulW9LuaG30F+dyKbNuSjt3RWSF9Q9EXyf
bnOLVSYX+7QA1U28W+UrWL3V4VmBW70XhI4R12qhLWmDgSg1C9+d7DvOSOFZQFUe5CfmvRM3YIp3
ITzikL78V131Y33szEj579ejv+UCurK6f5afoqMYM34VnNfU5j7ps2HJn1LRYo6BTtFUYxru37qd
amXXr8U1/dZvU7w3D1PXcziqJK15HU8L+1YhjQcEQwDpIbL3uHnyNN813FMfIqSzXJw0OpKLhLRX
BD++67ctVXD2KSuyPrY2rniQOfAHYA7QaqFOSCAPjdqQ1IpGBBDRGrdy0cY7O8MBmrqPws6frokU
6jF/nQeCzMp+wONrmtVlYMGSQdXOHlV/rSoZc0IZXopPxb+g21Ax6/jVRNKTHKvyu/5KbcRAskM7
zlyLcYukcQ0Isqk2EzcwjnBOG2TcNiDDkSELvQgr05O6fg3vNjC6TIgWclDCmFY2DOax/NuQFD68
N7exYdj1IYuCuoMpV+KbL43s2tuZ8/CN5tdm+pFXMrXYxRt701ZQ2vLG2Y3klIj5C9yetE92p4IV
B0ofjSTzp2JoxiO2cI7drfk4MJWnf1YeeounAZ/RZdMacvRFJqaGcUiIxa+0Pmgg/o1Mt4avpkaZ
Ln6+C/yj/mmJ+VHGCSw1rSHkplb1KugAG0/T7X8C+CAqLReama+qjTnFgczpDvmCGtTJqsDZF9W/
LgbesMBl1Pw/Id+1/l4s8l+O7qRE3q6LgUQHVEPpvSQXhbcynIjCJB10kZDtndYMxXcn4kMPrFHp
MIsLRAhUD+NPwK8vb77ANhj/30WxFXaBVQi5ZCJhofFshW951SeFcfhVpHDmHMwg2StC5/m5G6Lk
jNhQDySgbDlPCExoCeE4QhhpRAHwNO4T11GtV0vl9dpIUpzRm8YNPsaxx24sBYzgUvv0ewnEhTJR
kV8OvFZFFIPvS56reMg9i9T9t3Huy/TwC+IfQ1oqk42A2E5kiyoojSPzoeVrMLZ2Fw43BtpTsT3W
pclB4V1Cs8Bs0M0ec/fJ2+eBy3KN3bmlfoo1U4QXIH/T/5bp9c70UKMCR3nAa6u5SrGakJYWhCxJ
Wg9ugp17MpW+A2kREzaXVVVf8FkbddWnay/NHyxRm9fnIbWLFVUG3mrbiH1+0ePhkQdNREnMRlWh
e05UKF4oT0tzoZQWYaeiWtGAK8xQYF/a6OjTBJTFPV2Zz0Hm6iQP2T42mDz/EM/BiteIbP4xKvUM
AEJ89/b3Qc7VEqOR78HidWFU5WamFQrt64F18X3FHLKAAGhXBJHUIquklyiue6SRi5/Z5rwnBOO4
HnIPSa5lUe+T8pebqv9LwqSzlXtCN7bd0Kbl+Fnc+iD+b3NQgd4UIXA+uWE0kBKfcntXAubWhRR8
tQ3r7SZ5mtH3B8SBlgPm3GBTKC66W9+Jw8sprZMudiUOeF5JCaTheftSvUme2v1iuOFxJJZusz9j
3DOemWuHIVHj0rOx8tdIL3XYWrCA1diZBHkHKfGqWklPx/lLhUjJrSgtdsuqaY7uhcSu+gDt5XC+
psndCc0qB6r8ANJzOhMbEsLPaeNvIn8unNSnNHr6s0G43ju7kIZ2GcWREN7CvedOy91XlFYOh+s/
cGACNAYYgUIXu1RgQw83NoaBi4ir599EYpePH8Li5f7B9lwbQA11ocaVtcYcU0KSN+00NyehvqlH
ViihN6JxFLckCeDMFG2TcHVaYDxY5/lmVUSxmCjHLynso5+8gdndDvclrx2StMJPRm4SegScVYXR
WXSfQTpqBVJpn78SodHZh9kkVX5M65DrT9SuOFRbP6V6v6icVSKLpSSikY9egnDE0Dh4/CtwVfjV
08m6RypLL2nwIRO2eVduMA4tgnyqCtjiaxOt6XkDzg+BsJkrNe3U3hapBR7Ia3oWX+TYSsYd34GF
6+p7tiDf+p1IMp7BLPhiA17XuJBnkh39vtKnbVS5iR7EOnDSTplfiVnAPwNYymesy16T1tnAAT1r
VN5dCYRvrCRY8pADVtfuXDsqH3Y8LaaEX7B5ME8vwSlshHhUKeQPGX3OLE7CkG5bKNPhFV8gdQUm
jrbcxxQ39eb2eRZUgy+GocGSP3PVTYhB2OFbocJ/olEh9uYgTDxda9QTSxs6H4M3O0W89L+CHf23
/cz7OUOTHQv8/GzC+lnE5uwOf63eL1Lu8JWpuCJBSWunnjZAINpkgc6nlseH/Gx/RJCANke7Cd4C
eGxHaQ5fE9Sm9SpLjwSWGVEZK9UAgFRClvxkNrGesfVYn66cHuSXZUz6hl2fymjQQ2wFW5DR1ltB
d53nefYR4u9P00uGsyqMPA+VlS21d7pITAJShEX7ztpg8sRcUk2UHSxM65f1Md8Nt7Fk2eweo9W2
H1eO2FFAcjbypy+dy29mo0qvBKFJzWMbCjY4jh093DZazGCGiXDjyXjH+pWsxmVLuvRCk0fXd212
9U+X++G1zxFfj5MdC422hQKTnR942rIc1F9XIouyWVVoiDgV0Lxc0nqcZcIzS31QiP8uTS/GSzoh
ySlMDDB4zfdZvjUnBlm8X0qR/TNYqXJ/FDxIaS7MaHTXeV0siYVnc7sn9dzQqmLjhusjylaNR1ou
mwdsFG/VEGsfQq6T0rQcdxwKgLAiH2mHUGgvIap4eYEgw6PHfj4iB5lJ2c1Ad6OKpimCONVbWeb9
LqJ894zIne5e8BbMDf0C0v2ceX7tSkIfJkI+nTaquHrVEhmUcQdOWmdVpeQnOsUf18gPGqh1fpGr
C0E6qY6kYKBb5EzGJJf1ShTDBj+Y8Xf71tlUy6x+2S1Z3sACukVES7rHa7xwiutUGLdplTZOE2bQ
l4W+GVxxqlRwytkyI3Ph4HaISO2Txu3Kd247ZxyVf9K5pIJs0p2VJJF0lfY3NKke6t+Lb3i2oA+H
QdAsKECc4bYWIExASgISoyS8hNo/vY++Bj1n108WRISarEuNqESvQ/EkGY+Rpt7s2VdFYvsL58VM
u57xyceDq+JzRxfl6mhOUuk08jzkn6gPtaQ552rrT4LVb46bvFE8vtw7nXoSHVscmAs+B4o8DHNS
KNBg85XGizMcYwXWPj8HTXqPIL+dRGaJ4bk4yG0pRVuk8/LsCMvNy1h13BJXq1Dfja9t+PhDecqO
ZMbUfG0LfYUas+zdtFwX3xS/5Jg2aSmLLbW8HCpX3gOFyON7xLL/eAswIHP5rKmrMt+5/jhNzres
bvnZW5//H32MuEidlsR6Jhxzsss/vWVw9wlgZMpLmEUwNXGayYsqMi2L2Wg7AJOpQL4BjL3uXW4T
2iXLtZia5z567hv5WOyETqriG+p7CaSGNB5PCjM6NA3vCw25t64JO8Mk/kPI4mOW2CESF6Q8CEdO
pKmlRisLglLQOxsOh/qSbKtLNXxjnut7GsC3hx+++58jsi98vzptQRGZvyfaTs09BgXppmLdsutk
pPKOhnv2K7jeiZWxRHQ2/sTh6pQ8wuqixPuF5/9VVcybXqs19/ekqlHGr30arKXnfqvoxLHbN78p
MKEJIAweTONfI73R/LD2n3Ada5o2nqpg8F1G4HjbN6Ob04CY/fTFYDVu62cuw/WPcuP4DItcTnk5
2QH2YQcf2j2uAtEZm1aQ1+ZUwvq3A1FkvR0S2195zYwu2cNntd+TNjAlOJwwGoJxAyxuJgzxGsrA
M+IrdM/LN+nzqb41L4HQprcDscAAEjN3mPX8EHwnnhj7xJ6IwkfXdaIRDhT1eUE1CgpBwPtljk6p
N/VIqWwsJZR6u1IXd/cbpy6ncEiputqHCRkiprGu8hl/19r8kSVS7OQlykVegxSn/Tq1B1hTlv9d
amre7af0z//ZZOc+8udcfJvxDpqg/hftpXYs/eMP7fjxNAwX41Xn7vXYzU0p6RchKMNM0E7PIqT6
vK+LWb7Ezsz+3nitwMsvw4JXy7xyiqM1J0zQpF0tb7xW0GURcwwvkytqhB2EBMUoAACzMTuggwV0
1BzM/KLWphoiG4WGfh3lOQouYq2cG7uY8T2HHcl02V7tn9fTaVatRwcNmUPeX7kJZFIZpfU26YKZ
e4N3aES3mGeTJwLpXlIHh0H5ln55Qt6r1qF+rbdmsan34vZaIo/in4sWI07BKV3jBj8x0FwvrlEO
H5PAy6dniu/Orlz4fH9L2lEqgpPlhDl8gLrWsSZ3bslHFIpzndZadq8DXm7PJRI60A5gR8WJI1Ak
TlugyvrWZTkxewGzaEqxCn1FCsg3nnes4L3/P0O9OcvJQVjlZVc8QXJjbg/L2noGAsNe5rU3WjnS
RK0JTQCSCCTOiCPNmbENngqSFHGtYkK8g8JNCYl5uuhcur5wieDwniy0XLXCqkwpUWn6uosnCFnP
4N2rUwOsjE0POxBmU4/fCKUsvNbGRlIR0T7fwAqG4HkWiHRswXqJ0Z+Cx6y6aGcdkMcsLQcmWcC4
SuxYzJ76MtdA6AVxhUOUS/x2FqeWBm+wcml2DvLtJNNTN5glNSdJKQnlo/nYjm9/nsOuziPL53Ta
9VMeOumFTXG2SNg432ITwsgHq2S1Gw8WZsE9uWy9ABUx758VasBCW0NGgpzS8yrzOHeSCbKW/aPt
hrHrJo3X2LRspc+ycMVjEE2yp1newZcntcEjBVRk48xrd9IRotpSpekQ3QGYKqyGHG72dlJ6SvnV
kegm5GJIXMiswv0ArUXTKv7tsLkO7Wgin//rcBmSyWOeKAIYlW4ENTm+tNR9zhwt7PGj4i4bHOZb
vtCuwGZ8qQjNFqEUNbJk89iBx5O8yWGHqyT+B6fYwXgMnXkMLs73uk4i+H8vi6/ZPAd8H2Li3SNt
0NS4+0PoE47bxX53dy6Fe5UqN2+kKpVosfEiE3d8MxR9JO1catGgtp3d8tdvmH/0yKIozCrKngnL
+KlBTTqKEF617B+DvuWd9IQVTOwnN0c8axK+vqnKGsqp3jtjjIS3V6Imz5vu2FAeuewKcCWxTj0P
8m3879xTqwgvCdERvmh7Fi4et4vzzU0h9xJLv0hwewa4P9bPHwkMNq7Rco5fowv5L2aSn1dsFJg/
5mSE1PwNTD6PGgxptBDq9NTYmz+zaqzxyTD/32dvWneMvKsP82entXjO1Z1aBZxy1UQ3yC8qOgzk
2jwYbCncFGZlA4LzRdQaFopCks9E3sUSvGbf8hbRyaNmhZg7RuGAMZtKCy0VOXWNGPbSN0l7WqC9
pJkkBVcLnPYIPEnYFWzjmjcP0gUXoHCAO303ZbcOBB7izPg63zIWScf1y9fradXQXlT10HmnNUp4
FXP7S/OeuR0uRS1BkwN3Nm1ste5AWZYW5PhaTf+KkNuJSBXcoqGZ1djXxP41DWLx2NFXM/hzkKoU
wa5sPxpACObl4yjIM4XRzZ+hAJJCxacLyeBrWK90HoUyUWQ6jYuReqh33eTx2CeGuu+ZbpxWZvT0
ffG1d+x0OH01LuLvKEWhd9TmDqYjf4axBknnn4Uj0FyDO68bILD58sDLqfJcnyupPf01PXTneN+z
8vFKfz12FQaJT3NSg+hWJ4BPgk+9aVfsNJgIdFjPFJ4B2kXBEs+MNRebDPQfHXHZ0IhJg1tHFEeS
pWZ8xla+O8nJE14+V2eWErOSevJrHP6q438Cv9DJOZJMUy0Cxj4CkZljot1dMCM3oy3bqJBsbTA7
RG95pjERa3VMFW3NhWtYW2lJ3WGclGa0B+KdyQWSqJPMZpQ8BZpwQCY6E7GSDpdM2PWtrV6g/pyA
p7/R35v3tZ+9cz9ZrgubDIHBXahMYlrwPELyKZD5JXI3ZWfZdKjZo1VxZ+2D274ROvjAXl17q2NA
Eccx5kdkhBqveDMRyocifxW1Im3jLxaXLjR9DQpWGRiWGHdKX8hYWtUDhxWRNZDbuPOlOnleBI0g
jghkp/nrZDvg4/ane2Tw2CIBQoVGWNVghkrMKboYqyjlI8fPZRGV2zjpU4zg3u0pNUAEDWZVul0P
hkQ+PF1VxYktM1uys7iHOLh8jD9q0aLAgp5XYDWUgnfF1oKdBRwbWFDULy/2zXLoMuCIv3cqcJrH
uu5MjZClnRFgs2TRdzj1lTNkJtjBe6NdBPkPx9dNqu5kFGlpCyUL2Lyv8OImWRj0ttl8W5AsFFNh
NR3/VrURqXQXvBexidKej2/NdrxiiaIkX255lbgQOHwc6hujLv2ldFFGhPlJkDj9HGhiGYLPjaq4
zDVNN3cccOmidpLTjHYmpT6mDdevZl/53dAsBai5s9s4bslc7kXNwkNCM0NbjXIwGvo+UY0BOsYS
PzUeVgf8oRJVtwyNuH8oZkwNtMylZ0bLTf8xKKVn/RULbVh1AeUP8/HQFhHAN8A34PnWWURcoGr+
YApQkkzdlyHKajvBeWdqXveo0iWvU6kp4+e/210kk8Xjxd1p1W4RBoDNuk1XTx8OEhn4aZkFUqJ7
W4Av4qebqdW6sRu32ilt8OfdiNOulMyW0kMy5qpLGovvECRbMTNflioqPAfd86fXFiMKUo2c6wYY
Ofpg4hebDXMCS0OEoms6CK+Of3FnOOnzXcvaBfgubVHSPMXKAsmGM0SVg9EqiHEsfmp1NhhMFmdN
Rq8oD6V+gu/ekIrdHiph+sankIPCxUTzJwsA9UuqVzjNKHpngCt/BSd3LrMEpuRhQX1LZfOLrQXt
8GgPSSrWgekC7GupkOEUaUZayEtcE5LJJ8Wud3h5y2zicgDpEJzfAbmlC3+d93fUf2Hqu/IJy0yf
k0DN+mKQju09p41NF0oc5HtMHiyzhNoEg2ZYrfJL/eSVpPyqykq2tKLL9ggQNxR9nwkrKGwQWev0
iDlmhBlCPScwOtvp7FXxwVafMVwYDMeNAv6PpbX+1x072fkeNAe/YIXv34nMVeai6Zjwa1x7p0XW
3l5d239PoeahEyMX4pWb/99OGM3AFLv0vqraO1xmI1xxEzS3Eo7YT8PaGjNp06sS0EXCEz4qog/S
mSaeDR/UBsYS8LYqVK63UEEdOWIEyleukzMKvImByhAF/F0apGx/mYpD72sSkmdbsPNTAWrNMzJz
8K9HbamVd1TRmL6uzamCnl6RoVlxKEt6AxUVNMHVRORKTPAeyU3VlVctR36PG2s3oUWOuTziAHeF
bG8vis/dTVfXIb626ssA8vR85FZtBZo3NlrcUz3teQfsQwyhrN7nWxRivKwY/abN1hdHE2XPg8WE
gIhwd3nfBZvI22Kh9vSEhWUO4C0RWiuMCWwzY3osvz0WGQ7EDkTCtfXehg0dqjaZpjXwrJAkpLBu
s/WqnV1DHo8RNz1PawwmKh5TB+UnLxkCIpL1pv55u6e8C0yLEc4tIqYm4Evq5PjgCw+Qk3diBoxW
AqF5oxCjN7Ib8J3RqEkVCWy+f/nq4JvFcBVJxpTnNFMGa7zwvtW4ikO27pMn14BlS8IJWbEGjrkU
c9TF8wsK2r9rVdAl6PkPaCtB1nfpBFEbNtbADwbSVA9UNq4ry65MPRIRfEPZawHMHIRENolFNOzE
VKEnR5Fxznb0Oetxt52ADpNcSOVz4+DctWH0Uc/reql6+36twKGo2FXfeYn35csOZ1zX69SW3XKQ
L0FG+OZccqAkhI3c/K0n6rOIJxTzG6O9qNOI1g9bckrBXGMHOQUtst1KYXQta2Cg891dY2c0Ir1H
1OcPyjtrZKKIddQM3G5uZ37mqoJm6f/CHIbtFxLUVlwtTtkvp7xJr9zO+95NBTyNfY4xgJ3Slahe
mh5xeJzF2BVbVqm8F/UmL/PH5d6D1GQ5UFBdSLNuUocxKnmG/9EFYis+Bz9maMammv7+wW70eJP/
OswxcKsfaTZRQpnO4B7NXGoGcBd3yfG3WTi/lM1QERM+A6JH55ds4VECtXRrmPV59DRABJo4iSn3
l8VyVYkDSN/xt004H+I8/qXie381pntJyx7L70Q1BGPGC+F3djuvidDTDdtrejNgGLX8XFFqaOyW
NWrPFiKuQvjXeVxNIArl143QGQ82tmwyqv6WUBzvmmQgl4tSkPcRZLfLz528nLP67UD2uFxF3duv
ckRUNYrayxszZBBODLu10OVpQ0Pz3z6E6Pyr1oVFBL04BlY7vXvECoozxdH+Ldu9zGVQrLnYuyhV
//TIX0GynFWTTLg2VV/hIz+Ulb3QA1mzJCewnv/0XQKxj8QK5Z4tEWVGDK42pL0z3U38s0b+K7Vk
baAojrg0kyZBLy/+gf/yavUkz6clM5+GMsrNXH9W7BEzcTnVuzmsPUsz6m14Q6NkIjFIcomJXVnI
8RGEnqflBu+42R8L+qFLFqj646bSTD4lXtA3VIbNnm8payDJ3bFjjRfhkFS9L6NvE30fsMzygX/k
gmjpugMxHZRii4o+M55GnqPzU+L/ggqmLAQitgP5Z8fz3FFz2vXT8IXFZKjxSGvlRrqDVdJHs0kG
IBEgT7NXNRNraZ0lU2Aiy38gabtmuFGFEyxnTtVF6RGxvAxjx1ZR2b0zl2i3KDe818rbQN7GmqqI
uStz7p/k9eR3cPEgfdgRQbHg65KTe+YaQPYuOmZXp2yjEy7MScHLRmra1Q9DYhiQPpA0a4BAfxMS
nKCWVBfKzv6TBvzeUxjOXqfJ4eNBXhEOpfwqpd/klq19AqF9qcSrPsupvveEX3jog2JiUOSI+Aph
VFGqEGpVQxBxYSkr5p/5VSuBL4WMmSij6DZPx+PVjdPxOCsuMOSw+BzxkQD3GDEVCiP+/E1BRXA/
EpuRez5tyG36ri+Bp+vhPboAwVGRrp1MJZysGR9wvUTm9MiX2u7L2KCf8FfDGZ4qIOAu21fJrPwk
me7/i5NkFdCa1Jo0hSyPfmGbyRmOxq98bHP2s9gjPbOdJC9fC9XH2sVyWMKimnjV2Jz3Nj7PbuJP
9iAdI0D3mPbZtnVrGFf2PSacLupozbs5xCBU/tPORHjByVvDgI0k5IJC7sGiuC2xXfoO5DvwcLZp
xEM9Ht4zhpaBlIVlJdeg2amYMAdmUuCeqdFpSP+pjaCPuGqbBDQLv4klbkYo2YJdn1+TQ6QtvP32
BojXikNSAfDlv6TKPqniKMqikIKYyg6rFwxtH6HzE31oNDz1JkHLkAhSCful/dfX3Bc5RlQuvgyO
3P5yJoHbfRTU+j147X53RwTchR3xMkR/FfmoHmL9HFGgKLUA1KkwAlpurttS8dbutKecf7TEyitf
YIpX77qCKpQT2/XtwkfnVMPDH0JnTe1hQXgvrtrDtW7ticnmeE5wCKZljgS3awTamHHr1cNOy40o
a0JN1TyDEVuCKz/81ti/XdmhmNb5AjkeYijwkKg1S9j0WmquSTqCwNyxFC61ntzlf9NBvVXAZ34Y
uPGp3z+ygT+6iv+2TrF/iC6BEwzbavudV0/BIXIeB/xiB7dW11S6rJi/gfSBnjI18CjUSRYeNuQ0
IJganOjd8uJGuqkwHO2ZBaDq6dePITH6cQX+qH/tgm9uakhmf1q5m/YknUKsqiqIihp4ZPVMPtV7
833WchpJ/G48z2uO7okVBTWvL0dAD3EmB5hQHX+Q4Ic0mO8J0jILw8SIhTzabO4hHGTig0zzQIfw
3IhsJFCObVi6xLXXCe+34tvXWGyZvUSnfKnF1Z+isLxUyIYtPmU8E7AtC1Xv/rixEWaXwJ6f+dGR
qqZH6pp0yKI8/TOXekUTHK2OJTOzknQ78Opn11SLAsyEcIXRAVcVxPSrKZdGbiE29m7IN81hrMnt
ko4TL/iyDvjc9iGugOmmDuQ3UDl/jw17FfQ2iu1t0rbOtqYRK2/nxh3MBJwSn/EJK1d0ARcAWtJC
64dttaUbaCOEczXUPDNtiObwlkyb2o89qWGuVVPNqRlbUrOB9RlnJOge8rV7mnbT6pEslCReHd/H
Yb/bAjHZAg0fUS/sfoG3upMPsLYrOgEDPGlgzmbFkjetGsofKz+u84QDVhOmXAbToSpIdXgRAOYi
tXcD1kkXAPmoFbYlfdPjBr2+oPgcDjexFieli4J2HaU8TqxueE/sU6mtsLjkCR/oN0AtibK6+16f
zqXRw5O4oG4xDRTjYReZjxVkCIJpXxjpniSnHiJuaJoBtr34y6F1NuruOpMPnEslvZqfQ1aPKopL
rTkqdPH7Xp2ANGbCpq2YTuua2I043q+TRXMX2LbGsHdZOFpFYlgpo0/swqgi1b3G4NfUkQmzlF0j
ea6vFgb3YVYMS4BqJ2wTJr9nL5nBk+tCWYRI16f6JmOVVYqjJJGwtGp05JlkvBm92YW+KEI04QTe
pbyhBeqmpI7M7wmBkreKttqE/Aa1fYZ0pegfLEx+0+TPai6IAMQpZY11QXDoUJlcf9+dRxZG+5Vl
a41Qjy23v8DIa0x/Ch4GqXfvBVWO6/uqPtXGxo46xkxabLn/EthzuK/6JblH6QvKGBNLXrtQN7Id
Asbm5/d8hu1OkHiZUhP54SrOK7/rfioUdmMDVB3RZw7sErJ4bO9WkKG/3Zh1TGam0gvS2uGW8pbC
EgsoCVCfLb1mVikMtZ384scpPlr9s7kbSzSvKzGvYRDyUwM4EvixfWq8bBtsrgcUKCXjswc1dZi4
cm1fwCVW1g/veWVN6PdDhrvpvAX/HaX77MuBdbJmQNqAN8wTzh7MONw8eFoArr9HJXAPgF7MZdx8
O8Z5IP1S+iKpcJaHGffZGSIKj/f5qhAg2D0V8mkTh/nSe1sJsLhR4xoLl4feGIB7+9rCe2P1w1E9
TZNIgD1YOrqAad0t5ceb8qS/ZH5a1KTuEa6mYeWAd9cFGAHJ5lTdYlB9OpyeGGH7iNUDxg8gYfFc
HegKcdi4OVrKBtWMsNk7GBSBqq12+vIZe32XgyOdCP+X0OOl+f+08AyEOV5qAlWaalrla0lD4em4
986ZtPwAzbifOMOBB13m/QUzkjk9DBXejAioup6DId7xbTTMvaT8v1D1MdhDO6LgeQAUIdLiB78i
3qoG0OBJkCOTadZKlurejO4i7Fv6P6xgOaFeJDG+zTxvVKDTCQw838piEleWGh03PyyRxCLiaIGl
xJUr6xemgXA6sgXvhNQl/T+fyhy5YV94eF6jwncI6PEHcJPPIYd1QFmuzAUJk0UXcs5R237EKxLC
Fu4V+ykGlPXGkCKwI6DUb4zRbnDNqONxuSLrgqcDMbq5SrngwTRHP5Hx+0I5uij4HcKcAGX4h5PH
7qLkSVJ6qzwjRbnDKQlvM648rqfY5CzVAbxg2ORp8qDoPrpNrOR2llR+LJ2BSIboXPsfTrejGFJd
0BTAAZSSvJWTu9XG8QYP/B6OvRzfA4x6W5E0agn0v8BsCyzYDFeohc/zQpP/MjpU2wD6F9bk6KM8
ZXeK6gCfy/TG3aEc4dLOyPrNcBVHtThzXd742EvNGLclYNhYElBIe5XdkhuYHp+m30iZCTwW7qvd
Zm87qK8FtSj0FfXFk6hEAgxhSpVqY4ISISYk8VrYmCaWtPEh2ffGJQmhkoLfDMtVSLuTIiUmmwin
vBWvYSkvFuNohkN4rSOvaWqKxctycD+jeHUF2bCaLjJ5IpcFGQqNqLBcEzt9h6ORD0ikq2j9V3Mq
w5QmW/snKdHY3qbuTS3Dbq1b9eAtjKstFhV+hP6df9S8SuFdDuU4nVaCxgFKKjJe1o2Bv+GGP+wn
37bakeS153tp0scoNQnzpGZNYoPB4Ltehi8K3UMuWXnN0Db29J/dQTeU4Ji2aBjm3R2Ft8CzdIut
4XApcMRDJN3SwXidt3638O1TDPnMlOWf2aZS6+VsnXNAxEGvamvztMDZANcL0rgUe2NMJUeaa3Gc
TLyNXJ0kzyfdFMjlUQcUg09e3ZEuhfE7bkXW4F1Q1KHDT6YvjZAaiY1+va6d6lO2gw/rqtEmAA13
fxRU8lVjEcoGBqkxuwrFG7PxdW+F6fr0jSEqs8gZT77kP0Nk1qLKaEQivzRW88nL3vmXjn1700FU
igbagxIdpioHQoMfyi2/mWsxUq8lTSSXZsYxGF4arxWrTCjW6XM3YrUe6kqQvLrwt3Ve5zFWw4Pt
aOYS4QWwUXrijpbHi0y9hXVMC1JYetAOcnx7yiL26fJNdnC5xZ6ljafmmSr2dhr9bvln19QS+gIc
xorIeCL6VKHV5QzjSHoBhPxWtZrrw1sOvgNjQiNZxCA45b9JK4dkl9DKtAQBJSw/e+CrhGDK+rFd
QWTdYIPhcMNUS2P5Keox0lbF4SRSGamlCG1XtUZW57O3o1yq6ejknt1u94GEXtrHhqpIwVcw1mBF
f1PNB30TKLfrB+Ncj3fkvZHNAJ5NpcZnsEUZX7RZPrKoDRA+WY262nNT2Pg+5Yek0WjUmk/Ca1k2
tyb2tzVpbfjrZ+5AWVzWMRf1R6ofrI9sUXQfyvYJcaDnD2zTShkZ0AdBGIw+PQzYobsyeV8/O6Ch
PKUV1ac1QM1UHsyZitztLuMIINgNb09LkvwnulsZ/RiT7xiyK7YgPPcPziIqq26KPFRyEoxOD1BK
3l8dw8p2RCjAjHhQLaNPpMYL2Q0DSIjhLoed+XQON1rm38Ty7UZUkNkSDsSeHuvLZYz696JNusYt
7pZb5cDvJjR9Sl2XOGkc91BvGOaIM/Yx9mHA3pyijXqCsTTy9EwhPOpxg7kFsMqsAZY0BqI7Hdyh
J7Xs5NaJ7x9pwFPUIA6uGyBjCvCqH9E7sNzqtt1GV2pgbiaR4IXzV7uAaYpo1ddaJ6gUEbLEm7b5
m9agfBlZ2hkJUBtmXp2alFhWf8Y8GR1xTJ0aVo5DV08h+HheiUTzSKDfw/pjsSnBRDMrWn/B2Ngx
QFhO9fA5U7ikhK1odsDT8jqrygGLo1J/uxucFOIct8TAUmAxHDs6dIiHwTqHuDDZl6vH5Xmd5OA4
D+nXQ2IjijOinLDOHSatmtP7PxFtnap7DLLBPHHa1SjFsxYT4oucPffPFRuF4Kfe84ppaO4G/3J4
c8Ld3HeyNtPXmvl6GyK7Nu34wI/bsouWv/M7vmehzbS5rRrSSvtgWl1EmhIqu6hGskW1Ma7gh79l
omHS4Wq/zjIBc3OLLKWtBJeTJgkip73/YBOyBmTBpChJnlyYNxAanKzeUuadb2Btzxtd5Jtp2AOk
gaHijQqt4v0YFAPCWFvxyFVeYZNZar0vrVpCq3ptPWZXgowt7hG7J7PMk9WGyA8iUmSMXb5JLsVr
4KaBI1He4RZvyxtRJMF/zwdLr3VMBQpsO1wzRsQA38NDDLFeNnDg+xeGqc+Dz/t0IX3xTqeQ7nTW
oLeap3eA3tJy9YcG7rnPPSx0eQnzLOT8si9g7+HnGdFVkoCqkdNMdW1qNOYv2ZN3qehgK5WYvAmD
IO316Q8nPn63eFfd3Z6d3zPNDzJzDIYJ82ohld35aMq/i4Ke9pqkVZT4KG92NjxZVoF9p6uh315t
0cw8ePdkmJng/DpBZlFo1z6IPfU00tmpZGxvZ1nEqJHEXl0h90Nu0eYb+mz7CFgqI/9E7ndir/Xb
+HyvNe2RcX69LiLaHhzl3yfYZ8ThjGy7/IXebtNuN0/HFjLHWE2rAcvrWt9n98+CPh/cVIQ2LLPo
vr2n7MBeFuhw339ir1yWjJZn4jjdMa9cecOCAdv116BhhMkK9GcW9EGiQ0EPBWFchmcBMlgQHR6w
S0EbSYrgFTI9FmtHFjH8DEH6V7wSFsB4wxBJLCYIxpQbeVHKPmnpKWTCycaJDprGnFdICQV7EPhP
JvxQ7nUvy+Lwmjmo2WbVytR4ea9KUcyFfhV5nGaBKqSuBRE9E2Ry17JJy0QS70ok6DkjcB3GpQfo
ZCwTQZMq0bHqUwxIP7jkMwyE+CTyG2vdyxdfN+DEMFsAG2NLVpbdnv885NmhdvdygufdjXqHKK5W
CiOPsG+Sr6EJH3kRGhJJ2HXfln/uYrrAHkGyeO/W6DwM8h8FPWNA3uCQ04wiwEM9O5QuV0Op3ZQD
Evnd8c5heGSp53aSXkQalECcAOiA1aqw/J/qYbi+6malc/h+VB/vBsCD+jFWRzKmDqhSX4PYNMg7
AFKvmNFaD8zZyS4XwSnJJnMmGgWXhEQLq+7qa2078/arHBjjFVNMOg9YUje8J+y5L8FbQLyZfsiu
Ug7tIbNxcpzhj1CIF6xYy5y/RVfaiBypGZvGKQ5qeVuwrHXySS55bZlUPhVtgn36VY6pjl/GqjCC
5h9bvU310sEqJ+K3Q+AXs6FPSqXihMRKEf8r73dg/k1vozNUJfknaCLNvDyQuQgaf2G6hBXLCJJ8
1Hc5gF2KAHNexARzYPo+3tooECmKKZepiq7/cUJY5brR+l3BIfC4B7DPhVqPIA0Q2NcXqQEPmwlH
twEfZ7KT2GRkhnP/AwqJuMNvtrrFm1J6dL7qmXz4VQtnPRnkKITmTU221MDitMTTC1yKmZKVrAIv
aZCq1jk/vttdSfd7/aSbObnlgyY+Rpz1+reCwVel7klxkkGx8rDslLpY7B1blLpg/1RCCqG0MQjq
hOJl0lNZjZP5aVSdPyRkZ9U1z4fQjL6cw3vanYMsBfldx/qA2t1ZDn2Rwq6MjYam8fGEqaZW/JRa
nKvt4NqthTafoUzQZGYsEc0ivdbZPu+m6IVYI6Mt2UmWnfoon2tYRm7J99ULxSFIzzDED8kr2uSJ
ntqDC2SRgUanJln3XSb+GxnlwcqIBUvyUwRgc2taG0w2N0zALVZFXe7Ksulg/n25ZFt0bLL0RUOJ
YAfr9AxN1KN0ZE/cLsy8NMmo8ZeMG02Q3YFr2oQqBNtgy7qNv5jXnF1lxgW2ubUqYyy3HwGLqkrv
58Mdj+ebagfpjX+ABsmKqwix58e9NK6tboV+pjRBmhA1uuyTzKZEBZfOEyQOjBOfk+1Vg7+VbzA3
w7qeDIgy5fEh7F08VqPrVUfFNyJ8N291M52feEmeWnHNlrvg/g6scw2t2ScEKDYZWvYDAkkR2RZw
zlvG5NNdnpxjq92mB129teQMKWSk5FzC55j4KID8MeMn8XaCMVXUkgZ6++2mU/w2o3U0UsX62Bnh
uktycq23s+4kKi5D8l3J5xG6hz4lPqGDx4IqTpJw+UaqA0bHyZiNgk8dl67b/w0RLj6k/jfl6Tkq
q97123baZYwYu/RC3sLtvSUm72v5Ay0BHFJk7GEoCD/jNj5MUrELXFZCAaoB1z66qitGagyY97BD
CIRHwAauipxXZ0wsAwYOWCkZZ053dWOfojxeNKgfDX2OmIsnljZCZNwduFYCnW9NG7jTFLM3QI+M
qkAviX0VBUD5dh8y7sDKmTwOFqzFCPdtlXjNj5+yTdTWhWRGFLiAFH48V41MV+PL7ekdSY+VihUs
eLbJiKjv3OHXgpGO7XvnCyehsVtVB3yVPMJBSheHrSDZfz7hn08HmRXazeV86ZLx7r3vncfYeE5Z
b0WmkhZz52sUrpCvtvrdOOrx/+0qQJ7d0huBcPPYDYJgkhyEJhoYA2Izs8yqDLz7XATAIw/gqwHF
8P17vCAOvCrxJDiR7rhV0ZIlRVYgvaeYkBcjKlgohT2GXYcJneu0bKaF+ph24SPSF5gsBLLD4Idv
mJpFWmtjGIEElXxCJyCWQ3fn3xAGRPAF4+GVto9kiCWeFrulxZ4P9U1BMot925eZ5X/Uczn9lb0v
oD0KxcIyo3ql0+gwmWglY4iyQQqoIMCyUzMwn+N9mqNjwGUmee9iKXIgYCe4imDebs5DRSVHGFTB
f5+MxM7rUZkhv+D0E2Objo2ECq10yEfmpsYj0n01ZJBAGgLjYgMxg3bRWL4C7dkzZEp8bH4Y9VG+
FlzWQfRdO9+HKF8bKF9GPwuW9ng7Zmxuob+L9IMuqHNsgGormP1HKZBByZLNkWU+tVKgq27qKPJu
SODth2TW8wJjOH3KBylHtUqyZNXHByVLa6O5xKgCVV1/uwSSYrrg9/S/tWz6E2EtmdpaP/4bdUL8
7bYcQZnzFsdM+T8Uoyg4w8FYQW15MGCjIIXQwngty+E/ZQOOhY7CkrfcymZvkaqa/4bwcDxPR6vg
7OhsOleIv3PNhBWEfN5xFAmW+RNEttyqxQM/495GQ2upiI7eaGLJHxy1bQEpYHhsF4AyOolGILjS
/cFk1YDNCFu9UP0F8RhVe2IRoG5dww3BLVmjrhw91kDutzUvKsVXZPQsAj16gLO+qk+/sWOqYOcB
KAQ9gtU89aQsnR4ZCYe8nY0XOA6TsF4nIVgVQo/EcbSd60ztYGYwi9g4I1VmI3/Tm6qRABDVx1yr
eQ0CD70iT9n6rXD2vJ52lSrWR1dXTSGFiFX6S14crBxblDetl8kWIEz2G6DJmia1OgCeV8TCj6ip
OD67zUvfxwursuMiO+hloFUrNkVwR06FgFCDhudt35pzOP4sNNaLz940ood3VbiFfd4Cvv0N6yDb
7CQGIFFIVU1GmeQSuTXWcsuHgXguQoZ/zdXOK9qPVZwkusgY4z5weR/K9P4IgYK1flyIA4Gxg4kB
LRNwIS3vTeoVHCQS+4ynK79u0vXM5tDkVqUnyB0TVJ5vVJjlyGBjAM6MjREMV1PB/jQ4Bi4JI8OD
Kbu5RTy3V04TEwnf15mix7Vv/XRI7nTYePiZX10kahX3TiJfUsaGL9cSsEwbO9ePrWNB5lRA/Miy
IRx+eEQD9akyWpScaBiFVidOWKnFUCLUgUyebMeb3v1guZ5ByPD+nLQuDSvA4l2CC7o2d/lgp9uh
3YZK5nF4ekedA7fylah6je8kdEGdUA+yZXuE7OOJa9Htk1EBhcqxtIZj32hk/1QBm+cLusS3rmHf
tEoDtPmcDZ29CgH462XebGpwETHOH6oCNHa/tFJzuxUgMmTRmFbLVcmt6l9vsSsqOVU8OGiHIMNF
TuPmHFN5SwKu/U4vnvu44+9QiK282Ormvfg5UATz1Z+kvLyyBpc/jCFZouTmYWBPPGF4EQNRh7qT
rL3jkMafaujtD0nOleSyn52mDz51cVqRTmloUwn0GExWFcTvF7ocNitr8fha/yHacEIpkYRv0BGd
zQi9uPkvc+ILhyM8Tb9WnC5ZAuUvpvPtQZBva18yqk1ztkrQ4QhABE9nhWCC9u++CszMmKgHllPg
cGgK2ihqQ/hruNbbiOdzOsEFnTvLAEbz5MVa8/vQb4ANCzae0magG1inYX+XcpZ7gnNYepvWF4mu
qDHxHHzTgPl0jAkDXePpgHu3TPfXogG+yLTBjXxCXvNCXQ55Nm0SMbHR2r8ulOr2C8L0SPsbwdHK
npUIELzIetfPrZ/idTxuRzk/QYumOP4kBg3MNFfO1KKlc7XUllwqqRSXKXgogp3WJGeHWg+Dg5cI
uGuMS+xW8Je0dqc9oCd/koGQbPCA5kVPN7c/MFP3g19V8/wNHVGCO+Gw7n1ws+EL6W9PsXe7YIVn
tpATtoPVlkPFkahHA/SMO07Ohmbly00CB4PH7K1Xn+VOeBFRGaWg8CcT3kJNGaJtdeG5HldT7GcU
6MNUJGAFdpRD5JLhqAroAGiqnwP7SAbffA5/TNzGEnP6Z5OMDD4ThEjUC2sf4qBs8w4dzky0yRj8
eQTFSJDfjpYZ0TcgLmMp+CzNNZLkZ/uV5VG+RuhuXnLTtBYd79iXe1SFKbaDx5+flQ3fQBsArrOv
yPjAfHghyCHSOswyfmggK7V+C80LlR60kdtF2upwmpRQciYgwt0KY/ykdOTIJ53Ys3hRNIigVTl9
UZ0wNg9t2o2mTWOYJfovLHVzSIeBcFVeRR79VoxqRgOk9XlWLBD7HOQljbnE7oZcKCx0klzfTtKm
5eCp92cxdBo8v9UpLpEQip3c4l4xGd3HObm1qdQlTwAFioVLHVpbQ8XAeGVqv4RyK9d1Dl8/iXmr
SsJvCi204qzyTDfLnB+vgiw5sd2RMoQYa4TJJy5K/VGnn/lgF3lBdApi6TZqaN64triuqjd7mmHL
wklXkAyZTduvC9QSFliIVGDSDO4YSuuy2il6mO7p0C9JDCtI7tubnO+nlna61w5yc0kex3kzHt4s
91y7Z3Ld9rOvNv45EG8KyoNnl4pcirjap+0vW1oNuXa8SWq6LGlsUd4csTGCe7WUtTbbsKhauNPi
Y6dEBCXhmyayFi1OxVkzZxIKASmcag4dgKXEuwseW0U+9EZqXr9MQQkJ/IV9pgonfn+UpSuVA3o/
EfuygZhh9E1juUkg2tzBVCWQSJARrYo9XsnKKCy0aLjDlJbimUoN6bJlgDL3pzHJDwW9gNIXjyHV
uW9Y1YMNzl7C9fx57+vlZBx7EnTaBxLN86JKg1+BXXMBjzsO/rFYfL9gt7YdTo83Kf0Km4S1Wtkw
7UNR3YNRPmBb2xXnQATo/PnIWWLLGLaEceaPM6NFknOcW0KX+Tc2POSBsBss6q/imyquX6m3SCOz
PgkwZB9HfuDjKsW/UmB4ZFReEXor3SyQhugZfeD5DH9umc0beveOZlCTi3QaYbWD/IeEPdnOkxrg
gei63pyA05Gu1xUhgv6EihHuvCEqBwKQVR60jjqHp0/sTwxKUwnTQ3i946Jhy8kyegA7mGprkiJo
nfO017BXUcF313VCQFZIxA9kIyW5V/nqcFylFdTy9f2EBO+ZOusEbHUts1mY3fjTLgxvUXZgnhAH
DLeUrMHnErJsT1PzmMjrEZ4aIChb0Si0maPOeZcCxb/SE/pW5ZFDWdpeo2yRkCLmEe/7kDE3/8YT
k0IkvKMpDmZJ+AcV/I6+eNefv3I21V9x5CF4okbrfiCEfxlYrlcDOGLYVoGHOFWaueFgDqdwq+25
e276G8NfHWaoeSuZ9rP801LfR7HuXOtSQeuydyMh4ktcjq6JHuLtykUjChLToo1/xTT2DWVQhIg4
PMZSd7lMt+XVfswlQQrkMTjJ/HJX+2mMyKc8Ola/L8nZKUvhWC34ZCNDuBZtdlOC/Lm89eI2SmHy
KidPfzsECpsaBkJVcGD91YcvrPZ9BZ9C2uPfSFPjmMyyy0aPw/eUply8FoNkWH29UXEPFUkBpIny
9Og7mXeBhpuZ9z/vkz5fPgHWYXYmo5hzIO/m+vZH4YS6QHIqLw8ZqxmFBLUijg8hUGR8+sOTCcRv
huDVc/gJ3CBR7+jftmYKl3Q3o9+SQY66jDxZv6F6PmjP00Ad7byNNiGSPDgKHzabtC/u+z7ICWD2
+vv27MkzsLoiDqPosCckY0cYKrpgC9ic0YmJvpE64CtKF2phyjnXWfT9rRhmUyrJSlhI919GzbuH
bgEBXCXp8zeZAln4P6kC0divSX0MM1Azna1GEdDKoz/P+aDatXhICCj2LnOj1xM1blAGhkdAKvj3
RPnpvF4XVmVRfhek6xeknV/Inr1x4P36XuOWXUwuUfagYr+xYFscCToZG6gVxi7wvjy8i3LhwD0s
b+9SaKEqA5Xz5tljCvDiNaxl6LfgYzd4c+pl1301KpKrjQ/0uQeXDNLQu+rAFWKsJ/YgO2VD1d0h
g3QEx0P5h0PVTx0UM//voOwWPyWg3jX1150T6RhOoy4H9Efn//YtOzZNWEfOX76epiQDhVsrn2K2
N6jQP5ufqWJCGPf0VxEmioVjKWDTQzud+YHm8hAsF+tKbM7dQ7uyhny0QkEbX/vSCkDTxBvN1h5r
xgIRc+KTIDTEDvM6U4ahMusyj2r4G5VYsdc6UR/WWjCVduXq3nC5oncd+DULcTS06R95ccp4f/lH
snr+LBm01qhNdMEFV9J/DHxbpADY9N3VqWFffhLkKkkfJeeHjORW8AMJEF0H77sPSI/GEi0oZ41N
6FZNe7s2Svv9ZliQow/LDjrmxVhuZoWF77PRMBgJNoEsqT+wlVR8Y7My58ZczfNm7WxoXn4BUw53
+9gw1x2n/mTrrxn/sugUlOMVzdrjKJJLiaZ2+zWGkpnw2CCVzM5LiREpU62/dTOETuzhKptXgu7m
TkrXzNzalQnMC9XTxvKpB4nEFJ2lZR/XC8RHLkID04nHbtQQPvkf6UFK/Y77r5zN2T68VlJ7fh+d
OpNwrE9krWtpw6DmPWRmAKN3s5Uf0tg/31e/UTX5wckcCEBzQVex0bbN1oVr26q/D0azXvajl6nf
wlz3dqYAx4whjlt/BWwhgoWVb5vG7mISBdl5h4MECD50qFZyJJCJBnr9ufH/rMr7f/IF3hHSnden
vrtHQdn036TqYhllwe1CfQhluuSq3Gpwz8zhZ+JP2vIkgAJViAMik4YYn8/5cs5HqukpWZa9sSDE
7h4Uw8MEcxOtg9WW+ZKIkF7kIrvlhUYhSVqLRfMi+aVuBrRTFCVCmBC+Z1eaeiWwtyEDlL0e5gqC
E+uOQBXbyRNwuQ0QjciIE0bm2UTfc4FyTKwy9M7eCr3eR//LqrAQYa+Rqi8MSvoXstPMf0keiQsg
xQgQGqr5yupS7ZKVldbIBg9gkb8vxoERJSq1Xu708TQwIQMgK5CGk64kPL8hX2oerVefJ59cgMsq
g6FC065l+3ybE+aZJXcOfRoyz1VMFE0cn3S7cD/ijMMBKaKJpvKhYn4UDQdAQZi7TJwYG1vy6k48
gFU3YN8mOsm4WyLMjwFvbnUBqe151fNx+p4QT1uKYst44+mSofnFJtldBaatyLvcSnMVYH0sLmGu
0Veef7GpOLvwFOttgqYfM1nSluhFo5vE/QfLkwnp0OXnfkW45p6UmjIpKchE/M7fSYPH58IF0kc5
3dN7Zq96r/NN92m9zr8pdJGVK0HSe6YVtOdZ99F5FOts4JIeOVLryTlEWwJa+e6QrL+WoyzaQJwl
JpLgG6qftgNzbofgx0bg3TKqlLp+azRTARN98l7TgrIF2OCSoxdvfkSSp11EX9Xl4hgdlljF7ngb
einr8OPmPiauPR168R+vLglvhj5Z2istJ9UaURVz/M0mi8HnkPXTa1H1Z0APULHv/gQ/BZ2A4XFf
YozRBGKMwuhWOEseSXbkIb1PcHJWJ+/IW7S2uf+GV3eOyUUj8MKObbSXSXjBbZOFJzsEnFEUBiDi
KuYYAYtmNFvHJDqvjnNNdEWpZoTxRCAikL8l9GSOXxgC2imITcDPV+E+s5trduUcC+TAKmiQhjkm
hGq1QOzP82rOtZNwBlXzMQfCtLDe3QCvTQ1B8oD+JQGVF3a0lyiCY+jf5E9ci+KQxMRLCieVJ64j
7AUOnDdoN8ODFRdM80ERQwm2+YVsM+mMp1vdmm2JSHws+Ypq4WTg7xiXTXMxypa7lvhqob900tyM
apuIdIN0jtDRkLHA7H7TrkYQQjhCtWHJ9/J88xrJ/ST+ITrgdHyJAMgtJdmYSImvrv3phZRIS/B+
oS6B+2RpKQ5CJltcM5Tzuy1YdzRGGQX1iwCTV3D5H02UnDH7FBakXsJ2WHD4qzsc3y+nMj6ZpfpT
CEtRYOqowsGe+wV3dVQBBmngi5NMvWf6Wg06ay8WqBWd3tB7ZGtO/jdYAgLkljhYf0e48iOb/8Hv
LPBxDbPztHuJgy9Y2+mJh1nZvmEoU2tEUQd0CnGoXpjVxDTqH4nqA341dhFuuUP5XzcPdbzoLqzL
2b7WkE5JewpPbMTXdz+HOP5ciAKNVtYq58WegVDoRgHDqC5oSghX+/9brq4V2MSNKey9Ase2RHS5
sNsBYW0yUbfQ4NzkTyVTlvx6qYjSk/zRq0mVP+cIgJw4IJkwkkRyDRbNrlkl0/4wvxxdEdOPFAc8
XifsHNBNrPNoYWrYa0SCripn7H0zn7E5E17AiD7Drof+rNcMwIY6ZtavW+Hrs1rW94nY35ZLGr1N
9/MjbFd8p4wigekF0GWtA1u/sCyFNVOvjqbLLQS8SrmhgKNPXgE2GAxsGVqw9TF3cEhxWBffWuZV
NeWzYHxxDd3G21ERmme0oKtcWzGNlqQZWxsL4kb7DenVePkGKfFBSmBkC9I6mlITyGdbLRVk30Tb
zG/77llzTuW0pDMpeuCIsHsf5t6CZt47uGu68C2OKHNlDJCHKurDGD6ODEbsQC9lwiQ140djQMFF
XNhTJ4Mi+3yqB4WuCD8KDDGjOdWdeHpnDqjy0DJcbkjDqnqR6ckIUqV8ldPWLZYUCK2L69aOymaw
RaDyz+gndIHp5XRjIyaKqcHbSnXDnsh2N4sH3mQFJDEGUcAWLePaV4Lg7B7NZW2uW8k24gsJt9CL
6aydkSNKxG0YsHm+LXZ+kjvzwC4ocLQcz7nl7rXeUiuicDC8M0LftDFEH1ReARM1iCvhOTQkXGGz
oiGLWgsQT5n9sYLNcj+RZRBSxp+pPQK3TalhGmRpkaFEtuMD5T/ozdBInNasKzc8fCbAA7nC9e6L
kYDPD2YQRde/UyU02SjJhGfFNGriWYXpA2XoSSeTDSGcXwnqxL+tn2meG1Bx5soIUvJFn+hL7RbM
pfqNlh7omHZpPLQgCRYGNMby0MLyudbCnqDjoKyhMK4hQhdEvR0BivEl/O50zKNxzyxIqT64fS9M
lmOuObqZ8YplPkFX/B3sVCEzDcOHTWNzoVHzHHZoacVujbFPTN+CsPWi37+9mi5M+Sn2YIkA4MnM
AxxvfKFgthhQgRQQE9v5dcz3YgZNJxWZXEiV3/9zNV+subP3nGygeq/VU5vsQT3mP6dKixg4IP/l
jcPWqpJ7TVTWsMo4dgLjMRHzyswGPXYE4gr4E+30Dblz7priuDy/c7wE+2xX9PVg2fEpsGHqkOg3
NJAQVU/NdP1ROOPFOfFi2zZwy9iutaZ2B/3VTyItMpbEZZPf0maiHBJdN+el0qc4Q+vJMvltOswX
YvE14vNLkOOePGYVqPRwQlixGNXSR4z0MWN1mKNaoa/Oq+6YjLAbOs0lh8Zql5JnFMBsZXvFTT7e
BAKrKS1Hi6EGSv2Ast44Y9Q6lr+trQzzxt81kzg0DgJUYS1ClDb2eHJcD/46jF3j0TXbEa6W6MjS
22p6Uyd92i+4NL7Wkp/XBNLHXTVzZdUUCMn+bedtP/a74pyueQLYMBB/jE9yAVH/PAYK4jAhxTmO
LKMaJbSZk/O3cdpZb4yyz3LvExlFxeaJ1rEiKtIWJvF38Mvs+wPrOy+2agqqRCh/wVSWn1FsikVR
RWAmroxN6fwETNxKp6pqAUwf7NVHptsS031f09LVHZIT96s0QBIb4DfQNOHzeVoFDjpS6RMw4Vcm
YL2AhKeH6vPduK3rUavuOB9OXSx9vkQsLyOQCW3dwqanuweN8DoYek/7CvpJGFmMGaZCBLlqG/Hk
pcN7daham6ogYfTzOYQJTCEGqnSV50o42sYGKhlFOUBT9/9EvGZFBrJ5XeGs6wrN7naIcr3+OvXL
EcK94hFfqhKZHQwwnc1tlZePt3L9QIDma8CBF/I+hK2dXn+N3KYgKXG9nSk9qeMo3AEpMIIfoL/j
mWMbk9eRHBBlEdM4VD99r8N8oN4CJrENvFc4SesJeXer9oif+ePBXx58dpQKpm9k1l9kzR7/WCbM
8F8HHaMhv7cH9koeIIoJ2SSeFmLnQGCKVktDlkuvfhdtyZT6Rbye5istjjg+Jhzlm06Tc3Jzep8U
fR5BInZu+ozeOsDbPOrcZkdgYXW1CedzmeilzSVc6isf1MErjFmjqYMJfMtQAD/Pn43J8BoGQ+YJ
uJ9bD3MxzsrNaYbXz4TaWN5B5UGNxvYAeJrLgZooS4vcZ0DnDEgbmnk+mmNKlm2sBWbZFv9kK3mH
KZfyrb2+SAWS+K4dCrdEavPu0Oe/NaEXb4kX/SbWgSEcsXFJsNLkeVEI1yipzppJTZcszXRIGYL0
iNvnXhJvXw8VmXhTVy8Y5HI4Bz7EEwMeGAGgF1KAUNV0Qw4qss/cGIf6ipMRHfaZgqde1AvFUkmk
SKbgkfWofguagjehX1KI5nDu1Qxkr+NidSpKEam5AWwzoamgM8+pzxtLpTTvXspfYmohIZu43+c+
gmqh9l/fMyLq4DLKtr/tsKrTR0zZlH5Ku7DffbHa3w0ZLBB86lPJYHTjIRaPveCxu2/muqzuxhGt
dRwATY7abJyR6wWKYAD9LughMlyo0+Nx9hQ5JLpF3r+l8sP2tuKyVf+/WJ8gVQaPl164ZaHNjeKd
MCK+LXjavrqzjTuAo+PWJuoGFWGN8t2g0V20n3GUkSG3uNVAssMsAoxdtstRr5lF2SIEZUF7hWid
jI4L3Ah0lHTqu/0r8NZ7/S8UpgzsJansdhMaHX84bWX8X5z/mAz/OyHZF5UIXkkegvkz5/tl8cU0
GLAP4ZV9V1r9zPMco9iDeS6AMl7a5HSY1GvFqWUtQLuAhxpzw0YqE7F7n/ibRpBlsPgtgkaA7Bnm
+YSHJM/hV+KU+BKvQhbTQh8bIcKZIiH24KSbmwkNvPRhqiTumjW+HnMOJGS+xt45VOk+Vx5TNis8
8Whfg3bt1apciTOsrq0FzguHLcQGGIdLeWmdENKUKr0vEPB5EDk0qd5Akih5iK4fg+P7ZGOC2eN1
BGx9XIZazhXJM1JnWYVpUGcVoUvEejA9PK/PHO2pzS6QfeVKX/nAkpZAYzMLul0/geMxZl4DhXPg
300Y8LIEVPc0TcGb1DV4YwWzya1afNnkP+ReXvwhqR97TP+2OObx183Iae9HwreNJA9ACb2zjT1s
ef4n72OUAszmtZGa/e54tbm/QJXZDPT/wuXhfHJoZoPBYJPna7oOs7Xe1VuMDV/EzPtrbG/P0lvb
Pbf1lSeEWj6ZfwehPiviPUZSlm8pkHCTbyNf/xgZj9jj0HT1VTIy5jG72EAR4IiHtvAM0run9+TS
LZkTcEzuXskXQHqHSDSvAfFYOvYG2ad+WHUSrA82KTYLCTFsa2oTZ9A16cF2Jg6cGK+l26qfTcoK
n7ed/oAZB5JUz9VBrRhskNQc9io7nFa5r8m39YQJHeKXHmfSrZYjnESF3oF3gmkwDe8ohSxm9Gyp
iwjOLy83HWYZ+oq/XApflKJjCLWFGpke16zMG3NpnY5qnGdTnaNhmwl0QqxcbkRNvsSn9tPFvg/N
NVtJZmGyrL75ylMifz7mTB3ZgDwLSujBAAGgqAXCmO5VwBXlsE2ScYdt9kWrAGHg0h4m4IuHAXoA
jDMdBR/4l1cm1y9MyI3vSZEKvqUPS26M1fzDDHD9Rmp84IoiLTwAdYTixR/84MOXFpQntru8uNBy
v1a8PA7cFxXD4IXajMSLIxrxZifMLQqfbTMDQZ8gEDrVH7G56ZbE1TFdsVesqdA9sW1hXpTO70qs
jCFHv35pPwqW/gYIJo6Vj2Ktic0M5J4Uh+b7Gw58aWo5tJKsJ5ScMc3cn1tO/l3+eFP5GESsaUyq
DiSF2pdWghghHnXOKTNoucsU9m5lrBNTUWidDAfYb0STI8ujClhFC0TzaD0dCnJnF4ekhZQ8dL5I
wGzqmxNj/q3i/L+8TOVctrMkR3Krjri4vR1ZTu5jBVc4TgFeZzKatG3iGNXu9jtoPyt2j1DDdAJH
XLl9HwNOHj3HIPqYVQURBGgQagICXsp6mpHkFbxSL9iSt3FS5EfI+Es7z0h7Gdx/Ju3oM+HPzKpx
lrbvtkH8LBqpupeCP8gD//Yg5D3iKXlxxe08IbTimN5pfhLTmlv+ARYFUpseGbJNgFx1OolABVII
I5NjQQyNi36WZFAMLzjbQ9Q2YXak2YSzZ/1zSlRPLnUHBmgKHe54SyQP3IlQL6tBX5qj87uYjzii
CqI+J3uPO7o4jQY7zJJ2ATVfybZu7S24mHKhOj1GgW0iH6uRmJj8OOGLteGhpKcjpFcHLuJg8Nch
FUsYmmYLMKMck68LaFh7ImYYAn517BdrhAWp1Xo3uswY7NU9ej2VkFU+TyxXNAJPLk76wkai7hgZ
vpKByywNVKoFtzPWIi0qed2wwf5TzOVQTvvem1XznD3IBNv5nf3Lu6UbJYhv4Y47x+9PsSRFKqMS
ofE8BMJVJXFzMZbtxcQ0/1SVKChonjFCWGn4WDMTmX2h2fMbIZ5GNvscHe8GAtMaB1t9/7NxyXfq
dZ1osUv4yZSGypHv4VPO0KUiXlO0pBITMFkQ30hlEGXq/Ge52KaluqUIsiB9OJB2x6b7NYZRn51z
OBSFruEzFLJy3476k6en5PQuTOJhdQYcBDwBbUajzPJzNHkicr/qOVZqji96lLBGTuDN7ftovgxP
iCzBr18+6VpnKu7+hQ+iuTs6UbheKaxZnx/QkxvMBINCAaN0NdMo4PCGhlLf1jzIA1yjUyPIQRuH
FLD4BxNZgbjZnoYjn9TTrSPXiyG4mFmhOevsySR/xqKd7YbvT5tivyynmxRU/mJOaSMXKIc91Z/5
EkllHAamxvLrr7gt1Ti/jlAiLE2sVaxxXiDrXxP+zAEiy1PrrIDQaMLaCCNJ5IQ2H8PkhqcAbb7Z
+s5AmoScqtvK2Yjh6G2vhpq/TjjCqGEXL74DVnY/00nASpXqlJBEPZ2TgTSR0zQi24IwJAaRCZ+x
O8eXwlHMpT4KJebdSGaFJZM17lzc26js9d94Kn6OwEWb8s4lBEA2jcTj258iAEJy1AP6XA5VlPJ0
pbWldfero+4/f24+F0kUcmSyWaKsIAVlBSPqA2ezdanbyg0sAch/HuAPebg3NrtnbwP3om409elA
4xUXgUuk3xeA3MXeCzX6Dqow72Oj7XnUwsn+shLyNIBZwfnjx/iZ/w7NswwpU/iWwCCVS7t78afD
MryYm4CQaM7HMEMaofOu+DvT2Ix0yfgIz27GsGEkGUblzmIc9ZbXCDV1KMV/IQspPHz7DkFdtzbw
XbUG7DjJtpocyFPv4GsXsBTQG0lUFe4NecPPk1ET3QXfMUxGrnngoRKVLJTa0J1y+scJVbD5bkSZ
/cdY+875VGGVT7vFiKDrJcoPlWsjKIfczCKq/lWI9LuzVE/GPAHDuAkZEjgeoOqV36NdDOlnIU15
YOrj61xGQjh5BIS6gXsJ/bt4LZFum3ldd28uJUjuFtg27rXythTQv8hNE4qeqYsBC/nRCiuzMai7
UhFX+wOCOZh0JBhL/MAdgbfnkkoOeul2XMWO7NuNFppzDR2tzdJ1CG91/JuK5wCm05J3viVs9+wl
abxyddzs3Tjh2Fo6VNC4DZj0lKBhR1x4vs9jcMUL4nl04Yg5LouDuNtHPJpiZZDx9++vU1U9V4xr
kwzkYfiUgIJOwqZDzjG6aBWd19ckdZ16QfqgE0utjgtn+e9H5pkgIaXb96ifMzuJfHDSBp/2dqt0
YPDgdXMKwnQdTR0Va5MUGEW2MTN1/DJXh6cUUVuCiQP4WVnmgWzQNrRTKJOtx8nMM2O4TqJOW5k0
mh4AhB7CV5tijzsBBb+W1vJXWPFtGbdPWKWOKFdX5MaOGG91rccLuiiAZ6Jjy+Mt+y/rljBqxKvb
+86ZQ7ETTlaWLgEjvVS5Faq99a+P0X24gLfD9xQZFO6dUXwvqlugaPfkXitAe0WsPNrR/qS6PE7q
BWYikFGtXCsT4EDLUv2rSUxVNR4DlBZ2Xs5eY5vANnNsjFj2Jm8W6VtYR8/QAsIGjumPuXSqyZSU
iPABa8Er9/6DvCu/VfSy8B2PfIkt1nrOJCyCbi2Zl0X13nn/O1YpHfFkEmDu8Of//hYg+DVQiN2F
JA2IBEWAAvBNf5w5Uz6QpPL5VohKzvFGVxYLMU2dQFi4a1w9Nt6N9/KmfOWsiZBDFO+8/ZHVcjv7
uk+Sbyp6vS54alK2WKeMyQ1lzu7LJht3hkPUNbCL0hC/snXbKskU+cZiH4EYiF3He6Ko1uG6MBKH
yS4c9wdNcCbcIvLoE9HkfvHXHDTjQFzaIw5IDxrsG+pAUamD6Lzrk7+49lh4C1WG9fEAqh3sggbD
9uon8WbRFl96wTocZ6Bcmfg18u1ELLm/oSBBgFkFqWQaE+tB/oUB3konl1ZG9GaE6iuNnYDflWun
ubYLPHIRrrG6SCGYZId1AhjybBbqRSiRMKadUzRsGlGaauNq3XOKWqJHJbjkf6z4yBYUv2QZy66A
NZsuNLjYa+N+KUaqJHsGC1aDoy77RRltYKpJos4IYwZLStozOC+55+ounx2fglBDJgAkulikkjz5
7QTslOin/wv6R5k0GYkYr7K80Aic5oEHwnTV4exYjY7Vk+XNlrUuFn6VWQjMms/HzysE3iTlvJ0+
eXpuQfeoThQXslZapDT9GPfedT0AfId80hc8xm8WY3fDcanPcXCMWijQ/UoPv16lZx3nVVQ+q4sf
JpLwzpHkg6AGQwcDzFfyQTJaLYmvwUrMmBHCB8+iBIilG52k8spDf4f69e3x6F2b2q0gbs5YMpxu
FIHhZYy4l2NwIGLAxgBfkVNAJw8TRb5ecHsZEksbQgHn+PnSl8ZkzgJS1Y5lX4cFcYW2zpInr9OA
1mSCMjFOsYzoMDQkn6u1wMUiJFpw63Q+w6VMsLE4+ko8zz2oz4pnEaKYAVgmRY6ESL0a2FE4VP5o
oHNZLFoxqZH4afpkKko6Qe6AXMgu5jBbktzGh/NTfvHN/jK4o5moePiPHVHKPUerOj7H+nWUuOlN
MUQyHJsPU71cWsO0/ru1VCgDTtw7J9HuUToMh+D0/W8MSsDXeOD6k3pU5Wl+/bTT1hTrSrx2+kB6
BiBXsJM++2OqwSWAyjralpz0dfThY5YGmq2h7rSPpA/yD+Rb6qaMFaU+HX5wr+5fNrqYJfD+ESXT
YwnLQpQlI3mSsZzBswlBfque9Jgib0fUxhT5PpdToOTQOJRBfLxDUOyFW3PcNwpm4XNKQWyUvjnd
IEgS7QN2giuV0hadZL6IaRxdOsswyhKjHhrkZjE3WeclUSWMclJO7CnYxPOQF2pK9PWrOv5kuWFu
gCv8TekbntoO4lrsg+VFQ8hCxmLFyQ6rnipOsrRIbT0egPohZTblRJBftCDJzbT888rtyXyjjAlF
Y2HIpq8qzkopC0+3VabqE9pQ59Wu4PF4wQBOtt9SdcGVYr6CGrilxqIueO4w1cL8xGDeA2AZhOtA
kRWat3b3s7pYhBB3sRIaH4TyVd4Trro5Yae657xlZDd2ZXup6usOPHn4CXueUJIUPYX5ASqMrKIn
/C+58zZNod8dN1ucmmPHH7pAaqH/sGB6+OHTVZ2/i5KUr2egUTog7P2ruA9sz1liCtbdxNYodE8k
JY07ebDm2UzGUZOLRi0+TMPrkmk7iVcb2lNzV6wK3f63O3quCmfvDST0VbZyKT7TRsmOamoJb4QX
durkqt68MII3AG53KC+B14lbOzQn2NG0Uc6JoGP14XNHRFJPwvkBqSUt0Gb5wSpISRz5gFdMpQwF
h4KGRDmczcEZRrHZTlHJj+3mHjLcPLq1O1BWRmG/usahVZokTcMb2k3WRZcXVnZ8mC4rUg6oST6S
ZWdkaPmMp0amkQQBeq6ZBsb9ivZJIEF67sDZx3a8rBC9dz9xhB1Yg6vRK4Nt9UABGREEeseWIjcf
01aNBZ9Vw+HVP1FXEo0gLK3dtRtYGGu1Q8zTRZ0kzkafAVCIYoPe45RoIEZJuAfp32rIjMyWx8Lx
9aQzgdp16H3z8p7WXvrI5eKJVoWNEPQrOfoRjRAq4yi67gHiDboSwtvrsnUFtzTazrgbVZwnvsHk
jNHHvxCnz9vC02CdWJgmRnlr8wKH8ImKoaYoROdwePUXVixE7Haw1Mt6iE/ZEF2G8oTYbD8kaf0c
C0vwKp3VbdC/L7WvoIQGtANyH1iJDIEIN9yyKaIl+wH5wFCUDvAdUVBcROQWBCssXK/ieb8XCuU/
BHmBGeYwwnC4z0uSPHvn+U4sOKt+re1epj4n8JgKmj7y0Rl2nf8bZvpZ+hn1WFL6soAGEaDMDsH0
asmzPncEPDNWvsKbKrr93X/XqZYDJoHE9tvoC2XRaN34nVj0i97xdxDg4Sfwm3JCH7I/0fbmJKPT
dClhvtBe+xo7YxL+gKfW96QJow2Exf5LSlA+AVALS9N/jlc+XALVwPR4wUrWs6XkQKKaF16q/4uo
pfsgdIWW8sr+rxB9aG/cKTn8uNug7MSncehWtNJhhcA6dkvnbRSbNjUNrD2iyIf7lDRWbGoYsaG4
uqLJ7e9X/WXLF9sy5Wxi/OlJt9EWcrUh1iBg3ykc/3vO/iBKLvTMvrDcW6lmbi4gVlDoW8uASGHo
J3zdiXOxor2RdzlDsxRps+qDN4lZAB2fmUkvsktqxIvjTmAnmI6OTikkr0/+CSzZqCx+ZU3Vx0JI
5MmPdyLExew6ixMSJOCD3Dd5AjY3Fa2lgtAouwM+4VsWWJkVTRQX67NfGUIECQA/3+XgwGi2GYOz
M/qTIWiFocSwTohKgmylriESA4qMvhFJcZGqRW2Ej1JYkq2es2l3QZX4p8SGJbMG+k4T6o1PnH7b
mlnmREmJdoA4votfSIuaXc7o394h1j9UB1MAiOq9ZJwiyuU1SF0M1GsxbVg0IzoDFhwnM3qVeQVP
Govcq97z2HJCe7gV7zj8wUGrEfg2+I6HmVeyProvaXCM73AxWG6tfpedo5/Q4mZzSAUlLbqVrTo5
399FNXMBjhiByRBKS1tnE9SYtuS3isu5idBoXe5LXO7C2hdNI8XqLrHUwDnwZh4c60S4T88/4CVH
/kgSkRdK5dwITpUhTBpdCLQkxhvBzTeXHPwDRmdNZH5AyyDi7dobUltvapgSaXHDsjsb38H85GbE
lyHDOIfNUG9uceLtVFpM7CTtRPCYCU8L4/h/5taKmbuGBPjWjtnZYwB2MvZUHlA8C16IVLogBzIW
kHvdnypJUjo2MOZHZaTgsXnF3dfv1Ouq+gGVc8epVGM2ZyBMX/p7Kf9zDLgl14dhqMYIpc1elcBz
gNMEGeuViwgz6zCMRLv+Yc3kowmUiQ1aq8nM5tc6IxG2EADBe3ahk0d6/cOj2h/w6fe2GG9G0G14
RmoSabGYqNFGuKoUdTWkjZ/ZcvkFYsZuM06x67qinjntELGcRBZXWjpsBhP+H3K0XANk5q4vrfdl
e8rn1JoP9L2KyE7RCEEmHW4Ng87UH2HTbzz0R0V1tXGNRrU8PXRcuhuYUaxtrnwoeiWqflsL9vfj
MoFlb+VW27kcrcx/DEx4m++6ppKb8HOqv4JPjmmMaQ8fwqY2PzU7L6e+D7A49wzbkgYL9TMRX5Kp
YwidNngdilnuvsurNvMHMgEgIO0dDx+XU3zNHOcVisHNDrG3Cb/RhCv01q6D9LxTdixGElXijwWY
fpQLrKD0YSe7tjVJyNIYlYvzvterJ/9fNzUwncKunwC8Bl7pi8LOfMCKC2H/noMRwK5vS7gBGwSQ
KF1FWZrx7fQE8BAy6dl5BXDEkWXWDCsBoFB9nUtfvwUfIEu9iYVAiWgXcixJVceIMUVqro2UVxCE
xJz2DirkdhA+3aPvp+huRG4YPJTyLXNg2YHu7Wb0adQxRKuCEesr/zDJrrtXlrNTl5ylHlRgdqWU
/nv6BN4LKtkPkIakIq4NHavrtfk2yhOC1pZ0tOX+o4iZFetz9TTCHTqGbkO+004/RCxJEiq1z0lS
TL3FAvTUdwRx5PHdS1rWd/gFs6BCJRKR7tVuJwVJ51lqncx2GDItx11ozwkEo1Pqv9xxJm0AZ67G
acq8GghOw7wp9YNaioXbYcKFeGCo56VnSQRYLQ4ISFOiUEFpsBg6P8CQOpg3NL+Mv/PFtb0a1S6N
UDrnulYPaKvLFVR+NN60tIL5eeN9Ko/xEYhwP6Q3kqCjNlDKOixKngv3+CkyKMvE/NLlclnK8N37
YT+70R7PEPI+7Z7qL8pSvT/Hq6EfaXptR3tVXfkkl0dcLHITbtR9Y8njwHfsu3Krg+Ze6q3rUK1E
pQvo+F/jw2WkJHRjheklZ8yieL4dnQVQ2zEz0Snr0EiFHLfhSslWWJuwdXOClywqX0h/3NhFkyUM
iM2EIoaa7a0DJUcvLLZ/5pjG+j6pDXfAnJRQv4HcxQGxBnxS5+aevjUKmaTja9bMMKbhMi8lcO0t
hxnD+FigtMALWtEap7+VKJ0q3xPZi+VMUSZHWIDqG+/5++JA2KZwMu6YpKV5xDmnaOPFtD/m7izb
bTLKRfUQ/c+rGU9gAuAQ82I+rwAYNM/tWyJCy9xOisrjIzyV9zY6O1WpIkWDgd1M47eun9vs3kcQ
O/1iURlGj35VeNu5kSzc9kB65W6sG8nSr4kCg4tPdsPN1mWgqVhbpLzmI63VYxjSV/buqxw2eM6J
nWiUg9zikJAoL8rovH8uNBjevY12G/mwKQ9uOFkyioGAU2/K6qiYsqKLNwTBVF/qz9/Nd28ETg6b
MOtB1unjnBwKUgXSLJ+hFhksv3wtpYMcW/RR7R1WlASy/V7FZz8HwEIsGiKXBDMc5gheahAhEtPT
VFZyoJqIDn9T9Yjj+mP1bnoRZJKecstQH0yU4iMKqoxxMV8cZsVZrD5o1S/BZaNIKr0fBrbhzNPF
gmoxes/GgFJIVu1FZa+pBVx5qZNXhptZL5K23LPEXh8p0bUDQeg8X5CuOeZY7lyM2d3ahVLOIVd4
Qp+WV3MWgDM/qa30+m2Sk3cIc4vc1ddkm/JkillYwNQgnMMSo89Z/sR+wBWMFDrFvMtJV7TL/4O8
zKwphXWxPEWbWvn63hqUf7F+5rOY4PV7y3gGGEpOvGHS4s/rMXbfTqisqlSO3EFpSf/z5V89wkFL
pv73ispmn845lvGJLEIAsTTFXp4/vKkOgpSmYND3lbUIW9NJNo62IyvxldaPnjArNKWEw8GQJAUk
0ho0GJBca7oal0+LMmsgSQOtC8rh1uiRXaoNOiEH/SaiETO+haoL/CA1xp8blYCxUjf+JlY1ydSF
KSe5HbzGzzLhnk0B3Z16Gk2welMqXeiIu7Pl2PhG9yFCCu9SnqB0WquVNPDHX/vKnSHnAXrQrAgK
IX1WdiYhCgyygKOv7OLv6WvXNFJQeZzVhDNnV32K/sDFcNkQWo9w9NeoLTDucOQUZDcmeRv8LNHd
2Fqm9v8kdhQDLvNvuuXSllTYcjMh7TihfsCqSavIZuZC7Kh/d/n9rSwjQNrey16fyH+yICL6xmbL
kESEvOyJEACLEsNJVs71LWNMFAJdbnKemCkLTE8A2YL63pCPiNWEefEkLqRiYao/N84IXWEInLBY
KSfySrwqdgj8Bbdy5crLsOymHIwwJwrp75pamdXnQbVolSmeFZtUK4JJMRApcc2yo/nNqf1szQDt
pvu9tYYUV6uLFEIt90X+GTFrF9GVXrzoVvYhXD5917FpGVZPxNPzAiX4ro0fNv7bUZ6dHXW5xpXs
2Ta9kGeRQVFyjRLEa7X3YfvoNym9MlmLhKZ/1TOxc2+pL2B2F/Dv0oBCK81n4TXZPmCAETK0JOWg
LjwpN5aPTdRsBpoju/GMvhY2+okDtEExWEYUzBwddal6AhsIkkrRT47waL4arALqDcnFzj+U47B+
V8SDEUGg/IMXi5ieYYkQkj4qSVIDs9z130hw2RjJXfUBCZreOru3IaEexU8CNXJJooNheZm1PnXs
HN0JWq7RNfts1Htz3x6O8kq0yZfQpkpOJigFlJsyZQu8RPabqkY8K4fK0oE8BdumFq8/CTLS7U03
y5R4wOarvs25GyNzen8rC7aZjbQ2B30vZYN7AxdHTw3OFOxRD0JKYGCJi1awcCGq3OBKbKpM5zoL
0P35clm68ugdTXi310bilGVMzJhLeD92WVHNQdKC706HLjVogjDhDjaD3K3XG0bDQ84qvO/nfJ0W
zyuQePKftkkD2oclgwIzuuhRWjzbMFSFIXjKPersIjiF5DSqf0H5lWLV4eOQQwo5oDZxGTwGgNx4
SKmt5kehU4ezG9ZZnkGz5qt9V6/3enZPsAFS3yIxdmOCTiX2HDIJkmjjKA8j+fRj/zrJJJZBMTni
ExKs/fsyvInXGb8hGS/vh2uEuvfs0FV6vderpRuFKXVjD60SPhfSjc6uoFvCsUiQP4mzP8O8NvKl
lFPDdDEvk1k+SMXX92Hv5VFOXqmjeNolCTj7k5GwmyTlkmMWMIodibncRmIzPqlW6KWq7zsGLW+R
tA4mURi47pFnvATnGkwUtkKbKRwXtQhywzx5u4tX30O/9KKbRKpbrOZy8Re+p+e9moFKR1C/OJrV
aT/eQvQl3zWo0VBXfyDShmRTeFUUCkRvBmZSA1JGsmHAvW7DnGXoad0gL95io2I8IP760M8Clm/K
jOiyzrnjBwjiWgxHFm1vWzBXoHEzogJAEfUdVA60KTgSE9HJb9EJytbSHaNIsls1q+3RNaenBQ2q
odTa7YwLOClCuKPmCknePvZrMgGOy7InrWMo2cBHtu73cPTmz4A6GO0Ta8MnqEy2LofufDJqdNZc
OGQaKCDZP/qirFaqv+qChYu9TwoTNIuOkNJtKoKUzwKqJS0Uwd9BnyJMYGqG49Hw9mrQvC6kIfPg
dvsKcQK7SzydTGQ+fQOfRhKMGSZ8CBv1f1m4daxrqA9RqjYKL1K/r4SLZX2yc9HIm/0fXc5QPMmu
d3of0bdq5FFEuHZit1sgSD1M8TKFJXbZGBEk3NeR8YAVXaBbqTtTRld4sDUNeF8E+rx+sxSIzu3E
w8XxGQkuFZ1JuEZUhHl9GRBgF0dX38yQKQRNk++Mj5v6R+n50Z/tMOx/zYg6JyzRVak+XotzTJm6
4Ea29WG46GlKDu9Jdt89OvLfGLOeT1WZ91x/MQJG0ZdpFYTO/HMtWL1/AdQ5CSAef1pqGMrTmlk0
ie83mOje8IIx13qOsNo4ApAySlFJYWLLN5DBDl5iOY/U3BPLQb5Ed6oHFx3T++j+NKDuuyQXDhQC
I6j7uA2/DoljyRwjVa2LsbN0fhVfIsMvElf0M8iG8KF8BtvmhNwJJ5YVgHCY6FCyAKLV0za0zXwd
I2oTZ4He975/rpNjYrwlXVDPjVVGHgeVw8jdpB4iuiyV5RTmkDDWi9tsthgz1F16Lq/1ykhVMY2V
UFqTnxKaFB2RDWDfqY/vd3pVK4mf0Wg2/dhwlx/TRrqiHYt8BTkGHnmNiDkHL6fFmSaQdpLuvxDr
Ijs51k62VH/zNoqGEu0U5xFj+cnbX0r/I1QnTFmnAvcOF0t3yEjLRUpqlTsy3NBkzaL9RLZ+BT/p
/IIkZpcuUZ+dv5LquUo2iFmiCiAVgF/WTQ/xF/ocwrL5F+S8/BnyxW0+3vTJSBSnKHJmOqmmf0Gy
z2syoMrwXsg4CvEKS1aEugk5XmOyCrze8cKwalPHzSnrEauMyi1lNpC97I7yacShNnXKLFW69/eK
h3Xx6225H74mj2bdmdPoizKgpypwcnFgTqwARgjXBA5g6MT1CQg+lmWB48zjScYIKPtDm+J+BPHU
YH7v77p7uBgPHL0Rg9JfcECQcV2O9yv3x70t2mV+nxw+6EoI0V4yRRoEfFjOpm3hlmolDkwdXCn3
Ybjs7F+M7xrLu6sTODKJw86GKsU7eqBYNuvIPkBCYoSw7tdi/QJFVJRRgofON2Bo3R6ta/Wqqt8L
QSa4DeTdThHPHdJ/p2UhS43bilauijJ+8US+rroPPFotauOWC9tPpZovdkIwIWwryWPReeVJHbgL
hDwlgEh7fLKA8uba2zAXSUnqdhct2aoSavseqhc76KoLadzKBSfSWWyhW7Lk4JKpnQ5wtq4hWdqh
p7h6xBez/j+ACXY3vh9pxJU/b27D0wqeRSPmUH/mx+tUXQbOhLwNOBxNGl7ZstXorxjH8Ru1wPe/
psxqP1w5PzxbN9Sf0RBRHqhcNjXbV7mGNSjHktoWuAWAKNVVb6ax8qHunxNjw09CB2c+llNnZxnU
hn9BQ4gPWUF3S2CB7Thc8aXucdjU6Mxb/BQrr9hcco9rmjh/DxOFSl66bISgH4xyPcSqt911g1IV
a5pSOoVxHwvha6PcX6xN68tNqTs2WLtwA11XwXHupsezMuLoMfgmYbezetnufAA4MZB/jW966M92
p5bOAZzAaJzMlN2+wk6rNrF8qjCjlSVb/GGCI5/lqOhgKmVoVFd0p+cEq/7e70ZBjR4glVYFFXLr
CuM1OJ/Nb/mFiN2rPBkRRgNqQ84R0ztZCOCPc1AKmo6xUQ611WN2/M/90uspuhxX7GqpUbtuv5h3
FIaqYvmZDt0gnbD8K8vXEdWs0kfoTgzPh5VQxrh1GR+zbOrkidmblEwDWeeiTKhmYgyO2EzhoFNg
3KejLBzZgTXkXqNw4pcLXBwSqwVA2yBEwu3/91G1Q1xqxTZ72hfmSlVlUXWecBIgbXT+biqbPqCL
AtG94jcBY1ocqFj+LX1wiLOH+IxND/rpl7scl3K08IbWytt2e/dV5OMoDHDRKrBfdqnH23UVXG7w
s14KjGlej5LJEp3bKUAkzT1NNfQQDcNWNqmiIONnV0xwEU9DB+oTJR/lz/r8WCy3Vv4yz5OiseCP
+hbb608hDRtgTUKJGzgHnnnQy1eVT0SIc+uWOai9dw9tGeieVdl7cLLgsl1CvhFD2nll72XdKqU9
OlDY5+oRfEW5VauiLx8kg8deCWqOGMjQrrkzFQwVj64osECPXGeU1ocD4SJdd13lys8/F0BAhZIt
+rpsCjFYRnM6KtvExSkpr25ASTSa/JxlPy2pPFXQVFGTNWDu3+FjsdlGIKhdhr6EKlmbIywKj6nW
XinQ7Oh6/xz8K7DQpparH2llpQjuXLXNrpE8kiGdMtq7/X8qdEgj7BZ6bLdrpR2AYcO35EFiE99O
nHzD4kYgiBChIA3xuVBRjdzxB4f39pQMWHg08Ymmw68mvIa5I5p/ctE0IvnkvXcsjx74DTpKpRCp
aWIt5rL92Igw1zCaJNJwdxMvOyGyocN2AsuUjUehp/p+q0NLL9hJVmyBmXZrYVtBBxj7Oqr3sRvR
y5zhas2pu2nI+HRc5/8VBjlQmiAMLfWHqZ8AH4d5fK/yqj0rCKDhCObssJ9DuvkMnkko6mbJERX8
4bdLtKgzaXCCvnw2eQZ3CKhKqkNhCIPpKvepaH+pEtTsL6gs7zd0uE7odFQpIAmQwtgQ5Qgsp8/c
l8mUpcsT7rhd3mhmsQxZuzpmS/r9T3lM0GUo8Z5ik1FgRqk6gl1N0evOZuD2i1ByCZvYtS8DiGDx
/K9JKUdgeBITq8Ar8DS4pe/qgW+cHQN/2HsLRh/c6gWNzHonwUTkoZslKfa/FLpVcf2XiY8qHJ2h
FEmgQX3irjO0s66Y1LYRQA6rwRai0oR+jtPh6QYNPSCPLYY8gx0vGNqDAqTbtzTU8dPTYM6ycF8w
YsGlxtA42a8IBRnle6nHjNH8BvD5QOrKq8L5Ay69ysKGKx0iIfZR2q2GxAv/3cQ1W4/0dThM9Y+k
F0gN/zGt2XMzBAsAoTWIkLAin418QNFCftvPH7GAjdcMjWt/egFsOmQRL2loIR+706HZ9SslsD/m
U/rj6zF5qQZLsqj5jpH81KxHGzj25ZiE1hQrgq6bti5INse9w/Q4isyT4nANp2OW2e7pVJqeYct3
17E+aQyRD9/GUqpBYk++z+QKywaB3b1qhYY2q8X4gShPKZ6Oqa/kX3MCFgliDdeDzIZjNmn9jqDs
HQbA2s1iecSdjH8B4xj6vTZQ91xsfsXWH3RqDOHdaLl2Uk8oid8Mmzu1FXoa0VTFuDchkXTmJjIt
Wnjz/sOtSbTy62gqmy9ZtyXNIJa6h+rsi2jltP+NKz1Vw4k/W3QE1jh6bKWZZAOR5Q6O0buQ8SRB
KwO2twKpuanLcdSRVTDpBupj+U6yy/Q0sO43DtijYCZ5FQlBr2BW7B6O66TOIXssFO1yQzgKmsb7
oqlsD134l3+r/GtMQyP2oykTJf1T741tVmF5if/4vgaHYJ1UOnD8Ocr/0e4Wq/+0EsZsJrQ+sJKD
bywMofbSZglrGzrl4xgj2S3HkJv41dh7/lJxAdimzhy6VQMQlN8Xo3ED2s8DQmOynj/kw2DCPi2q
Z6eV6pCeEO8akBCRHo1brmGk/xoyP5efMiWaYMHa9w3mR+ptfA39FQwbTkDWH6meM2k1RgVnbCu4
DyUSdsQaLsSDwO/HXcabHAs1QpVvnSuF7LJSYB9LOs1pia1/8mIXRXxm/0bsBQ+Fo0qYFBZYTQCf
1slTlBOS42fSEB9V/S6NfPemlADH5LNeiQ90K2BoEyU03ZK3y2QwwX/3PvPPYNkRmpjplIgDsW+c
SfGLXCHFeTpyhJ5E5a/PUnL02jldPNlJtDYGdgVUhxB3di+Z62doBIQD4e2KhQaEu0bCZO54ZkJX
kHsixMwWdAvaAzsrWbdBjCtYDCB7/4mMWgJSsSUkyBGPOlXW01Bg+/sMlrXvwtTl8zL5lFPV7PLe
QpA909KB9/q94i9mtv6wHVfRabUtt7OnjHhRNR1DOkL3yK+180O2h/EJX1p46+L0SeftmBBS7gpi
Cz/kM3Y0WuASc9Lq5qICD8k6K8WHNvMRJZUXP3NvbGjSFe5x9mAohGuPAkVtyVsIdolq8QWiR/7I
tjNgeleeL7Pjo2QbocxBbqyRgptgnKKi76FGk3igK0jeRwZeVKxr3GuKFjTw7dZwMgptJoIjr51H
715WGbHD5BW+BFqmjaeLaUWktQDmjhOMKu7aY7koSqxDoMlYUeY/wBVFAjnAjCq0xq1s+SlA9AmG
vG0hAjEUD+GZCJu+0JSNbJFLsfCK/P5uHuQJ/5/8CZi/GdbJMq2T8dohefuyIqaMwNyip5M/2DaL
i5eTOeIK+czd2WsjfGt/IyBwSszbh5GWsXoQDMN70ZQFllwUHKvpejgNXoKOnpkHtnYtl7sVS7Qf
PCHNUxS2CzNgGjsmj6GViEr8rp+X85nn8GCQg+UrausFUtYbE2lEL3zRiaFsZ5Caq4f4yJ9cY9FT
ONqQSRGiSzBo6555AcUbSANDnqwUnbwb9yb37/C6dWKG26GrLpULvR0kfbsWUnCLRRRvZoWyGu9T
KOj+6hkPwkIvFI7i+kcE4IkohP6oFYS/So6xQ6Hu+9vr7TidJjjQr6Oh8aabUah+swdPEsqOcaz/
TJon3Cm/xFLvScuOl2QyI9ZKtlFn9Pg1CA1Uk6L7g3h2+3/EXZs7MjwOsXKyXDqGGa27wDXwY3za
Y2dFoKEXe36tKaCcJ00TOV4/urms/vnjZNIMxnAGLHpaSmu9m08aV55CiTv5Yn/Hd0onhtxFYsH5
bPWAAlFUb3dSqFhJe5csmgneK27BB3yXHWKLT6YGtAjthGYZQxWlJBzs/V0cR/Az6RqluK5lHU7K
CQ5BSvIY9Ba3q5KK6df8uvC6luQM9y7Tw19uSspPv6cA8Re1O3XcK8g5NuHTk/UP2j/pmzUq3Jsm
Vr28sBZtyYVX+g/w9mOqc5pBYG3mO6aemF7h9LYMIMZPti2cbic+/ORbfY1gA5Jn4XD1D8qxL5pP
SYMsj1CNsB65f+GBDumOhiQjApxETYT+7P0uAEo9bkerPHUQJqQ1zlv6TY/9bVDfFejXTpI4IRdV
t185492XPvJ4mvt+1zX0hjx7QaNU8u8dsRuQZw9m6M9Y7LPkh13OmUWNm8kWSAGLA6YOZ2RWNfCf
s/r2s6lRGR/UxQYsoVw4PQNBP4tt98td+aPa38g6zC5jrFcX5RX8jYcjU08XoHS/MWQruG/reIzg
CnsKeK3ILuuT7tqbsB8JExZhlL1fej/H6MAZFGlavPrJg4h1zMebsId0iYJqiKReerkjvzrQpnHr
RO5SCoUGprSXpaAVLwOPhvxX/gOpw/ub01ghNEGriOrHRYNa1XYH9Xjb+Vwz2WLJEECC3bufTHwv
jq6d/vlQHeWKwe+joAmG764sKaW4oTNYZPJml6pywM+jfBY6mND7jIFGHKfddbua0p4+r7EVj3p+
+KwgPW3DWEI2Mq5/mYB37QAOlHqKXH3K/VydmpxDuufAOKEc3VMVfhT/o1NEjbRgNeLUqzaXJY7S
SJ/l85RbuxrC5nt5B/u1YdAZtZoyFA+gSPYRY760KDeAO/jfm6Wzc/egKKdpxFGs8WUDzkjb2Nm0
CPQ4cKnLx85ieQ2vDBjgdY+gBQYuaKRKtiXobtsff0wWg2dC44P1JzfL3kHANpV0prlqFDbngiK1
eCPvFwYhNp3h+YcUbftj+Hn/xa+Z46SWlQ/1DwjbH4Bs8z650/V7/Z5NSy449NOtYqgTN2WJoLrh
G4k8AQJQBWNqTd/HWu3nVQIjPDuo06ExNHsy776OsicnuiLlyXJB3HpHQMunu6idXe77vUmJvWvD
0C9e8ywVUDHnAp8tdG/oeoWQV4mSQWHqg38z/H9EKceG7DgYPTcm8UK6X6YzUBP38/Gv4DkK+ke1
o9KCzkzQnPyYKIJJdJubjJRvjKK2xbT3Ib299YsuElWTqGwUR9We1Xi042CsI03Qx3afTpZy918n
0tozElaKQy9x/1TC1/gctfT0cIqdOagnMMHXqr/+mrWv98YoG+sBIGJg/0zTn38vEZimNBhVOUx6
RXqpobwUf1O7LdK8DhjT1hWYsbWS0XLtAyQgGd4sTGdNCKFm4RCiVidkUPP17ynkMiF9dqROJfxv
hajQZ/NNT8Kw4lZ5Xs0W/bR6Vj0QsBX7rAlkjgKec50NJRTRQipwAwUp21hjBvmwjiVK4psM9fZ6
gMhQ+X1G4FMIGLc40Pu5uwDnO0sBX7d2WozkxT9lbpqiKFoDjjoVDIfLyFWyAkgvh+YP989pB+iL
TI/P+YEESXydo1DUEqWe1SLr6G27R8OnpQkuh+Dz9l7EsXDQ/OEwESJMINvoG0rGkyYVDYvCK+Xy
NtJJ+pvII7WUoIu7CCXhRWNfPrkQX9ZNCa/d/Tx6Yca7kFcpD0ykqBe+s7EHb2r4GMdoRhWh20ND
WiwnW9DX4bH67U7cHjA7GsF7vDk45wKXNkWa1YH235NywD9BEzJDJjAVeHxpTktfiB0sVi2CHY8/
+bZCIi8SMirqxcCD27akmrrS5JOYkVpu8qII4/WhepfRtbNPx4wGk+OG3/KX3CCHYHtXb0GS98Ev
WanY3AZbh7AwZ6z7H9WzVQDNkpMMP8KrVxUqFL2vQP3uG5sVpxSSW4876elFPY5xVm4tHFhA0I/6
2hO0oYNw4wve3VFNexR75dCluGIuswMb6O8xeC5fiZAsEOxCUNJRK90/P73KEkjZprfUfNQGbT0t
9ZFbEsxvahxCIW37Rl2K93/CuvTJ06j5FfmiEUdSbnby55tDL5Nxly5vTCQY9aMzBbHFB4YOcdQS
TckVcua33xy+tQcDGrMWTDHbElEwQB2UiPn1SIgaTnCqIkicFReZOOzfDNU5ve1NxCZw+B97cdFd
ZvmXyAdubhOaBXIsUD/tjA2eePElcf2Z0Yk0I8ZD235UeuKDEF7LdcUvhJMMf7iOglOT9HSmKjXq
ieefzyn0F2XVZYzFM2ehmtiA5t6zISyrnCVeXO4TMd74wrS0Tp1dyqLtBSpLMbMG/FTAHfYuIlFy
+9bOWVW+Ltr/RsaSjW96t9wxqpmGBSrPPwkZJMIxTFkYPbbDyyCqZf4MEaHcP64/MGhvMB/OQOr/
bKmfn0OgmzrKXNdaM2lLXePRIjAOv4a2qOAKv0lp4C9AFQS7rvNcZcnFX226E+IME7ijtvfnWZqg
Df9ISNGrWrcJX7KEBfbaQS+hUF3vAg1hl3Xma8PO3y6c7CLwlyMQElNqrEfwRmUOZEDi/jn1QS3L
K5c9yu+TSDWQ9cjmgYj1BeE4/FzJ6nio843MTOTFrmsNcUWButdAk3ny4We8H11MoK0IfWkk8mHa
rAnOVQ25UVwNnzfSmHKqxzNpAnOJEVylX30KyvX+XgjxhrO6MUY6XoYy8HqLcPZuQuvozcyO52Hs
PLgbmfNXAQ3TJgc0dJpHW8qG2WatfbRcOodeXuRX7qUgUSGFFjgX5uzok+eMELGRh1KA86IYQxuq
vixhXeWAQG3kp0KY3uEh/Jd7Ckblw/X7+HENX/RGY7oExI0k5TaL4UXQ2sjE75ARnJxBzrDxQ4rz
Vvrk5pmW1jy3NzmIYYX6znU6JH3O7WJBhJOp51uv4v3s2cc1P2pVLb48LecZ7kff1w76FHDVKG45
K68nOO5Zg8HJ5yEeoQo5SNXX+KaQzgYb0ToNsl4mJQ0L0g8KVnD7FIf5ytykismB4v2C52P6SSt2
rV344T0M05+ZkihzcKmV38BVvaDUoSahgBElM/axQ/aFCkw2Sq4XobDBpzU1bcyKwpNHioThk8b1
pqR/7IW/0ikEsDpb7JJ1NSSFF81l96K6CuX2mZDQSoNmlh0GTW4hx61zJ7sKnwdX02qiTiJSHQ4i
1e8JeaJC9EIgd1uqrM/aiTZNb2sJPv+zDnSzDtMdlhDomogtQL9Jp9Sk6pca8qp6SfZf7CjBYs5O
hmknJrd5IqZF0qXzu26YWBXNyWcDOO9B6VWdi+CGf85e0yJBZboV0s1BGjGQVSl9lYVLHQ068eSA
8Hz7quo6IdoRsSE/nsv8F7S3ACrheGHFg3NQ5MD39oQlMv+Q0RmGYAjNoNPH/JkJ6oHA0+RMg001
Zh1aPj3iwIHYpoMOeycyfRbHmmzeZd9K04hkwgsEp2H2CWaEaOiYugrc62ubOLbdYDW/BYiS61zD
0F3+1nUGRwsxtdyYNd2YcneqmRQnxbmd3dF8Uzb3IO1UUGRBT9IPFwswWha6LaPfefBZ9YpurVZO
+1M76yqe2pbKKZHgAcg5rr9HU/cELLAW8cO8849AuzgpPZubEPhh3hisHVLrM3wj4aEcu8nMAti8
SdwmuXyvvzmKiaqOIeyOvDwV8ULvCZTjcImp0i+Tly+zsDMBi+hgMAhDao5Lh366w+ZCYrwfpJ18
6eZKKF4BOMEM8C8ORxbzkxYXqvOKz+FTSfNsMIBckSq/nFJwg1BYoj7CykhmdicXQZ/keQuz7NHv
5LSScGsU+tkGcgU0du10L2eYryrIosr7dMCVT4xXQI3YfNVKgLGQFbBPGHM0WxEwXtfbXm/+UI4T
iriO5cyv2tupvQDX6I+stgml9p7b0iNo7PTME7qaF4Z34VaYBnxaI4H0/r+pFzVEWYRq/NK58+MH
VGa1mAo0Z5jkojt1rKhKJyI/9CDkjRG8jTz8zIM+9+TRPb7/WpI948eZs/no5ERApnEe86Mlx89L
tcy+yImTxyJgbycYTJ2ryEfu5fwurF55FUPZXCjMCF61aSsPuKvv5V4CzSAw9Mq9eUfsMcC1030x
4CMoUFGbgcYMKo4VBo8GRJZGc0FaDlxIj7EtCib7QEoh0788nssSZ2trtfvnDvd6lWEo9QgFJwkX
iRclwtvxjDk1QdViDyBKwwNFrX3G0VYXJL8iVrphldy3JZUPoXKhXyPVthp9N3Vxy28DxEkWaoS7
3XhJpKF0zjFEm7vGP4N5lZMj4NKhtxKl7PVjKkl7tR6TfcTOPyVe9oYAmV/tw6KZgt2nVbgdG3kn
sGc6BYIqWxKKENqR1Tu2PTjQ5wGefUv/NkvbniJQWsWySkMXaWxoCKd+nMppi8VA/OWtbWkvuXmk
lZlnEXghfLbCV+0O0gbOGSLDEd8bZ7wFYkR/RpgdSk74cmibxcXfRC9t7Bo58D15eanvH3Oq1bfP
6rK8mvtDXL6WYU0RJkFPF9+0TxBhzOUdD3OjglTV91V8mWfSJjnOV0cKgRLRZXUUhFcySIGxCTe7
QnBH3UciXOCzU0V9aD+G2d0zQ7rh+TTktH1kxO/fFdZiU6Dux561gcgGpfghp8xVqSc3L4ZWRbS7
jUGY6IHoMWUVjtiBblAqd597KpRAE/rXr7ychFlODtUwIwhYJISEoIw+3pUUmISvDcVv95rHpO7C
OyL2rBqFB3dKCPM2V2lPhr3cHiI+kG3tdD8tmjmk56oXaKigyc3su319pvNDQteKxAHwXY5vKxdn
VZuUFtyA84dzjXT+/PQGrHtiAUa4Cov6i+7WE/aaZmJEe7dNJPx/BsyWMLmDQcnKgejQhqJAVfgf
5D56V7Jsw4afLXi79uIF86z4kz8fZGSrM/D3+iJ/xDx+7AcjsI9Rbveg11CKlcFXLdGnHXJfsuOY
/0ofuZ1pJSPzgwKw6WfyjsPfI61f4lTvNFOGMjWza/4vnbuQsqFMAS9KHJWUCKoI7KQ6XrJxeGM9
dM2FtdeDIWIOkDIvto1/qRQNU96vSXfLvaplmCnO+tzIm5Mdxr6Y3IogcfH9+VLgCExsEU6UMmzH
CSriQMeNtMJFQ6866AfSA+dUBcLiXYXWHk6PyyeG6PfXFiBk/0cY5f97I9Irv/HltBdmqLKX7N/M
hf1i4ol9jqlNS4ToxeX8BfnI7oXFjJsu/hN2rEkCYmImLFjdig1UvJwk2wNEuDPIY5Obu9taSWjD
S+rERdJaMjpKl6kkQAfOWwLYfbxpAiJsoMakU7AKY6EpTMBcghMOF4ka7gVukNBHdOCFxjRVcRGv
E4OMjI1EfaqTklzXgnN0Uyoa1Eg4uXfDfJwhyaYsftL5viw12FuJSKvrpjjaFcN+45oJDckXIunq
ZaB82OWYKyWlVnbAXD5ka/c5Iit9vGXOu/vFpgfJ+TSsZjqRVsJPK34JkyDGmvESSwmjw74v2Akf
plunju6amvor+Bng5vXqcbs6VBR3RC/ES+kc0qTzb4ZUzFBRxFFh6NV+MmMs+vvc7jcK+xhRxGRm
HwwSL2ZihEJQ1dWZlXhLMKpW0nT6PduBWfBrndCCnfje8Y26kylKd3FzleZ84m+Nm/+GnXx3YU31
Fs2QLGr3WRv0Xgg/N2bYzRV+Dn5kD5j+9Ge8OctrI6kvHHbGImcOdPenD6NueHQKRkuk4dae7exq
kwwwVe4DdSZesZGueFBEI2c3P7np68XgIYznahVjIxcUisCJQyoStsIfsMXWE3KGJTy+uRM+ikoW
rgp4T/w71OXsbJttdXo0ckuiCynYeo5Ko/mu6hqooLNy/4KPXO+Y01T/BtAS1CBAX0Ice0bZvtW2
U2WsgYAgq8gLIHXyPmgCB/ifsYHma29TqopjeeWy1EXubP6vIi+IqNyZgA44cTN7FB/8epGI/bYk
7kYl04bqGFqd+vhKEkIqtn5/D7pVhUOqkt17BNTQeg8UB/nu1XEI+NIzxx0JuFOAunfNPZzBAqii
Emg18Mgqp6i8XfM7a7zSfaPWyeREmU6h28WVdyZ3UClpQmQN3Zz9lSkBlZowQlK7qRQHAM699b8T
cKPBBnBeNRNYxT5zCC2OfnmfawVCYejeiAvre4xwDOo+uZwHTPcueRqaGNc2fdk5xLyfbQB0QYn1
ykSfIce9ks/hyFfVoj/qUhw4w/Qq9FExIz4BIjR9ESh3/zMHCB5fGLI6wRgZfsOF1FYqXYY24I9y
J0SjY/s+zyq5wVgzVzcEfAwenwHVxiFMNnpotLTYAGFey/qZxsK4AZ7UKhvgd78c195ebiIEJHud
4vHawAZNuI0YaRNYMKvB7rHP7dBECANMtabIMNJ7cLeD2Bv2pp/NRr6KhSMM6aPKuGEK4wAGpmYq
V6ySQ8pPsvcgZ+6iARdBwMUKTC0XKZSPnLx9U2Tlcoq3BbM/KzCYSB55QdBopb1yeQcgZ3vC4TFX
SR/DBQ8zHevyQMRnK+4rCRBIWQpvj0oS+8kfVWo72LeKLFm57piOPpFgljKjZlD67Fy01X5JJitX
qbezpSD7RzSjzFgBqKkxSRUhLKKISjmismSgFRr85ZKS5yRokY0AilPvLSTL57oWinPHi9gOM4Ej
QZaxE7zN3yrbEZDRdgJObhJ2UwiVLOrxmAwcBTxdIGgS8CNqqYJiDhY4wwbyw0EYrcKrbHxcwTxu
1nJGPVmQ+5WfY7Qmeqg/P8kvErShAo39l1hjIkaM8RZ5CJ6tC3zchTAbxHR2sB0v8F2SawCj2Vmm
v8iYngCFnxb15aLA7X4bgrWv90DhmeL4pQN0xNGapik1nAJI2SRwFFfH7M0csAF5TIpdm5VhaCw3
GtLtCMTV4phbHvIXicqs+kqmOpKqkYjBXzalE83fSFZuCgJB7h77dmWGmno3ZDQzqYY6fx9nsB1p
PaXs04sEHcgytWV29N9B1WjvKKk/cWgDXp/hPzK6C7+bhbKTRX/B6qli6qVAdlsKgb7tZCEHr8hg
vciywQJIRZI0iohcdW4jePIjZkD8gcbSEfZJj3Ybc9KgRpf5SwjUth9eVK81W+cm6FMvMnruJOI7
qUWaPUkjLikFzcRkSK/YCu6pi/0kJcRh7Re8kYEFZsgbioa6TeR3BQ2sElnhxKW1ynMH35ywgJjf
wyeAvRrHvX6ABV5qGJGDI+6dEMI1TheWOP1b5gNls5l8o24uCcB7Ftch3WgqBVvzzJ1Bjo0DzyiX
yxuCdIfh8Kx9HWk/s+zDoqmXOvFd7Qk8YjrAnzJYPTyPirLHefdHUx2P420HNlGg2XGanaC8HR2o
uCwptQ+8ZoV4Y11yD9wtZE2Q5qhTuX8hfKAwdKfvGpDM0iu7t0oke748jiPiprx8E0fS3xKxK/Uz
MDi0tPC9UAqJUc4u09NwxH/BQxW+zNE+J2n7qVCoAukgsfh/r+iIa2zhfslFPDrKAqmaGm9QCzjL
EuS5ayL3F8DlEvSegEYDfgABBBKY/nssd0FxkD6Q6Wct8VeqQ2/ajN+/jAwSMACU7zO/vfrwQYXe
IjWV8uFVVtPDuT6c7pHf/Rw/jqE/wPdcoOhuYuJq2fK39IZQorw6z3r2fYsFg5eCfsYIyeVt/5NE
HdjcEQtnlAXa4ChkdmtcUK1JkdTGKuVx3nYgDbb1+5YeXupppCbm8BNY5+biEUsMBSvPvf4zjYB7
kLa/DG53Se5ku4w+jiGGKP0NV5X6zFmo/q7kuOnWOpSXgzFI9mcJcqjEzeIia1o71GdMr107We9S
TCsFuWunmWZP7o8pKwUrByfriad66NdSFPBorv5WW3CHe7vGAzvmK5XtPQLDGKKS3Buv6dYAR8wK
F+o9uqtrSF+k2ophv+6cu3SBQsO6h+tAP6kxm9BdvwZNh8OwNrlUl3qJ604r8tRja7Orqx4GDaqm
Ca/xhQgRVME8Z5LoiGFG4RGDtrWioAwHOL1RCojslhgzSK0iPUN6qlzNfqqWwclW9nahWVb7J1Md
nyoGC9FXDM9lOW3loSYTXARMoiFq9q1f4Q7oO1sIXTRFr1kw5TJTowmJHTxnyYqqMhzNh0dJphKf
9Ph2DLsm8sVNr0FbNJgXg2n89BgNaLr8i/fPDqKq2aVvsYd+0lJLCFnxj8kouiDUFrlefq4/3dQZ
yqITkzeydT1Or3hz9muHxH7GzcVjUH6evlVMG/R7I5TJ2qKksnrC6S9MMWXUIOnuu2f7F83SQQXv
8WWIl9xEqMC78uozhoFmF279AY28gKVEjlr1laEyhi3kQC5MnkmOGu7vhHsJks97QS2UkVGk6Y/n
LxQwiNuyjGoiurnxLJzesYyCtbiz2K6YPTDN18YzDBBoSThnvUEZCMr6q8mAduBl3GEycMEu8S1j
/jT2TCnUMalsXdLkWe9/CvoUm4OVrzGFRA/mvJovEt4FDe1T2qaaHYKskkOlzw75TNJEVGsIPvSD
KYsdhtdhlG4uj9f4UCKAy9bOxnpE8PMBqBNkww9VcubEzuW95UhFekmdrWiwufWRUU1qS+/2CEMc
gciaqG0ebJmWf9u7C47STlr6wcTmZyfGatK0Z988yMT2ieqdzPQZZMvHuzff92X1BVY4XV8rMMIC
DXYagcqJqnkGAXAwJdqwtm7LzDj7KV7S/zE8Hq9aU4DyjsIxhis/pozhMZKWJFaG5aVowuhqBKTS
vN56PTLv2QU1cjvdoOdKJcXoAxmIddBI9fIUHE8vMPDSTQWsduEUQcLGOga30zSTlYCpDJhmus8M
yJzMOZc9/kd2g+dygDT6+L5b5indgLwz83KtE1+eodEiskZc9QWq8BI+tTMlKCO5+7DrRrPmxMKg
pTiaWUkN65t3vIB8B2G54Oe3rngsGYaffFKUsrSjHYm+TxSBWU6n1/z78AyCTtsrhf6Rs52yPVYC
ImmrZAdG6TJbi3YLfpy7gx11+vpNOLT16+VeV7KWsUsOBX4S64zaMf7mc9edzsRYiBSubuG2hHm6
gVs21nC9xKp1B+/dns/C96pwdB6sB2Mdxd79gpbC85FFSfEnJw6I5ANrYAq1IXjSHCLJ5MtD1NO4
bacJ3b5loahGB06egR6U9261NZzjVadltXEV7cw0rf0GNGN9cf1HYTGSan5Y0Ra+NG24gPfK6hgF
DVp+3/mtQp1HatMQ4ELgVskl2kd21g498okPLgGF1pZ7YfhLaqGT+3IoxTJjsk8JeUE1fn5qeCl7
RSnwtMcVdBGBspjJlVeg9cqpYjF9NIRCZ1DiGOySR9FAzR7qog9VWAUmqCIDTknNwYBPXXWlQMWg
LoVQKRPlztVIUHX7WrrjYqs1zafhBoLT2EV8JVN6kjk1YX9VbrcrDXFRQOsp9CGGF1AelrE9wAbx
gOhw+Qff1PigzkmnAwxGu6RE0t9T5G0M4X5l5wTgMKpDqNSH+2d/InM2mWyXk1mFH6tX5BRkD3Rp
Ti6HQxvUDuw1XJFRqGZptMM4l/OPm4XKjBYg5gbeyxi95Ch7Ks3L0u71gGZkWhudcimYBZnzVxuM
tX2pNgzY2JeMGeid17NfuMmsH+qQuJK2BFAfZXxm8RzTgn7htFm4nChxKQxFjcH132ZW1o9Ogkby
Ji56ZBUs6j/YizIEROmUiBhlipqwt95vd3GfDrI6eXKnvE+TVFGBd2CRQtVXCTeltOr4qQlVttL2
vyWdjsJEybQol4IqvqSgM2JPj73xfyOXFLmN4C7mJ8/ciaDAn1LakTEqj8O81bPGRH5f9gA/xnCC
Vb/ulYjw1Nj/DfvCGGUEbmWLBDXL5hPdCRhm6p4lrro7FdryURpEOrIaNKSCWn0MQGNgFcLM038t
Khxt7n16U2aEK4zBxQgc5KcsnQWOyk/dN1Ky+tO4z+S0pf9Plq6mUSYrcMdkxeDnLfS0bFhr4JOH
oVwdo4aZ6PtihuoQx67FKQkoR8+LhaKv4EqqrpWlvKymPGie2/ya3DmSA7PCPArIJT9xgLiZwBb9
An0MENnnKUSVdqDeviYExEkc+5uMJrHs7r+O+G2kKwreGyadnQ+HS9hGUeeS32rH72tBP1W+/4sg
h4TX25w9JduddvmzZ0DmJDegpiPt8TAANyVe1m7CxM9VuFsWSpxT/xE1aXoQRpF//rHIXxnCokll
nvLt7lizVRVRVzt0oKTCtbbJB0grmUuKN2tR7C1t4wGRu0xC83280W9MbQw6x8LNciBoqdi3YoIk
PRUUs4WYQsrri7XoD84VqkprD3y6oGLhDe6sMRaOQ7PZiUM1kWmie9U1wuKiHTsW+s7gHzj9EIsu
M17LY9MozFypw2HiOr2LkFYVRhJKwMFdq1xBxQgiy23E40sAW09jIGbPlNas6bssgWDF01sU9nab
OHBnbUd9KcVsre36GRnvMjIDIDZaCIsQ7fIlvmom9T2uTa6svGxJf5xhMQRWgDeYVQh0yMkFYgk2
KosVkCvOEhAyaAjMLHuFbTWO8YFiieeuj5GdMWRDCtH8DQ1kx4QVtoCGCONehA/Ax+9xH/Tv+87Z
Wliu01hYgGaiQKkR22zsLGr7exhEpqPo7ulv4CbiCI0h5lm6QCfZBWNtKQxEFcDBboxwkFOd7218
X5QNVamCSIanxYNwECvNoCHN6sxMlQTss3vkQwtE3NwCKcfOeqiGlRobCiuUPI2yZCjrkzvps+fo
x5xYQtcuSHh3UfHpckSOQg8jNL+/PnlI7iN38TYT+ixlJoX46UokPlQ9aVYMjoM2oO9tFoK5IzGd
kjwcp3OGymwS4G5wbL03B4pv3WzLF6KUf4E0MrR1yGI0/p1sC5FjJtW88xGAvLeGK3nMAjgR2Jpg
5+W+OHb64lBuJVyd0Npy1aJ8VOSkgV3BtbrPrxok8YLS6NHUCO7tSddkW1dBYlokU0fJGxqyJet9
RJdDCZMPl+Hwhx2Sgf7LdXsA52FBGZ0Z5c2DQZeMOTTFvMeVZBR5aTpQzh9YUYr9UNkma1ZFofbE
ezsrlMALnK9xAjgl46pjgOTUQgNcfi94C/zlbGrrz8KzhOE9/MmcXNUvW289C9NDfHRoV6MOvhyn
erO0eBJmY0GGhfU9HSoELvq3N3xA9SHGn48yZMXntH5Sya+CAwljI15M8mAjw3dOPOb2RpofVpxD
2LQMdCjEp/ItB/j4JH4MlX4bC2pTNCYKOgzJDCj5GfzjT60SOBvt++GOteUq7f0ZeyVkI6516leM
aN356FTQ2CvUWCQmuwUC64sBKEHBqv+mBecvjGJBWcbKz7PCyT0INr7FdSnCtA0mTKYpN9isNoZ6
9rc+Ulto2z1uF/vFSe7CF5m+B5dnLghQW8qlL7yNCy1i2ItCZXKrtEwpxfZdzqI0HB7NE1tkj89w
nFJxA/W2aEQu1ev8DL6bEsg4nV8efbtVb66kjXtgDoIKnPlMZROxsJglWbbihoN+KDjEIsRsVDKY
aFAvIfdNi9jKF5CvKNMNgOmJ79AYj95JwGAuaKh+G+ogWWlhsbluVQwAs/Rq4g0XUmR5CSh6jGK3
AbY77vj68hFZd5rK7DXooO91iiMg5YzNLqIffSAXhZtqFwbKMed7i9yP+b209pn3s4ALk7gqOjHc
Z1gen8CEANAT3e7OSDuqfJZkA5na6QMNvW1PPRO4aaVAE4yxxaFBJQSRkXCz66joW/jMh7alXsFk
VeeuE51n91hNXr2EvKyt0Xx8AMh5VBbTMJ6NzMmaMJbX27oLBqsaSoxxB/Aefoj6l7r4fdcFRjAn
Q/J75GlN01Kqsp/Cq0DbRindbZDA3rQQbr4WhXSfszcGcZF0Jei4KI+/YTA7Cihw5l9y0DTjHZ8Z
miHaoY8wJZhXlKugaX/0j/KuPBr+JQgev9irulaPdxTWkxkjAC2yCun2mFTSb1dMLc7+IVJS+87m
i7XN7iuJK1Yz9zPAw+apYIrOqVeDRXFHYqd5ydnkqqukkMyssn/3EXViUI41hsb287XYFSe70wnh
OTPuDu+nkAwwolLMpZVdPF4TNlLVMj5OdHpQfYudkr60mLo03Bu7XVhHKj4WB1WwWWITBAYhZ+MK
yc4NyQsyjNjQrg3Kzjte8znvqEB3UDTB2yz6AB+ql/FB4ZsYZQENVB975VDaQ8SVLAjkFTt7D/t9
7FIVzLBxTrPZPmDQ/JOxNPSwsml7EkE78nOt7+KrB6evYeY08dH0nvEAHk/kt/W2aJCJuZLPAnGS
MAnWAwgEyT5XPX4xtQ+v6ENlAa+YErEv+Yy+V1GTjjatU/9IakYT9FaUYCADrEXGbwNStC/lAQXb
G/b96TEuAAa6Jn8qGLQrpWbcpjjBvKPC5/dgZErma6wJ5qn6mE1xB1U7vfcIxHBUGg6hVaNPGEFE
5zJEC38nIOpIlD7oTC1g8jsGJ6oEyWgjjbLBoIQZFKaiNGLtecWzcFyRiatws2+DNWG9kmf30tdY
4OwnJRxEKR3/5fN4C/BHy3b++6S8U+/9sBVY7U1x+ZZ9KN3ZOuafEH8bKKHK88JVGIKQsjMfSTop
fphJJ+qgj6FVMUBZwBhqtdibOtfen0awvdHPR1At1omsCwxmvE5P9YF7/GLyf32AYRrJ+fmMJM7u
UCn9fezCAlBT56lHDFj1Vkc8iow1RW89giJbwvzy4+uEs35bY3dhH8oRBBW+EOBmEPcVshbsCeRv
MZr+NBpZHngahxfzTNWXP/v5VZgI+myubY/2gHi1bk0zJqd4YTmXBUalWsPKwoMZuyHaoIj0eoAU
HSqdz+fFVopnhFQHzXr8fq1/BNAE+dEmvItj5kxu/tuDLJ4cTBd7mBidI6WXhFvezljlJhAQSSNe
8hzlnfDEf6jBAzBJV6ib+Jmcza2pK0ra7nHgWi/lOvAPxOxViiyWI62XQRdx5Qc6sejjGGhurAhL
6jiB4TAlOEg5IMpLjTVuRlcG0k/ZG5X+/jduQ5w4JY/XFKVNfiOChetPxON9pjlLukM+debO7tMw
UFTVLlyEc/qNP1Q+dd0nwU6BrDwzny1UaXuGNF4pMtCYn5gYAqwa7TLRj+6GXWplzKPOfu9rsjZw
g+Y+9+wnA2n4XSIRLdiVHuMXab2E2ruQGmzmOebmsiTljuGnuysu5tD9vJDyqudcUYwNNwp8gMyq
F5RhGsFx/3d1s6/bTTMu5ueN/ZbSIiEV0L1MxHmdvFvEJTFBt+fUUTaKFpMU2j5WI2E1vauVqSD1
THiDbVIqI41d0GvB/XI0DSLyayOKEkD3r/e3btVNXj4YV1WGul5J/M4SE805lSy8uuU2k2ynn5ZM
kWPy/qOlkmi341WEhp0Hfacv3u8p6WUhnuRF84xU+EjTgRHnZ6jbTjHtFToyhfWpgxNKijxj4C8b
y1Dn4kQh/UvVPHjjn5ufOs82s9//5bCMPw3mRzmbtQBm2moLPKlZ7nSmlYQouc4hXsIcQJoRA8fj
mk/UXW/WYwVbEYdc4pcx/9F0TzbmeyvLutnYpudB+rG21R8YrWaIR7pY1RBsyQFwdnU+VD33VBa0
J3j4dyDWr4eduODcfbwudGuygDI0frufzYorlMHopEG5qtckziHzdVFVHlskw7EntIMVv4L9neRg
q9XV0qNpCmd1hvF5dpZSbGaidTClc37yHJDmNnnqyaH/VuNILd0cZP8twnvX4s7xTZdbOorGNZ8m
+THb3P8ehXcP8OhdMePiBM1SQ6BLlbnb0hOrxIX4rK6xc5yjATLehpiXPdWKcicIOb3RVgjwrcOs
/YIz0Ox3sCTwl6wx/yvavU3NUWtmophb2I+d6FWyDbsxZm3+3snX4aGecxyR+zl3MM1Xm0Oz8i1r
1btxDq1SYToelgc3Xw6zA7YExiA+ONC64Lf1+hy1incLiJ7qmv5KC7n0ZpY15BvZxe9UbrQh4JpA
hKX9zAuSdwSRtkipKjj7c+LbQQOW/s9059bBjA4xezwu6kE3nVt7pq5xK7vUfhsQ0NTYUUWeGsx5
h+1JtTqJd3tbil+8WIr4PdK54MS4Kll8Qy0VksP10qYqpBWnsLX8HDY2xWOFQUrdMOjKcGgH+e/Z
Sm2puDmYWmyqT04L3Y/SezhY7taqXNg5UWT/20LOEg2Yj6cOiAJXbnSLXwrue3900VzR0vKRd2El
cTkXcmNxZ/LzBdNOBlBNZBtppWm3VhFpc6HkGy6FarCdw26yGH5r8ZNNHv6+AmaA8NI3aOZfNVzH
e1gNgr+D/x+/R5V2Z+gCphSBBACBV7rzfgStiK0naZsSUMFJx/bEpnzgJytGgvcauVPY0vwV+NZl
orTHhw+1X3TXYfq6bm2bhTVGb9rBHoQ4VBj6zJhZADbX6Ps8hY6icWT0oRJHwOSA0sjujjC9aTt9
fW5Ra1mbGfpTxSq5jbb9BjB1Y5pqfpWyRBwZLZ9lsgFzfOnG2BYEdgoTO6UPf8TzUtkwpbPUXrgp
levrmmDDR1kF+0fgMvzYZRBFcRcG9cV2rPhmFoGYRzgVa14Z1rK9qGj2vnWrGszVyOnodcp0ZJY+
3nu2/hCQ4UNG7p+GOA/bDLjPpgUG1ZbuAZMol/ly+U7dUXt2Yjkmbgt18SYV0CJAmoiCWBk+UWpM
OvEmIqRMrdvANB0Dn2dHeTWzZfK9D6zJ/RG+u8qfm1WJSB6JDXVz0E47/4+lO1FeZJA2sNYD3kJX
9trhBVCcp3sk2qNwAgO1ifH+CJCUifLjzFY7dsSMHtX0W0HEWoO7gLwKB66TEYtgBMVr5e9AIeXq
zZDQIcOIz8B5cjImDj/Gd2o6LEf485yMMVQd038eJ3Qzn97wSJ0G52QuDizgnvKW+H0WCUY1nApU
ttfOeNdJ0dPwD7V1Ii1Yq6+3bqxCzYXWBR9hdUuTCjSwjAbEOiVDrADR4LWZlgZ8KuVUseQE0kas
SsWDmU9rG6QidqrVhamtDPqJLJAgl8NdOAFDyfO8Hqez35MDoMSNirMyi6kpv7Eo5bHWrMgLAYlQ
PsGJEMIuYGwoKJjxeXuqYQFo4I2Got2N1B+IbiBNNVGhRMXJ7z9i1+RkQOr5XzWU4n4AxBEnwBV4
tQFEZAY28QwIT29OkRR7adYccF2E6C/+8SdAgDJnXE/ivqo0H1/uhxe/cKjvsJUd93LhCmdc/sXo
29TH+3vQdTrQVYB456E1a7cBe7jFcHo4vDDAMYzmeKeskfr/bRwmSgOJq+HwtDiHicIrJoqnk8ne
R5GOR9e665qayEagcDRdfg2Lj8HCE3Ncy9/OxC/yPZRoQNKMTMXcCqCVU9ga5QKUKLZjqrG4t38c
4LpfxxtnRRvvIFN+SVLoPicgXZl2zFC601ZIWiz0kh9N/wJFod7CxdmP9Lg2fvfPk/cYj64ECmql
v4370SuTacWZCo6YoRI4CAsYITH/LnInzwJB6D6oyn7q5LxSmtH3eFzk4QySQNj0Pl7VxnVPuQcU
biGNyLJknfjT13LJiQoOE55oqP8QpuvYkz6S+XlKYeKwxh5Zfp2nWDHerJiAs7Lxbuc+S2YX1BKL
usNBQyYaJeqyRg1SgW3ZRY1dDeZQPNEsPsamHFAf975A9iJS3gJdPrmAmvSa7q4OP9d9frsBJC9J
pmsy5tPXRNQ8LCEQtpaj5Dd4QuHJi06fOfj3p3rSMlFcQU992ZobhHOFkBbUxnTWuFk3qZQmhCs9
atRztmzVywVG+tV1qsBRf5BpGZ99FhQ7as1dgesw8UI1s3GN/AxJM98NLLCoYTdKncpXoS1Q4J+J
BqLhdco+HQRhmnXtxxfA6OHGPQN8PPpSWjF9/YPtbRZ0RJmQJEGe8PqMupk9RUroUUnXR044YvH0
vkd++SVNbVTd5owxbsOwyXl1LeZvqO/FdLDZVPJxJXro98dFd659REG/rm2Uh4fFyz+JeAbldkl0
AEpMhxtAOTT051REnOldGc0oHXDpR8fP6sNMByrdm9RB6pqv0LH2o4xSBTt/l5nGSZaxfNzD08o/
Fdh/x07IvfjhnVxo11N3YXoVUaPlKx1MgFN7a8f7UqJ81xJ2CGNYsuLnnMuVa02lwM6dnd8Lm1TO
aeyXprNaibOHkJcTQBFahTnxwbsjjGGYHJQcqiddY7WtuKMBtXtRFZLDVY06xHBuO4rGb6NjvVob
xosp6XCH5LJ87Sx4mEpT87JNuZZ89tSg/umPJNkqW3KRQsHwfsG3EDmFCuqPvg436kZbsZpBZP8E
zHP3iZ1iQ5cvsPGSENAy+vEejBG9X21pZQeRJNg61SLJtRXKCkrbr16YHuDQLTCB/xfcJllTB3KN
C5MTmTh+kMatEHjcyxBkcQhGFYB1PPRrVmZTZKUun4LRspkh/zPnh1XsnqP5f6Iqi+ltBJTXf1aH
Z94FxDDo5XGFN8O46YhaDhuvpsfqdyAh5tis/t+Lm7FOaLLz67Lit4apqVyyJjFWr4K6Te2Zfn/g
h4la2wtD2FTxSkDM+PAm5Y1BuZIB1HB0hf6DeZGqbXDCksNlyH0xfSbWdJKjh3iZ6g8h1m/Aok8q
aH4PPvBaOgTsdO6zFRpJydAF3fUqbrtxjQdp2GYmAhF/4XOX81yzxPGQ+ogLi7iuzBF+ppAkdL5C
YMYva1hqAbowchhLkASmOZJV7+hSyA0jHpNGESefNlPfWy9nnPjiEEcoYGv78qTkS0L27DMMVul7
rtfDFg04SwZ7GgOcsJJrRNVnf21wJGGxpMDLqCvQtHPmYNVlA//18ST46VJoj2CBP1cRct+9JMe6
UcqwSnfuFQzIRgyhTH3Aqq7HNi1tF7b01neEmGAvR4/eUuRqkkDomIeTjK17hgPsfyhlu7MjCJZo
Kvy/+voBiENwwulRDfV4p+/MSyna25BDWbCf4IjLDXXkEyLXm+yzcTItHVXPnNNr1hevJZQi3ceA
jvMrxAxPE8axT6jhqCVmU138ehZu9q9ns4BOyfMAx8VgpdmwEs/cDnq3eazBWIECoG7o6TOJamhk
7kkn9UhTRifce0YG8OLOBylxLyrCp2hHIXxug+0IPzhaQXgwAWmByaSiFevs+z5XvAgyq3sFRAbA
8VrtTHevmOHuIvFe9o6G7OO8oyYOYbFQLCzQomNheIecQsEeyFAGgdZMMEbojBvVNE1zND1Us/rq
55RBhRq+CV1sXmVk7Y3dYjxc4YcaX8YOaDDZNZZz/UdazgjplmwO09iVsVZWNBkkyFAAQsGkKz/7
95VIIL2lCpeuU31szik+VFW87SIoIGoJrmYiAnBvzsMUZ7APR6WChG3mJCp0qt1h1cLhZ91mBcKL
xuZ+nzJYTb8kR5hKwZS94XcQK3e0/wim1PVDg2Ua47/4JkNyULY48HzVHA0r+YSaZ/wzJwe4iuOg
NMgf9mflaFlKY2hlU7hP93HKmbeDsbIDe1SdYG+gWFwggh7N1UcvUl3sf+q3JKtbeTyyeZSxRFFn
CFWy4vx/2SiT744T4iwiLI8QZpYQC4SmHpHOrg9GQyvAQr3qsrc1wYN8NxX7ua7JOqNgJJIBjAF4
LSnXDiWYFCVyi5xAlMnj4V64LlySfzJR1ZIajc0cA0gx9r3Ud+cft51ZQX6rDOI4ip2NsCWdJ/tK
GsnFCtaXMU1r9jXN/TT3Iphb/l6imWCV44LwHF5UcmxR+Qqqo9uVwrsYuEbVCwag4VZlOUHrnTvI
NwoJE4OD/i6E9Y/HbD/gpjvrJ1CpSxS5bQYx9FO7obByt82xi3c+/MoAvjzgaWixlhJXaiv7z6It
pNeSxb4+YzxeLWKIA1b9SqtaV/HPvxU4RUqFTvnphIxEFLgWG5hKA6u2wBN+wSRXhsBRCci+6bBn
eupKHZ1cfmCbGsDvOA0v2FMB848/N3cf1uUholySWUsU5/pSRWAWtyJvzFFDSj467eBkkz5NjjSq
7MAEyEvBdi44xHM1O0u6nZX/Key10Un2Fke2VE9iZYO8pqH6xr90jpW5EdwyqZtfjFULh2YUUxx6
w4949wwixm7dSi3BAZRscuJ9BCvcKTdBaMP1AQjsE8rrTNc1xRTo6X2e6nH0A+8UCUGNp+DoBzFE
YGv5UwfcYmuprr5BWiw2HjHBOaCFs9v2vxNEcTD3/NYkkEHjby7weHSpD7z04n/abAhxfhn5b0NP
YiMmkNd5E+xAudiUrlIJkKicm2CYOn8nrDznc2YCy+NfAHxvhbJndAibqSXMEuD6Gq9Lbv6qtABd
dtyAcWWJOMexVzZm2KpIrXcPZAk3g2rauCpdUoOLxkvvpgNRE2j7OjyekfP5DtSbuINKleZp0CCa
IZblpV/HJJhndql/nYYac05eRw6kwRvrJhzlf5/lhI213djvQgDOAJQwLpZm5r7H/94hnwrHjg1K
JakgUxaI3MlxWyiMNZTsT8ifUAuHa+JDa9ejn3v6DnBUMBoIMaDVbxiiAVdbx7i2OYVTPRPzHNOe
N9Q/XnGPu6790nXtHGDaClP0sU89QPE4by/W3Akrr+yhoSpUQL6Qs5kuqvQnauyT37/qRVvVCT3k
LeVZDJEg4fGj6eyfI+0Eu473IgwjNobDj7123ob8nbWjjKAhuPL11kxKsaKWqWdMQJPxV+/+dAF1
AwK1/kMjdw/cQkCVHP5zIaTdpYRqFIAy1NKaNmNdhk9eZ/qng/WgPlE/u2kxx0uDWHqBSsVFgVZj
ytbqO4EgUShX5TLfm9ZL8MeTRtJKWvs2cFkme+1XkpCzMZSjUmkGZV5fmSFzGnivvtWYo8C566lo
5oBOCjEnj+iRO5b3RJXaxjr7k/c76QCSpT6DEBqGU5dWjxJq6OixjDz+dFxZJK4tNwWOpuMoBUta
t4OznJWzhP/0CnnERpT7v8NS7byx+3y1wUMCTza9zkvLR9EcT9wEWFoTGQ3NN4qmDAV39p8G67GI
v5BpN3CtnJy391lxcIc7rW00qu5wmn2gC5JRJmG7gWD0vKGv7sqvi29qSM4c+dxxH0dPMkBGo72o
TY6zyLuy1xQ3rdqHtiK3/U9CTWZ4+54plXY9lCYSrls0eJvnUdbFr6yp075Dt36ZMb9NcmhPJGIY
p9SLK50543EDC+tAAxIs7cFf0M4MvXzBATwaGDJy7ftPHNp0TAFb5Y0WyYQuRiCapugVOM7pGLeI
gc+InVXv4KjhzJEAVwvg+wTqHQpRIaRFOATjnIAQ2AWA92Ho5KA7KIzSXG7HH93m1xjyGTX7EITz
LHuSGwYlRzxJMi3AivK2kmou2w6LoF2G6Q1UdlCHVHAvgPhjhfuqGfuCHrL3IwuEPQTJULktvGpV
jN8SjF9iTcsUz+fCxK9klVUPJTP/aZMO6V2fZ/o5+7tJCKzOQB7SA0+Xyj8ltYT1EoqQFt7K4N3q
w4ItLWCtjAeob+ZEzAqBnEg2h5WhLAzXf8jaSTUw46S/yQ1k4vQpOpPZUTvTDc3uucgp3wDabYmr
ZHd4s7qBUtR4NqlmJwjDlRqPxifcH01eVmyQzuRpAOCiAR4YoRFf3biVbALipKBEXm5jVdPcF3ic
eWHE2/ZIcWAJ8yIeCIvnOhR2Sjpqd696TbEd1gKzFtJdPi1gmQDPneBnKBaRSn75Jk0vE3gA7xJy
BME9Ab26psSX3KphXI6JZTiwDtCw1W3li58BA2wxkYoM9Q9azWKgF4SHmJduNUbIS7qPmJg2WvI6
Yh/RuxJzeAfOqjeJrWSLNtWL8VHP8dvEnCOGvODpEWnXYD82hUnIoqUsOtQ0fNdWid/nxz0sDuzC
++txFK2UvoOSFtQPwi99sdHzhA2WVqa/stF7ucT5pX0wjxhZOLXlh5UDJ78bPkfDlCIsAIGSKEB+
Y6TXx0zhpmG4Z79K6YqbRRDbQbtRw5YmR6l2amE3WZpeZ5OwQTTkfjNY5AIpz10cExksX0HwZrTg
7tqQWLLCHJB5KBjTBwbPnZOdApjSVkcK8sewvgwkkIC5tPAztooRWXGHhyomnAtsS/ivDARivJHn
8LCj0Xgg2Cebg8i83oDQNdgTtPM5hqinYVrPZWT4rVZI3DRK0NU2h8C7pjhob7hRpaAVIoWAafx8
XPEQaVq9InKl4B6feechkgiss0XAqDxnre8jsbJd0aRVjI04wMoF7JB0tUUfFKYdQFVLerdhOuV1
vOC+a3+dp91/6mJEEvvgunSe/JAUub/Oa71JQyHEDD1cy/yR5iDHk2S+IEW8osWbb5nm0qTQD9F1
hIF5A2kgr/zto9prsIi8amMH5hGZrhP65amm0dYoDLT1FGM8ga6le8+NcAzq6IX55wwCiRPrWz8A
jFSNbJnfTeeTIl9CGqg2Az2yhd8J3ckg2rbs5TrKuQOPUlHKvJ2s+93sv+HKbEq+/F2wN+wgXX9v
N2MG+JJOESIChVY5ghzOF+L+Ulzt59c5ixwtvhStZOOuMZPYnCe7b2p2d+5JePEoQvv1XSrMTmMm
Fca57lSEqBI6vipP9LXUmYXMy/gSj13vryvqV88BceldWQTs0pSbybCDtw3amo4Zss0xB6SyBlcZ
dxO0kZa+d6aPoHjEJu60YQ9AJcC7amjrANNlEI6yUU7LIaVfDpCYxy5P5h3SAXSp7OMlc/1WfkGn
mnp4hm41HeM7sY2qALPrajxpOcI8OlpMCAMmmXEXQYP1+C65AuiGXqFr0fEhfO5aD20XMgEW8xc/
wQr2BB1EfFrRzPvDBQk/F8/ZNI0KDZMd78uqObyN1sSoSDR0lmAMpnSdskj3/77L/ZyK5yjIDA0g
tCjy1kvEwe/yVnFmMlMisCUSxx1TOG4xiAYWvyO/mp4j0A+a7aRLay1IG08jD4VwYy1rZhIOSze1
Vn+o5VpoXOr8oPL7rG6VpkpPfnFV6YuzYltNBPwRwCKnv6+Q6CpliSVDW13QZS9GVvZPxMxpNteJ
Ud0pVklKnKuvJ8eo/1GvteEdwwv5bdU9Gf9CBbmL2cSrB2SnYToH6HlfyDKCC++wcPwOYHWLkZR6
95G1codlU006S+YplxcnawViW1/H6USM3haEI5XCJ3fBrFGyHgec7amz0DyxGCGmemwqSi9waUm4
FzvfLkRi4RXva+wlD0IH2EmlyuzzskRMoyfdCgD7OhF8JhaP7fzvEvWdeqnJ2RRaSOOk5AhOu6kx
RH2NQ9/0K5TCe4NevVAPgdbIuS5Ldfmwh5MZ5nSlBvdIpHFC4KAqsjTBWCgQY0lxxBJJ3BXpqmVh
nOuMS34m+fOpyK3Nd13oBd7hpzmzj5RY1AM0KtVlkrwZeU3Vi8rfm3eTWZZCHoKFtHF0+2B7BrXI
KMuwBGffx4vofjaiZup8crqJ+78lql1s0MctQAmRfpT/2G7LIFZs/x5jAOD/FF8a8UXpVsgfrIm+
14+9EUxJ86tKFFErJp0/lqs2/eIdv0TgkaPlUwtlFBoNnkspXBn8nRHd7HlXgqZYMP8EfvFmuJKN
8tLCObvm5jyhUFeU4YorDlTfP9YXOxxoiDee994RXMKLVG92nlClayuvemEqG7F2xF/n847eiM/g
70zDmL+xf0m5kH9MmDj9q0ccZc1FFnNuJ7lCTBBomAsddmSA8cZiUPDka9YbFsWkbKGi6CQ4jVdF
wuPAmBxYCNShJz3E1mCmFeARcBHMZq7s4qQNj5NWe2CCANV9Aajj4iAN5QDozVnsELnuKasnmyho
MC8aQy5QjwsX8o09t1PsT9RPF7gv+qpQpfqMk/p2x2+fwr92Pj6NklNj99bClcaZp8V7bVM2Ov/X
bPLylW5InYujZy7blnU7oiXlfJQSLjJezoVEkis4p/NBtGQzLvC0/xgUZ57IKpfBgogXzJNzF9+P
OolurioqFqoEFJz2tSKNSzQXmbnG3NZ6Yba0jV6hIFp0/PrMkWQctNH7lSBH3b7iMxbK97Rj9L7n
7FADHepRyvBJYVzJgplBTUvI0wQFpC0C03L2mxjAsHXVsRxt/4XWiR5+kDEJ7pyVDcAkYA6mSaNO
U6lG8rnWMuU6YxzOBX8Y2rydSc8Vn9t4JG4izEJfjwJzN0VQEi06ZG9LlPjvp9ZrBzt7gJyPlyqO
NoIAwjfS6WJ/qlMrODASNofgO5NEocHvIi8Y4gDkKdJoaUj8EAcZ0GJ6uIjamKf+qSdRKeB+n8cO
sat1+V0lI13GJelJyj6t30sR+8BFLscGpyGup8das3v8Cu4/TLQlhEZiY8Y6msoYQwSeblyMqZdf
I271AHXTbJUSw684IocSa9v8oVGipYDMP3IYCJ/l8hHolg7hicSWmg3uW/H1zZByYrJlauPvs6Qn
Qe+bvuDyBaQXIEj3lIHn6R8eI1781722A0OtXbb+WJ/NG5iBkHrTUvv6owRZl+yQRkZ9nY9StABo
YTFFBPdFuIWaLi0jIKt/yqikOkNJhGtBXgi+rPvjgRh3WOOIpgQJZrFPExAsMzWNEBsMe0L6/rVE
PBP7+asiFjLEHlXOapzIinw8NMB6GRZaeYqDJh2OHGvlahyaUpJ5bn4j+OIRaIuiSlHAL9UXYHJM
nBRmzSJgVhwfjoMrTi5KZk13d+bZhckWg/l7GAKaGbzm6fR2itNhG7MW0kXsxX3b9JooaZRzIwAf
lO+IFVM+P5CXBj9mw1Nc47vIwRiYAv/tz9PuKZcUzsLkTSz6BZEIlM5CXCbWV1JWXKiaYuf6eIMj
vjFMzA/QiIcISFGOciMUfeC2PHjE93flhufp57PjQY3ry8tX+RSGc7TKZYBqE4L/VI5hpUox/2cx
OYSijWE+sawmff6JHqs1wya4s4GGxRTSt6vcXZZzEEGYxEJvn09dAISD7++0PilhqWYSwBu+Z8z+
fNjhs3WhTfi1R2MewSs0GKqLlmW75r9qdgSTefHlsbozLHxl5xuel70Gqm63SbbohcxJKcOO93y2
+XSqg85IWV/8VuN+qSCEIdGvbBbFIW1SZpKKkOGmS+xllWSkrC6WCDbt82ZlMB/MJca+Gb4qNNWs
Q+Pzabm/ybwk4nQh2uTgkQb3aKWsugb0u4bZmfKWecmOCsFWe6v089kX4/UM5viNQSV5nwTFxqSo
ZAOg7MzTxXq4SOaeLTZH58SK54tz5ANrIiTpIx9omwaIqaEZ5W9Kv7nwxUbPtmPYsL2wm5U8+QOX
Oii7rljBWtWCa25Lzicf3Vr5SeXuJaLixCD84ft6cjVUNgzwTtitFooinbwr/mILvkfeI8N47Mw+
YFarIJiuykOnZZHCdCXeNFJmRp/uE5OVzGLuzgIklNyHtyZ8ktdWUD8ekd8hdkm/H7+2kpoGkFQ1
yWYqRqY5Jowa846FQo/DXqvTaLdwP2ST9hzey7QB84eMyphQNyJY1is4rFBW4+0MJ35/jxwdLY5Q
ne977IFLfWJqqNdkcQsnYKcsNfPrF5Kpb1mLY3f6fRyN5CFGJkaRhoY1ewNDqucwHym2XJQa7JSx
lwx7MynUQjsn7sB/qoUPG2hd8qohxjnRYcsFLpSMhSYoJXVW9GvhhYRS5bXSBrzka81YjMc072xq
nee52PoGgNvVC32znEMMjaQDLf5x4F41nTSVYfhJqPnCDON77OUK/HusIsL/Bod5AeWw/2xpRsEa
rDm0cbr31U0XMsxYLJQfY21Azm0W/eWcWLeEsC2S/ZzSFGD0KY03Xtjt9IT15s6jNBAHDWMAQdum
Ntq5QTYBTmeyVGMWuyDMjlRyP8alud1fGlDCyR0D8GLXZP/PFIyfmp2lDWp/H0TF8vW5hTi08Aeo
RlPIMueDy0YaH72XHCOWPRdifD5WXzhMgR7YgAs54k+ttfn+xm2d+W1UgYmRq300YdAdOUl1EFYb
qAJqpCRP34maeFdsMOeoVj94miAr8NMxKpqaKJ/2tkI6bxSO6N24gj4/VgRAIyws+jgH/Bhns3mR
OKqqf88K439VMWaoyvtFSNiejjICxoPNPnffhmb+FeHf3pUij11SHmf0EsVaLOmeC45UGSbPNcHM
Cgu2vfDGk9NIxV3h1qALkI4mkBY5t+UWMBZY9uV/0dnUnvMQLRUttm2CMDPVVjAa7Fv+DODbLv7W
gFPOX1h6QxspI4dTaBdtcf6A2W9tY+kTWgXgJVmfv4++ZWSY1NbEeGw43G3Eoehn5Pr60JVwkVnB
pSdERmCsDIoTe8Sume8/xKOwnIALMNU70DBzFADDIL6LH6lmpqzU2213SkKcqXpYKqqUo6aht6bv
y5gcJDNNZZndzHrxiKpIBZLjeX/16oNiL2GjOoI9i9wapbC1jJz6dKkMzpNxc+8mTTEXisFOLlO8
Onvd3YDMKr0zKsLvfIfhwa1AQIP72t4m9H2d4q2paiPihUEVW7v8Irn8x8QBFE9aADvs/bHXykxy
uTxj+fOVzD2bBrO3nw6is7tuW0BWuY5myRBsOy7BsFa/d8nlDfzauX2rt+MZkT62Be5MN3AJQL3v
D2dp/953yzA2Y4lukeVN/0Xzzc8T/3BiWFVzmWAschkUEafBybQTCBELrgXwjf2hzMn2zvdJgVqv
q4mlitcRN86pQihOEF7YaLUsszhLfE71Itf/kZXxJwwb8cKd8kYVuonheAxR35lzqKsIidOU2xEV
at+ynU9gTwHJkkMFtjf+5FC7xpZNyvtR7iC04NJEWgYVmDdpVT8hnuLLQ9j/QPRiiiXywFx9wB+u
+PjXTmjDCJEh19llDqipqcdRADE7fZcN9LV9PUEPvtTB38IptzNFJh2ltHP3WZq+GrDl5K6q0GH5
DF7d/2IjvVqrycU7XiuCXc4fCI8NCmkVchK5n5B9NP9c/WMHh53eWzQtTGHhiiL0IQ7GDOPIWHz3
ZY+cAZVpvIGhfAD++rIbQAE5UsmiU/TyStW6v6I1K3KeOPMbDWbuf3Manfw9GZfLhWGVe5KnHN3n
UZKZ+HPQM0jMse5DHHx3048Jt5Dn5rB1ayBiUEuSjoAUnnIrmHqC29tYsu5JIpPZinSDLmorajBF
/YZXQRQOnW9ClLcj4Y01L33gT9xiA+K/GpzsoLsjKNPRnA7IZN/R4r1tghe935RYxZBdttz7uwQs
pMWe9PyaSPNXhc9AN7eGu7SiOQ3QuymQyyp5ErntevxjMNZqTmaECNT4tovgXnF/fzxXnXwXA3o7
cihS7JShMj2dJ/TU5VqoiEmrQ8TG62AKW2sBF+IqzpW1rPNwOSYVOND4GVigWIGvCHw/rRtmHde2
nM+Mb8vMDaivp7BRp9LUkAuwqpYL7gLG+rcJAYI1t8zk5MxzrVY5Km8qHnmigsc7XKAMAuu/iik5
NZJEvFy6WOW44XEErwv6hZM4jiKHjfXjPOb+fqpS6IGNsOHerc7s1e6BaBRVs5ZKkw1urd/P9ks6
5J6vV9Ied3vKrESxwbuj64N811hys0jDq7E9pqCaqxkaW+8e2y4A+Gt9A+16yRvI7AKvsepzFbzn
wknlIgAz5CUjQOTSltUHbG2L6DSr8QKvoV6cqd/25jaV9CqgdFeYL4jvCxoqfXn+59Sx3hWn8Lfo
F7F9GNYCTCRN2+lxUTULVN/IZjsP7Gql/6EDxIB8CGeD7SS568Pg+vGQTvI6ktk1TJXZEisVE+7Z
/+ouQfR1iRTHJcd3jrlEgGSWuo90/hT/AH/2JhjyMxa2I/Pht0SmqZAkpJaJFU4xweyUA/CTVKjz
qyTe+GkPWdtO8KIDJnlO//vzIjjk5h272Ff17jW+kujm5/Szp8yDIZyyefLk4N/2cCtpyL92iHCf
PeQ3OWdP5LtYt24ODUmBNz22+BH8VKPKD7Q/EmHoQkpu0AXHvYQXVboBAF3UJLKxrrToT3TuZxze
7mof8PRqyqea+q0RbEvsncqNkG9hd4oiWS8d6M2embp4t3fkt8DGEvHbA5Vb1SDWTmBOyd5ctBCG
Ck8RGpuXkvNBX5/vcoUIZo4TCb00XGwJhngUyYe+ClM1RaElcQ+cno6mzkor3VpAQ5W5PzFRTA71
chkJy2JlhddknIaoSYXE+lkcm6Io2PgQueSHG0gXtSf0A3y7lhPPyOVyMBMKcGE2VcedS/WlzfL5
3xTLTNj4jfjffEfvCJYgLfFAGpcmvZAU1Il9ZVZa0fp9QaGVNQzdrZiXUikfD+mSPoytiCe3scgC
w49cocrclhlWyeAXBSJrpCIB2PiMVmok6afnOXxsQ7WwdBq/zqeWWRCkpDlbRgCyCpssFQOI9Quc
V+2OJkSu9ktJEQUgPYBc8FbN9gZe19hg1/yzLH/YqDpiuj3no4iLkA+6HxpXdOpPO0eT7V6fOHs4
e1da4Vt54sQ3U0pcaQPrsLTl8iH6vXaLhv7QT/jXiKZOLioxKYFsMiismO8ZzIk4OkJ47dvREIz4
vJXgSs8c2fLSD+6zyO4L8OBA7mbNh0vGBe/Lw+m9HLghVcBIjxRZXyWm+A+OeVbzQ62O+JvryDMQ
kSLWSO6zplhDLmUBVLxuKpSZm9IZKE5CF3etuTYU3KDWAYhx7M1vEIU8SvJj6qNGJRvGO2Klm/0v
Oo/QRfngf0ykOJORFhUZ+c6W0i9ec25rwdlN3eYMSsdGhtLPS3OKTmOBPyGWxWEm1dthCnIcwsnq
nAdCY9WnWffd3uzP+guSOvUq+LaecNr3E7MfmSv/y1xoesMswC078rNghxgGb/wu2MZdxj8CqpN9
Dfosykqo2rDuRHOOjKWjhn8zjQevbJbXk1IT+69gI1OONiHwIP9WdpK7zbKv5CHIPTRQy1TmNLgS
zJ24SVM4Rl124xG7KH7f2efX71x00FxoJ8TCV7pp6snB4JzGajJdRVQRHrprTFQiyiEN5vhWlJj7
u2rnGAN2En1XqhXI3G8ALnbTiZt625z3zmQdgvpscS5fw4u+SdxyJXuPLAN449dMnPOPY7IPp947
lycoFC848p/ozz/Lx9ae5bCqQS4WKRuQ0D9Q1KtboPkhA8MDXr2Wf4+hq2UMIcceYQ1SOI2sLddi
7RDVmWrfIfjAVNjTTjps0vwyfjGV9O3ZAW8W8gHwaNt2td3mnGrkO+CfXUcmVBE6jXRfABQYnQio
WbSNxGaQP8gQpSwb+dIISkKXURd7ICFA9e/T/dBblxR5hbhlEmcahJF+Zda8clXcMypk0kJxjLEc
QhvdLMMwzeyReFcYoW+F0/UVltiRsRrCLXl9867cDtZFETu6NdG4nuEIBMvCcIDCf4nRawIIjQHB
ya7gK5pCGjC9VnrTNOGklDj6v3hVWYEq2KY6rjpBPx7aPXHgTJuogTxvG+zrwJf4eL+v6/ix3lnJ
HmHqymAlqTZEIGsQlzOga+SOW82kJ/dMAwxigmGl2tI/J7LJNgdhUOidFu89lcWer3oXBiGWVBAn
o2nS6b9/EkjJA+nO5bGOAWY857vM9fejju7B9QyutjbOgh+fxUHSWaYmkU9Hc3A+F2TKyiOO32Hg
gsyuU4nsZ20klUbdAa8q0dhv1v+0bt60IdOEaxUNEKqhB7fM7Rf+Sp4Elej94H6RT6qLkJKbkcs0
JPBOyqCzXXtT23jzX2yGYO/MjwKWBlaiq7I703vXndcLThr18dyceUd9ATbG3ZTiMicAy3MMgqQG
MgCRDjHxTp158ovrA3S46nBnIKojPZjaU7r4gZPffV19Hq5vABBsSNSoHFzC0+apRfegEQyCTosO
XOqNnp6JI7thtJugt+2m3hf6DltRmfpiWnO+an46qb9Q5jDcw7kdx0PfFTwqFrSexd85NrLRVUF+
S0ECt328jxPY7yBoniPerbRUwwwAsYmmpFvZVFGSiyyFG7OTA3bGGLWrLxCstfjuZ945aNkVkXVc
RsliAmI5EYR5XbKCTHNRmkA2K36dkzZ1USWqLB6j4DqglicQCARf+M2mXLniGxQCzDw4KhJlUkmT
Pc+kM+uYnKn19WtsUSKnzSGfw63G0qQL4Uzje5rQsIRG+T85aI8XpLjqloBejh24KB8MzlND3dmP
5hLCF2NMfQqU1j10gVrNVs1ulHPLnigqHKFQw8pIx/lU9RFEyHmjYwBAzKOVF6PaLXzHjRgCSVt0
7RkqqKzCPRwkIDj3Ze9jUgUulM/uTSb1u/H6RETqGbUf5VCRID4ciNYcgt6cpT8ocWY7s9M/FsKK
36iuo0PBK22OZP0s0uj0GWv4nKi0OSORFqlQZaE1+9a7A0iGNT8cuOWMd+C+E+2Ajc5hyLcwizZ8
KfBNM6qMHc1j7fc/Z/4ETuyAZ3ODfyjYi0L7R6CUZxa+RFBD6GUeGkRCQLXhdl3PykeO3ln0eLWE
QQKx8Ti/uQG6Zra2D5kqMVh5xO4OARKzSW2Cf/uY9fxLLwUvfblfSHH+DRQZHU7UBXdJIJ1rzPDP
TqtXXLg7aPFzEL1PDY0qscKl9+Q/fztWmwe7OzNzMGd1yEqjSECIsgkCqO5Q100SJcH/JKet0d34
Tq8efNpUtttlp66+bFnijqJU3rRFfYnZmD5x8amagSJrB6WkpXjFM0MneePd16hv9NMkcO827Lbd
A8gup+QLuq0yuNKTm4PZhMVXOJ+HpgW6Lo5Fszmxt6jmtaCp05ivnSvPTS8UNZp6pqNOelNJ3NzV
IKw6HJheICNncmwXXN5borDXEVgHtvT2x3Wd9ffiY5AzA7kzoBaqDyTpMKQwcLdPV7+xKIQ3McQH
HB/MLF8yDmSAJMomDv92sZlnJmADHbZFw88htybxAQJCo30JqHOgv+KzBCWoKPL+ZVlZ/gmyQRUe
heTjvEBwhyazTZeoypCk8limkCOHDD/FRYwlkmWGJx8aNmSs+IsCQPwVs5Z/YhmWaWiGIx3C0iTv
ZdYuUiryTzelI25RX5Gg4utERSN58OOKfT8eivogTUgf6ytxoRDMC8mjxjXCz0AtQdZ4mAsUL0pe
8hG4pDSiyIEIdAkXyuVnITkeql3xx4X/tCTcrdTuFto3+lFONtzbnruEN2a7XeOZKqK1RlNJK/lW
8l2erGClex4nbcffgEKO1Y8wW3eNDTHF/PEckCiNb6WZVXkwEe+1RcpZeqWpchwFpNByHFNDLYrv
aENGlcFzpOasxVlQUibCatVXEdIWvTPJ5RysUmT9xGn91Yy4MKdppEC0YiQWrCCzEq0fc0NPn8PV
qnm3lgaZkYPvgXlhSDqaK22X11XG/dOohkrozlRZ6Aom2kzdJD49hA1ZxL88UgFSAVWtVgnTnEfo
lWXaZHW9Q8f/RRMmHNte4NYFDMm5pHy+QOCB1Yv+1vfMcpfntgfCAdmb3gmU3nS68r4ivKajKvhk
dXqNsvYCd9IgMBAt0+MlzeR+EPd/Em1ZHha8h5L55ExBBo663JXrdLjvduUfbr4w0evqCxF21oZa
vcXEJDz5/PdV2UhJPmLbMAFAJ9K9I5muCAL0dJrn5GDJ8013UYOx4/L+9iCxAfJyHz5G9Qv7hlcw
A0x6pd0yFnmGFu5lwiMzzD2QZHpNuu2bLDtPaW7KIZKYI2BEeDd5EmOZgM/LTLDfZI1/3pCd1P2f
bQiRmBMTrfPn3HsnqxEuidUFflo/jLBzfs6wSkt3VsSRllcuiTMMffXYv1xL281S9kjWmA7tlCe7
SL2PpLHfQlTLKjBlMAIScP3LEu1sqILqmt1tHwbncOsw+rRh+mh0rnY3eV+vU/kVYS8THoyd4htr
jCL27e0rzRvHu2s1iNiaE+czYn98zU10gcDOpEHVZAem8CYUvzJ6RS83Q4klnTx5pl+NzyzNE082
bcKUw/+WFtZVrA+BS1O+DWZo83Efpo9RlpxF9ehpwGs0+WOOLprXiuXrM261kDlakyGJU34QuAYY
HFNkvz/3koTD6+ow28z8WXkN0fFNWdBmhthBJezcfqp7kqtsyCVHP9f5CHtOfM4ZWhG1tPgSImj1
qKZQRBpn9yQVyhvZrzkVfnnlveRAFrV+KohECCwcUqS4pwKE2SVm8YqojpdPK0VTEh7DHqFmNKXL
PqzELX4qqmMtHq+IYSGNQPSoFs/jB/sUu4wnDX6vsEiVwIX6hR7c5eTPYDHyXiq1D8FFej7orDAE
wxiyPAo3V3f+7kDGecQxwhYSMC4AaUU/kv4S3h3FaqNwTh7TztKnTwbcEEXDJ1xGAvbIDT4tgtf0
j8JNImBGIWni9RyYAa1tWJUzeHaH1eMJegB+yr39WOMY9DRoE/iMHKF68dfHlBYMlJCsiD5lnbWW
qfDrWwaGwqAC+VXfCClEwwkD7taKGzc5AqFokP4VNYD+BuhV+nlPeA8mm20zhIoOSoi+oNnJHHm2
Sxl7/UIR8A568QIM9d4h1q1pY7BD5Z0o4583ZDKBNrnSN5AW08ceiREHtIehydZpneGDXQ6nrBhT
gU9S450yFcHToTMoV6MXjqsmzYYp2YHBssz1hwQKeARQrhZ1crA2szax452+D3z88n0S4QvjNS9e
D6GjR1CPBaeSK2lD+fcdfr1lb7dlJty2W3jVIefXe4Sg5adHUk8Sj+pt9NYoE/rPHps/w+zPTy/R
vyKomazCVtbMae8FJIz4YEoS6askM5HnQWBdf3nKkiV2tWNn0MzVf2bKcEqN0l7lx/SDTsiPOqU7
ZacT4CVcQdEPSgAZIFlvLAyqRiQzZxg/up4m7Np56uLLiOIVl1Vp/U0/30jRjGh7DZ4yh6rV56Ye
M12WpwbIKSuMhjqN3+sbW2ALxgVFQd0PAVEA4OHFrwnaHPon+dnVpeezWFNVupu+SwHlO7ShBbte
z7AgqezM9nLxuZkLya7ezL/62CAMBxRhPcgrsaPqo0GNEX+h7kJ2YlROd4iN/YNRIpnkKkqO4JLo
i6gulk40dLzEbO4tY9l3GDdUYt+yHhRywNjYKZWa+pLBy1oT1wcW4FiXh3N2gTmoydD04ayg16rq
klFrmWjMKFXJ9EyU/2PEekrVb7m/edRq8MD6Y6NmYvZddU+Y+K9ZNUJLFdFc53AkMr7EM81qSw8C
IQ8rEzslYZ2BpYi0B3gSc+M8HhJIvZ5tA4iz8aD6sObZlPCAQ2DAXsQ/jr5hXeWmkiCRVdPfDhso
/8errwy+S56MTIfSpHVR3jYnN+NIn0kdsmD4rjcjxMfKpjwAynGt06ChfuqWnnEvyuq/wq42Ly4c
rm1ZPazY8RDlp0DYeGMwlcmGw1edCNq1fYJ8hpCraujv37I8S4MbEHLVqISI63aSJMwXkCKJV9nt
aukjjDYDQlevp6OBKSE6BMDbyQvpvfQK7b1qD2zsCsaIfGBC3dqA9scjLF0s7KwCXr6JSO/NRLr/
L+Zi2lhNQ5IaXhgKyRS0w3aEFU2V36VZFWzU4wDlkDos/2EZHVcPCYzTC+drYWyTF4eRFU8sd8RR
4GyCl6OgZqgrEzyhYNYxVzlDpQke0RgJadnsGo4KlpWIUMPPyyRy5wNUXijpeHlKYG2Jf/Ui8CcO
pf8eYFx4bc/l5+jwNhOx4yULixyEa5aL2/dhMOtPbwxQN4OSixsODVPUo8lTaO8eApgbkLtoO4Ac
xX9o0l8F3z+1qD9P4VUo16grHX3D+JKUnK2qCsrbwnHJGMIfQ4fHxDBhuZEakpa78vFvL3FNsptd
O8YT8WG5+h/PJTb1ns/6aSAbHwzkhqsLqTSROAjhE71h8QP/yBWt3VL8I8TSZjUoakkLwfky7iBi
6qMVcHNWlSwqRkId0Ehup8ow5tDEKtiidAA27SV1GQNNUXwMMdMgWq35rT0m7ZZPhiN1uKJrPrf5
yfzRdZ/Cw+FU21TePR/VjdHlg/MUVgtMydKhWSE5073819o+pWyzz2BId0snzrs1GJBT5DGMpajd
R/yFqf4d41YVmyihTAUgMLcbmk2p362vxS4oyE/sNvCDB7sHAo7/bgonC2skAhDISZrEI/1OUhFs
n2E/zP/Glq7ANm41NDVQmub+BHTA3W/8hUjeh3uHc4ZVGwyP8K+urOTHRIfXJCzaOnx3W2VXQR5M
S4jLcHBt8nKymTNXdKHhT0ouYUpODzEl96atbdq5GH/CP2hJG0PCHWfHvVWSn/pNJVi3TjfrV/iV
QRkNmuEbzQ94raFhoY+5zS82T8SmjYrrgwKUchUQiwBSwJnrkvDfNGc1GKR3v6sy0V7ZVnU1FTxV
qRPQrLoCv6yZIzgTU6VErrnbajunk1uXVpob6ioEER1ekVgeaScsELXyuMbZDsXvqoN6/X0AOcvH
pvYya1R9b5ZVgVDefxaquBE8exjCKMlo7Sf/sUICSUckjzdA67IceQCaU76KsN1q64Q/wFQvxJXI
3WRYW9rw7IBpof87mofdYbTYJ6fSosn/k9tYLRFb3icS9MD2DZ6x+upE3j0ceoQSIByp98Ldgjki
KmK5N8oDi4c5qch6erpp5fCY/gz/Wr29AXmJVJCu2GO98QdI+TT2aAfNJBE9gmKJXFrTqmaz7v5U
nQauaODTvqS12GcCXFfynfeLcwzCm3VO6u3PQDOXWio5EpNYkpPuIB3M11VcVCrMUc5YzHEk5cTP
pJ7O+y00+D2pWmltlVeYWeyaYe2q9jQbf1QaHi69Eh88Hhji4WH/NcgYnWNIvpI34x4vsGaRrRv2
V8nQAPafPB/Dt2BsxUTXOYetWTjWXF6zvnJKKGAl5A7xYIlFwdF1tRnxi0dX0vYroh/38MP6TCMS
vWPiGvWd9VRv6ncabmCw1RyrjQmdIUz0aDzu+WPO4xKDZpMoTvyIlaiC2qgoOmVOeEX0mR00OSAQ
xlvMHKYk0v5mFIVpboZl0v4swWrdOKWo8uynehHKCh9cAeTZmBkzeHwAvvVQZ+ExTwjbYOHyNUY0
ZQfAk1u5b/kjxfnlVWGK8NL4EiIg8aEH0QT8OhDksTr1O2NO08Jaja2dyyFVqwPJ+vJKIcdmn/Db
9wT1p/YLfADp6H65DoyRCRgphFYA8fRtcgYGnUD++h5OBlsleKgsMq8jmRMCfPHl5fMZGyHI4OkN
lcJ/CurjBhhzOGq4+AZNBg52OIhUY7Ilas+Gg/aCvdyQJzhYTy0hgVp5tmWVTxGHc+ikOzdDC+Ir
TFAJirbpIEs4PEquEqC6NwoRghFSqd0fZS4nwHbIhYpFg9ggmvGwAd2JO4ySh4WLrOFNp8IXWz9O
A5so4LTtxDg1XdCeu3yuD6BfjV2QLzqQpffY/lZk7EgxdVgxkLzxmXcNwD8LQH004Fwi0IzhIGYa
hQbutzFq9I4s/lRuyZ+/sf5iwltDA3fN8WUmYT7nbJH0vkkLBI2uOnPSgZMfiFulgaEFBrYs8WZu
EqsN3HHPD+7g4nAmL+0VUyWHeLa8UQULswQThAthf0u6R3cYpTyFOTHdZtFjes25etQvOl0c1HOe
RCy33EWsKbcEMwvWCT1hotJkMYGrX+Dki0RKO3EKPWVWg7Hbc9ECGhCzVmG3DoOE8xZTjS/pjmX1
NhLHPR/Yp/EcrpvqfZSGgJPNEo1iQ6L19lS7H41QiLtTgMmooq17WxhGVuD9aHS84/RAYCQOuVpz
KLmNtrAxiNSR6bjKJAGC8hRxZGcoJlglqYa9NIgOWrjm59iArV8YD8RYqdZ8CnLPc4wjMSMWnoMA
xPevnGLobva8E+BQmOtnaYSC9g87uIaalKYu3Ks17enMGfAZtbaMy3WLf8j7XDCtBZDp6cPNWTnz
IU3heh0XCSmckiKdyD+IvhCT+MbItc+tIiNrMXOqs2GEiiGZw9LENnBNSVz0wnovMNdWUXtY1CTJ
u/D7ogtqtsl6MBHsiMCtp1iikSvu72oSGQ6yRSRti0Hk0UV5XmyRsLIUcVCU6w9umCTw9yWKr7Xi
v+/ygqT0b9OHb2TwkYkMY9gpTcGoQCcBhrV95n4Z0VdEVpKyzuup5s5tFqhRoahiSrAtPsnu7SFQ
JDp8dwdOjRMp3WY/MfAh55ZP11QnU/gEYq7h390cTm9KVQ/QY25Uw9aSBTZoX3IW3axmC4aavYPu
6qoXymrewo+Za46b6v6zlGleiKMmXiU6s2SeIgnzoq/7UKdbgCJJvmnf32ND6Ti3xOrPWjuvThxx
9W4zoRBzEgy8+6M0YEzNxPlFIthhMRTULp2D4Z/Zh9he1r77ofu72I29VZ58vMl8MPrHI+uIi0rv
2tlKFD06wGZcTD/X94Mq/O+gus2s9rG9MUznhBsBOslQhto2wVjdCYZxpSGaDvCabYQkNueOBWY3
o/VntMBAnkfD/UaJDQsYOhnWiyPfN3ZGEcDitMloDF4KUfWOIZMNzQZqJW4Zbvlal5T+eNFnEOv2
0OQrK5WhaQyPRRkTnDQN4MTPg1h/MSvG2wSLZgDV8t/A/ii1ppTX4m/2EYc7YwkWtc9PuzYO7UAm
voU97Y3Zr+sYcQs/JXV2v8dpao9hJ6UjQ+DI7m/ORGbVen7LAyz1LMaUxGqP7pm9wGmH9jVKW2b/
rr8CPXB0tE4PWDmJSsKIszZLWn7KqMnXZFFO5kBa72/7+ZqzNuFoIrgzTw+oKYYPJ8Ub0XGWTwLl
d2eHgYe3DSfhPEqx6Sy+fO1XEarIsiQpBi5By9W7EsPmHbMRiPQiPBy8pi7A2u/Wk274hJu3KvLB
HNJcpII4HQfdA26pBsoOEbwzWmFQu+gARPQvdDYdfvaMXW6WB7ga2/VaDYtuwQ2uqKzXJ7AnFl98
eJIBQ/NQ541q63O/umO2ItcsmCmWLfJlTirRjpDA50ZAlr0txo8J8iWuA2ykRtqwSG3wv0cajytt
ew7OTBjtU3jAOHRAvVcI2o6pRgL34GPThEDSeCoVYzndD9Wj6TYtDp963R2m8C/xyOhUmoqGszX8
LWPDBKAvni4XYIilBaDPHIEePPyhU59+zhdTQNaqU4NcesMq06+9Q8KcWHPZ9cElPLoKQfMAok3f
8ODmDDMbQZCuqTXtyPf/ygU0qiIyDzRnvdll9FDy5R0oNq9IogAZnJM8IBRVm6eR9iz+X34Cl1qz
yfcApQfe4B+O0UtQeD7AxOeZXDg7Db+9amT4zEGs9LBRfobbIxkpGC8s4zEa1r/OS85tfx4Y4fUZ
8EvDEQL3OIOFbR+c6/IOIOj+gZTQQiBxP+Jeovxb+z6kj6Q8QQUPcdhs6iyo/sfDesCELMhSyepA
ZLAO4Vn4XHXuuuvm4t7pQrAdl91T2eoFQtC/Pm33oXvw+E2cLMIzA4H6/r2IjGzsCovaIS6XvtCe
tuBEsRdZoBudfftFBbyw6l8GrJ1C22IvOcVEJwRHuvL+GgCA1TOo5hgUHRLh3xpDyazAJ42piiLx
PhQYOTMxSMbDXcv+X/iE0L6toQPslZOrWrcJKQ29ufAHgE1Gnu0vree1XOD3HdMtyBVs7VCToInX
Rxn182HuumMUoqv3jAf4etMPXKsK2dWGcsQY2PCdzeUuCKlL9eoCsdt/t9pz/YCet8EgjP2XU8+N
Nnq03eTl6pogmFo372TesN2lbxPiHGygsyIItnazkAcelPpuvdj7spK79rb/eK5oOcNB4iJny5E7
zuhcvmURa1l0FV/FpvMPcFvfqFHq80uR3C6xJP/DER8H9rO5/zC2YpUtzHA3Y0b0TMMhiT063dqL
L9zeSs4CJN6PpgzWHOAfwC97v4uM5LKHy4NMjvPjLoQmnX5DaAbHZZssrnY9rxkDgFcQh+tRVAtl
Z+1UPhaWMsHiaVGgq+VhqffkWqRmx4srLf6Ta26rtyioSlbaaV8qsyNC0EoAwHJB7a3ZI6/KDp7T
fim1NOK0c8P+MpsfGLsaaB0MrUUU99943j90+zMytfFFMGHvo86FiQL0XG0+EL1KuElPfO0fkZGv
l+y8BhUm3xXRRXfUhCje88glarVN1dznq6UfBK8iSKpfClR2Wawx4aUCs96a5YR65QyHbH4bbsbv
FZ0ZdAaNcnA30sHbgdW0ZUx78hlU+muwKEfZMAHL/XLW8rsdZDP6HTHZ0ZuekLkkCDWlyUee1cbO
zkUxWHbgFPn03NjTAsPwLJDmRWPitvqaJHIET9dNzeYBkQl4TzqPGWpwKtUO6ssHOYy8cqM8IBeq
HUmJJ/K5PEsl8P7o17iOpcDEth0JG2vCsGpXtUCS2NIYynuLZpVkmuv14Se+HYGiMmreJ+YLtP7K
XFwRrIU5fJc8L9p0a0+MHDCyjv7QOLNjuJVJkTJw6NpmpMxVqhkiVYz/eiXCw1lBzJWFP33/9hG5
amZoeIPL1lwo0KYsHP/I4FVRj9Toftpym3B8bbW9B3ixmWY1pdzCA44oXbmGMrd/3FxuSqywYyfy
BuvwwouOKOnkyQXyrn3SJdDHgoJg8h8/GwDA1WwrLjtfhSh5AT4XP9kU8MAntdFprAsZcCrcHNI3
eFJKhDgaTzYAhzqGiDqaRqYLHp2r4WGN4eznKujzl73ofLExyQRrGillmtvE6krO5pMy5FbT+5A+
rgtDm3ck883vrh6RIDD+H6krbLyVkD1VXzBdWpSCzrn61TZNjSny4OWoQHymTcp1OsmMgoSJ6eJS
RM7hgz8EDUa2ZT22lKBLTsorxYD60cLMUQFhrB75JU2ajFHJuQqaTIWou7r8wVWzHqXG0+yJIuvX
Rfvui+VO5bzGEPeyk9P37gIU1Xz0Fa9hYHS7ckJMzTQ93LEYEegxaBCd7Z6saw3a6ag0DcechETf
JH6WeutGDRPbH3QOfdgeTPaIxqtGVQQ6fLuD8suKcWEcnmJVvxVTLWwCtYSKsKKY7UmDx0lsvLgg
1c5INB3BZG6JLP6f4VkBTq5/CQz+u9NP+EXQbk96rIVGaKC18mw/5PkS8X3MWZTlT+nEuPMBUsnb
IUbnjMb2slPVPdGvu9uylwA1Hf8um7AXl2pH4ZB6ai9FrJgKLbA143CePUkpzwK4XE8FHXyYEXih
f1P/kBzvhX9sMm4fIPdMjIOiNXVpXxE4xhsV2V2u0QP/2udscOcJ91MN7Is6s5vM4+VF2KN8ls1F
aC6B2W3RcYPTyhx/EShfCM19BQ5Maa1Ek71EiKpnuzXbpv9QKDM8+cnVye+tNi/UZrq8YUuWwYcR
VjxgMFtutK4QkRuyRagm3lEVF52CziYubPAoqTX+8POHrgUv3W6lUz7LgG+lxQxkCKPsmyGfe9D6
cKeEJrrsmTtkorBRyZjzhVI+sDPyZjDa8kJL6gY0KFotg5N5+CSP92p1NmfLqS5uElEOvlnvA3ua
7V7Qu4fVDreySTmNgT4M2IvbGy6EWEQw4BB12ecpvBSIFT2KuMucsvRqv/uzA0Hk69Drv877BEHS
7jpkz//WBz0OGi0MuOr/OtQqZ/KmWA8ICUZCQof7H8FOFEPnW9HqyUGiwqC1JyWeBSkLzYJNJaR0
suunHMQE9rRxCSClTlfvnH99TFvHEb2bUKwxSCM/d9pOJUBfmWk1tYyvR8LhkSabXu8iop1QNbSQ
AqUPIa3F11xBcmQY8lPWxtPTi6YJtTIpQdKM2QgmB6KRgvYwqRerCdYFmcpgG/aWd3Z6J/W79eBX
eUNz+2xbY4uCSZl7hBamnQUJM3Uls9U8nOW+ZIb/uJpBpq2+BtCHqkfR8af0QVjFlkCAX4I3VvFJ
qUar7si3NNWD4E6gjM+CNzVGqeudN7O1Ilp7Cp0og+1+NLLabYDsHxDWVGydIbJUKUUrbyziEMTy
MTCFpBOBfb5lBCECGDiH7Dn/L81iB25pfLn2Snist4H6WSyUAPjBDM40caLI2xyJSpa7PqZmOTkG
FV4VdttsZAH5QbxuST+xTgEJoBLX2lHCh19+S1TNe/GS+g1tAHJ2SzBIQcrtZHmPWNWdRjF4mMnI
eB9Zqobn0eaFzjjlnFxVXpDDj4lXDQJZJ+9YYFVyPOnF0WBhBgQlVf8Kw5CppxLhqitvYbbwxZMw
fK9+b3Yzjpk6z9OjDxbxVVbVOO3ZNHtMKm4zzezVTJHRM2YIE4gV7mHiKQ9VnCeM9YPkzTLRVSb9
f4cvtFHQXA/10H6lrHL4SDqDmAdTSUplDOVq9VQtk4/4jByv5hW7W4T7bmImBQfFT63shJ+6b6zm
6XNPm96KXamakwpgFgwGStDqmMbDw/cOACzNioV4UDlBHrkUe3d79z8PS1ZJicF4Qeag8L9Sm3Y2
9qgkzvMEKd9yB3XXtnfRHZdUhr5NjtJkMXwbVVF9jd0VcGEB6VDXooJupwGVlo/o3pUilDsB23Zp
48x6NoHePUA6z6O/4tAt8bE826VcTEFaYwYMYVXIfkAX8e0hkCe43A3HkrtSmHpWTMMh+xyDk5V3
cz0bNDYoMYfHJXeo1j28Ayy6q+TpB8En4aqP5GD6njL0lEvZ3x6gXUCQpFUjfwLaBpG2AwWGTE4O
t/JuOLAhz2v6wpe1ekGmNuAECVB/cqWHB966W+pBCP0iQGbBIGoUbbzdXWVe6Kvqr5w2B56vsH11
9SUoZwMflV5paX20PCeTG5OTkkLRRLIZ344EX/23pHMBq7ODkIzEoxti7mbuBB3+45qPnTSYV/b+
u7DiWaiIUDCykWChcbdD7oC6znUwOaxGP1ZvnrdGrrAgUn2JdFw9wJf7bA2HLtyxFeY/8cKxvi64
cCkLc94ecxRX5v/qMFosOeVwbOD8DmwzXOoPI7vFcwr6Z7LsWealuiiOR5A9p6iJaMgiBzRICIHK
Mwf2d8SwxRF9jRqXEThZR6ym6vuT08zgXwJ7PzGPYeYmq/i03N2Nyf2bc79lx2Ghl72KguS5DU4K
CYlg42/z/Rk/WMFdeyWUM/cB/a+5WOAXVtPrwbhWPLRi3vpe1ZY/+rpp4lXzMaG2i8fRnBDAMCxZ
2nsJIs28NazNo3RnNjKNTQE0qJnwWM5iOe0EO7nkUTQZy9vTwiUvUBP/8kfIwYikSuyqJgQhlkMJ
D4jaa8dT156Bj13xLzxnvgs6J2O1Vg/AEXCPXEggrwRlivAU50UGjG5Rm2EyKLbr/7FL6dfGUX/W
PXR+GyoBdZagPOo+W2fTwLSlnmnAdkC38q/o6GOWKQBGb/vSKhL3pH6OCsBwQZQ4HATOnDaAfewg
42IuPBXrTNpj3d9eez3S4mLesFO1N+CtHXKSI4iRkxhfJ3HeVRl3cdJZ5tqPK6+R22BW9hnVMFzF
k/hPBelX3CqKrjEj77Ow0HepoI6XTNpcBCYEULd5UWWkYED+UsOkyrMThZIap7ay7/yBven9Lter
ClSJCQUVkJ2pkQWSBxPAgrVNwB7A4r2JGfpQEZcNzqBJRy7tPiWpci/ciCuc4121d83Wff/PSlSo
NMMWBfKOHy5FSzBuHEqFEZNZwsvczTTiNLA64Rou2ZRy4Gamnil3FU47z7zczue7lvGcccdROX39
xCiTNNPPHKID3pyqGhp1gn5sBFia0WU0u5Q9FRQIyC3M0BxRGY6G5fuynxMogj5AJqR2d6ybFw22
yry/H5L1xKK8q3oTaNcialHbZnE20bMpwZe/vTy2UupZP4UQ/GLO6ceJBVy+ZYk3+XdmgsKmZ9pT
u6rSvmsLreeernJIFC3M3t05u0JG/RupJEZgAtQHSfzxQ9FTslburDDf9hg9xRNw+iinEx3gz9Na
Yd3dkqy/xWNbWHJc7N2t7NJ11IXkYkA6/YopynFw3ezMTw3W9D9SZoY63BLjyNUSN3uRpJMziLDh
HlKSynxYiHV81haTPZ+YTddmApjpq312lALR4mIp1SJTgUzjih74RYLyNA0CeRSogGrDhXuHJm/a
UgVuHCC3ykVe4CQNNl2FYLH25l9Ee/p/GFcdhdZGcQBp6zhhSKb0SN7E1gzHfaMhPjr+IzZ8ri41
ysBLlrDriyH9lUNroIuqJ9dlZ5Mveu+/JQDjMdMK0B9lgT/mBvL7smn2DpQWNeXXzDO4aFezVCQz
i5dUWONTdZCSkHAp3eQOwil+WdwsyYx8ygrJsaWBQt59DQDXhZImPpkDdvUDE/xhHfft5RW0TzK6
H3cMfBcpV8mkRMf1wYWFaUzc9e9/zswkWERs7y5Cu3C0Vi/kpFyVTLMmFJQY2QcWoGvD3vZ4sUki
BLiyyrQjxEF0u0v4A3CZpT0WotJWdJAbJEALUNXggYdHacl2fYHDbZSPIOqFC7sjk+oRy42YXeZI
TMG+/xOaHSA5rQjA+jnZ3iOys/eYmUKnYD0Yfe9Q5YeYdErkqKc7HvkOTBxJWJjyqmcE4M3S92eL
sNMG4I6SI4oDq+faorlfghIp+7VA9/l0G5CiVaMUI06ahcj3xtkMDWh+fo5ztN/LRAbj+y9BtKiO
HoOumPmqDXwrfzP+gyI4LwMDCGcFw+dFERf5vnSZ3Btbn5Nguov/XLqix4IJ0QlqGbh8pcV1U3ae
jILuZvSbCCTJN3ycYleFOBCdKUKJ7QvUzFvX2wzxkcxitkyZ0SMWssrrLZ97W8SgLAIXBSwHWy7Q
ZHG0eA+cRmhdIw5p5ra5yCrQz8I03EvRn6kooBdZ1dP/zUek7wUgWwM/ZTZLzbU13VvRDYFEmkkx
U6F+CrguqhSfvILrEjN7ovFXZ3YWmWyWaW/VICGi+Oo6b1zyaQSfJDlmiQl7JO3C8yVp4MJglTiG
HIHC0JGNKaM3SIB5J8AH+BQk52t8WspdQ3BgQIlFabN91hIEzGT2GVLyXgtiAVuKEN3AG/AmUcqH
t0yXPTzn9p8BBoT9DIZO4kzNSQ1kXTUGz1CuGB6NnW9mGqEAOew3JeEZkUvC6yBaDyiZar5U7STU
n1V6WPTahuVQX8d7kluOyTjGrDw2PTYnz4Fb3Y5Ym0EUX9EJptOJvKfTq4nNGirKScbnwFWkdRPw
gkF0cBPYdjkvJIE4tWCHO8ObQTpTeU+N8nKxaQi7XEDZ1KUTNpsUUC7j7rBwESDGxuOUIH6EndCB
DIvkpui13rNVcsdZSSlOx1gpvtTR9koNJZdnCC/v3R5oYMhgnsmnZGSy3hRrVDYAQOu7+UCFH4Qx
3XRpPQSxBS6L58PeTfzasKEzIicdJF2FxSnO3+XCXKhz7VJEjb/rQ9v8VV0n8oAQTmGKPFWgiUZt
DGno1LGSEWgmFI7Si1Tc8up7lfm9TLQMWr6c25mstaPd9A1lOD5/6d1yf7DdmqNnYepHE8Udxyc0
jD8udsYvD6UHPn6PgQ/KETyxhM+GHHuj0R4yg3Ii09AeFRb0GXAfbnqq1mSFXN6CUsuvwiPbsKFG
e2NbHop1h6QhBSRGOR9KlQXFA7zB4DbUOkRYgJb1UxOkGn01XEs1RYwZt7HpTTz2crgEWk+aETo3
eH8yaLIFBadh6vyBYPlT4I2yTOe+vyVuqag9MkzCrqaG0t1FoRSj7mVZEuAiDn0zam/k3vOqpvw6
WIlwNdSLYxfAHpDpA+hHyVT/hNqYyg1qFZlHH319LRbAGez5EroHKO1qynwNWZWlwzykbSsuMI/Y
Xpnyfac+lF4h9Uv9d7sCPld5WYUTXP6Jr7EQVHxHjafqRsO/QomKElkhjh48b/YhXNtLcpsXq5mg
WIwWrnYUuaKf8W34j34tignjjU9+bJjjuZZGP1x9XOeusOAvTr3JbmwYesK3AbhRmi0XWskLkQrY
hKjgWxxuYAQYHBrhBkgKTayEJjbJbjh5v3YBDzGn2PH83yq3p8855Z3MgQyXEjUIQdEjwfnzJA+r
4SPDleAZ+6Hy29a1XGf3KUnRKi5A+1DTjiSbp8KxGe73Jo5lbXOIqom107wu6/A+5Zsm7A6yrmnp
jaYPx+kdv/q+TcoXtS3v7Y1UxnJs15rsja5zkurWBZHvhYBQBOhRiq5ArG5TaaSTYXFDLegyELu0
svFHh0Jcq3PvMYVfVNfFlQ5cnK7RKr0ktslaVphOqcyIuFOgiQRKi6DCbPD8RsR3koRgShCHS/An
bP2AuOUzHn7xC2vYK2C8UdULlYonjbAjjz+gcKPbDyNIt4L2cT7xT0hUAayRs9g1eHwltqKCiseD
ie39JXOU/AmgN/Cy7wAVFgFjVpoj4EJOXKL4VRVtnkEGi9k75zPyUas6HSmZBhlN8HTpdNCXj/Fk
n0IuOACxUKmoLMjhQGsf/a6tEwsuLpkG/97eubsujVBuQAGxBVNVYQezLf6Ph1d77L028GyabRf3
SY1rUnIu4EWkJyYOq9TsPn5QRL4j2HLyDCSxovXutiMEWw5xrnd0LE5NjnW39zCuW3Ge2AaT44n+
d6SxkH4Ss9Rxm0PkpdViNvDRnTrrduLT+wGhiuJqi+V/UGAWtcQVxoNYAiVfH9PEpxd9r8qDU8zX
GSinjTPGQooaQQMAme3VERcSV36oNI7a4usblPJPoiCiEI6TBEAijBqApsXZLOYtY/Y4OCYjAcA8
zOC+LHGRSBvt7D/1jc0qw6rK/vnEDkzLJyXNQFLgLLfYRkKPLRDH0dn3BmDllXHoaoN2L7RkwrdI
pL9xgyvYzNc9bTow1PSSx9z+SdFIQO4dCEzeMuV9PsYATctU7mYN8cR8vK8vRFZiDZbxzuzqPRTf
U9VxRmVqZcXRVkbyTP4/CJuCjfi9SyXxq9LAT0W2tNcbA95+QrZKHAWSZ2hVLQwc874e1jTUsvvt
5Cr457JW/VeDwvOyVGumqh+Khr0Fdp/J05VIoQ+soUSivPJ5bwSzecF/aTASPQrXM/OJRjwx+OXI
z3NODDmdMXbjS/ZeF1LOsEV81+7ePnNXDLoS4/NX9rCH+5zNdl8fQoDr0Yo6D26ZaQxdtGiwiSuo
aMEsj7+czIPKF89G/zmPPrt74dWj2fpVgJnLBYgwL/+y+HYYIWeDSN6TotuLtDeZssQ7Wph5p6eh
6FV1w5bAq0u8gY3WpVmXx+nv3ZwiEa3ZfHD4BPN1PSYV8tNsHjEAi6U+aYoyNDZcKmdFATaVwWwr
7k01eGOAHvUlfPhTczI94qKM0qVSSqF5ItZNJjh4RACGd6tfaxIyfWh5Ztmu+BSpdwN7Rd838/Na
TCRSItGag+VXRSfzRTQoI8kqoAffQ7tkk0Gh1LINMnNtXcZvn14K4VngknTOLf7FfetAroe+jf2Q
DVe9LkPL4WF6kJBAG89TBgnQgl3SEfF53vXZhA5BN+nanIA5pw5Uor3EOCXPVM+YzZ9MEVrjFivu
tBIjMGY/5H/H7eDX3NPcRSDYnyMJ28191gHdmCWSAeXM/SvEPaSJJLcJEQ7jyr1kmFSZPR1dhsY2
qGLh3aLGc/zJc3Y9DHC3gLofEq6f8y6yywwE73V3FmrtxaCFegwhvnCAUr8gXqNmcyqhunYw49dC
3qCzyipkvyRTs2/ciJcLW8pcjkDXNZMr4ViMl71Btnyd4oz9CAXbs4cMmz33mhgo52q9wVoVxE0n
8fAf8kdbBobr71nW4bMdgKwd1+pf6GfN/dzIQieetNBp16V08YMF95wVq7N+yjKmldpMObse9Xs7
XMCl0H1kgVhE6eaVh4yBAhT7OvtQJK6Clh/Z8o2oVDQpUSc0bA2TLB84bFqvkXE9oQLfGmmM8N1m
7mHzgL76dxkqe7exwTH0uyuoc5FxAuuveegM8peAL5qCJDpIqotc/VPXeOJbxP9ItZTjRkvFN5hK
47pF1revnEHLnaaMS5AVUNO1seqiPBx7r5tMsVHupNNJH9aIqWVt++nauUL6VVCXlET88lnsaHOc
4exJb51kYy8T3+Oxo0NqD7XiPxOWrEzkjvdBOTn8F1sL3gBPwyWjKNqqedBwo/2LaErSVZ9/2r3E
FIrx5MvDYVX55g2qwOTsakcySq0SeoEVx8uXtmXODMpjZWB/JW5F0cyJxxU3B7pz7AeIVwQWokNX
DxyPq70sVQMy2MFd/GASwKVwx9eoqYVjL+pPAFtv9tjEKHWe/z1w2Wd/j5V9VjxcjPbklg+P/xkO
ANe1OLOon8TNPXbUHJYIOr5i9pLk9C/+7Hg1zf530TBWd95DecwW+c78Ck7pYanpjsPusYhNF5Nh
Ga2Alr4gAc8iRjLJ7YJaG1eFDTjYI+42q4NsBKB+9yGWuBjAW/bLPvDr7MdD03g1kIn4ElBEkOwx
TgJFmP3qULT6VcIeJJeSsc7f9AJlBCSoN+HFlugNUt1dyOZ4f74umI3u9uH5MO+tvAd6I/kF7vtG
tei9UcxmTzNyO6GzpOvHZwyJPMmDsIqNqrW0nKSrCfXJstM769FYY4EDRJ7m8sDlccsIHDzjTLpQ
jl6tfJb9ElUtio4fv1wviI2HsoVIPJWF0SPaBidrE8PdL3g2pA2w1/r2U23LH50PM+qy1Vsm/22q
Vll5GftwG/ByG/YNagiyAxCfxK+F/UosjZ4C0u1Ld+A0o55QOZw2tjbZlQzjj/FYTHmaM6kWTs/B
0AD7oyz/gp+jKO7v+jPFkj0/BwwzQdcrAZJcMzujJzNO0v6JEpEd9yTjMvH35Zb17e8u4DhSPwzD
LWi68Ss7lvM2Y/jgpVAnnf4TNsyAUsscsoV0zgSYc0eYhjJMwAYbl6UjA/6yWVTIWpRhi0v6VFVf
KPTg1pjKTFeGnDTk8rzONRgTlVJhRAtQJQbVryjbpK4pb9PPlmYkrqGO0p38lXNHcflRalKvP4hu
n9yhxPFk64RrREAnkoL+mXoeOwnwiZXsKlSjH8eO6GWBHUVPviz7tFm7wwqdDynInq+AiqMVLAak
ljeoM9zjTLm+JS7XyHAo2rOG0baxKmBa2FeadhGAZxaLAkW+WSv60d/s5qimUxfKEivGeGde8Z+Z
nuLPS+qf793HIxykdgyDaISvfXnj5yAc+7fADzKa6BoINRUJ1rSmZ9YeMTWIaLFEJLeOuzS4DEVJ
zcaDph8T3Oew+YM40hULbVrvcuJdvLBszru7ehKdY8EOy9kSeHJ3hjmPnIY3yw/5EMOUbCTKW4tO
kay9kqr5Lz7F1/WIsdsfFhbRYFPiJYdeDrr4/RHWB8sBEkeOcQ8brgeqlzqjkC0aIizV1Juxjyuw
q0mslicUIWLOOEQIzYl3i5TIcNC1fflsVjGebo9zIMCqlaH9GvqydoJi5SIbkWpE4w5OERoay3tX
DwxSG7M1CS1NtOIZn1zo4xPtyUOEILMZ43lgfBxkzuO6AGUnW+pmyhcnWFv/sMDIngLBlY3nHaHn
O28ZiR0LL8QtfpYPRuCi09d9VMJoAPUtii930EeDNDFT1om+0Crvk9MfBtuH6RTjr+Q6c4yQuIQE
opSaHgiuMA08rt5cAI/IJtjGmgELeDVNQPINquvyQ8quuFJ0XLkLPvOz7ppgIDLoH5mGoUIfeFUr
ysj6ReJAqRCPY2TArdfmWXH6zicbfkhKp0OFalRHa2HccoVGT2ZHbzs67YTKiTo4ACF4onpUBo67
yxisoixC5FfKAORsYcIMQKs8vCiY9HhMRCOHOdtL59owEOcarCFrahxVV0SPE3p4epWMChnatEy2
TeWs/4Xn9R+dcAZa6F68CgMci08ITxxPjttx7sHuBzl5rLGFptoLJzKScSu0YorW3KdKlvza3YVX
NS6RTWyC6ABQ5YRzklAalAXFIuooAJFwcAZ8hX83RUSikCwTKLhXG7rnHTSB7okO0OJCoK/UbI0i
y+Ea9bWWMA72KlyESctT48DeIqh+ub24pLD6LXTbMF7KXw6gQqzdKALvQdf/LpJEc+UwQQ/PHbma
vnR/WinA6DrrrNErFJsJBqD4AuRC9vHmVCOCQdeRpiJj7SnyRB9UHfKSnTEcZ4lO9e9t3k8bAyAl
o3DjiOe5J4rPh/eBrWgA4f49eGaklLehbzOon1c6MbYSZUfEZXmw4aB3G8T+36nHxyVGYkteZJgI
5IYHZmkqlGn7/kbMV1NFCPAOE5CEW4MuPzzzydGgF+HE9jV4h6i/iytGXogwGJt4Lfj8T36g11/Y
zoTzuCbWxId+UH0FSUa00YBz1va46o4uQoVKy5GNQogezX22Bh/cOb+Teh/PT3UnmoDGYPLD+Gnt
wWsxf3RSQ5E0aC5bymsDCmNqs6SGU7IcsdvSy9ITFa7lCeeDAIjIMaynoaXe4APF6rQhl5yGsc/M
hCehuzLdt4CbwjOeDruP5VNvcmMPvlB5u29iJGXtuX60npDzcMVVDXZ9Pa60vhIAFreIbjRSQTXb
zWxAQZMTa5MDZofzs5vdgJ+/+HDO4kCdwsN/Hirnrt+Os7NaOo27xGqQN82DELH08U7gi0dPWKwy
fBzG0eZ5zL2lYD/2lr6JAlVIzi3Iqxghtz0sRUlRp3zHcFfdi1s9Iu0aaSyKo6htZgdX9YOzucwM
sEmIth8kNIC7v+B6L0OcilYLdmuar94KXk5lzSVmEQBNL9gcfEHzIRJyrRj3UIWFiDsrcbN1fDi8
/zS2YCsBG9SA6YSbYoaPcmfsASuOI/vt0mz2B1are3QqJsx0GN9iaODhnr86rK0sZzqGi9V/KqTY
ql23lGFACFE55oC+5vM7I7vlSK7ZT5TD20BmDVtvux9YLa7WwuIbv9GwaUCgQwZ+uXjeu5Pl0lwK
MRzFu5zre3Mw1sMPne77u4+SdM0o7KbR2BVVoI6RhlnWjAJuzt6UkhvdPpmgccR7apiZAPJ2/LxU
J92ZOL0NYgZxSQeXT1IXpdgjKNyCuNtHEaIcC1iHP//gTrILAsbt31qwzVU9i61sITXlEgQB74N4
zjf69+5GC/sPSaYacMvjwgmbln2t4uBHOk0C/ZyvCvxnD/pb0OWX5ChlqvOfnHY8icYWuVGVJrbm
v2Zn7VPE3iceqRWX8yYICW8NqPxpfzqV53JuJgIu6jboluvK9v+IZCr+imIkEBCbkfuSQ6qAJCBf
y7xbS7evl+cMmDrLFoh+ADTNvBlFqu+4ahX1XrVRZj1WcJrbZCVE5Imtx1/Ax4RSxsUsm0ql60S+
15s5qzfH+Ke6DsfbRZduxAy8R7wuFk0+Di8piqH90dRMVWOzzhqPQZNAPK4h9+4ELez9OgqQJwVa
RFtHQUrRZIGHp37RhWY6Kqz28FpSnQy6eZVt89nDbZgvvWDe6FVC5GWt8/ZVI/O6vkmMExciEJZJ
Nimbde07s6yZWMIUq3Ya3CZ965FmjcSrqWXVh7p4bmdeg+UUovCQg2j3MsJvX1Q5vu27rUlNEXjR
LOsCAh3aEOfPkeFO/DMB2dtNzjkutvSUuwosLhqcquM9FEUd1RPs0wqtjGaIHkydSKp+WU/y1swb
tqpKRAfHMIYA9DkM2sgIZxWSvY63js/gGWLPpSHlrvbUB3EBYlpYZxmHOmjrhORLZ09Sf1L0DBL4
Gy311jp7GMj0nq3SdU/KxlNMMMKcFL3O8Fl1I03cRUJADVae1I+LdoDYRw2W8om9RWu+sQ+AL95t
w7NDh9Hr0pGqDKziIfNQkhsDBmU3kSef4HH0UUrbX2CDye95y2Gp3at3a1RpUrWrLT9LzL+UXzld
7DzvTYy0KToZ6Jefz/LffMk960Vx3qBiiZOzPallz7DR55jkZ/DoHXTUMy3vI7jZaBevf9+S4fBm
dpCe75fb9EwHmOpv7EgsMar0xdAZSPBY0fzsUMFNhHDYJTT+0tWH3KqRz3Anu8nr8NObHl9mNIxm
dXLfEXriU8mx1m8Dz3KoTkCGDtmjGq94v6o3Bf6RdD2U+WnHZ3DAFrU5vO1tU9PJM1hbFndB9brc
GP+GfnP8wgYNoYXvu/7ObaLg7JJ/ZA9miFiWNas4NAs04kX/l+oNfXL+Q5PD1QZ928gyaFNNsTBM
Vs8Q9D2e5FVPTWcGq4fZLf+E+tdx1GQ49byssPkcnBEW0nfkY0xq5aLcB0GjuyMTQ1j8c9YrGCK8
vwFQ+12GIdrKL4CLxmEg9w7YiV2yWxZF/708+xpj5/2niSmXU5Epk6iF7wkLZIULCsHGq7Poo5om
WH4upSBGJfXJg2/ocSjmIJV3N0bijKY2p8tv1uWbMysG6FnCprlz0Oof4KuroSatl/Bb5zu3sjfX
m/s447bnmyW0i0OMRGzgsbztcerYHHTHWxUlE8VnrbuTj2JBD0QZRLUnIz7Ugsal7alTtm4BYAVT
JnPYZLIrOtZ1HWQiTEu17AkXjoZX5Neqq98eMIDcf8T3ch86pgy8eQzMmg9JmpjeLsgP7/OVQOxr
d0YA7CgUAKiRDgx9XuOMc6sVO7orK2WTH7sVvDn0r9/7SjbsnYTZSz+VDK5vV72KkdQ5AuZwKQ0g
yZdzgFmkSq58pCSH2gV2K5zASnzAuC6NMog4ac57ObyfFwsLPK2KgtYLDeba1B7s4h8s5v4eDW0h
UosG+XZa08Bu9Pu4aI30i4ZUq7/GtGkU33boWBwKIf72kDJDm73CWwaRdessawKGkW218X12FOGR
g2qJYfF65y60Vvexxcom078zX221uUbxOJyOkKD31yVA9XFQhGZx1FlymxRPYZzuHH5BEvGpoq9m
vdDXF+wGfnz54FWurYq4+h5XToBcvkCgb6i6yAXLE+xkIkgRoVhXhA6MdOhXbIE1QoN6E/p3UwC9
epbjqR/Lj94Z6C9x4C6RzKe609NcKt8cstuQsxEMh9aicIXej/k6KX4QgdqI5IZp8wgRYzh1pdsn
41jVAusrcDzt5gpft6O2PCM+PardmgmjLj7zXWcx64RDw6RQgWeLyfuxaTe6x8mO3Dcls0E3qBnD
vmjpefa2aNR+mpSF4BdjocCXwsF7Zun6aCCpQItTftBXDZ3RUr41t1jEgOumjy+aqugYfE5qe0FH
rzgbQm4zn8/RyTbt8EOxniaq/2vWymh4VtHUyDsQ4v6P96M7y68w6Z6YaQDOHN9I62uWwLFBv9uC
jbUPat2HZN/k8jQH3N+8JiLg2aXZ3c9M6PQPXkgGfm0jBsi+vXLzahITn6F18cjrz2PATCl8YSAa
g/sxyIViubG2TMCRCqrdiDZWtGLNCJlTSKqVC2QmHlB6lieKsX0XODXtLFJG8IsIBLGDcW/nvCST
rljEtC1wk3gsyZkc+qmeQwZciNeLsxI61Ch365r1JTIKKPyHh+qf2tu3a10xfC2utncgFexXP9OS
GYxq86ZpJGrwGM2kQOE9qxZfJE4NLxKpyPjvoldhJXeZxK9jOQjM2uXgZbsfi99fHmjVJ6g31eXJ
JaDNknFV+Uko6qVhLprVD15izW0M6oqjlHQn2tID3hZzRZk7LsqKgQKN2pv5usKS2TfUmSC6opZt
SYkd5ZyM6TP/Ohk8SyEFKV6gkq6n9RaH5i9DvRBFpsjGkNxTFCLR8ruckNB6P4KU7lRotX/mqdpi
LtfNmv1NDvTDgxej2AwA18jUREKvPRlZAE/S/whDRqJyZ3GtjCoEnYyR5vM58VPQghxMV9Sec7co
ZgGdlJRNcyWaG/tAqoMIZ/yp8erUh0XeENc5FCYNImyRSan8G5AmcZpZ5wr4V1LirU0ZqPEDeH5C
TYUS13z3M4uLLKcBbV1KeJdhbQGJzXqjKRJx0/RM18Opbwpazn9Gcn5Bpaw+HI1z/k8eMyyc1dKp
ENLjINLlmBI4HY+2QAXHlPiXypzb3gwtjZN33qzc7QRZWgmsGu3UVJFFOLlcCx7t/nv0fOWQQLfW
C7hIHFluddaRJOu6Jtj7IfVh2/vv+UBlw1sXEIHLmfEAmV2OrVe3rOPRmvfu6aPN3GhrcGa/34U/
aHvjvMPwizisiD1gG/pU89EyOWUzf9/FHIkxm7ulCj82xa8WAoA1sUFfLvtP7rSv8Q8B3ZAyhbOk
yeIP4haMYrds6MVvjMsHOzYJfD2dm8bEHRq8qOBTMFSm7h/trf1kFUDGxL4FwkxKegNTkQqX08Zv
+UH2JE/gapSR/WC50TGJpt7Rkas7JUpwXtIpjVymyc+3rLgPcnTvyXPmXWhYPAV0a/ke0d0npky/
Ju5z6XWRQrArn+eyzxTCbqQJfpWD9Ja/QXeAi+yNtdo2plpf80qAgnj5Iwkr/QXtkoia/6Hz5GuN
LgovXOABpAJeyw2WzmHOmjbIjLt2j0lgoy0I2+0I+EdRjuR775Q/u4T02qKiKibO/JBRr0ltEtEU
JUyz18tAreJIVBfDoDQKFOU7Ov9cYYyoq5fYHMhQQ7HCLxo8+qEKz89tFMozXylA8QXXeZvcoTY1
nujj3GZwDYvzOWFDr4SLvrKXeT26zbY2QEyvNKnpBjJ9Xr5+4UF95BdYDLxK+wt5fcKOPmz9v3rn
e0Zpv2paBvgW8RZFnFwr2JFALN7u2g0P+wVMzr1j6MMQBOzlY3hiyDDg6mNZyxPoGu69M9hyR7tF
7zTwa7xK8VJ/YCMpFJfsRyLPocHwFnveXlXuHsayIZbSR82+ki5BDuyEdHQvgwHQ8EZWGXR9GYlv
2teNqy0TTWVtN89GmZ9rct5xIJfDfmhtqGW3rLfzrENzcLswYDNXuULLWDfFnyqi/tXk3NgMIvwW
f7jBwy4aOj4GabO0lWMXCg3RlaqmvsUsU3yNMh5XPB7e9/1QD29p/BaC2I2sybRpV1n8RMAcRqLE
AYQxe+h5xmR/3wVFPPZmPUqgEzq0lYh6wiwSmCsY6nevUlTTJv4wRbSyK3tNutpasOHGH4wged1x
7OTN6lqeJbPsLoCPG5Xm8+KR+GK5WPUaCw9DdpLPRZ187nKOQ5dH2JQOhfNmkZ0C9XZuUU42JRdm
EvJfbzhbI2zP7F/HbWnQL8lsfeeuVhe80xEcFsOxn+QAHVI7JiAlJlCTDv1G4+yDqGW3rXZg42EZ
lI50x/IVw3LS9s4akpJq4fsm5rODr/HV1fbY7sCG1JiH+jydExekchkB3auAxmrgZC8gYoJiu1xs
ICvds82CvjNOVO7nyyGJd/4CCE0/Rxp4Gy5LAWszS4wzH9EerH13Io3Hbb773VqH0c40Nid4DPHi
xeX4dA0npU7gTRtDp8E+VcF24ydIO3jOF4sSSzu6BYeVdHubIjKz+WTgx+j8+iQjxdH6yrkn7blm
NQfOEbqIyNVoGgWO/GEUp7rhRttjeaci2IDBDMLTyOxg8190RnryHGVTT50s0sihnRc0w6WVDoFH
5XC124eO68KJAWS/YxSQCsTEpED1G5JzFE+SkwxOFIE3ZyFkGRPUHREn3zjPZX0Z2RkahcLl5efI
+Mj63Lri/Pu8voXxCEoZUuDvMnuZMD8g3Mukb/vOMk9ISmOQSQb87kmFk8noKU9qjbMPayggvEgr
2NGIcOOAyHNX/NCGKpum4+BqCWCbhwkb5CWWSdLImc4hkTE0yoLV0SPbkdebnKC57YX6P33Fxt/z
7aQxJ2xv/7SU1wHEqMsX0OimZ9eyNN3+n/soEJo9SIwIkSPM9htIsYvFg4CIj2nJiNW7yZIVMQof
kCrAFZn/CuISm81NoS9HFoz6o0TNVnnns2IyHK0k8q3pqbctPfToS0Y472yWZYe3f7C+HVTpurMo
9bQP/sn7KhGDtIVkstVYV28VwTpGwlBcN7RDc+rWLvrPykZV46czKy7TAbQOgmVjWFtPbUQlvCqx
JubLR9sJVpgriY76VIIo19kc0gA3HSDZaUiJbSR36XvzMb4x7dlhBGxinwFGHlBSWl1gb9rH3iVp
xJSrr2M66iFFj0qKzHO38rjfCedckQJ1n6f5rrVXNENXBFNwfzQq7PDGj0TVKBtH3FjOxam1ILgA
tDnBdoTjnqydfU8HecrYMGLHCXEJtOqtj06zy2lxD8lIclx9pjUzqX9U0i9hMt+vyRmowO45j1Fr
mRC+K1xX+LGCGfp3c8LvfZ3ncJUjoQjtqDmoe5Khnh7EN6D4AhH9WUsB6kT1QIGf9hrbWRf7gvBl
ffOU09saLgkURVWB1PUVSyFXdXxDa2D29zjOgA4a2zcZMDdbJrL77CRHoKkeS/6Op6hnDiRLLf8r
npO8aArlZakIIurSG424eet7kPaJBvDUbgm19w2+Km5OWGY9GNPvvn81J37dQrCybZO/zQm8/KzH
CO4wqdyYi3V6F5Ip1xx8dAzjmZBLdxuT7CY1XJPk5PkUyI415pD/F3VauT/yaZCbxWs4yDG+2bkq
kZLOtW15TerrNJCHRnDwpTMjH6ZT/jtqrzRwCxPWZBVqY542KDrErEj+0hypuw0VURRDn/2rQmru
Eu1RpWyLFM7Doo4e5ZUzSAT6MUq+nEhOR1KOfhdwNJxjA62FmaZH7NZo7P8tYwvzxrWtb6wPkW4v
y7CdgoS85XWzmoTAVYzqHvU7NibccUzJD3bC9uQ0lrBn7rdyBgjg0W38V7ygRHLuFOpbRp0SMtgH
Wwo489kb3RjsIipomIycMC8yB4AjqdntuOQgGA4/BDrdg7Yin9RHzqp04wiLFkE57B0uKqrzyvsc
DRT/kH/FwCR+GCTQlDB1MAm6xaAov60Qdwga8B3SD95Ol3JE3DVheJp1xP29C62YHgmDgcQV+UIQ
zfJiXZU/DwuEhx/OxwzJHjguoH09xtNgu++5SBDOu9WMnVhipAeTmSw+TnTpez73cVi+iz1E7UiQ
9gRyZhLUNJTrE3yYVdzYtpBvcoG+H51myDS6AP6k+TQJStKuRlEee/M8Jxk6WW/7lrzMS5DnOAT5
GaSKzuc6lnpz0UOT0X2gilhQQsY7M6TqrC1//urfEdaw1IuHtzyRyZnFfnUmQyMb4HOdRIfQRsKH
/kflyLbQQSfTxa31vDl8OrQKwKsI1WhCMoOAI3qUAoioA9w+It44lY2WsjQoxRbgkFzexSE+5O9u
+TjHxOUfGJ/pDLb6U1VJ2kPRSRpGXLiKJP8VNC5YSxBknnbtrMybBrUUn97mWp6h1xtmbXk0C+Pi
TeRhCtajgok9uV00exYn7rZ/QLc9wtbGK6lP+PdYoUHRIEr7cFk3caaPfuO+1xLC0yA+/Pshqj33
vtXoCA6ZNIMZGwnxsAYCVUWf/7j/5ZnU+9OST02pvmEI6VL/k2VePTYbZkwcFm0O9XE0upUr21dk
ACG4lSpKrJ+I/vLz3A3zZLl4RBMYC7guJwaAba6XlrQAr0weR8Lw01sTwIDITg6jAe5qRZw3kvDC
bb2DPiStOAn+5zcFRIyOUCgV1PplWfDEiPDcwmK5UPIfq+SkjN545s/tg+OxnAUIlpFed00soS7a
74IIBMzFdHLvWDxaV7RCtKMc98zRBaE44PNioB6rzEctzNQTsKWkw8+kc/5MYtAf5ZLj7Uc9KtuM
QZtmWU6Am6wOfKVhATh4d1mKgDvIuch53oGAKJ7nOBPdnGzQrSEsPuH0/+shFLB7Qy07eQfSn+O/
h0MLvPxdfCmmPsEWgNlOdlcHnIDD5XtYsKxSK5aA3tZ4loPXUCS0saKBsx7r/Zurti3GIf+RX7a/
l5pYqcSnE2kItkVjYStwUAQFVwOKktf1OhW890hciOtBO3ksAzeo0rmepP8ras4VmAUzhfeaUm6u
FT2R4vUiLaeC2X7e0z7FyKEGdfvYuYp5UkRPTsf9l4yJ6++3cp+cinlTFk9X/22ZAWr8wGaedbQC
qoO72kA44cAO+IWEtZP4VXHwc8K/SU2zIHZt+bMzs/gL3sGfv54n89RFDjEOskmjH9np976onCQC
o90XeemYy3eLw333Beun5WHOtH7TMRD7pyGRKRQdhNErg5G/O4DDUIkSns9dyqPQrxNTNsyM0mMI
fisurDNL0PEHpqyrjn5MYqORP4lOQ07Htcaobjh/05PI0Dn01JN/iQrwMxDUuz/BcWeQ+C+U8tPI
bcYJRyfvtvFj1QnFXpdZErrzeVwJI9+Hw5WkF0Jj4VHHt+BnqZwDP/uraVK7YMAcsXhIuNFXdzLw
jcaIpizUrV0hqyuyeOKd2r7Nph63ZTr0RzEl8TRuw30sc1uJePZaBnqj7FKXy7M9P5NP5q6JWoR2
+q29Jr8dx/dONTSM2aTt/vQgMBpxKdb0yja2/zI1ujxWW+6ib+k95COTSh82RRE8A+I+zRCEioPh
3FdkHKT5gohZP0Q4zx+yLMwNkIEERcwiRkYkN0J9dn+vj1e84/1vgharm4A/e6lBZcbRpjtA63xX
O8osDJi66kDLPiw6O0uPoNBOZIiaEymZRKxrBCcQieq10CouHVLa15PIxmlwAxtKkIjhkSPp8Eja
RMdoa0EeFfepj7NKCMT1y4e+u4t3O1YD2NqEhvfy4fWhd3/0uL7G6L2bKWRuHE3ac1bfS7xnHlKa
HXFrsDz+VJWlpSn9mW0cDnpJZpczpz0fs4K4F+YYk0Wkg/7Friwn3ODvH0BoDd5t23uB4WMbI4QD
gExvmtk+ZYhghMrsRRGQN5DXic39EUOLoQAEhe4yPnK4+4d7vK8jdaNvFd1r62t7Sq0uBm5y1ytp
0YKVCRECq5iBXwCAcaGsL3nX5ZjtbNj8BSg+5XXq9tV6jOQKhYZKhxD0Mh43B2eiSkDLFdihU+6e
FeKyLITg+RTdDzqAgWpzNeJVOo4H1jD/jnW83m+zdk4TUaCtCPbFQox+yKd7Mt/EcSHIuDd9twcu
9EpTR6TZ0DlLfKpjMCQyEKlTMc1GxpouxSg36W8tTCkr24c0rCF0kgcS39LELJO9cDa0fp3EX31r
Z7Wy4bx92hG1lYtRt+KQDW496pX0ohY6Z1Nu2Ccbfp2857nP6dgcnaUwObrA8mTtmrCNEHU7/WRR
8rajsXzvgmZAMLK4PAYbaBRsQE3TVS5RHoDqhGUz/H7YTYG6uYrleGPW6b9BjRqdrvG8SEqgUpFb
R97GSze+6wS+8Z82Ax7OteysuTENKUIXfcfwVuU4mdWXF2votLes90SFb9HnOPR4LFK9vCUU0oKa
AZCXZ1by9l5hQOJ0kxlP12Q1gupuaP/AtCWDd9thKkcNs8vF/4/KGhFndQCK+hPdOgxcNXjAajew
5LIHhuqgiwyVFer2yYXYeE84vgfp3bqgyHmBngUWgktanYXt0uXnjePahfcH4XGfhnZdAosEewur
vhQ3A7sE+nk+H3hMJjFxxKldfjuJf39YpkS27N8TtSfG44dJbgn+ka688SXggRFbyaCClIQI3JqA
P+g1WilFl0i0G1Bec5gQD75TEyIOtJE6UDxYJVcTEPqgzxzV/HHiljz3UZczW8nKCxht9YvI7vmL
scbCt+FA2vNRMu3Oegpq+PpmBaO00pEl9JqXXQ5H/Zsi86nSWkSyehTaHL9O20sUT6HYrDf9afVU
n5k0GEUyiaILHtALSbUgvZL4XqpZbOScOifsI3ZQuTZIhuvRTrdRRNokeaQqDn+smhg+bcWX3DzM
xHthzEOgECpcQ1dTKrOZgq05JiLfWGnonXPm62PaqYxGEsaEgINjVeqj53ot9lSQvtbkweL7rcli
9NJgMTsw6ZtzxjZwpcB2xFL53cIXFchF78NOEfwEEWMbrdakb8yMIFRCd/USnzk4eBdtEwjej6lk
67MnuEiD4sewAPz3A8tRdNcbU47ai0iSb6TjzOQpIbr+/Ga2R/6bcoZRN1pyzcYjjsFBEXVXJMLe
Z3DK6noFIqsZMPsPHCzWQG1dxosjaM0E7syYc+fG4dj5wvonRsgGhG2iAmaEzPliPnN0hwdCQfFj
K6IAtASC5DJKe12MJKBWda1LHSV+QuMrrQd4JJ0spa3tD9Tf0LcTKnmOdOXvvzC45aT393vzY44H
wv/v/VodNy1B6DPvxwVo/Yld3vfiz0b459iZNT4WjCyImZImIVrbKDeuuvOIZ/0htwnr896AnthZ
cg4OUjbOOIwwRjU3lqJLnpKHatUeS4hZB2U7MfyOKaSKkToMzh8VBvdQvZgjALIgsg0B2Z9u2VCd
SM6I2AO2pG9zqBylAYgowhM1FFaqT/+nR1VUcmXG/2DZ9auAFIXSMEzG0Vp7K4k46qX88IH4Lq5S
xBqUhrspypxSeiCUCeLQvcx6TiIm10LOBguEfjV8Le+7osuJ0tr5pJeCsEuhUeVjwOjbdIvwWKtg
xFCTepnJOKD2RXPiZEbmXxFwHO5M5DN4lRwKgX/N99iu9nmCtWaj1VQot+jSKwgj/1nxESpTkqDP
mKMAEpduhxb6N8JbvqgxzxlJvemf9i2cSjb7RP8vsjnmAy0LsDPA+jJiwFxQ94IU/1InyjYKj2yW
52CFEiN8X+7CFR0eveXFrdjsEhLJP1QxbCqfFJ/h5cJbBwI3oiXuT7atyDjB5QhoxBTEFcXT9Glr
LAaN8VmThaj0kiawJIqVgUoMwVooshu21L9FQA4BJTHp9eArqAD1cRvEQWNgco+zRU3VQspIHytP
BzH1fNc0anUASkUt7/MTo/BMj+PzrZdTIraZb9q27DpnHXpvf0Tbw+x2fJE5qyz9aiD1/E8cuBtz
1pGgE4nZJkcbhH2PIzsjQ+3YPxTuulI+gqYHGAA6fd6WuIcjiRcoDHo39tw2beIffd9BRdBKGukO
T8VcdOeaDmFD4J3klvHnO4UnRe7303L05O3HFmGJjpzaSZUcEp0aUVukFQZ8SKeQAD9ggClBGCKI
WLfMBmOuDifPQ9yDHKMPO/OSqbTNuESxayFMl0A2P7Go0JK4ROD2LemZ5J/Pqd9nJkGjXtzqU0nI
MLiTAWdCNOhlnp48QJ5yh3PYjRh7UK8cK23vsSHKBbLi3FWe/M/bHBSfY26wfZDMOZV8gruHtbQp
KCKTqH9VxhF6vgtn8nD6fV/iopwjS1jEHB1sYvdAixet1EBvmRCzdbjHNd30MSSqop+F5VQkFb1L
d354HOWkbNGyNiyzOc62vT4mFfTonVKFkTyE96liyzT7/ih7uZTFJK7LnQZj0wVVbcTKNJzHO9Qx
oNilBnRJudn6mWbV0hCsIQFSOwOARTOjqtt0WBss4ng4nVNdCJwjM2dpzfzqiDQery0t+OYuYSle
fmYPXh3NsS8miS1ztjP7XErYgsX/RIOI3m9ZtHhZ7TbIwsyaJx1d7B9IqcB4BYSzvmBpdefbx7W0
QACuM/91jHzB2vBTGclQ655c2ZS1+TpCKJgHHVP/3noX6QYvgQs1+uEWkesHVZup9swK1YwwIwo2
xojXwCAjeVELhRJPt2CB5mtjR7GeeKTyITwdF8xFmvplPfj4YjSVTqaSxklEtJK8bwvG2lpi3oVq
JxaOkxjdni0syK8+mbZ5BCXYrkWSaPsAu9zGLfs3+z1UF2YxdGak05W2vHQCAR7tMitKaIgM2KMT
4m6vn9c6hm4nRVlW3apM8O8jWb23IcDoV93l1RecSP8+g0MKfoJmVLt3D4Fj1YEp1BVtfbiWfQl6
XWwgZdfygM5tIpB61i22Fq+eVPwzbxAhbbhE4F2eNv8w39d84Ofn9bwwIR/dnmW7zoV1DfqsLxVm
QLTQWb67cdvT/Fzq06Ychn1mt9r4SaoQl5PxaoS4vAdcI4xEp2vYGKkiGGDmMh5c4cBp1hZKKmem
AE2T03Y/3bkVSGvt2tMFY+OxklU4DF964mBX2230LCR/+nEoyogonx+qX8HLThZV8jy6jblsqfpt
a8jhZHW3OEjl9CVpoak4iImu4Xd46CM60bYvpkzvW2ub5hVQz4qm1QhlgMRaLOqz9ODYk4E0rC4c
bI8OM3Pxz4+yNXZglypHUtJJ4bLOupQ8GwzMvcOqPaOyjxtUTAoDjjF8lrpP8zUXBfCEl4RClDt/
ajmjYwevDie7bEnIJE0O8YMUn4bsnfpLoC4dG6HrW1O8sOiFiRO3AAg74+XbzglKmEq7MeCnZ6Hh
6O/BQ8leJLEX6Vp5nK+c5lgJ3FhQk1FXJPICSS2LwBKwHg4LpA2oD12iqYj+2KyEkQzs5GTIr1bs
bl9o1sUlRpnRP7DQ0EKiQanTQYcTkIPUhiqFiiVAl9jMo2IXS0wF1IeudLd3e6xRmn+NpuRqInUH
+K+ybuMOA1ZqT3DLr1XjImJ+LPnCEnhyk9UdGV3oETgqS+7oJ6fXHwmY0J09IXn94bngAdbo8TZL
WxZZv4AMS2xrpyXhkzPUndTKEPIsLcTAvFvUPvKUxMPJYLZq0q8YpdjuiW66DGiFA9B805wqwxaB
Uix02P3Tq7xKnT/+e0MB0BHmjQe0P+x0aGSxgD9RZowHmgLhIpMqmb6TByHd5HerM2ZT/23sH+K9
A60Yv4jHKOQzprwFuHet96JoZ+wRR0hOlNBtYGoYpxJbuG9uReKfp1WPIFjzll6F5o5NHVtnQIUE
XsNkBO1f01zmpHlX++cwNvp1Yw5YZxabrxsN5t54y5hBIl8eWqFXX5+U0Snbgwt2dNRIzjqtZtOD
r6NpUYVZj9cPNWckFKnPlQGWMLHidSibNUt+flapJ74DpCmceyiEEWUi9r3g2+H8V2DgBBtodDiV
7ab1gFMxf3j0t8NuJsSgJMX642zrRK8Q1hlAHO862+OHxqt3m35U2ASqE6tcazHmkzk/PErLWxpA
NgtL/194THdmn+nI79vssbrW7pNqtULfQdTIUYZlec6BlwL0ghnGaW+oIPN1jpvOicmmHOy64OXs
WzgK29imQJWQJbQrFORJ0A8STNKKK91YF0SzQ8fE29Nl9mXufpTTRxAnpPpmNXaX01h7O6gRhhs6
xya8Q0mB3k1VmOu1Lb663zSjupX9km0eLt64TtJ9YJtks13hJa9UGwMrs56/DNQw7uUZLu1mwlA3
zZDVicGaurWY3F90lQfyfENK141l2CB+csopRAibVlKdQYuIJ/VlMzVzXm+7hAjktsPt1FO4v+UX
DjPc0fPpzNxCzGr/a5YAEi9w6YJ4KkQg7jYqrkFtMQuaQSftbGOjSJqVh0FbEQxr+KxchC8+ZeKC
GEK2hpsI87ysEtJSVUHXQOJqwTDdoyr/wrK8/39k5x04RTRFy3hXwYE5ETfjuGLGUmYgSLW5QgVZ
Bkg2HwQFzEjdONu8o6xgI+f9W7ynTNyqRVHeMKJKEyG7o5huT1o8BOG+lhQOyUMnGZk0sgIESX/e
7s/QaZyghhV+rXiDKWoo7chSj1KWjLlEJmutTCpcvlsUUTBJBRwmGaQZ7PLsOBZezo7IQ1Uk5EGK
kNGeiOyviBjdaK9dE3uTyuY+kgIm+EU4I++x2igvJqLwzi4YrQLgrYE3fL3+JfbdnP2tbpONQH8E
Vk0wSQhyjJv0AjiidF7YWGtkEyvKT5AteAIdB5zU4/oJqpki0KghVD8P+I1bOqapQoEXHb4JSGvT
Y8mqGwikfVveQT0o+1lFy1OBwr3GPEBFVLUlhtFJaGLzpYhM/9J0Gse1UfoGo/buzMAqos3eJ0es
dfXFXKE6AcoXF1pJWuGqgfh1TBlMpo01L3uQUfFMozb8P2po2Nc80DQAkB7d7/uPEO5fDZ5S4HE+
lfSO1FbfxizzKlFJqbrVDewD6NDBx+bk0NbFPuv6ex00G4YsdU5g7ENI/OT3zrUryN5i/zhQstgS
LgXTE+9y8LrzZEGI7y1uf2J3z79zDb8AAg+uIwMEUbO6GIGYDJuyPWEAZk8RpkSaJsVNLaE7hsR2
NEvuCNvR/VQiICAQzo/3OiDEL7z6V7h7Vy1a/rbpRH0Gv6UUHXEl/USQDB3RQMYPD9YHgjnmwyKB
ye4Kk5rr333AFfj41Wep8LbW8B2/jJz/UHpgjpu8S3EzymZ1ucRjrWmTSyZnVLoYQ+f0eZqsqs3t
XOefurk2fLr+hltyQMHaYmwDh15xWCh3m1jZ6QEW+4rBs28QXCC3qU68wbrEy6AOZ4ud8HINfeG0
5aqW0K/uEl7gORLiI1EztOcKkkEYCF3jbNN+jCZjSP7Yhm9H6FraY62URWDo9GMDRlOySXwfiSQk
i7EnbV+HgebZslO5Bo757tj+Ck8pxuPluqRpvYaPe5wAp204Hg8ndDbxoczXJRbDv7ril4tuXdaI
KaH/fYjHxERgFKuj5f442A6oQ1+ixbFNF1Yx8Q6LIqtvLZbvZsoV3b6y3a7pJQHjux9kv949wWzU
UMkDJ14PST3eb7FjyFl834BKpgeYR/JqdU5D/rNAnQdj5zr/M0QP1XwpTnbHiQ/BZzFOaixW0aU0
JB1hqrBK9bqxPo29PFUicBoupuTmxBAUwDefYDhPozI8cpPvtjNWhaiMETbfZ7x9YlZWQNk6aImO
DYB1QDq3Yt2Qi/fTNPnxkwmiu5e3rWR0T0l6W//K2+p+fy12vGIO8YIfDhOcS3qNpLhuSr9YMJt8
tclzxZxH8TTNreoSMpDsCgvA9Ul+o0u0+k7axCirKK1ZT6XqOtr9b6rDHdswHWXBsT40nLKrAf61
RvB27+tDCOsG9r+GHXBpQD8mzrC6s4qv8oYbIdkx2jV1cah+TNscGhwe3ojwVGIMeNa/TPCVkkdP
bVi2DuLQfm7zPSKm6LaTeMrdkdAALFR2Ji/S0nfkXY/LZOB636uwG9ga3JiyQCo6+2mUTgodCZDM
f7A0jINAaS+SYxbF9GzmmhAmCbvizqKZ1Ca38Ls7q+xCSUp5C6bjYjEICYZXlfmefvVJ7YZvRR5j
tecYYSYnctWMD+WnXe4Q4BR4kuGmoAWC9e9X1QllFAc/dZeHrAVnRkxiYN6jCs1NQ/Lf7bifCokg
rpt1ari5IrbQ7F8V7OagAKAez7qQo5qdSruaXlgO/DoF0QzdrLmdS9Ski8kMmLyoEgnq58Ozez0F
MqKfc6enDbgOmeGGpE4mUPbSgAsiOXgQF4JHIBjwN8tugPGh5KB4iSijxWhyoWoZz/W9CVcjKwJP
3KJvJVsKW8C4V+tGWJpQ5/i5zMIIYC7LkPSOMlMK47Q7jNjUqotxlzV+fUoIbJxOVSiEBUu7ECRi
sjk0ukdjfbXT4KXowuvP5AFouicDjLspCs5XYsdhBSyzel3FSKtnlfI+9ZcVB7X7oHIfkQJRmU4j
j5gCgjVjp0a/uOqlHN8PzwApkQ9UeIb7kZ6ALj+tuS08/YXjsR8sHtZ9qfVKay3RVthrN4Xrhq1R
O6b2AkXBC/hJFbeSJV1bLZjC0ss91ZXqjnDchrxE+tVyb8O108VVbvU6DeO3YIlp9EASZU1N51X/
MaBJi5h+S++VCVM7RvjHdh2Ny2KfPstz7TMPUnSPD5TYlt0RKbF7IWTZO2I3ps/SMVPeCwWi1qZn
7suG3AHPVTKUcQeoPSlgmg9SFGlUybFWjqCz/yzqcLv6q+YOBqGbg70mTI6nST4fxqlbN/5an9r5
7s5SIeeah2hMaN6H4gxhz7y0tw/pRJZ43gf3Y2S2fcsodCEplR+mRajWoX21mfkUoUYzQIvYe/Xm
x1HQ6hzZ17F//FW1jS8Ixf0jCTYsewmPc4CBcVM+7RRDcvndfR/qkgnOVNJoRfgh8nws3mVa846c
b62MwovpqcJst2pb6ASBvkCCxkeKpK/6nuYa0upVUumI5f/qqEZGGKsUsKDHAhd7WY5y8amrKe5X
rUfWylQl5kf0csrYZ7dohygnxE/TyEsgDH+aWjcJEKKlnyaVfyIwqu0zZIhF0ARZo4pPSdLDDWFo
qzj7govfCZim3ODmwDDuyWZrMfwxrujNV9fGA3i2ZVsiuBWdlnJMWeYCxHERH3b/2wtd52LGRg/T
Q6n/glfaHABQHP3e/Ktp/6sBCUgv18cjdOA2DqOo9J1CD7bRL6Mh23VuU77EaLWUX6Rfqs8UZmRn
KEEFN4/Tk96XPc/ZM4DWKnNEkBbh5XQoGcBS0Zh4kiuwUgxJIw4zLHw/CB2kWjzJ9aUaHm/tdLDx
ziCYMx4Whqn27Xat2eaGvBXbd/QtsW8YZQInpQ0Jtxp0NoU65P/1mrjn09s13xNpW8Gwd7BzGq7y
KnSR++pv/jhEHUHL0w36lPVF1TQawKNBZehOUaXluPZ7OexmNEKI8X+SnkINfnOanSMwQ3b3ZkkH
Oig+0KPy8Cj6ugY6OJmKVR+k+FlWmRKmcYG+gRNwZbt1WnCypEL9LAUWe2efL/hCM2W/wYIx5KVX
M6xNnHicTZnPIrquA9qzGwd25O6yxQ/o2Cyok3+0Y6T9+cX3QbEvo2BL/IsakmeK2f6TRKwI0JYb
0EQumYU5CfZwzp6g9tNIBh7ht8pGDurlqqrm230gefQWbsNTjqspH4d8B6nDdbA6r278ugF3pBsb
KuqweJqOJadUavZPmY686SwknPtWHQg2HDWA1FsP5cX4L407FnBbtQ9wLrnbHFWJNyKLfm6Iac57
pNYzqxIcDVM3Zov5wTH5tKBPd8B00Sj71iyAsjr0J86Do3dC/SXL2LBTuByCJKplJAi8BuBpN26N
rFIw0l3Uuz/49Ll075e873iMSZ4Em+VSkGxeUFy6YBlhzkodKHMqxy5JrkveyFLjNfGxVHLUObcT
Qsj6UeqbIMVCY8GSDoUruiRziUf7fL8emkg3nsWjmGk6q8PRdrJzmwNNpoTeiomplo5r0M4885p0
W22dlKv6XytvrXo5kiHpAtbP5/QmkLC7lE0aEsVgAPe6258IOgusaWWu/7nHFohmshgycoHYb2ba
scKz674YZSGqttAHjmPBhDVLQ0UyaQviKwx5KvrWgz93L9aAfPkrMPd+siibY82psL2XPG3WT6o8
YkuFdRAozHxjLu2kg8+cnVpAlPqtyN18PF4ghIrzjxM4wZfiwrW625DWOQoAVAZ4wI0/h8ZtoEqE
avQKE+LEHKlq20XrhQGWwiEFfjwDkyQ7flkuMIVug0I97lLVSxK0QZdzvGq0LzEYLSSQgiKRQ1oF
rTMSEZ5qesAfY312L5xS99OAZPXRxgJv13v9vUcQk877SXVF4MmHCrK4lyfRPXhtLdhWrDGc05k/
lQh+0QiPYkR7c7f2E9NeR7bOrA2U1kzrRkllydPn2L+vP68ktXldqgzNktl1+XHUlDF4m0CPmgc4
6n968ayhMfJo3wHyUwxtpQkzUz0qW3G24UlInirtgpWC+p0yWX7qjAcGChA0slm4KkXgR46eQ8Cy
E2PzQhPYgaLN3WnsVHn7LUWI/DQC1QfU+SmcsSlKtrv5b0LS9JKK8mcWmmko3LUUkxOpKvm9buZZ
+f6FxMHr2OM5Gy+UxzHksFCUYfci0F7CtESJRC0fLETzpl8/tIDk+D/+vFZ2maF7bxysm4vUHb9W
5yG/hGmouGYzN/gFfvE6ClzjvbRcpntsVEkiPcMp0KaZIlIfif69xn7HIpqqzWtzvp8qcY12I53E
mgeOivkNphACokGYjfnpO10IBVzM60ac/d4e3RgUKZ/8dSVHbfdNDnIYSZGiAAla9wUYyqOpmUlQ
73+6kKF+xj9dCm+83IJy6p2VRFtTbNPNazDfuX+rB8wVqkAoIwbzTjuN82TsfUbQkBm0phjCH9oL
HbftXzdNMPN3mIEz3Xysos/WXLBDRJ/ShJrJO5dLpKufGB8B6RJlzpvOKohiVukfY/iZov7O1KHe
6fl+nF1H+BqZ8Is0pcdxWbHrVVS7y39PLjt1POG48Ezu5ClOTpIEQ3tZIR+nhSnQHzxRbTGct0ly
M+godhIIs23AYNhY8W2ujuHSl1j3FQjZxSoFI1BS0drEx/7RjrPDRyvveMACv3aN2rrigd77UnE5
SEsJ4igJ28OYt6LR7n1UwHijA4PdEVgzWGfDdF/UuyeSbuqP7y7ApWOfaLjSMyKuZER9tizI29v9
+Mik8h/Rnh5+LxpfKEsgDoHbifK08NZFCReyVmPYpxUbiYm2ZB0WcF95Mx0MGRwsJlNaCUiVGVmJ
Gk+mPuULueNI5PUycDiNnWWN4FAaTrVeKchJ433q1shCifOIemA2l8Q+KSVH4TIAjQnoxbg7N4Hv
/e8pvbV66g2hUXQwCAXenILiuC9awV8rdY+xXVWquIZ3ZgZPaRu1Uj1AczQoeFtP4azuZDR09d8I
1wHiu0B0AofXN/Nt6kebsy8+2SEMIPJpivlsCQ4v31WSWMDLQ1qpVvW19lHruuQcal/FCiCBYtDX
TVrwthr7ibjTQAtT24tvXBc6+fB1hDQd/9awlJW1XMxtn95M+sygW8QV9R3NIJ2krkSF1fYZbdnL
yfeR13mx4p5K8fd0trNa+qHQJbaen4JNQZZsY3RPjUtqBNLUCx57K3RFU4mcAIWMthYF/PGOYL5M
Fun9krM+VLeMqajvrUGbHTgIeHnBTsygwDL9pfRHUhXLWCBC/smDUZZzdpkY4Dv+xswiRJHTqY3s
3dFqDC5ByVXad+HascFoRHDSlFq1F2GR+aqJzW4ZUkeOiSAiEe+Va0HWJ+/xRLk5ScxMP/Masz0x
dxT7g2wKxpwIMVGBtI3H19dAFFuqgqsvh4YmiSnIVBvLHPK3w6gsKLOkAo8SorS36St6TIk+x3yA
6E8O4qLGY4N252yRysexPr9UVKTwVBhl8M4IWSiGMAp9rH1KTvoqU6UTfnJby+GviefAfrNCJalT
hWCdFh8kqjLmR1wkBqXuGPjaQPZkzH6G8VV8n2FO60ulyOC7cPbw+Tf9yLZKCRacelGIzsMeISpX
6SotXAvQ4NbX5pLg/sAzn8JDCEa1M46iJFRJcimqwDSd1yFrr6b+PmWP1qu025TQ/0xpyKtqE4U7
41IuXoHRdZO7+q1YeE7md04Hbu9rojODxXniQf9J57ftuBR/x5MVMimSPrAtwb9mcnmTZ4phlll7
XCm/u9z8I6ojRgWZdFfPIssd14MQl1y+RmtYA/0fTCYXxtXa/5VpyLIHb9Yn/r/PXLltMZgZqrtC
yfzAhKK+WaMuXoD5hASlCDkgQN39S1uH0Bqsc0zsxRgdrezUJECPZtHxVCsK+BTdSltpzC0Vk94b
rhPtjxC6xtlVQKxWkVp+J6tszi1VNITaiCBxFfvJnn4YVzabZtoj/YniWi4Y9GPVmH3xhopWja3m
DooFvZtD61BB2rkI75t+IVyj9Nb0z+TU+p+r1YerFwhgCXPoJrPIJYnAl8poMYGXxnq1FAYgfUzZ
kJUr3p6lh4Lkq6aveAyJC7K0Y8/ULsnRDnn1iGJohKfs4uJjqKdh2EihRJgRc8xbwD2LPOlDuxFl
HY95VKn899QwBIwYxir2uKU3WmS8LSRs6hKIKDmOZpR5mTbNAB56cwrrNbakatgoi94zsI4Y816c
PX7SaB8wNR2L1D2KVlYh2czbABEWfsxA3gYlic+YaU7byKrmyn08ZSDpnJqbQoljis87kxR3M4QD
LHnsrJ1qtvzk/usO4IkOb5sACrXuKcYdHzkO83oiZSvd6b3tVLXR6HM1GM97NCt1s7DVX988MF0A
YvB4Tj4NcnZgemuLZya3T+2Byz9glkMWaH3LeFUEyG5HvLR2S/rHD6P5qOiMXqR9+m4UAtsUA1ad
DlWQM3qRBlPoG6djzr2IVbb6+yA5F3jJUTrtaQ3eUpFRy9x0FoQVdX13bb8svhhPSX9aL5fXWtQh
pmV/gBYZBukaMMCC5jEmwrWrG4VwXR8mcFOL3lDYQxzczP+goyFAFa54dUY3hP4r8MURvramjLGo
OBOC5AQrk7iHlQ3NOkI5RhYcpAQE3o1DL8Qg3mqQ6KX+NwdbAAvkdhBisF+zgd4i14/7kgWezfCB
xWBuTClmBKkvirYZ5xDxsX/KnHhVUSb3daFPcxv4tMk7c6lwvTtcnBML7y8m+eZjCf/Bcku4ajji
3MxnRgsI53wAThl5LUZ7S9cLo9cXAcJXpcIXU69qMXqL0u/wTHYkjFPUTVKcHKFtCOivv57BZfgO
1c62ORBtNDImq0WFmsmjsd17+vfV7jz45ZRKjrux8hlAdZ5guGuSHq+KwL6JRf04nXBTFbMWojdW
y0M+p0GDH0DTSOVrErSMHcHo1pn8Hak8MHyO/MORUED6CZZ7+MKJsHZD79HEKWJqAlRBv9ujRZUM
D/ju3NkJocCWPh+KkYfBSt8OGnQpAwlyDFPa77zlPXAcr/sV4RewrQmAmouznBsXdtxMP+YMd9pK
vPWWdqOLv1UZQlfVRCp9n2XYzDMibNe+xcXOyrSjwqlyzaoUXDnBzXKyyRfcO4BQ3gYmtvo165f3
EZMfQXb0xOpHWGihEK3HO9JRsEEc3DNHhUdSVMF7h8SfYdg9552pTYoyxyDVNtBQg9hmjDeqKgVP
1XXknSGPEIeClTcfm50LPUy+Y61Mw5WJWYFB9BgtKkJCZpbU2xNsaWRMkkyuaxIFBU7OIo5kOI2S
VnljFMXJ9ER24gwmwVqCqUgKQOYlebioeqS1axLVC0KW8mdXBcumYcIaTaLmNUb9LeLgGLxkoqLh
J8qpEPXnVTGpED7QfXIahwvEnNaFCd5OFIz5pqBUwnl9CX5U1JAfJKK/Bmd8SqcHRl6KBAQRPbn8
4UT7i4iMgP/tCTvBtEzzvG1p2V3sR8ZpOb511kXD6aqGMWdu+uIY/rThaHgFaL15h0ApHwgTn8ez
uUx8rez60J12wB3n6kyJZH5/51u8NLeX6ptzySkOlmyGEmGNx76dmuqZcjjoUVyF+TxKGKX26lx3
1nktoGWiwqHa4oPVxFJ5fuggpGg/XETn3zKV0lvXs6TpbQfyhWwdMmDgfMQWfUtzFoUdYaqCcuKU
ENIf5/AT4h8xpOCMBgEjrDlJCmekbnU8Ql6QCObbkbmpJj3x31gz+V6MPELK+uzOf06gJ5MP7mz8
eX80rJJGvzRKtXlEUaXKHFPIVjXcYe7HQ1zaduun0uRYoA7aHacPcfagoYwJjGgt3sDbvCUM7z76
RZ7QZvM0T6bUeWi9NvBwgsshwQy952Gk5Ok++xgJVMLTj378BgK4P5JTKpfqma3tQ2M3nCoq9Yap
CJgChZ+aAOJKUCPY1L84yqcoRGlv/P7OqgKZIqTvT/yluxnlKFtjVwm4ZwbId5rFlm3YaKrJYMDK
z2JwLBTlNe08x1iqWQT2ZmZDWAu8s0QTTsTXOMLCzmK/mQXd5XmqyCRQxhQhH+DfvPjdQHDTu0F8
p5t8YuYP+mLw41wlLY3/83igSWVKzwxLBHZyo4rzbUTCK0uBTdhl9kuX/jYmZ7WVv8j0Ax/O+k1a
7LPukPepmo4PhqJ62xHZK+kOT1CZR3Idk0O9odXVP4YUJom5jsjHWKWVHQyi3I8MrfDyi2V/URmE
JRPrbk7/oMVDU4SUtyRocIqEpEwY0/l6/VepNzopmxe+bmiJKi0lYF3pbWHpFA9VOFNOoyNJKKhU
2flghOc/ZA201wBjoW/Xg4Iz5lHjtlDh68jW7l9iytpBB/NHrlYUfv546xTxFlLOU3e7zfCTdXqO
itCJ1LA5ef95d8eP2LF3daupdZOJEjEHWh8FSNGQhxWbGoufB5Y4tKVboe5wikWmLbbC4p7OVwLK
O7hPUBbmcAmpZ1PLU3hFL8aHrYMyRBGf8WBTWmjHGW8v+j+vzfQTLz+Ilincujp8RYja3sOEgzr/
cKilr/S2S/g4K3MRHa44Fcb0b5MPZUFv+EZ4bug6XAa8A+dLBI86rLLMSIgqkc5HEnve1D3qI0Oj
O7qNcL1c16XyPkazn+U7JhDY0zG5jayA34R9N/lBHtQkRRTkDrZIblVugan2P6sufYrZAtqWZVYA
bppCi/VvxT1fSgE8g4BMqS9uZp9aSyZSax5UjkUyQPchXwlSpY3h8oShZQixUvF/hjrNqcDrDgCz
Fh0MJxxFwUwJULE3P3ckGeq309gD0ABr42e+IHqzzul53Lm+WoxDtzIObz8JRoVO9Ff6mVBpoDft
5TSE17hn7cKaDxRYgw3NnJPXbF9pMqtizIGEymL/AzpnBkivqz0CLQiiRP91P9izBdxuG57WyOlV
x3TnWv8+XSXVprHKZTLsqAcErTfMNzhcJRdWMBVzyaKFtlub0mN4mlclxxVJ1F+jbfIBhzRrQaHt
2Sn20oZPRpVGuLQiyeDW5OG/9TVK7yfsw0TT8/qnhUZoOZUIJCLzc/VWz872MRCPqpxZlQh+xzfz
pEVKYTM4F/lz6Mq+kjQe+grTuXwYa+YQ13XFVdW9/EopStW06iHvPMoOIzseIwMynUl/qnN/JFbE
y5lKep4O+7z1flIs+CVF4pdtbWQa8d86xddopUR1SlU/yYoTwrnAuD+l8Mu4fx7yyjzxHhd4Uien
/ZCOtOGjcu4wGf+fd3qJL6U/MoxYuHm2Jrvmiqs1vKL7QFwm94gkK+j2DR11cDIcjo/o9JMSThVk
cGzDfvQFGw6FvRZyG0o8Jk1jEJMs826EHU+I55Lohp27x1RMmR2p9Wvko52TjzT3xw3ELPcCHRTA
IIBY9XbZzBxSkUnxNlCEtaIwY5+y6pI0eYDP9ns7/5Tw5K3x3MU8vCwbAzT2Wuv8wSBGknZKxhkh
zAm47SL5mFYpnar4CFXMXr3LEnnmmauIH4wZdJuVZz2q46Ii0uktoO3OONNQyec6+XIAs5qYSgRp
knkYhmRqwsoDDKE5kF60rGMrkWTyxHPSDWRp/OxNZjT6j+TQHEZTGb9EzsHKtrnqG9/mpKo7QSEa
1JKO2qsQCiMUI7quBxnR6XLYHgHJg87GdgUfW2Yvh83hbsxVZxNsavi0TVf28JuxjoppD8DW4w1q
R+e+B6sQyr66EZ5REYtc132l+t9Xp7iJ0uyoz55iDKnUXNk5ll0bJeC5dEXYwIHxCE/e5Fbvj/S4
HUX0qbu/1NmgMJydkRNz+qIbAbO5KSA//n3UGQDIdzQTO5SeXJbYxqu9X9MtruCQkBcYQzZBXp82
uFgOsO2049praTJPLYahQ732LWYzh98TaXF9A9F4ZjKQCzwC14o8w2ln5oyzDR6C3sl9gkg2efqN
awtpJDSbrhLGsUiR13XcDSc9VCIU0qGjueV/KzDZ6/nkzx2Z5b8z5CUEvgS7/R6CpubApyN4xjUD
uUULX4andy9/0OVvxQ4zyVrR1Phrq1qHqo2cVvzkZ/RJiFpSyInfSTvh7uLdGvZ+QQY2rNPOeEpP
Nsg+U5KJGSpdUEWOtl89uWf/TR4iVW3neDfPb9tNORUvNDq0CJ2PUM18t44uwhF+rAzVM1nFTqS9
0+sn2z0/Gl2KUpy5+D/Ua7MOjYo42XVJGWJaTfvNhbD28+HVEWSIrJDLquGorMSiMpWwmYst0Xz7
bA/bgjDvUcjUUU85rSlxpgf6OQIQBm3qeK11D1tLsUMpoe7uyE/Ya8rx9RPvlzTB9f32vknKo5hR
Tpq3GyWcsNO640yc795trUR1nEaNf/JD79hJE3rYc+4jJranngEuiJsQbwpmpdVH7smP6/5UVQaP
hoQkg9+pByKY19EmchW/AAi9qjRQdPX0H5cRPtI7qpnR7SzcYtjkO9toE2kcGq88ZjpA2j39Yk0l
CWPdbzX3mYlin0GX9EmiMOBu1bbKIHDbL9cFk7DL18S6mIGDC1VroD4w8X0sbASXSF/yNKXnavsZ
wdgdIfFAeaAMRJe23RGKVm7Cne3o2YAAEk9FaE3mVSL2oHEfsWJrT6l/3Y5SLK4oHHjqzzgP8C0x
0H8FaRpGKEQ5VCAF5h2URFBwkHQULHRlejpyiQ2BMByxtWEuty9x+mAz+rk2yX2XJ1tkTTkOoTLZ
gl1jCzt/LX5S4INS8RuBFkfSRxACHmUWS4NbUqBKsTZAhan2LuDzceDwOZYbZ8LKXolcIZb6/r/F
NK2sXdlJhbgqUyf79Qq4uPnHcvhVQhtAIxMHb9Vx8+U8TaCSfdQGjdEu0B18LzyoH/c+LGdxZ8iO
Ju34saIBGUE9qhBO34A4t/pIu2iW/1OIKDo2C9fVDfmgUC4cknpb8zNntN7mPqKWUErIyQkU2zgv
mkh8XX/G9NruMG76m4r2l2iemYaS6vEstUUaC2Bdy5fqWF+XWG6PhazSCY9lFGEX0D8sChHst9Nm
qizBTQiB3dnXf1YIeJf9xq3NQulbBFTUvZWKHU0ZgnGSSg6k0vdWf9hIluau3Z4DVN2ITO+EU+vL
iKLLHxrngZ4WzTpgTanZlZ68Os3Vap7cGcDO5R/tBs5me2r2Bhw7rQGyZeJfYUhIpWCPaoQ0cRSA
E6ka/Wh20Qh+MkuSi+aWylxKCrFRpTXO/IkB5iKJFhIh7ZtWy4XqC1khv7cQroF1tOtMItTIXvun
KrgYQHgndEtP8eOtVIB5GvjPFDdYcIiq5msjHw7EQ57wGjDRPkxmXCL6u5jPoh/d082XbRQZjrRp
caRfxBxXzC9W4qRNyygtAsY+dkHwkF7oJTJo0IEbUk4o9P2oi6sb8wdM9852cRAgjp+L2gocRLNu
LHVGLGp6dDgDm0qxgyH5vxXJP6BZNmtjBkbNZMM/JMb7n4S4j2h4zwW1d9P2XeIPX2F4THSuHBvT
aJEncmWpFIlg0UtPFKd4inbvL8EgPOTszGDBuZbZ4MjvMAa8nHCDkfp1GW2yqc2PtPj9CsqYHJ85
38ASioz2a1VjnpL4ur9BncfcrCp/Gpb8HUoGMpuhoUF0NnjngqPF01mSKqIuHn1RpniiHYJK1Cdo
MiDiZ0y0cvslVxkTEBe37gQWnn60+U6s0nVE94s+dzh9e6yWDwAMGPDuhnleIFQJLfvQe2CUev/v
kp3U24PNtvFBoFxrryUuPG2TeMUzzFquvQ9wtvGFP4iZg3NzfLiyrxcIMz0BvU9CJlikD/Lpg3Hq
JsnRfbphf2y6pIInxxnjB7tCP7KpmvvoSjIHPQ8TNHNR4Xu471EhgZDSUYes5J3lQNTa/ar+/70m
gpstvWR9FmtppJs4ZrJRLGkTMPm0NEqTw4tQVW7eD81otxo7g0i4rO5GPmV36IOcuyyM/oh6+au+
sc/0l7HoJarMLgfJ4TnCUtxulf8jKhahvHWzQheOtYI097wTJ7Daw+8pRlzXDXb/G331Dh93zgZ8
/A1wdCUtiXWZRdFZzdc12nJEHfzNEBdCoc2ZFpm6FjlPR80pRN6N4adz1Z0h1hDoo31dV4nSOzuq
XUyUnNDAzgRmUcYPpvvW/OWA3T5h2lTqEnukNsKhDkWZd/h24gTgL4w4mu4F8DrHZT4/AnOVrA4Y
5cERf0lSEtoS+Ifh24Wp/rDV5ls74tehBur7k6RHVQ+QDT0LIzdhGYtcTMuhR5RnX14sDPw3Inuv
xjrJTSk62X0gGB510NDvXObhcyrZNmeA9pIIG/6eR098pDxc+EWOXgUy/BJdzFMJeTcRqLKgH8I5
LT9yGB6ynxW4uDgUu+NSBAbEh9zmWeVAHIgRzpy27zPf627iataU7Iqyk+Wyr7SIo0FbCTRQ59GM
IWcFdvQCt5nb52otzI9cCllnDf4YWoch43PTNtrONXDqqwk/S4admkOB/kyIvZ/pGboHOhU779bm
KsrjMuxDanoYuuADq4fdSpxdBdVHp0pu3LrqpSNM9+I8ICXlTK0tOJUcUByvKKRdCj8EI7QpMmsE
+JqmFFR7klfV4vglQva7Ihk9gjxyokMjYfyP6mnbHrS/OI7/WE1J40of2zJ426Dv7bCxgli2ritF
rKY6Y6Pb8DKlo3usj+lpLn5kxG7FIKI5abEGjYBNwo56l4gksfIXNjd+b3cN3YfdiAG8XLeGUm6Z
QpI++/GCrjUJYB7W+qHT5nSElXnK78lB1qkseuz6uE94/zCnHABBt32iNMetNsQ4TszdCkvy3RXF
LJj1eqV7J5v9TlIMyATMI3qtLnfw/5hYOx+Pk76Jab51a2UyXq3PrXmArF8c9sQ/BeO4UWLeN7Hu
V/F8Prar48u2CRBo4z3QZK58ZFISmwCuJqSI8hIlaVk9GTSaMVGmYbXu0dTHPRH7oPo/y+9LSxCd
ZuSZgo2gPxwaJ6uB8xUzNujQ5G+QSxn0wG46HMLxUzBHpwm2KsP2DkQx8uMQnwOukvjr0eVRxbVg
awfaGD+s5LNl1OBCQuElmZb6H2qX+oFzgMW/bnbNgeuGjMaaUUJGt1lrKMj8XDGWs8w9+xHEN6/i
q2e1fbFRn/VcMd0UvnDOypGYrXQ+YI299+FtRHwts/BwbDxWmSnb/psdw+xzq81IDQOFcqCZh6Zc
Qhy7vfNJSHwtK3FT7E6UaSYj/jNl1wlp28B61uVERdgSGwKUmp2qXVlTYoTMlzaIJpFSilACdIIL
rhfUqcsfa0fhM9FU2KEhgDZ1r+27zPyHYeVJfwjYu7G2w0LzAcTBUEFqYHXP/Lsk2e4QisxH26bv
qHPOxAIKjJixVx/wJOpOpTBQ71WN29cWiLNgccdoHbOhFHwvQVvEBQUR3m5xOrTPKSnthF5BopbD
T2sXlrSNuld5SNioZTFaB+TvxvaCidR7cJLyJXETwKNzZuoHy4f2Bne+bmMI05XySfkAOtidwbgX
2otleuZcPhgTUtGF99FGhkLhnQDzeKmR9P1thGs5ltydfAZYrZGgAXEXCQd1NzOSuRAAXnOPStCM
XcN9djGQ53gxwoNkrrDVgGot8Fnf2heSIVrt/2dcJo5++nIRsLmZ/GbrVpQ6ExC9EEyvK2dStmTa
X72NPWeRSBghLXGr8pD6GFhI2ddWYdOjhPVYkVApIHwBI5H52xRD+p1d7fto8Z/iW3qdwrhJqcQo
Fe9hhJ1MWK2zv9dNtrTxNegheuWu89ILdob2OZCpf1BuHxW7YnaAr0gIZHFrjse8reF1hdaFmKbY
+JsAO70CVr63H9PCV3ljPVb3WB2XjY8MfgSwSEHITnZ94LzGjw8pwFYnQDv37Wn3TDHWwZ3M/+0p
O8DKDii4JNiysN57QFfXocvlzOB543Z5fs1tZOaRhdzwbw03PUXNFOemskJVHHkG20IMVuoBvfUq
UJmXbJR+STln9wjvizZi8Eexe0mJ+5M/OW0r+/DlIdUP4vDG6Xpf1J6b5nLNfJnX4pDRy+8HXrYJ
UYgdAfs+ktLJopLcKYmPeYYvHWhkDGwsxOQijM2ALSQkALjYmaQKSzm04teoQI9P5iaeGP483vZ/
dEz4fdSo/K6gZB8KpYPKw2+49dKmaIpAdtGwpng0J6rYQPaKzXEUv1ExcmYgufBCSAjr58KPHgas
U3E8nTS6uYx6dg+J+Xv06MJkxpBwNE9/Vnzba5p71GEfH6dZTqRaBUdx60jKBKQTDXR1dtvr6XZ9
7TFNcTIWaGdM/yidl/oIgbrJ0/x/FuX60eZJs8RgBIk6cGlSVg+pxrlCgQUfYjQSIC/ZRHx+y1tw
hlw/AKIOpegOqtCzbhQkOjSjz7EKMLUzNwSqyGrB+ve3GUJfD23jB7GBpCwcl4DPd9tYtCRrRYUy
iAKVbZECfKnAhZsi1lOYCQrYHPueEI70Dz4LvFsQXDC5FfcEnQObygjKh4tO/pM0TE+7DrPXrV/D
Tb6Zu5LcBRkXCftpWnRMZ6uMbSW1LNcrEiv3I1sdSgmQZKXZld7kJKjla2zDwb/HayTH5u4McN5U
2qYvWbSvZ9QDIBUY2BPLof6Tl4dZ2z8P/EglXlJ859gdldmMvH+Y8EVLuGnhaUZ6gkZPxTzoVydS
Jkt2+rhfRcoUVAl8sXlP3EGsXKPj8d7m6/QXAUzQobR04YSWUMZ/xJ9JilEOMaMOyvsbyZqsczwW
9wg5gCYsptTCVawF8aQpnQwSsbneMoeXzmCVDXngFA4hdKywlWWBdzB0V4cH46NkUe9oBPJ9uhUj
25l0DvFvqAP6wbi43tJjQbQ0Lhc8FtmSUXf5dT3pnCUZ8V8ViHhzfVcTGS5ie1L1qvd37jineeNw
hLO5eS83D/WX8eqxHa19qu/pt0shETJUWyPSW9A4LQUj6sCESaeb1jRucvcmoQ4rllmihwLv2l8L
qfATTCricBHpTyMwVuF/agPhSsAZYZAoSQvFMctEO25uqmI16mcj7Ux5O8sQGspXaOpI6gw+Z8Ra
8yTFQskwPSoypQq3IYsCMYQpBptzglWIvz6e3w0IqNiTKjAsx2NjZ35ub55sqwrPof/AkniuVY3A
oTvxbUmlb+d/mr3hOCXiCAuxowFiyTDCBmcpXECjFfhDfgBYqAQaBYPMor53mUEZ+CIVTOLeKn9h
zQzr1FuPmzebU2f989WVIAGLi4twnxy4snKScnjc74NtSLAN+hZxhVXSzGsfWo0MIcZGTBO+pyPx
/vqJCUCz14O+yFY4G9RcH1sMu7pl8TizXc/rdFQ0vZhnKOxnF8kUzLZ3O/FT+Uc20bP6NR31QSdJ
diPVAam0lPSqTg9T1TeLrCcgO3VIe4FU9y4lG2vNvURscEoRm2Abgzjkx8RmQGiFLEZNJ603k++n
5k1AzubY8UfLntFNU3oF+g5Km/iwAkyTSQqjnfxGsSum//8bepdyRBpIrK94FEBUCS4FTpDZOJKV
lTxR5WgtyNXSbdJWm4rILne/F64aH0tnaRS+MP76V2pIMntUdGZwT/lKSosUZ2Z7StFo2IH2/nWu
xNTCRPSnZwY2juh2XaqTBvWYSsDQM0vwud6KIYF2HkERJZHWWw8EfX/xOcsSxEKW2p7bGt4ebX/6
pmhBBIVXdskewVzQ1MJWC3G3ibfLt9ZyY78gwnumA833gGPz43wgmOU/5S/rYU4z+KX/8xjMIFBo
h0gFTe0peDYEdCZdqcA4Yaw7s1qrZwKyl7KKrAIdd/A2ayRePTuRgYAkjaCdtXri20KdANrGCi0+
NrucIniyndQLuG9wQ1SgqwjK+N1YWr+Aqg4JQEeqSvngTgOmALIPE1EJu4V924plzyL/+iACKKuN
jZytcZyiMk4CuhV1NghGe8m7Tzf+qFGrJsFQ2XCdzMwGuXKIW9KTWp1QECfPyGA9lZ346GzPZj2h
rFTVNNBd/NPOGjH2wc/nhVun75Taq5xbWcAB1NFinyLzEARSXWZJS+YcFc4Ru5W2MUwo9z2422Oc
RcGsxZ0c2PiwBeebhB18GLNCNZVSGU0+bRNiTjBwBg3UnOcnT6AiT0eyDnt0+qwfCZ6FDJakt3mL
7rcjnvWwCthaxsfzcP3ws7WMYTxqF4Sw43/qD8Kpakhp8SeC1y0e2Ut/XIdCff3KKGB38x5vlmky
Uwyts2ZMtRScZ73xwt0lAqTSXX7zbAgsC9jEHqmwQOb60KnOADWL5LH/ERjjYmc5D8FAlw62pIs5
OZO47QTPJxAdXLeg5VYxHd5jlyXV7GiGbBbwsZHdhEg69mXtHRS87ifgrahR1sT0ldzYawKEa9Vm
S4VTW7hrzOgN+2qHn7EQtRNTfXTOsMP68fWa7EstP5EHgw2jtgo6fxsahjtLl7m7GiO9edroohoX
YjxBikCk8rB2wf+LJnuFvgAX6oeBncFI2t9SZA5tbziqI8bHwlebWUo8bZ0VXGksELI2qIP2o0Xw
kEn7+s8DeqViW0WjRrmHKAdzbz+ULKQX/Rpm5yAAnzIVF1DcflaC6ZlG2gxB2lJNp6k/yrU05VQG
fFI3OQkZMqC57an6XO6dIkEuu9TiEL+xV3efjQAKD+ZALZ8cCcBr3ugtTXGnuHklV+MnYYh6a3gw
qGgxNR30ukSmH1D924Evl/03ETkvgj3JjqHEOcBsrBdmob/cXgt/37Rk9nX6r8Ck2CdbNij9PK9P
iE7UTdYJiDnM+JfwaF5qDkNW2hMeAaIP4UdNT7qYfkDh25Nuw0n8+I61LBWAPLFMJneuQb5R85GJ
IIAZD6RqSrar0RH0gNnefOCqyPJnR4i8bAw7nFo7OylRDN2QjQihv5EsYfnPBKbjZObJf8QfO+Tv
aHibDWfAZsaj31SqSY6x4IQn+sdWv9wm8NsHCMgvthdtWoxxX5Wm+JVRhsbSBFAXjsALGf4w4Pnh
y0BGNUkTiHyU9rxsFtrVfgOFi2wXYd/lFQfmItvpc3fO87+Jw1BcyYNl+j+IpyX3rRtECRMaLzxA
XI7D2Gl1m2Rm+ftBDdY+I9IaJNE6bgJiBJZIvEgVwZLKAaamZaLr3EFIoQQzkhsf/k+7JQqOPENk
rO81d/+1yJlUfVcf8mOXlrGHTKgPulwRkybXY/o5Py5IHiIssmHgGEOEJ6kfww9wQwZKp+qdzBf9
CuBna1cuwUgwATsRNof7hB0MMvVOLqRc9lht+J3NAIKCrLB/Wmzae0F4hki3AefRtJSKEB3wy0pk
dyODCMtlOVMSFNafrhaVOzY1lqFHiG3ZWFltkS+TZbF7uP03UxJLpfxMiVhfUwHlANC4m2wZWYNs
D/agXSBA/SIiOqPux/i20749536cxjdIyvFPr9+0rK1eSEL1TGrUyzyl9DxcupU3Nci4RuVC3Z+K
a2ZVmt2DespxPuzoybDw28/H7ADkJgS9JhehiRm5sAl+U0U84hEAQw1r5bmX7bFdJ37xJoZjEHpN
nFCKgqzFsZKWI/uwCIqzXXA6FVAfevPHZQokX77VKjNINca8iuobOzI9rncC1lk0J+KWZ3nxX2k/
SfmxtrfGJ/srlTi8u8a1Knjwe4c4IPJNMda0pVy2rp2KrMf5cbc6Ro6d6+ZAsiOhqKavbqruwv/I
VPZ9IkeoSoQ63xY2m+izGoxe3bCFF8dU8eQ4nX3eR1BkOFVg9Kxzvu8PTf5TiMOQQZzmKS+nu4iT
d5rVJP3tI0hr/Bzl8SBual+bdqcUgZR0ki/z4mpYHBByDbhEhLGDsMqZO04G43bVgEmi5m7X8bLn
Sd+KJFO6gC7Th3/dGJaGfcFwt+KkJyFxGWUAzRLvy6olGhReN148xCOPu/ae0WsYnZXe0gCWbpGv
mDR3qQAktqigKiT1sFJ3ZH8DcLSNFvG6EkeB63f3mSpO2m4/TZv1zeoaKfoloAznjGA8sL0TKshq
StMzC4IoL4+Xgvhd2u6z1NQOvJn39NXtsCFloWmLcD5Y3TeaR09tijH8+ZUqUpLOMnIwYybwHD22
ARFrmw91LY2GgpHwOKrOMKeVpauuFWxWn6B2U0tBEzfliB31QmAzDgqQZb99nC4pXnjOo9uXZa77
aBfN3ZjDgh/cIxMncKTh3EUKV0cT77HBZb3Yc6MB4n9i6tHyqVgvpeyny1em4g7dZ+KzvzlQoloW
wMWVvXf95Dxh6AINYf0FkRGV7+4aD0zvS8xc8crI5IPIAKo7XZjwqCxGe00oDZLWLKjddxzrOKw5
xH3MtUrxp2XzPS847HuT5crhAWhCUWygAluURHwiNKqifFoOZBc3LnNHb6ysBUZ2J3F4sjzdYivj
bdYOIHN9+CdY4n5wMU5HvZy7aRn9FS5mEDnP6evNkleM2He6oXZc4bIo7iFlD0ZMn5MwPoCSGVLQ
plB2jpS4nHBd7Y5IEsLBRRfaRcWc0iyh/SFDXgCaf95L35cAP7eR3Rz5JlcIR9TnrQUFwrQCAMGF
MqkgunEhPJik6wMjCjs1iQ5dfKgL4WuBQYzCiPy5VYM0sA/clMFwK3x0L+MC2O4WLrcXRkC4PwMK
78ch6Oea0lypdeypG7ldg8kJogSO8agzv4fePlpdutsibS/VCekWJmAAkq8G0yfPRTdCssCA16BN
fHB3uMvS0L75nd3wwHexGR5Bm+4uMfWHLecwWYqKn/FPe6Sr3rzOQsQ7l99TxUkxw4w2w9MbdwAX
WVM90XWwQtPbfDIj+YBlKa1Em4v+JarIaycv4/B1eIuQF01iZcuBvWeBSOKlIGh2hx8sqamOrg7F
EyTxqrKjjX+Tq0i+ylJlggaDdRiWBgm2b0CPCV5K2frzNwgwcjuiSlE4hThroVR1Z5Hj9jYoO6KS
/8q7iajjlXO9ui8l4q37j5YGNe7OuCeRAzm9gvQTQkF7gISnLuZ8LyUBIo27GmHQ+TuWOiFE70P/
caYNxT40ngSleoHlUDZNwV1PMnVR6TxAOIgVbpmLQyQ/xHRH0vv31xWouFOmrqmLac+/IyxydKuC
FUW+HivISrcm0D4Lis8WTtp9ULqmF+wVnK8VDtJjfmRpaqy9hcd7E31loExuLbxShZjbrJTa4y0q
IxfErPvPoTOLSa3XNsH/t2KCZeehxo97qgI1E7ry6z+ipt1cEV7h4C5TfIC5WKQiwdAir4GN6UEm
UiiWsspEtf3ahVDERyh9iy4qZLmXyUupaJWqtNxmGf0iYkXok9fCRoItm/OoSpu45SZzCHPuim+R
xAmTw0mIXN4eJQ+y2EXOo0yOMf6m/iFLwsWMh2mqKJVOy8tSZPJgjECE6VTrWMlVGr0eHl+V5LBn
WwabK/uAnaLk3piLpmFvlGgo8qMSM0PuMvcFilZl8YfMGd5TLhyrxPAW6dHYj3keicPAxgknJtBC
ITuYGHjiofKaMmTvUH9cy7bS2GcNN/U4yKJh/aabBz0V0RChf+0A/UyMswoo3QjPrk9yrwhml0Ga
XHzFL02MH/Rx2/UIzMlBHhZs4Jq7g5UIZ/vbFH9/hM80uGtkHAtMUp9NvhXyfGq0Dkls4QG04/ah
Yu6SU2pWqjDo9p1sjSA3F2zPc0qUhOxn2PvUS668P+1NeE14WTd736J5HdYtRJKJPA82mS7a/kTA
tKJSnT3mFzCNwQ2pgE2MvnMbZ1s0RLeTNeWN+TirF0V62MwzNr8XtH+ldSIrbtaOut+moLftLfWY
0sOPJlJvfAaQgX/2swybTkMKR/3PSARHQiF5TuO+fgoFOCaBRGwWxmMuaFDVxj9x84ZHRHKpgYfE
8gKqqEMdyxeBD4O4WOTmalnbBNbOSSApEALpGka+AvcPMh2QIEWL+ur9RAncf/4VqNrjpDGnr3hR
Yhf/bOcqt8OdBeNUpOobPSi+ehuXB5cG0ns041pDJQxmkDFduugYuQ2MGNA5ynDEPmnP5mAUBZce
l1b522SeUyqlNrczS2PLc6ZhGxxmD+ZgyFEhflm77xpAUqMBT1C8c5P2BXkyu8+t33w2VHGPQW2s
ytVhlU3NHJSkHAdL5Lz7KEdTYqGJ3ShLS7WXE4/s8BG4GaTWN7uNJhpJM18pHUy1/tVHGNMbDJaj
RJjSuQUoCvOropeOUasx60V3wz4Z/3ulquelOcBDO/9MTYQVpo/1shHKGezyKsRXLytlBjPB5P0/
naXSfWaRtyf+wOUkWus8hlgJxXRelihBR9ekPathJ9UztCEMoN73HbPFEZ9Av9zpYFRYMXO7Lec3
mjIH2cgmqjOJ9Q8wK1WqXwPrwxuoTItKSkvXE/kbvrEAmzOTUMcWn1tax9m/XUTinqx5vzClTi+j
xHfWiiclMv1SGsL7N8NcAHTGsAtjERvDE6NAAdIqbwcGDOhpVBLSFksbv3NWO7eQNzErQY2b8Mdg
xg2wdc7Sr3mTNm6FGkivJ5cr7WGwMvkiGk0EnJd77djPpQ6czaLpUtlk1EskPrJ9uXePPuz3hS6b
w0A36b70Qbr+Ea88fU7gvaxk/tHQwsRMZ4/aS/8obQ1ueHPJa8yNYcT6qKAN7XE7X+yE0nvXErlz
u0WrM2eL2l+zjYyWFr+/ETWt1faeA+HAO6pjLMXG9QWMJTnjys5NFzQiZgUXZCYA1e9/ruxAok7v
Ak8aw2QHKDCRtuiuHQ+YdOzmEaI2K49yxfsbGkoiuZ8XxaPeUsy6e498Vcc0j4skp44FJc3r4OvK
TyAxLBr+BJpF5bDCEmtejxIccyZ7VeYjVEHvhwxJ9s/SMPKxsFW2EoDpEC9KYZfYvkAJLC3MaTY9
M5gHOqubP2GBdKjyHpSUKOXCI1NQPnsjaoaS9LoirRjLJh3++GiMTA537bjnuHblE3cKQYfdcSP6
7CDDorTH9EZptUfoLkjS1yTkhRYW9qIgVtXf0eERdXrdTRipMuXFocR4Aa59gD0GsUUDz/KXPww3
BOXyBNatBYJ8VFhrIEvP/qd9QkDfEwARxpLR+sW2x24IAW3GORyT6Vg87LsITd3yXb9c+l+Y8lfy
RKXGyjfN9h0uvJOHMm2hbelhC5vxg8I3YSidAn+MN7Ma3074PYGjHNVbG4Bqmd90zCDHgkBFRwuQ
16cwzlLB1d7VNtpMBNY1Y8PZKQN7HzqY9xXs90C/hMhEiwmePo1ntMm6PahmtSoNHe8DPReOzo90
Z3z+Um7lFTrAFmvtW91qSG/D7+S1gGM8tXsVd3a7TaY+udNnQ1Xord81C2HcUEioEYFGCVz4uO5A
zASqzd5sTDh58qjnfQaBlUOvq+g+ZqSVGnqibFxw3I6ICBHGz6Zr3dniaC3yDf5v1Jeja914dRqz
iAbmFQljVd6Mxj3/3AnX6BgAlMGCOCYb5clUd1awaHXCp1M42l/Vqp19jIFgqNUoMKuSnHdts52X
1TcOIcHUWDMA2T32RsEHYhC1OLuS1yXTtdYT9nqRBdOzNnmAnfamZpYC44sPeDQ+2n2GJexAFKqj
C7ZFDICnz83uT1kaqJfUOdNPuubbeLYN1t1GDzB3QOyJ3kRGDzIBTlEMTxfcdnkrJZryMJr3Noh9
xhhD7r4eYnarJHNyF97IfecyZ517Dhe4lRAe8NelPh48DS5Rd8Cy9WcD3E4GUjq9LMXsvJacfnyp
+1RWL3D3ZPvaAOMotwSvz5CEkvjNVFaELoz3XcpBfJ170PJO4N3SweWuWwtSZZ78Ytx1/yNwVZ6p
/6TCAzvI3SJ+lcpxdJ+BjNRqO2OEp/57HSJFKkYk0RxVUAZeL5fHvnAaGaj+4LCZdr0Siw98jjeQ
id9YNib0BUwI+gG7nNcuLGCSHxw4h20XcdqSUtHX13TmZSaJKORYoZaRH1XHI72mS8xYO/6n04Qk
Fe0wsSVnQy3/3DScBo8BsxUAxklzL7QsCzkdAwr9VW8W8Zx/8nhAtzzCJU51fgaYKoP3cYcxdSiW
FnfxikVGI933fz+aydN+AhuhdIb7TLA9O1UB8RZ2ccp9Aflhg8Sr9SiG0TnvMS6Oz0f+Wf/GqaDe
6q4OSQQzDftbTo1f6Aw696Pa7JNwSDwSPbW55iUWWkrKFHeY4yclfFJ//15l3BR78pomKo9W3Y+g
/3QZoWKyHPAECBCmv4CHGAxsk7qfa5+e5ohAwMUSv6W9YcQ6gHibZZpj6I6FVv8O6aYBAyJYTMoy
gXwXuR1hIlPpTdOe+uXLO0zzsBNI3ghePpF26a70mN1jTWLio7RP2Q0ZCX2gwCOzzNjPzU4LyRyd
1p/iyI+iHsRTtzsioHZQ1bEtixtyOsVtZXCve8okho8XESF6C2lo62bfGT1wBqmdaKxTcgqHI92d
D6XhdAxTVzuyG2hjHbzuBWP5VDshGSiLKkmJLyGuqi5rL1jfhGBW6oIcNv3l9nr9tp1VlY2uLeVD
KIytL012S4wMwumwvHnphchEDy9ONciOw/jb5efBZ8hMBq6vAdnb3t9picafW21K8GnaXn/TZhCx
xBufFVVn1ciXvfnIxxXyl0lfyL3zqF3gL0IfATBTycapNSQ8qfdEz3HnIxJmBy2V4wgqMxWmfc2i
pWc/kTxAwvxwTuP1uJZd+TsGwRXzQ876eBiUqutjg4+rtJIXCe8ciGb1ie7YntWNfUlzFJDICBkP
dAAdSUhY2W7UyTTYOTp6fOhGMsuzLAi+xYP3Rvmls8pdx+R8gUOWOegsQFP0Kv7H8dpkmrXvgy1f
68wCkwdCiXxE1PLtFYuAqLZuKA+Mw9IXyX6bfoCESND1okab0rvJ5tK0m7TABykapsMawhxOLyvG
imC4VS9h1X0ItRUGFo/oivMtr3dpsA0IU38vnK7bobwJIj1xj2QI3RQgSDD8QqFP/0a48AV4nQue
4de/xR4YXg+flSM7yLJVKkN4//JXjMRFX7jkFlx69MtoClUT8XWY+fHkqK+C1rcPVlziKBxKfzA8
Lczv2Z+IH7PLbjVWvTDeNQwBJ7LHRTZES8fOHbHP8k/Ai7eZn4N1vqdrZgnRyMhuEXxV2HPjhywW
/inGY3yABCapHHxsyFUUdWojoGXuPDjcrFt7n7JnQbwQrCfMyEedDyFJwUnfa8gi4kEeGYQd/DvA
OOEztOVR31vtbV7RNvQU0AzWe+6SA9fOViH/X/oUfN+Y/Otl7CB92XCkkPYfUJeERdrPR5ZLxPM7
HqxLQcDKOgeJfZ99SRS/D3qW/NSU1niRT30twqpvqGZjioibc8z8ULGPz/+OM/3zGAWl8fMzmcAP
cxRNX+UEjpwsEXPCdoK7oKMh0z6THa9ZdrWnmaIH6j78x/NnAgrNVwUkpXb+90adLr2Rk4rTwbuz
YPSM4VjYmR/2o3zaP6MEeaE9RBnubcU2xBut/kAyRMCAdSLVVm6VxVpq7c01m+WuJF4r9KvW3hoF
KCNBYO3f/qJpvC4p08VFwuqID9hrr0p0aRmTzzlnU58WCNYOa/xKuAEPM4U4vAKTId3o4WQPopsO
Ut9uVxspcVPO/juFhYvL+iKD/tZKwOYsygSHxOphbNg4bmM1kqO4Tk+myJYzHSG1ibHXM9TyRCez
pI+4REsOuFBW8HTLjGzUKXInotADN785upwD4HLCA6qpYWicSWpEVYOnS2ljtwDMwdHmnrf1Jrju
LzVybYTlcOs1bQBqSqC5g0PQL7+iZzYy73IJnKtDGd6GC9EsKscOgA/VQ2+2WuaEyXoOX+4V9jzm
md7dNgZhoj5mm+DdPb1ZtDCfKO5ldA/A0JrVlg+lTmIEcFfB0XmJJ6W3Q3kQ5FuQKrCvNPvF9oga
oLROo25TR541AcKCQifd9Bs/JEmsHrYGaMgLBBegw8wTo7Cp6WB6SY5KQ38lAgI2RQ9fgnBbZz5/
xiNr+NWoMolIb0tC0W+WnIV4Amhhr4wX3C9i+0sBrNNRpvbkLyDttxVr/5uFWTssyQOccjnPBU5I
Tc1DP7IdbfguziqaGRqPWjUn7xYTqiTAC+WxVj70+NQPPyNo0rLJQIvIeipoDQOdxlATjQmw354k
xSP9nsvJASH3NsO7+NlfSc5nF8XvUlkcxY0ebeR9HrKy9Vnwtotvx+vkU6iRe+U1ciHd8RJ5QZk4
VvXWhN6F6tIaWoq1WOqH0v2ORhSysF2U8WmViywmJN3GwURAXIp+QTZyamsUmETb/22k+Ox8atDt
e/DB+hUkADY3sLkVxYTAbMS50BosEMKbU3GF8nww7FM+DqrfWOx+6A4EaHBYNGCViVe0LGOYDuDi
EFbbi1FOch9gOI5XNaXUN3fpq2DRZoMNOWD3FNAIHlJp1Qg9Zur3zfp0VNXAuRLghDC54slZeAeg
kR33uR13cMZP4FhK1jZKEC/SLa7RsJpsfq24sfEkS5CZYozjtD/sFl+LJl2AKLd7MR208gH2s3hz
MMqKYFlhlQA4ngO0GwjLBOtayGacJ546fUoYNlfzl828euEuUlpBwW0ZhlwEq9KrX3PYiLwM31RG
4KAV7b67E0J0zxD1NV8Wz4ZlpIZQbbKEiVk1hH6gEHpgKTfxmbWBPpP+Ow9TCNGg9+gShDOH+roR
qOslNFtn27SgT9uGKcCu9MwUzXfbyjl9V0Soi28WfydGcZ+aDaMd80tGdLcB2WoOd5AtL9Zp+UpN
AwLk3JI6+9R9s0i0iX25dZAPHUlnW9ORsOxh4ZEkVzqFgIip3po2llNbcA/tKuII9WguYMDorTiK
y1ymRxvCQbPJMvOJvQUfr14GRoyXwcxVz9sFQumB2F/EqqH0ypeQbF6B5NpTpWQoYeE+CTy72ZVK
i0y3UrFU3xOCwvZ6rOjY67eiW96XzR7dezjUe5Rt1RKgLTaJyJmX4jAKtHCil9aekcsY8YKbYyK3
ncRYQ8WGD3JsB16+AVeql91/UF/QvrqqOXAFt0e7Y/m69V1aIFgSdoqzqD9SlNSa8QmVm9aSNATN
M3Ty19eLCVYMdcb1XhmYsFtETLm5L3wbXT0YIlTSSOdRzlDaGkBBB1spcmOfcMjbBgjctigPYTxx
ekvoj/e8HKJmt9AJKuwrucBTkow4VaHKtMaiNiXWwqTN7qgtctmyzDhwaxzUe4UBNkflRQEKvPJb
RHThBAk2BsJJEbVoZK5wWLSRpAY73LvjKADi7BHPaLfsQTE4yfnpVArskWpsbBlxvw5s+Z6X867a
EqA/h7wFfGudrgFrUT2qf9A6yeylWcU2hvD/vQfJYQEOwBXXH1m6DHY2/WLcZTtkQfJE/Uh7kZnK
TnZF3ADGSAsCBKqUfVnD9w/Yg3MirGcBJ59HjdtEz6GOjZrz8A6cHfIde0EgGEKdg+bor5438oxE
kVtP8bxdh7Koz+Gx2jn52RfRh5sGVRF4SxOGjzrPkZBUMH5WQBWs3XTL2Dj4kY9wtVAE+meWjE3R
DVNLw4AouATDStLZujrDYYi7F3l9WJld/UZ6m5N+KuS8cgCuBMNxM7zvc0bE+MdcDCVpQsJUdbqS
SefnRlw3O8EE8CI4oE4w5vVndWbRVF7AIq31dvxjUX16yKi+XUtHjtPgMPFO/xRgLEWvMQ9iSKkj
OG2bANIqQlkOha4LpDgsV+lEUAhH20WblqmOkC6btfW/wxHUMXJBcVhrBduGNCJj0ARbSyB1YYYO
isIBwMZLvW2KUumoaY0CIgiPexCsShN/Y9ESmkfM4HjD03K2Dex/pTfA0/gyYZndzwut23b6NYdx
RY5oAmUh4b4tJyTcZa/2xrYm8kEqC58WdXwy5URnX4LK7TdWnXIVdztRzZo917IjZzcFjpxZQr+h
nnGNtSMoIKP2tcuLny9jque0vbkUxUWeg4doFWL1Ody4MJ+WhaDIW+3B518ivyzq6bN4QjUnMixO
lfOEQjEUcArsAMKknT3RDDw0G9FOZMyVEYk7lx7u+Z+RUIQouOh/KuDOx3ecW9IzGrgtb8TP2fOJ
zaPQHvDO4xINOuEppTfNl0lKLq9pZW846gU3Xb2L63pl74rbefMCgPnXDHoohaCrdoP9rIdoaHqS
vDkkKFfVSqCbnpuXp98qEv/QNyX3iM1CMVSdS0LvzxMMpnNKK1XYY42sqYvuasF5R2wi4GZEmOR+
WBJf9zigl8e7kbKFl2a90NcUhgjyDNguaRIBMOT3V9n8rdqFTs461x77V9BwIl/N5ybW7sY/H4cf
Z6zv7g/0RTwuyMLaZhp9/blHPecT1KseIVo94MOKUyWHTi5cic6EdKu7IFoq74CVQK8++u2McI84
gTDzo7LOfWwGbWCSz3/CHOFfeivMXBInP6pJbuD75GUZW7Sje/oyH+/Zpjr98j6CeFMfAZqYhALk
zs/WGHJLdC+Is/cPGkL6kS5GgVZsIeML8hjNdbgmuvCXDepmQB1u9wpNNMWjGV6OybeNqiwcS5qG
u6QjDA2uRZSd4EvuWZu+eCKgsLyxXeg/s44nJB1ewSMyxwfu7jAvPrV+CB9hO3gYJnaYqqY0/1cv
6yu3TpZlIbVm/dc8JY+OwHNjlv6R3rp9nfvG4qt+wvXLKrauWbk+PaUug2BVFu3RWxqJnhyCQuU1
XNs4ldoMAs3pFja1hd7xvpAy2l2tn/SAS8MuwykwBiNePGEdcQd/WKjq9R3jd3P/JxIQZ1BLC8et
UNyNmay87xOjeDLVaMg9qW+MxfJ3gRzC2nVkwMy/5jFQ/efhk/qLgMwZJ6cXwuWIQkeYNuIxQidN
VbmWV1NqDxLYkaS6N2GQMfCs8og6G3rqz1ucAVU3mi7JCTZsFsMK0BGYPEzpLHod94r1kNHp7xGT
TDx2h/6JJFw9Wx84ULNzq9QAzMi1KFWn2R6tjt3YIvjjvKdJv9RYNRchSJPjSgkuuhRoj6EXBj4V
AqwufD6nGDFcK13gZmmyoqCUHkOseBgmVqUeg9HV2U1f2Bio8NEKpuvwDnwq4VZvfzv+e+6nuGKr
4+5KtsInOYTDWchKl92e1I/VOlNOfavQ9mQ6VuMpumWm2zGdtInzZ4pc+5cGulLFffvKKSaex0X/
dkVwD4ukteKqzC9LVKZbVK04PY2SVgUHKLYOAuEdtU6H2Sh11KS9K5vtkMLXTzbCuMU+pJxMAurW
BucaPtjZhpjVitetdKPxKA9VofcNbZG24nhoG0do4wbvFNNnQiEjiL5EfL+U+IjMWGOTgLQT4ePV
NivTxdi+MLj1q8L4yZWtjVEQzIHNuyRIuJYRtZuqHiajsTh+aIVC9YVXjpLKwucA12C99IWpkrrV
qKWl4P1DWm2Cckf28iMeKtELDAD0yMR29BRHGkdcnc2qWIwGAFZWwbYOlt24iln47AuwSo9Sft1s
hPmNJOfW1eseJeLbIJDn1xNCGZeoi33U4a9xGcJCGmPvIodH7ugG/dMWd+T2D0CUUehFJMx8m9f9
aUkMmyx0EZT+HT+j+x6tuym4dudUdZ4OCsvs42H3M0BhdPXnyJl40Rx+SMUdwzwH29o1AD19QNN+
+YTfl6KBW10+q13+MSNfcGDOO/a+V/u9xhNG2ivTZg8pmesuHEEJMIpKAFxJ2zii/GHmIODR9PNi
v73lpTBwFDf3jfa3DoBfXsbyjLNQ65drCNJEYdYPn7fH6vBKedyLUaeH29kIVxXCgx2cfZ+CvHrh
qpmi1ImPyUbh/nL7VWsDKic55JSepmAvKHItnTlmA6RHM4vsy4WCEBA1u+ELViaUNWJyAyz5ijnZ
FWMzeZaeD8Gvj5dbLXWvb0aFYxCkscc6+/oOu19MnbThBZGG40IdFbIzugd+LBByMfnOlsgtBkcb
oP0goZth+szxeMrSYMToiLa84o6h/yc5AcgCz55qvnaSONBqXl0DkFPORcK4DlMf+/tuG6mzBgkj
jR24z++VvYMAN4S8gC792jrgj9hgqTbzHwTmqKk5lfeBohMiVF0ebs59oADwGAQyT/GPcrR0FFoL
e5iVqmY6HdKBo3Pua2PSxcLFNdz3MMbNPoH36fAXbaUwAhBH/uleeYLRmvdw0dlLbWZHINgC3vq4
JkkFwakSokhanZB5D1uJrjaAtA2xKDwAPZCuqxuvcDT1NbuKhZkzFAeuyv+wo9Ak/CxI1xi5JqPA
xpjxt2U63DVCqhZWtUm64Lf/ME0QoJyvUx4njwGdJaxlkZ7gxfFxrbcVdYMPudG4WRPwVqoaO9uL
gqQFZiCFmYAVADGns3wCn79LEuZC4rSfefefa1LeU+8Ivg/QFJHihU1guSeKDZg1DnNG3nU0cIX1
z/FLNOx2AondDXmaieN0p44lolQWwWy9HATicXyFpYzaA5dlXmYAytTDyeGneyUqBM5mJ2mVIoUX
4g9CgfkUkKkLhlI8Tv/HXDWO1DjmWLf/nCTRDhd30PpnPhuidOhe6JhrZz7XLNz023NB4KEgxv+I
Y9IXEIkM+Lf7IonncRcDUt6OwIh7qLza4vmEwMW3Y+4sM6adEuSdKqG4jdwaX9Hzeuu/w5oQYIxS
/5BSCpJa6IW7cKFGwrEMgVFATCZ0FFuLwN+iu3F77I665WYGTR931yodbaCQC1XQ/Hkd+4PwCu67
Mf+G5UJk5EuSOJfi/8u82K/hGGAGLv51QiyJaKPNDDwd0eRZTUyuEcBe7NVcY1OKYFh1kT9PaTdI
nF03bl2xS3/l1+IFzkx9ZJELJmhL/+aYvL70a1aNBDcsXtCHyE6V95yA5vjE3Q1tfrPSegRrp85z
yQkqB3NbPFRkuBvBNqDbMvJQV3CUQk/gHaIAXpS54djXVbbhOXjgH55sMpUJKGoCPiFHm6Pg0PyC
5B/uwNZiIqQiQabrKFjiyYnq+1UP31jdYE3fF4/m0KErygNJzH14Np+LAdshuukPYM27QEhJkGu+
08cCoz/JoZ+pYhM6gdX3OupMWGCsO7mcHYLpS4HxuSpCO9bMZGX7KHvCYx6odu7JHE67IRpZQj6M
v47od0vOU7Q33cXPQN/r+mQpx4EdP6VgHCIPjuINLD2bYRtspkPsAaxAyZmo4Z3udqOSmLCHuapD
/7tXBcGD/NcmYX79LOXRM7ABakp4g26HmKqKRqEfgK8lUms0k/J9YCx7IcOuZ28DNGCnT0AAw4Bo
9YS28gE4BW63zJ9lxRz4DDKeMOoU0Ld73I3E3qHgqbOEGBSkzGLNpbEExjnfFmo+XgC/C7pUO8z8
+4KinjMySTCrNyBE1wo1ra0lyvoLBPDE4MTFoS0RrI3ZCxXNhpRLsDHY5fZDlaEtokFcstTeUTVM
4SYVDHNl/HKJ5XD4Vsj6pnwTLDuI08nOpSew06ifqx7ph4ZFTh4NJeD3CMLHmYiZ+1Z9Owa+V9ZD
N1KxFNcbT/LxqrgkG61u/KcL9rbYGZ0g6GOdXX/XJt78BaqPRXWvRRuN2jaxfBvAd3htEGmlXen9
xEJgdZ/Qq5odZis651mGqZr0L59Rii4s88ehnhgDXYdKglU57t7qm2SJc390hc+M/CoNz4CcAt1P
QhxKYw864mqA8GFVPOiiUhAV1N5hhe+rmPOC1qT05X4Z0zb+ZLHyK5tfth9FxqKKsKLGoSd4BTI3
YApNgv81oB425SD7B+MV6fcK1Q6LLuRDjeF29SujOO2EM3m61rqKN2czOk74pIuuAJ5WU5XX0R5L
wX7PYNztcag9TPu+9Go3TMFC+H5Yzze1K6XWFu6C5snXLn8rzyXkhLur/SaT5wR2z7MIONHesYJr
06MtIbyjyUZldOkpRTocBOW7y8ftRxtC5MUkyx0MYDPM+fm+RNpi5VTWzwTUa0yaszhjRZKvTNor
lxReiSq3gH2rDBDjvaJC0UptfY2jNacTzUmQMdU6V2Fi++sYwEvJPwU9cmEJz/mV0nVFv/BspenY
iZZbOtA3Yyk6zf7P7Z0OANDXx6VBExlf7vofIy+mBRYRKXVn02rOZM+xESmsR8NHl+HMaUIUKLp7
SS6TqwoLVDdS/XndzY0+ZQQ1DDMEskqyX+ulm7qIlBlKLl3q21YnknUTXZMGQIpJPpKxoJU4XDG8
fgpUEOWA40jyYCGClRYIAmbEzA3OTBtF9Ti47rKqcyoL/A4vihTtBvCGN4hAExbzNPI5+7TmbIg0
z5/glY6NzvySW2/8Irjn00oKkCvpgR+kD5rU9XbvhaTNe+zoE60gIFZpq3elSy7/lOvp1pM57qKy
bPndk/PpfJ+XgdwnBeG3yGcrV1Wy9qqDMw4t+ePI8XCxvKzgvBuGBUt1QBK3sma1t2UfrgU385KF
3Ao0F97UZd8hXVBzL6xia8FvDymKop+0pHfPXLeENyrSjzajc+OIVxk6s9ZVOfSdvSpmhzMgxF2w
TxLAou5zg1TDfhyyxFIbvxbeNuSk/94CMcengSo8hH/cSvlDpZgDu7lUavU3jybH+N70rcIz3l3s
/49pCrqW47Go9foYPClApzPrdLUL2MjSWtlouUvEcoi0BYlcT8qSlgc6QHgryHheIf631o06FM3O
8AXgNrYAmFap004IoHciXQIBHeSkWC8faXYAA55TNF7E7bmtPMfB81yD23Uml8LDX0AGqDqC1n1z
x3WODsmidKL9YEPrxnc8bP96fvlakZ0/+txopVS5J+UlrpGqZ2olxx09JCR+cxkwhd9/4y/XD9CI
w1YN+WWSFCT2Lj9Ii2AzCSr9r8FCJTzB1pMnlFeH9PplkZtFGX21qQI2h0+QostigZGGnIr9Nhzp
DfVoEe1pxcWtyVh0ihbYLBiiGjPfGNoccdvbaqTaLe6W7uBaPp69yPsNl7RH4VUQb5LLTh5+50M5
yrE/S3suKlG5PLrVn9ivLLQbbGVM6T1f6LLmeritmuRqiDq2IshmoV8vIwK0RkaSgW0kyy76ykDR
7yR3o0zgCweGD8Z1s2Ds/3PiE/iGyl4WGpZx4IJXyjpc7rwZ5xOZAxjA0Yy2Db1AHI4ENl5AuqDO
a6Flz5CF3vNVdmV/efI2XP0MvD92Hs3cSUtO/MFEcPDsY4DdUGeL6ja9uFNjllizbhA5ANm3oFH+
irQfca6tYfgwovNFr+TAfFw0SqJ0Ykg8LH/IaNQ/V6mBZJ29YJmPYh3OtgHBghqsfcOpYql5RQSJ
ffrn+5sB9V9TEwfBdCtESoB47dQnvG1xDppLr/T4jN0kw5hI0JmYWr9ILhnUD17jja8TaC3rR2ZQ
dOoo3VAZpn61Nwuo85r02YCv0LI/7qindEJPJDvCQVwuyPA4w5i6gZapMDZbmcRYwMeWSux9x5fs
z9LrL0oin3uGkUdcYQFlsNaJ9zUpVxu9JolQhlHuOwXq71vpBJT0fedMa2fgKawShtWGXHS1U4yL
sIbbU0/3nQOOtEGltzLhy+OWrIif0lwI962BT/EWf8WLYOZYZ7QsUioMYENN0zxEKTI92aF/7dyZ
lcaukwuMSfjRSv3oNqyJseYuFbOT+TjG9Ld+i9Ded3zuTYRGWP7oSSAdTpDjAfdby4pn4FKf8zgZ
BffGSwdHxwOnaQCUKPA6UWeWUrn14YLXYVAF/RXmh3CrWirKLtvdN/hWVFl79fYJFjzw9ASOBwcz
4xRQ7TXTj9MMY+HcHF4yknuDSRKbFhwh3RoIATss/jj5u0lAX+3tCZneMn+H9ntXY+CM2OGEE93L
JRZwfydjuPU2Mu/m5yGcuo4Ze6/wMpnVketDpFCDbULgd80I/7gY4+qsOLl8Wivox5SSEghmq8EL
L8GiHGb0eDwjzVyVp1B23PApA+tDf4QK4Yddduwk6k6nqJbGGdDwy8YlB0pH7lOZj3yFbYoWkiT7
OTuXYAlhb+PEAqk7nUL49t3U/M8obrQFqI+49L66noNu+JZpASLXfPBd1JZNjKT22dCxNTkcFkWY
bjREKt+ADchQJ+ObwNDZVci7ga3V0wTHdPCItan1bOiRtDtmlr5zSF3VwyELmxiXqfqfcVd+VqXW
jXsObyyZ3TtIIn8i8AQE057wqeYvWohdDE+naX6a4giv/ukQTi5T/27brhVRbNAMIY9vhv9tk83m
4OmpEHf/iYuuSaJWtGADnkw6aysLySOg1LDrSkaZrlnXMB7zvhffo7ih2GHFiiZfG9bvzMeMq3/c
FQL6mDLQu/G3xtH7vU+A0KWCzZlFzw6on+nfuPTeo4e+g7VdbIWjoepC7bZZg1J6kb66Fru9hFyi
g7doRni+n01HZ7uqFgMR7/0/2CLGTeTXtO7vpyn+zJKlLkWwNy3QqMaelDFpPiUMPl+QkyoWP6Hy
OHpFjA1LBn4NxBuM8gjU0Jmx3FUxebVBTknbLoWUcDuaRElDf0Q2U3Kt1SXUA5LDHTcmvS7Ox9e6
25KzZY6jTyoUq+cHpoJDfEwTNDNKM5AUM0Lhk2e+Oc/z+oZ+SeYY+egOTB+AICZGzqtdY4fPmD4M
z6Ay9GNIORrNtpDWyj7eWU+LPEJKvKZlpz8jWxOhLY094KVL/eKLDtSnvLaP41Fs3orWEEOkZSv8
Jq3fqwovTEt5JWk7OpiB9Cf7/cGOogFaSAfQpKgL9YGdvnfK40yRoYeR2ISb6dosEFxbItr7eRWj
psLiGdyFQF6VQtkS17Ov5qNO9lS9GyDUlWOelT7rfs+NW1FRra/OfGOOuBFE4BEe/2Re/Nn/WdiS
7E7B6Neec7rqaGLQtLKIPHdDIxV3lP0q6nnHuqIexuaVymnc7m+GQg9BhEsiewBMlzw1uNtFrsxU
USmPWe4G+oBtWDYKBtsuxEzC/E6Z6tCJwTCTxz5zYkbU3q1qVbR5u9VHqRKjrieZ5E52H+P/I6re
Pcd9VviS/WkSmpsP4QpWK4ZSgljFJULKRGadxBGLvbQBLd/qPYuQPpC7nc1PCw31WGDcNDEnU9TQ
1IGz4e8xAzyYTGRpNrRpfYxOr9GyK+tKYBqUTgxc3XFZOeodzazyLB/kzsDH0XIOiBrxWsKRJdpS
Xp47DT55okn5u1RZ3abABcGRx+DtjL6UXJZtOYu4b448qRwNjJTnP2YKA+Oq9lvxGfzEv43wQ7GJ
JmGA87CkCUONevjiraqXzFozrS0wAmZPvaZtDselHQpHR68B1hxEpAWYePaVDIifkzY88t93B/6o
BobPWqyLX2H9LxP6lQADmCHDpy5eidTDr6/tJkNse1J/Drcwp9HF8XcJgSiVrxdSsdTCo1Ec3hyR
H3myMtpMM6kPZqXMOiZ3E8Czat5uJO4YrYabKRW2UtCVHYl4s3C0kffyKhceCLkTJCHyXVlmWB90
euDlTVgoFkMX+nyDbEqO6zb3JRbVaIb3RiCAsuZ/w42r04tYlZaYRB2omN6ACnyJc16Zs5AYLgY7
bWhvYKZUpq2qlRqo3u+xsXn+gl3wBUyTdc3kVTATdE6+Rv4wWkyS9QllkWk+0jysrfVqUjEWCEAS
N6tCj8UL20qdQnM9fbO6Dkbish+hYoIQPKqyAKJZykVBalIQSDM0Bw7KdoP2SX0QcGwFOqDsaR3i
357Aq2dN7SygRroOvckCKwm4DHlwuQqI2WfkEecyI1v1iYHLbPsixHlhmJDswxlaQXjl3x71TPWF
BgsEimBu2cebufOzFni0gxdfxesqkcD0HKjrNZBj+fqVfqs/3eeqU4q5Owvng7+fDsBzISqvTga8
IFNn1S0/ANt2zMAy15xdYbswV4ay6Hjdtv+Ro8yYFoFMXYBJ2g7yZyIS9vGJVq7pbpNS0ZWNah4b
n+kOMHCg02GbfaVtsEqtXdsOS7r4I+MF8yajyA5ua+RRMofasnHOnMAiaLlGz8HJVBVSIF1/T1Be
Z9yzH1AsUX4SX1WNqXFsW7mH0GHK2vI3lOqL+cUiOm8sIk2jW4vhizIIPZQWMcd+rV3gAdUwQ1Mz
vkV33z2j6lI7uRvfEW/lM2rX4VPc/sFVSEfFgBEwJEdlK70ap84BvQA/L2xY50qhMuAYJRTH0rue
Dn4LPi94HrJQ12P/fyoDn/QmRR42z2CgGtmv5m4asu1GJVjxLPF6nWUNIR5xdCr10OVlru3XmT9B
amR9nJP/hUQKt1bsLtAAw+5weE/fuO/n5J0I9nqHmuo9nqnnpUaCj48bT0c1dP+1hbNqpfI0QUjc
oWImoePVolW0u3qK0bsP/SHbHBcLcVuXiXFcwWFTiXqLctpKx1ybMRizVYfJAgB/SG9dexFKd2Uu
jkELe9GIrErBMBz/yKV7JQlTsVCC3i+30FhBbuIpnPAhQyYRmNeK3zRjr2/UtqyGBNAZopDuUSIB
//ITQmvoAYDpnWQQr/LELAPgz1DOP09NSBkWj6/LZLwaa0L5H0mkEZ7EQ4HJsim2WMQuiFqwAyZh
ylbl8bf5dkuolAYmtR2+YuvIQBYTq+KpchWZv9dor1CQNVcJ0y7Gy6GybEjpbqReoLINEZZVHQJU
Xz0rNgKB4RrkGDAovKGl45GQwKTDAScuKSHuqWWiyDN+YibWyRLjL97wX2gEuzFJqjmNKGkK7WNl
4Cp/SH8+X+tyWsESsG2y1lmEnYSs1OkFSUfIBVTuImcB2pEmVLa2DRwHPP/IoPRHP6K56S5BGQNi
VkQ+PF8BWgKExxII9VvHKizgDzIoq8qH5VKrQ9m8iv1IHv28D8prY2QBKpAxV4OImDXbz/J/P8dy
8h7C5l4tYo8DPyrzUx5P20/yeqbiY1i7iV3QYB/f2u2RsxrT7Sj7b+BtyI/wPWvmb5TotbaNDtPD
bSHz1BFevhk4VmX+vId+AbXRwxJI64F1mYh/grwcNghdBTl4TrM6BsbNuMKuKHVfbecMAV5z/Ywg
yFzf6TqAlluWu5Q8swRx7vsPDhysGifeQDci+UCKF93+ztXGT/CnYa58+7G7v3rRV0YijgvvoJz8
ty5N4X5kvLf6FJHY7gTuYb7uJhtWHH/38jZO6qlsR1K9Wmvj+2+vg4t8q/gy4PlpNOq9Fd/qTQcX
S6t7BI1KTMQjcwIrL5jvrvu8mnrVfIcbhOioXBz5S1xsoQTksvQsISlQdbiZuE/A+GwvJwcZW7pq
sZVKOpL2n/73xiPnwSWmKO06YtxcXUZbNkKwa/eAXtjcyP8/0OFTL7PLoNMx2slCZma50AbUC4pX
DqgiJm79cvOJ1emAC7I4lK18S5nZH8dmrFkhyTvZkQ1MRPPLGpmogAlze9S8JagW++9Ft9pvSaIi
PfkWK8hqK0D2gvOvJpTZz5NhAdUi2B4w3q+/939iQ80hCAHNrSlvAIlzXQPtrRO0bajXQk8Rx9JQ
DP1Z4/AVU1Cfi6u9Q70XCdXExo6cIi3FHFppwLdUEsFcH03n7gOdhx2uKdm8D4y0b8eCITXPivkE
xaYVGrcj6dT/SahaiT4/8oATnang1LDkp3cEwryMBBMxID0kDnrPJckQAeruFFhhq84c64RtiJSU
N6b+YqeLCgiI38z2enPzbukrW3JzAgAsdxpcgg2FJA9eYoifPVcSZwwcViUezETmmOuSwsYut/gg
X626p0sT8krPvGsQ4jWWFraCNqVoYQ78SPTE+3grjA9Xg3dJYhwml3IUFv/MsdJoWm2NURXPnJql
+dHg13hisBBJ6JIG6jBXWPIRyoLG5RrMnczK3SXtTRfrrgIoIeL1fpK+ockTZaJJ2Zhi2Liw8mw8
Y5q5R3iNtxLp5JnZn5XjXcwSgtVsO9TOLTe0ecab8yqC5Ca8AP+eGw7Kgek1sWzPQwZwygbtBANw
n5NG2Hk8AD89/FCTI56R9Ap4ER4hknSLkK7QpkD/HHYpSXdlqOpGcVi1WdA+xpOsNNSTDhnYXRV3
fckv4+hR4zX1NmFAV9GpzQ8GTYOTpr58UbbDOGApvwLRSHm98zeSjXad/NA7+OBB9IXwZ8Xs5aOF
/C8pigjSAdr+srcFF5/lhfMmAqD6YEL8VyYsH/8y2bGvd/lcyXhkEF0L+f6boJx7bY3KWaBiezgW
8hUO1b01173mSkRfynN9jtIoNsUgpVEmeO9SDZFdx/f0L5bsZQMWrqlqGNTrjMgEKJeQVQSY/hxv
fVu1HXqgA98eILx03eYT7SQ43FD/+9hXr9DFFmYJPV3wWfYCoR3umLd1GeSg/xeeLiCkI47U8DST
zFNhx9vZ4H1jHRKPnEdkdygSIPdFBJJmcQOew2tA+vLuGHaVGj5fdf5Dm1wbGZyyS0kG1DhIZHRv
X8hcXLuNyOhc1Z7Wqlj/2GOJc4QLJWP0AxqGmxINWCW3CKtixQ2e1ZUlrx3E590XwNORNRkQvSFL
tDX+TH6NVw46Kw5Jbh81rCYNsmS4+g9Lx2TeSFy/v88JCk6nCT++PYMNBor6VTirIXj14WfGW7IW
PmBfnIIxt+O9MY8lWY+VPpeqwg8dsVHqO+pZNZeWGCDo8NLDPjZoNNgL7gkqGr1XDkbcRgr60QhL
IYWHJZJvYMvjrrVvWLAwHejhfPEkF8XNQu6geTgAP526eBDj9yc5pBL0rIpvFOTMZA0R27TRrwVQ
wKDqbt8EutgwPw7KTeih34+B/gut2HpP3Q0pRQ2gft94hWUtDZR1k8snDLvNVWobKUgwJHZgSKie
vIAI+hLANG7YlJlCBR0nAi869uXUZFbVlhj4S3iAB1XB9yZgwITrbGJmRd80qaeVsQ+KEs4wRiHf
3O8zqBX1mN9N+HUGtA/g8QZ33CBGCvPduHOo2/cRWxsFuHVgXGxaIVWrGWOvOzVqUM+9P5CmviUJ
GILfFznzHSwxD5gJADIpyXgXDrYBxdSifHk5uaT1C/78PtZAObEJMOl0syXdCjKvklOWJUn30rXa
4MP2+tBS73ECJyUUrOMUBt7Umut63j1a2lRtWH13Sc2Uodpa59AN82XvZklhqh9k9mWxaQR3CXNx
IzL6bYdWMb4wDbUUIbhPedCxBiDcXFDzISNr7dfykEuNw9BlMkrRc3yadzhukcx94cBfSrgxo5t6
S/8X5vOGFTrp2ST2ZmPPXIN8jupCGWosc6bk8+zurcgWnDk0kSXdWMSbTcPzGwfBjIZeFSFbAK6I
31Ay81kybsVQ1cHyco2bWwqtxNgqSJ4Uu7RYH+4iiAq+XBCWBOvqNiWFwtyvfRRSY00OmI62lmQ/
Vj06oAjbPWbNitOkB6V4YlRp/sLj0grL6NsUmMuLPqEWnjbHeWt03wg6nwFEiUvxPiuMjo2iEOWK
YmBHCWLx872+1EjQTErnN0YHmRua60OppMH6Hx99dk10Th+vF9V38e0f8W/yictfZQssJc4ZPqIe
BVrxBNDkb93qC5BV+LfNOyJZ/JYVSDV2cWXeSnjJg42thoDy8se890hJTneZaadGjOdqBdPetab7
48VKSidQlg7u3lNcP6t42pvG2KeVA/TBVgJfXPMJGt1PAltN7aOrkTID4QrxjBBFgeUK3TJhFiPa
9zxuVgBJ5jP/a3ROrppe3442nt5TrDgGvgSG4KLpajF8zBVRap0Vdsy0xw5di4wjHZxu1Rqa8KAp
5inE0R5Y7jZkgx/tjSjOydgL3tHNJv9ZTYVH7qzxU+kkfjrieSUFpiGcyqggWv5moHMM3Q4+7YJA
hvSrE1V1UQFwSMgLihzCsee3q9pbrnRZK6cRwYZJx5p7WWrMLG7JcL3Gl/951BJ1GOKUB/kLGbwf
HTBhGpZ7Hw18UjYo7+abgQZN2zgRvF0noCEB0uVMTyAhTPA/JN0zfxrhvd3kGCvBidMJEDyr6c4f
yr982i50mp53fakEEL5OKW4J6KLKtf1nriCidV/Mc+3L2RiJmiA/3tGnnLvNaVNSjzfsEjrWHAZR
Yv7ZPNb91zFHVN2zuz9GQbVBjgvNqEJT3XSKg/hY5RnOOV6xAu3LG3D4bo+5t7nJPwsijxO4q1/c
0ANnhjzLULSnprs4jNA+WNjUasX9/4rI6qgVT+8H6BN+0A37Grzs5pTDaVrxal8KM52e0FAmVtsZ
ohaCuU+xncZp0sQZDVU1jJCjMyPyto84UqlXzFSUB0Ygo9p3+BrGHmR1TXOEDX8b8vqvzM4gL4Cn
xZO1MqDNE86ozHZuL3a8qj0qdpag+mK2MxAHRn2/Znkz7N3LXTxBGdG9VjXoms35TTvnVvRx2U4E
PQUIvd+KTZiPr0L2mZK40gDWJqSUYboqcXpGDv5+9eTDmp9suG8WgdB6H1NRBOWas+IHX07nm/lR
5JYcTMvABOkENN+zXgGadwVP95wHSs1OuNLUmZmI0dWsVda2BbBkF8nn5L1zBq54wpnUFg4ZIkT5
cFq2Pn6P3ktqtkZD37TqBt4pEOCPqwp8WLScD8MpJjdBsQWzhMFrx+hpBKbATTwJA9M7algbHoos
rZZDmLPW23r5L2eW9AkQUaCqHpo2643BWfUrJBgNEBZIXfvUACsgMsKl6xoNDZk/w9fBi/NXaleG
9PcL2Q1bO60lvsnh66cJBt0Flo9nxg5Yi/aUV+cRIVObJhu5vqXl/q1QOPaeXFt+bbeQK07x1gib
akJmlshnwnXbVo+oAN5gRbYV1u7Sj/LrTWW61MIzJRwmWFPxLAlCvGHQxDn4W3F8Y/ZHrJ7NRf9F
GPpAKp+8rwH2iTPQ/O8BuZrM2JBgBehkK8ja8dUHfUABPdvlPCjE2QxDc9t12fNtBXkCQg23JR0Z
icGBTRbmmeoZtMQ/vtMBT5Ml8LgVxvP6AR6jikjjHCeWKXDXgzmNZn1GwUZYCc4lxEksXsju9fZM
YX9xrEl80NACYrlG3GjjpHYMU0qS+S8keZVnaaZGZJGKeMtrw/Wi6v16vil7C3l7elxfwaHX3ydW
gzOmW1epLvocqFYC050vDfdUiFPeuaSQsFTVu5pDNVJ2SXVViGvt1I6vSR+tsmJinVkKeQkZUiVB
mrXUlcczSN+4mdAPNZtr12Q2E8LsK2AcH9yrfTtvVVms5P38TBRZzl5E3Vb53lRRVCKtShnp363a
mZo1f70jGORDsRtLK5jxiNJymcwO1UrqrkP8aQbfliIwa3j5lJ23DWvcsCJ0isn+ro0QZEWYpUCS
sEuuS8QdTsjvxiDuKiAa0Lyo0k2FB3eHvzx/YxQuzKoC4WF0uvMua6jix7O+3I3ArMFEDnTUQnQX
vTV2h1pYXNSJL/EjCKFDArWDwgm/tmJqR6oZqcYimvRJhOgInMToo27NgNxTe/W2NhlD2FKw2Ep/
cIYG54De7bgj9rr+Zx0U8DWIKS0HOlZLAEPrZXvl0M3fsZtnGOFPpgLK6B4U5CPVkXHtKzxm8fbU
Jbp4lCuqaVgGOBgQotLVYIBEO7bP2YRrHGEoE2ORqcIV+GxOqKCjsCS86Yx9T4HMXWC3oUryqfTa
RuLfmNJBWvkSoiSR44DqA1razlxp+lvFBX6etrZvm5fy4exqjfVUOBAohhGY91/RjYeXnJMDZnhm
K2r6WxY8FuU5OFgBCMMolI3NASDq34fnIWtK3vTBK8w45up8J+efdg3ZTUWk2MaQA5g3mH1vXPHr
Tlb3fjV4o/GFKSJcuS60aDSnOBzjqDPgGw/iHOovDHlIB42e/sqS+sEdHtncR5ItMqEUtuQ0oFEH
lAflOJdQQkCwx0WWpJ5TOl6CDAA9wOj+G42FVWo1tdDcVUsAimId+DupcN2Rj5/0wqmz2o1HwvZX
i+1bWrUgpMBsFZG6msbNejetxA/4R+YeQQxVHk86erqtSevtGik1fKh+lsLjh1O3L4HXXbR9ztR4
RdFTVgg/RqMMNzd4g1F/rC+ySydSa+PJQC2r5pLFUZw997Ex8Jz9DpHmKG+IgGim3hQMwvvvk7hk
bkXL6LRn+xR0wIVOvDTzgD++s9uZUmExMY6eRLDX85JFtjsBGJcYu2P7X3SCmKr5S9UBiKGQ0eFd
IlAr3m1ep9sO0/0nbRxJ5gashe3QShj0csILslGaHrT6DDNozrihszoO66ami8vEsmZfzrlAi5H9
1QuKW108P92bKwhn8TdCFyqbu/Lpdd/RiAS9AGu1y7K1yAtNEWr0smUHWvvA5xpkZebfQAtRXzFW
JB/2gwyS8G8FPwRJatfc1qUc4CGStDphI66voitx1uyZMuCtjPre3j4DLDELcZoKXPLj9j2euc4L
A3B2Sed9LU2vLn4wN1QMQz9E//+BlzokQcOa1fjJD3UgZkFbSmIAhm7H7+nGtbfDoBqpColB3Bkr
Zo6a2dELpSemvTR4pnEU+XoIGL62UAXmBhRa/INCAHmP54R5htD0APjMM3aO7V8Kk/7jUlFW68Cz
yXlVwByaUv+Ugg07Ss1Wj0ilpW2E7NJvjK+Gq3RRxibtZMSBTgrelYGY83zlfS79CdHhBpQRs+F8
xjP/2KgT+hinAX5lb3rE/8i3dgGnDF4lNsarCmRU3mPD838YS3BdDyS1Y6VjSFUwMWR6bLDdBDzh
YKCX0wXvaH8WcRg6vv8Wsp78QpOYOKkxYdhuw02ewI/ulIy6yE17EJVhgbH+ofMBnCH+JMqwbz7k
WpTiADob6ipOfZL42NMzqapOminL+SwGu1ofBHmlrgt36X/fBOBvshXFgkGZmjLmSwCsIJh/XAl+
cfPgE08lfNDB20m3F/QBk6ktZCwkmeZgLluya6MzluHBtRGpRoqNmX30u5X0cia412GYK9L6ZF66
vTJxjfAa92Md1EpHZD6J5QZVgBv+oeqTs7cU+u3msfe5a+Dm4THq/i/AmXOwfRWHs7Q1M0+pajE/
0nvfaJnWr3LZCR+gaMsNFhB1bd9fNtZrJ56pR4EtSz8heqUIXFERaCNJyfpErGfvjBkLbCzHDB1I
EqRg7k/4SSHtJ0PDbQatCkHXeOpQ27A75Bml6CoHDglEnLBy4Tn39yalwztkFOsmPE8qF5UULAd/
fH38gwwqFzwu+l52l7rfSq9wTEWktPzxFtJfq0YndOLHpdtvPMXAm9+xw4vNsBtiOt3SixDa38Ta
nNSVC/3MFDsak4h3wCzK4rdheavgEPBcBdm0UiUhqZqWmMadCwfnKZc7oyfMA0WUItrne7CuouRV
Z6CUFdPw9yqb19OfdQiOsl+/xukFNrp1iFQd6OS61Vry1Ai9f50+ZgxI/AMUni6Ct5Y7KVkMNnKJ
69T4X+2dDAHB524koGtso5Vzha/6p9S8gp3fNHA1zeVPdN826ewpu81bfBsAZj/rQDi2bS8Lthah
XXRTdmCow2FdJ042Jtu9R3nsok+IP9VQ2VzIHMsX3NYA2XoLVh6aCUYnVo6/bEowm0gLkf9QBjX3
J6nPVY2P+Xdac0GkrDuuVoiH3YkxiLanTtFt4Yl+035ssyOrG5DVFZ6aQtVZYG+As5IORR2oedCo
nI1DRc2pYKh0KNj1aRAKQpzmZRO4tCicvu+AHXhDNZ0Gq46WmuT+AFWe/Cimv+V2zb5CY1mGWg6P
2FhR+lbooU63llYn7EoAWc2XRpyVp/VN7P5/UiuSEIG/aKje1P+d5fw7bLwg+nE5QOskbFKZAHSb
51ny3ZwQhXMGvJxl9qot/xf2t7sGoQqcm/zo7xKCeLvJopC9FIKF/ri+LrrvDm9HTE7MxGF5oimZ
+h6KA95dh3VCLBBul3mQWgS2pIFUOoZbYusXkr+quphHqzgGF4UuahIFCJumXBDp3ZGvBuXEEOAQ
2BttWg87w3ZfIaKfRJ+19gvy1SxVdwFsXjB5fmWcJsC9mFqNVzYu8GOBMVoa5uDcrdjjgcq6llh6
D4ev6ckzOY3Sgcgxeytu8j8YlN9Jo3uQAQANM+0QTQlSNGKRACxp/R8NDZ9/sPdRxAuSwwBDvX8D
cXLjryZTAc7k4AL4N9jAyNnoriVUA9F84TYdMdjozOwQjaVJgoxBxFVZZeJeCVt6qh5LoADY/ZY3
Vx8oJ8246p59lmEtINQLxFNV3xJiUzQ4EGpDl4nGkyiOi0G2rMj3Db2p7yb+nuTAMfHbDrzXfU0V
9i3uMpdc6G7Vy2u9hdZUnJy9/iYvh74WTgZIHcxC8JdqcL/0b7XJ8XaQuH+2TxmqB+gwBEhQhyIV
p3iwGh53bXLGBUGTrknJfa7jok45RRgiVoL7xqjGy42r719YzIP2B0uCxzKyqbJghXr5ycnq3lfA
2clucUkaFnEb/wJWx9BzKQaKlUdz0OrsvOK0KR1bkrW0hZgh+kUEgLMoZ6T+f6VrtLB1Rg7ET0aO
IrXE5F73DhkdhykxKfy9gAqKp8lHAVtZEYa8U2vmNZeX1eKsEs4OAQGsPLjBGkNN7UAAEu4uUS0r
e2MbJ8V/ayh2/+Xhn0DFRYFHS7vaQp20iSI6y69q+HLVTK1MQtBz4+tlgbxAa8HLkiS9VtSAKXnC
Xabswjz726+jkxcRPbE3BR0Ksz3/GnkRcNNAkyEi0f+55caWD8xNS2MetBjYgxrJxx3agiCyfCEd
rCXiYV8lAp5K1gKQ7MNU24wJA+aJH83Co7oRz90fmYbnryvvxFJJCNx+7Wxj4tqwPDxURP84Pcsj
LhGogHqH/1oVb9MAVLOiUyWVrOGTcPUX3gFu3e4K4IE4ez0lDecBxE/zVw2R6LlmlXdeSSJ0dK18
tDBGWSJGFLbb6rfhIlJgRVl/EGUMmPs3OozPnuoS8igX6v+xgo0HQATF9m0Rd+JGm0zM6N6iZpZd
0fG/j4Z1ls9UPMKZmuVOxuebFsvXBIIW6vK4znifwKCnC2cVEaUF9gd1FHP20Gtj6cBd/nYstzp3
0uJASfK9VQgdMjA8izwo+5Gc4C8Lumfmd1wdhu8jpYmwobp7wnNPtcMZ9u+lgb+947KkNb/KyAHx
i2ZxR/pix1nu/qbDjGIviqJiJZTSAv5SMtOotAlm/GunU4ohTx1CJWst6rYoLd5CrhmEOTSjX6c+
onrFnEdMso1u413cNlhXEs/GlixYvMHM5rNuuKqgRfjh1THzr5sM2IDjdT8BaPsCNYnzYWfM6KsG
CbPqjYQ2FXWgImHsoldUYGQZyXpsyDs95C6+VDz1JwEa8WrkQibJYm8srmrUiL/zanRZBJXcp/NE
g/obI7PuqjlgxgXobauCXglAk7oCx7Sm2WNUteQSYVPCqM4R7Cz88Mf4fvagTTM2QSrz2xgs9knz
hKnrdW7gmx3GlFmosehcbZLS7izxQhBc0jDdO/OCWnwUl2U7TM4juRC/dIBKCGKjUjvHk8sHJ8+2
TD7RfXJQ5Q5LFM4KdnGR4aKS9CNQK3ZK5yi8E2T4jQbSLi08PUHzCEEzeaf5uLCd+AZZ8lMpifRs
ZaPUAzgVqADq3CMa3pi+EZdM7rJ+3n+AVVgOmeJYN8208IVvcvQxH6fw7SJOLwhJ8dMTDDkN1zlq
+2g+N0OY0ppDp2QzhvwhdKpvGJmLHR0hgua3h4Zoy7Uqjjc60Z5zPXT4EUTGGC18byifZ6dX+Yfb
vFznAGs0FI5+8khjzxtFTBUvjohlmENf/4w5LqE/gSBjmfpdzDhexWcneFxY/FvQNd0fZ6+aNxj/
fHWlqs3ZAJZ83g2YYsfzzN5HKhb6aI4fhOLdYHxXE7JHa82oNNVOag9uxY2FG/6mXWKdaaNvPmqb
ZLpKDaIq5lG20b2YeyZjH1Pwm5Dhd0dcVvEQ3IkxrK2zV+GOXzidDk6xiqrerBhnvVbcmc1MP11K
f3r5sa9wY53BRiPm6x/AP484qmDz1Ylkhypz4yoc42/IhU0morCnFHBBhxNYD2JSd3kxHoWusRZ1
OVujj0b5810KiXErCf6KXRPZUkpSPkLG7uS9Ij13yBbU9pI0OaPGlHrmnUgtoOKJwYVLMF78Xs48
CNHz2IPNv5qnzjgMo0Z+fb19upqwfyiCqxOsc8gDi6x2C5nG8SgStPkJtRdjZVe8F3jfc+hfkp4S
WIyLId2WCupetriYwe4RFDIU8IG+wUeCMx1VThJoPpmoinyoho93/PuP/LbUEekrpHNQXCFKeAA4
C7PEHIYxBEKy0JXLDMqT7t8sVrMtZSIkoGLModra/qQ+FRtwyb4LnwP+BIB/eiRdWNr3p15RT40T
74Dgua+zIGCf+NL+27gL3tSy/S8i1w5gRbC8VzjKvzbV33E4HVHFmEMnafj4s37/dxh6yueXURqW
TujJ9yMFQj9JgSH6DgzldN5QNiel8SHOi9rEaasaPYjVdrU3i6kN7yk7sY+kYRyrXp8JZmcdVVAJ
Gw3Ds0i2XsgsWlpr+fyqJdfNpIvRSXhXalmwPd3QQ9WLYPXObCLTIrsD0bH+jszW2s5CweQGCexC
Luls8KlhsjT7sGqvBIiKc7iBumSo11uFh6Pd7uc05ztitzLBEe6CF7bPxN9UaxZyk92EUXIhM+AH
pEqrkgragPiUcmtjyI/L7UliDH6QkEwr+vS0G5IWW0xvWBLX1V7FYasQJqGS3xW4+CanRuFHcZ7u
/a7lDl/ShYrXMrqErN3bomSagDxSu2sUJEymqQmxXD+7bDJf/ywp2sq/0Hrvas3s4prGpwJ50TJk
J3NF6fRn2FYCZRqjgF8VvywyP3IUf+v7luN08tALHAkjO+DebzGidrJWqOseGGXzpZ7v2nbG18Yy
S89d/o/X3lKrgqprZcDynX04j1lxLx4yXhM/8ssfs8LcLIMudbb/KCa8QzfG2UcOjDJ/gWlpSE+4
C9qDmrn7XK2toY3F5AlHZvCOOikWfQn/kp0TdSRqkn1qzmqMtiBXC4QIm+M75aVY6C18t0G3A/N9
ELJzbsnRosE9HKGCcuNaPssvg6b5M2SDPL/Z8Ir7k1fU2g12G9icBF0j7iJenYM76eDjQY7wnMg+
c/kWr1zy08WvFFttwt4nncm0e4pVBxMLJ4Dp/nuMF51qEzTPJ0xnX4gos8URCpH83pit6I5DtOU4
aPyHiCxiHsVU7/CgAm9+8RF6NAVKSspybiqOWBInP4NnAVcqsnqBRruMviNkw+ipJtkQk8SGsocW
WJT3AuGjCI4sVx0LYYUVZNCzCTB4iSq1tPreckI/T+wgCV0ZjBTdQZDI37PevwEVZ8mbBVJc4nUl
sPHMhnUQtw2XxzU8yr44paUlsOYBJkz7wdlGQHPcgsZLpQWmRj5sho2Fp9/Fc8FryZNk8XqOJklm
A2Jm624XaUMXb0z9FY0eAlVA2Jtg1JeiDV1Xu7revcns2ILpbeL55Qy4m+mosHFDbxMb2QOj/2If
NiJJ4nEET/aQveY4B2fak7XWUVsrw58MFexf+HLr7GDLc9vep5Y64XzujebI4u4aSqm8bmHCqu/e
mznnLRxcXp0UJhSkmh/A0IlqI+df3eOdZGU1M0Tt0VfQFPgzpPjiW7W9AM9i81dyaK7Y95iaiF0f
CwfiBoVPPvq4h4eN0C7EeXT4OS8HFZFT1DOWD9D501145gHdkzdfARKxPGcm2HqFzveJNuVWq3g+
2j7rnSMHGI38Ofd9Ie5pVorVwQq0l/sdxzaabpi0+qyYWegD/cMde7eGKJwnCOKeQfcOp7EcjEkZ
7fdbA1AKGAHfgVwkHpOyJbZQl9Z+PZzzPjraYgoAUYr0dDHliEUdi3nR5wGHd6UZcNWsvBtrYPXm
io//b791vc0yQhi7Hoa8TLg+IELK5qRNUYJUiKG9X1YXdoLV7kFWjySZlkU/sfB6e5a4EC2x4u0r
i/FgPDEuVNg1Ug7Ask5rX7spH/s+9tUJhf+AkrA09c1ISSawWvrA/6N2hjAnE0WDlp7SH/qEvGZV
ZOonUYaUzQsKOW2g8x3nkA24iAZXsDO/O+Aqh4y/+3HgD39TvZGe8npNTaZFzMjeaeQh9XjaedQu
Orx3a1v4LlalQO/DlOxySVcd4LES6pedsaDMN6ko7hFSGJeUNXquwbGLD2UOY6EUfKAtJlbwckdj
QMIChcYwBeaXZ8Q569oBcEqzzK277E4KsLAIse4N3SXCc9xZI+g/3cGfIKavapTRb082uR/iFh03
X2Ir2zhvEqVU3sDo8nbeK6sDshB72HCne8ELDaKDIV3juXZ0GnhesG/RN1/OlG+r/Ke8pXrq5HNu
APMlo+wGd3edACIGIbWUw4mDGKzZ4RTVJWZAMIl/QsSrHvwjwPwSrj02cl2WSOmjd4DKd1ZmFOEe
yxR8dL9EMZ7mjk1ok4hAkAszgQYC0HxaYWyb8zpXhWxVJvqC+Fq/rsFO3DLpqHCy60Ch0QreGuj9
FdfCAJbea85MAx7HJa/IcTmBQm6jvLrNPBFS+2npsmHXtCKwI0aPG5/J2/YI1mR1N0SvJBG4P71b
vYcVFLcrOwjoTgz8iEWPxkS2g/EawcpFAG4GzPYfGuJpWWr/DLWDiLzl6d1buL+6jjQG3ljUYOXf
wkkrdBR1jAXLXCHbpQ8/QS32TFbQ2zQG2D5aq6F8jHzDuCIZczfJ6y4uqlTFqRR1RDAR+ge2Zmnn
z9lxUw+Q1Ey1NSWW7hTjzqqmvo0IyHrHFAPa9ZQjILYjAaxKU+ZADSk4b2pUgR5S2ANsf79WF93T
meaWTfT8NP5xZsIzQwsgupW2hqwowN2xZIVz3Qs8me4fLUKX9/cAD/hKWxb6BRF3mZwEwwHlR7nt
NZ1ev9UuxDrAwS99tWu5HxHM9p8jQKAd6b4RllFkU0AfklZmqAGWKY34tNcjBbIxfVyTWtQ8wanV
eO5lrjsM/aAb+4eU/29CxriEHJl+MiTlqTfRg1b3Mf43ndWJd3qfwhRkoROY0kegJNcZ7/JVyTMH
DWDdph3iUtQ77UEA3d95Xn2pwfPUVinRuvGZAtZJm7X6W7Kpy6iYR06LKFxgGoZCvUNmwYzgVGe3
d3g7mQOqIYLRchP+xzYoMeAW14NhPyLQ6BDgPchvgDi2CV9ckSBU3iE9tghOrizMmgGDH1FHprM4
+WWd/c6HtQK/T0+4V6V0J+T8Qk4AjzP6JjN2yhjlBFXByg3zlpKo4Vkz0WFNAwfmOmbj2unOPhsC
0wujm9RxtA35+AlwEI9XHNl1T0soIiuiQyrMt0vA+jffDh7c9oHCEUnV5de0LVhaR7L/KqmiqdqS
IoZzONE6r80nbOi1G+cOE9lyE0oJozs3njHsnlL1Dw3yLVy9iYfGwMA3GsBRkPhUuarWVK+SmdvB
MSbZiyO3sIqEKwOX9s7pw9zzf2ViO85jArCyf2rrNeTm/awUj9BEOgLQ224LhdlqBCZavKkEXG8o
3PeWfOpBtfgNJL6regcYdKO1y38s36CIzPE7LBnfUTkyyf+YXdyK3fxuDsVYxOmDl0zKP246/knR
knPIFRzdVRS6kAEtNlPb4RDIoOmwDmxgYaQscpkBc+mfBRGW9TSufwIapVLcgHS8NxyVBuIkyWb8
7XXeaGoWJjXuOXkIoJyZ6J00xTGXUwBMHhZel1CXOnOpVkO3r1OcG7njv/jQDNF0U7/p2R60xQ2U
jzC1Moz+znMkFUTVRNs5aLjq+d57yWeihA7hrVf2jOfGyK541S+mOahgBEVdWnj8ns1I6YNpq2vF
yaHSyarKcEnf4qh2PsoBWV2YOmxhEHaSkgwDuJBuTqgl7GdVKx+4J+cj38HnJObFuLVucqwolTIa
CyNHcN3ni6cAdUSD9b0VxV1m2f7k+b2l6GycO2H/PB5HFBvdPI2y3PjOZq0LSE2scPjXfk7Ibs3I
2lTIafxmO5DmneLHkd+zNIAjsRXq/3QXi98KGNRZ5QfdCZ0hynxtDcrZCcrC+hp/c2GER7WbUsyI
6S9GT2aVkzDt22Dpg/3R59K+CzAIaJreUjTK1NknWxYbAwQGABEJ44tFCcMYd6W4AoiVV8S8VlAZ
J3RgcwsrZjwqHHBbwH0C1+U1y6Dfc7NQ9+vgwn6VB6oeKNg9ufM63SrohPYY8eNSSV3C6bPbhfxG
HtfVCdwNeU8Fxi+kTOe8zAP2fnj38UzPXq9z4yRzR+BoOKkAGQUM5uAhusQihO6uiC1feWERBEmD
+5FHComkCo/E+5TlgzEzJUX51E7TpQjo2VbBDBExYmBvdhQo+Hpmbk/09+8q9NlE3xMSElhkEOFT
gr7IHE6aWeyXo4XlUGpTgzVBJXe2vxSSb2EIkqHCilnd2PdbyinhtbG/TnH+bd8+Ni/rDMEVzbK1
s4aP2/2qGs4Ckp4LjGuEldaTHBE2wdcwD19w5n+5SDOdvMMGy0EXbKXxa+a/ciYoCdy203XAsu10
BhFybqm4RykJf2KuK1CoRAvMtpZC/MMPJ3Ft3T2tDCTJ2a8gg26rAHBs5jaTHsdpudevubKWP7ko
JN3v5WbRaGr2X2jbu2OsLpsK7kSox0Fan4sGQJNHEa1dgR3RauOgFkg/wvOKGEqqRWsShXg6jlPJ
KwkKwFhoWbsY2TSaVtcCEtdxxBLRSXXkSY6cVmWVni6Jx8b/bkWQLaOPDm+Jr0cDMmRSI0cHeTUv
oORRNZkyC1fDJjdEykcw7s7ORj4wWTCWhVmeh8jQHf6iNAP7FA6MCtSMd1z1CfwAk1oyFpNB62qM
MtH2+/Jq8iXpi3skGieem4gWcwRbDix+iJOZdeLRUCPbezA3ssrfeYr/eivhjq5fycLpvw1DWpiP
LrrCAbz/c/HhzgLBGBYAVD4Eqtbtv6Ybr8J3PJ8OcQvXU6RiOac/KSpmd0+cDHt/+FEXSL+6KnGw
KRZ+l/pPkimkWUV/hrl57WMHlCdkTb98AeshxS2Kpwa5+QYVrE9TyKlLTDPfpdG9CF+Egj/NnJYK
JkKsJJeHmlLIiXF3RmUSCX0IAsDc1hUEoGQmgE/nlapeXIx8x9P+lfv3hemoyr5+pYv84/uaaPMh
F4IZJfcJCwrgATdR1g9Uhnrl24RPltm1pSCk4iqzzfoALRjjZ5DnQJbJDxPHgpgqL3eRIdmJtVGP
q34Tk5z2FBQD6iaAr2POxctOlsENX3VTDArddtgeswb2kvvNS7G6rZ0ben4TZc67m7R85Bte8vHV
mAG/cVfAc7X/ygkkt/QcNXCnENhyOfXLu2zeY5PWs9r7qyV0XV5Gke0l0vOEir+Fj5PDGJIUZlA6
kKrGcvHjv3XrPY5S4kIFTyTlH3S51R7B06Ah0EaBdZJtFrO88eg/uvcR9bp2RIG9su7RX6rghvhX
Ek16rcoFCnCAaJycp1Q8vAswmtdXZ/NzpHNumLA9nb/+tTvwMKFO2sOdU27JlSmC0icLywIFSdMm
jb87nOQACMvbIO7WmHWmr9WQ+T36JHHDudTxx6+Ceoc1VgWKOi3I2/vyoPrw/Ic0RNyuyP2A09wo
xcG67i+Qf1PnLa2phf631wqAq2O4uZP1aEWRkgBwHBxvgMMrcvf7wPqJ8VU1t1GjP/n66DpREZdf
y40Vzx57zH3qYZPKEAWmsx2EG0TTsw8YwuNI/YUsmifdq8vrb04De8G0pvivv68rDBwHHL+PL903
tMc5JXNx315E+cysZOGLRswaVctB7TE1NbzNH2UmFbphC/9P2DJ1oaiXwU8DP0tDp8f3l0hdC2Cb
DKc2E/idi1lJ4pw11xJPp/cFTo1Kfu9QTmHsqrjJlGu3FqVQB8QXomR6VmouY4lpipfvYqa6P6p6
krOebFyxXPHBN9oeCsVR6DINuQeUADPq2C72NVpW0w5W0L3NOzns2W0vvVu+7GAaMTNqvHrGfFJF
gco9nAb4eEmaBvDvqF18iV0987ZsEq+gtks7tjgo1SRZto98MTucjObkfUav2WPXyfizn9E6/Bu3
wsWiZhwZzW0LvLJy2sb/tB3ujsYmhdBM32bmMKychcsg5tVeWJT5n9ypbiSX0bwGPa5B2A8OIouU
QXgz/XXqJjtpgTVyCxu2qkVunEhQ+1QplNmPSd64MrjeMnH21PXCzS32FTJTXW+e+hn+U/XowTky
P2CYEScNCF2jYQuieSM8TaiUWXRvObTHY66ozA+R7zsx2eyM9DOHKNx9SCpQGF+t6Qc3MwsVT9x7
DfO1bfr5t4zLsjYU01jgd23ANBJlnj9lwQEj9JR2zf6GRsFUgQ7v+JjIsUpG4bwoGEJORDDubcfR
N0UIDQ4/GqJNuKxoQn2b/KWYyJMec3kE8YIr/rIBRNoOG1NRk9aiIrAUms/EUMLgfH1fvnYEGVz+
PIpmCtZdQwKcyzmjqFyXEdCaFHtL7EeitjmZ4tNt6nXoZx0tBdqPtxxyvDEQmkdcYGFKr8QVC9Yo
wRU145ZrrT1Cmbibx02B/9bDuOG7Ct4JyEt8N46od1TWfli4pVJxJjG4AoS3iWefehszh4NkNwIL
FZXc6p+ZW7axtUEaI0AN6M7FqqJ0URFJVptDyQntyuXmQgrdIZp6/d64G5Re+bFArR2lXnPhe+VQ
7f+wfz8pZcaDDp+8mj3+ihKMV8KGW9Sgyb5mw3l+Z//l5qFiXdUMWtJTRgP1R0toRsZwMo7rHP9a
LUMWaY2Cy/SB9dSJxGO3fXPTf7tJu8JUBT+sABtw5Vf8nO8gaYK5LwF2+Duus4JZjRtDPYrcpBqc
IDn58gwLRwiM6TBqmjsZ4osWMS+9NyUWE8kepMp4TR5fH7wrdqCPwncgwIaGPR1206LTGcqCefTg
ZtFe2UXBFnLjIKFcVzWkP4pQUuC9roE7ljMzmBwjmB1EajsmO+zcwEZr5vCCJmThYTVb8nXiNlpH
m84uLRNArTl3h5fvW4PT9Qluz2xLjDQrhyLivI+X7fbTgISciN/bA66q9QYQ4J6SGIa572uOoH5L
+g8yf4Y3f2332ZT5vN4A6IyEtQWJfaCPHPRVHP+D8udnxAedF2RTPFv4396z4Wj1DGHTgQ6OcK6Y
aOW4g/UBjkD32KtgoiMVcE95UQYTcVfuJf1LsAMvdOBkBYs5SsaKj2Kv5FQ8jHfxmKxPOdi5pkCC
oKOBw4JQQEroNAXsYNbsAjVgOliW0MdiI8WtgkB7u5hl+S+C/T3FmhHv1X+ynpgrgwA0/wflbeA9
v/jxlyDO1Etnir056j+EhFmNZ6HFl29xYjNqnSr91rvG/AbeLK/QYoIvThLEcZWfjCvz+BLryniw
32A5PpQrA2CiybfjzgnLDhQpiKQrtyuyK0kntdS7s2QClAZVp9crFUk8I5eforwSV36l/n+qk+IJ
MOvnYgzTZmTccCF8PHy8CXhD2yTi8cYy0UjFG+jO4xEMRJpjtXwnm+T0TUTC3rlUXXnlakOP1xwO
58JkT+LRxI3G6HWunnRP1pwLpXGbWaW2o2BV/VgSkwFZQKBp6G4YUIPBX1k7fd8hsgwEG+Om9pux
tGRSw99vmhf2k7h6QQC46KZb2jcQwj1OZTwUVgJIqjpaQI38YBeZ46f+MoZ7pZDxzIOh14o/5JVO
Pzp30CBqHL75sg7C4a2WZc8jcde9EA5KdDaTajmcmVqRl8nh41Y+VmyeEiqwXwOe34ePKa5WVcnA
BOsALXI3UOACtFUidRRxqaHyWZLJ4YKPKbcNme0OjgxUrWJb6yhoEuzZd4Tf32Wti1TZc2VV4qbY
SWd6XPxQfhe+GX8UpE0kDP0ZB+PfKptlSrjInZBYqeTs88uRYCC13M1iyAEMn0CzGkUILPdZGS9J
2FTM9NJPR1karLroRb8XQQhRLpASj2NJF/jU5O4zH7y3mFZ18RI3c7hmCOWKHB8FDiTgmirKHT3n
5sl4/dn4Lk1xxj0S8iOUwHV+TQT4H3xeaNNQ79TzHPUy55VZESfDgAvfDUKA54mg4T2/Wwi1ztxS
3ByX0jVHn3quv7dPaSCD8PmzhcJQ8KNfTEr6gS8qc/PAtZg9QwJDqnW22BsyG6TXmuwZp3x8kcfL
2pKsXQ3gwQ8OgE6qKpEdNvGCBB0pI+JmQ1vJTOY7OE+Xafrz0jZhKtxGsWIkzkK1eX3FZ5qdl5vN
kDDWuou7jvLk36T2TWLFo6wlS3GJYA5zq4pc95yiomOned6grY5AUjUizDoNUnzECdqh+MwUvP8x
bySLgLWdIStl9zjjRgwtl8hXdj/8EOU96uR81Na99GfJY4tdj3Hb2FexUvlW2lYfIOqLLARbflFW
QN3/c5o2RQZ80/qxKcDswIkw1dTuHX5HUQE0dj8iJM/INZ+0g/FjQZfgkaCZNsEtQwMCfZmHtylo
/9xZybA026jftrU+9bqccwxFr3WFNXTAtpOBPj5M8SAvkORljJTGDukAmH0tCd3L7GdVGht0rLZv
lg0ieZXPg+hVRI9Rhs3I1MJ+KOG+DAFVRI3WvnRJhaioIRDtGUe5nwPi2vQASLxXE3IUGA8CzDXi
xyDNXeZ/By5sJZpsxMJUqaif5LlECzMLlL//Ig2RLO7Aa7IhB42RFtTHc+ACCjVESOA44rp0hIEU
oJxL0oot7bTkmQcOuP8FlxP9846rqtbzb7bUH0MSkcMlF8VG8mwwFsdt1bXWQYwA4d+duwTw6Wdj
MXiHGn+0WZRR+x3Rl+TV0dpVR7msSno8SsGWliUP+KMOn3RQYunFBf3im3P3DXh9976kkiCZNphu
JQnF782rsWns+A2irBosfGxFtVQABfpjLvaCmOo1cYSS1l+ocaT/AfPz9eJPGaHLK5RpsghwoCLg
CQt7OZ0K5QsVNtbtEkFFMyuBBg1NczPPGEoWvVm858QBM7GVRdXw1z6xb4iST+eECnuF6lRxX3Nu
kl6TFFQ86U3NC13Q5wf2+JQdt46LYWyxj3jUQmbiMae1badU6JXspX5auDsFmXqdYCRHIBYUrnyF
Mef8ma3ycr+zakmQGDQruzPSzLEyDoD/T6BtKmw/YVvCl7f6shDRSVRBk+GF+jIdBqwOsGRCKZrM
WeAoN+bdUskd6/GICzu0YjsvjXyoLomiLZRHPqZRJ3/AxT4CqBlotvuzxvXfAuhmCAyPSGPnyqxX
fwBp4brUbaKofIrWt5A9tIIv0LQm36au8qJMXnGByYKfVda55xRp8XU9s1E7d57P5JqOYRgT6vCT
BLGyAHb79xLkdOs9XIz5ZmX2ucA7Kk4Km6Nyaq1LingBUYAAD4hitA1MS13QHcjpnfDbs3ShNRW6
+4iWABfk56jJFp776NJ3BQk7RjfE7qPKShDXK2dinAk7KKyy4xjEsLrpNKdqKPV4vtxSHj4SQzMu
lAMzolb/6IOnkm9zSPOSlmio8LQo/ydrZOD+iVcEb62O+KoTsuKgqM8CIjURq14YaQnbazm1tERF
X5o3AJMiqyOilnM9PCXP3jLaIXxZ8WBUmu+H0bcYxWpRKr6KrtlBlH2uV2FYrPUzGmwbjhDWYJpA
htaWTxsf9CSxr8qq+UKlFEOAb2H4ndgb/HhrYQa3mO2kB5OKpKupwophuePBrG5LVRUkRJWwiCFc
nqLBDgFG3kwz5geGAJoWvmne0EDizNOjf/yCSa9keRJ7UBBcwipt/6RCd3oy86gVeSNEYGXOUuRp
WemzNopPLyDLOe0aOHzpYwaulw7cIPaQK50CBcevv4tPSNAS2sJGTL4QoIUaInWIlKJ/wvKj4nZD
Si4Lbdx0BhZH2dPt6UbR7vtPxak9H0iwGXltHRoRd19KALYcg9LrmR1ccyR77bWSFdylMr0fHwJB
9GqTXf/BMA+2e+Q+TekRxTD0mF5k8kDnfnsS0BTgx5b7NyTtrfBsjXydkPIVlJ+iZ2Gd03+/lQ33
LIDHVLZd+cJ1EIsAR31jmamPvbhjeMtW8ofBw9YrmVK/SupIl7vVpzqWbsXnxR3ee+LX8ETGCjZU
8zVt+9X5U70C3W51gGqqL+kLmb45kc2pFrIyCHbtWsCruYTfCTJ7moHZ7br2Sg+Cvot6BOXqJPZ2
94Ftl8j4FqGYqlDWfUEgCFV04AvkjuhzhKtkuE6eFYUIxPfidacDC5N8012SjIrEtNMHOjE7/bh8
EPuvsO7sQSkLyDsZdCZB3/CMJ/DColGwb40jptfI0JBy23XByTS+IHVzFBPxITejHIHXwDgmbQrA
F3GhEgRIpNiQINrkm7aNZ5lObCJLP/TJHFFj/bRYPPhJTGbf0Rltc5xBhQOWDWaQ2lTnWf8Ghgye
hHQGKJ3sSjmxXmOfbkRcvk91MBM0dCSz/QoSouvEFsg0UEnhnr89XFLSR2W/s/u8893BzdMKiDfE
U/v75sxLYr6LW9NrS7JMgri+i2zpWnVb8B2PcHQkqtl2A2FXfTGfguAOSFMNDBsYfesEKOkj+V7o
/g6A2En6diGsoPrgivar/XNHzRc1XbKXg9ZexqCUNqoyyNQJzB4BL/+DUpT6EhP4z+9otgKBG72s
GzR1Iuycxux2YxgFy9UsEJQmmepc1DcI8CxOQkBpVg5jqQGOdjd8zBPkHUqNfLTyoQUGtGEdV3hk
Io0i1HRMsO7TktNWcwnMVusLEqDKZftoN+9ebtyJwWZ1/hgJx11upnm2PbZf5VntNNg5OHjkZmqC
iFfD4SMWDJxZqDNCv+0kwGHSD/tkP4kq+DV8ETFJTIxkLHc4c/dXw3FosBnyDY0DT9kayfg4BTd9
i/RUwFIVUlDcH38Vdw9YnLv3LMtmFcxre8AJlpgZ/NqaYhJsTFMnufliPoNECBd62FA5KVOBjMmL
O2+hiSr3/24sP15oYwuyhN3JTm6As5nkpsomTYD3y5R7P4Esv+CC4hnCohFd9BIxG/yw5J2ZTrFw
MNN+lNF5TYiBqtDgr2LNPLvLxXUw9G+blzRwTvDx819LM7EampwZ9NWEl+xOi/P035fZmWxtesZj
mQJW3Nxv3WTnZ+vVRjxAXULG9fu6uNqJU934iLwqwNI2bfuUpoYRQidcn2rPUiEkg6VjIsj0fB8B
ZCzQ4IIg0Womi3G2HdyCCpOuhilsOlEPqlukOTdzQHHrG0uO8ecPvzjqvF9uNwEl6jqaulHYQU1K
9XV6yXPDOmwPfB0Zo1zJ6D0I8nfF1D1R5s6Q3Zd6SgT8aUyhTI5CC6+xMYTTv/9ekoJDAFCbA/uD
HoWuulp4HJ3pcAUdr27uhj5ENsXp2Kbn02jrZ4by0a9Po9t44ywtbzZhRniPfqjeH70eNiXz56Ob
KXksAHrlG1M8HCVPRag235YFs0ayV+4I3UuLsDtPfblpy/hC6kus1L/IKqPlf5ZmM4c9FbWLGELb
uWi4kAisk6lW+ahTvd7r7Tf+PdQKex+dfdHwHP/zkhdQucTSyYIcst3E8yTGIzjOE4vGOLzJusuz
yhMr4Y64SuFsrjI2xp96HQQFWAHr4cOVQcahoeoovb0ECqiHdTJsi2oq8TM6KXxQo7o6ZuLnCznK
ELnZmWYXyLYTeRWieIdZtvdI+d4kgWNU7dZ6mykIhRLW4bF15qY8qf6btRXGo7GYLqvs7O8z9pwt
V40DzVwEamgEYB810V+OsgmZL1xfwyiZTigTqx8nTUPbhkV2ShWZPpVttwh8slQ8VPN9mBNQ/vOv
R1BEaP6hMJOM7AfEecohOqwBML030jcuMq5RnX0V7vj40+iIEhTu9iHeeSpICFWrDOjep8QZjrpa
hHlIjfI+owch7Vog51+9vWb0sOL7Orq1AZYjr/1KvnmLMw60pKwDYdaJ/sKFdfQn0YEowoMv0xIx
DSgnP1i2ON+jMr3iJulWniAdOydzF/gIkig0xFUITWLZUgLZ194EPlh2sDr0KYCMyN5ggpAlyxsT
5UnzNNpjmWwWbSQSIJ2iUQb277YYMS7RLJVbtPFmP47aTPDuVBVwj0Ck8DRhgZWnv1i6EEp6AmuO
Jzr8GZsXfNR05PvOy5MJ5lgXPP2+VDlcylLqXK/LsGBo1Wgwmch1S2s5sYMBLuOkorkNOMdDrBfK
HxbflZAcbBs5FT26R4bA/uhPjlAPSc3xyyPftPtyD8xrqBbvXNlKrQNrp6x6JYGSMOwSwtEE02K6
qvtEbvyoFocRdsnf1HPMJXkzwtFj8a+iyKPX0xfSumEw84YcAkzOwaLzia/azs2oSshV8Diy+arb
IXW/Kq8xhi/8XjnHLZw0/e4PFcTiL/+DBNkakN2U5C455FvoOs7TG0Mrlzz460dSjQumertrMRRS
+rE8WA0T1PA9WsCE4m2WR6V90xU0Msg/ynlerdkZrRkZznl2tLcjw3D9N7xfM0WHjstnq1J9sa67
Ja94heJfL36Z/kHXAMmExfCy6YfznoFISwwWe0ZFDx3DosX1C4PVL3x/H5igav74rh2Jx6XgNR6h
Q9uX4JgCRCfDzo4pn8VUI/6+l7x8ihZb0clmsPnGF7CJyqBGr3Jt3umpoyGRC8MKxKyVCyo6ycRf
mKRcAcgXsXrgtOkaz9wijyxFiaOlXIhFB7r/eMSaAbMOsyoReKTXfv7lkukwQUBkcOclCL2aaKLB
UIUb9P0cRul+L9XpPyVQ1rJK51YITfCSGS3ihhTczrukj2RdCFlH/uvcAinmc2JLUBeFo0LC/Qz4
J0W7M0SgD19H5dKuV2l/oOFr5kvCsklvrlHfhZ/tCJm98ZkhTxwtDSnHOJolkERN6aHBvTsELDHX
QRGlo8lFerZRaFj9xGa/L7FlUkhQKkqeVwakJDsvFeE/qsngAUpPhylBBLoTLJie7UTOUCYUyLis
dqONGZUqEn+wrNp/WkKPS4Kqh2Tf1oQDsbIQG5iUVeyoqyw0Wmxw+DxZ8oLuzqeFWGa+qaUm7p/z
1og+nsFHtDKuGCA5EF2T6H+gC501fQFBAgn9lVLmdIPl+CIy4td6V3ljRXzHVp+ZDeTuyqY3zWAl
n/BAHP5ncd2SJqEPqsTDA/si+/ORXC5VyTN4J6lZMG+g+TwQARioJ06JkJfrNxYdF3WBaCa0KCrz
tW4qO0FyvaKUxT0ntdlfgwYo9lQRrmg1opbaeNnQGY5kgnsNtEPpvWtJXeoK5U5RjoMZ6qd59xvZ
IEfWBypJjr/3F3rf+k5PfTDFUnI3ICjbLRt3TWtgbo0GBKZMoh6vjn8qolXR09gQKifMRJtTvjXV
zkwb4JMFPN05OCUw5sEyENwEsThnAAo4OjDQKK/ENjA2lYWz1ydMS4o7DiJ3c6h7MZqDjoDVqcfc
dDr3RgY6ou8W3NBzO9Q/8zlkeJd3cAhMn/DHpeI+WU9dMjaNTHqtdukuJgoLQv+yudmUmKJODY/E
5L2n1vYCbjOy2dtEIRDKZ8Vh8EzFmoEc7VhbEHgJTKaGt9etzfj8zMeDgixxUNA/eeVrFYuyVxwm
7O4E/twdWSTXRC3xwbuPmx8AbzR06k/+hkgiEB6Dj17eQNSBau24O7c8ZRrOcm0Ao16BxXuPeZAF
quFPRGLzoP7LMZ4TYANx0/aBYXgUELs9O36PzQqDWUBbLCcMubpnW3NKkxexA5WxlWGV6zsMMwjO
zLgMtdGA3L0Dr4n3owhnkm9CfCT76ae7mom1uUZkwB7XI3ghpMIDH7hsGSMU+oWeWxlQd6Cdh92f
t8NeyTIV4tgvto7lkUXyStkzzbnzw43RfmokrmrAgjUqd9I77WEW30phakAnvlw8vHoJ5ilmu0Ys
lctXLuz6c+AzlgKmn12+MBGzjNyXL9HT+thOyJ9T+a0ZHHydUTDDl5tuPQBoeHkVHlwGwXtiG24k
FPaRG+BRyLlhJCMqSXQ5ATU2WlcpcQh8gTYuBxeGZi0P/V+IjdRmvnd5WHADnZhrW8sA8mYyWAL6
Jo63hNah/kDPVDJCPXTibRHzPgtaMq/zJk5Oaxcgy2tl97De1f0yrrUAIviyA3O5+ymvZoA7XKIJ
sM5RsNv4yxmgDain5S8JknHzBtU66Jb5LoNXuAKldxJHLVzGix+bSO6XjXrPwYP9pkcJHzqa/ECF
2eAkONJLbMaKayAC80HPILz6jXow/Mws3h70PdqClOm/j2M4FHwyhzm/hFptqmpBka++aE/tTF4z
4AanqIz0bugM5c+XkNRD36lcH/Yd7NGTm0Ve13HuR3TSfP8t/1Ici8VGCN7qJ3KiqLahIZGE6BpC
8DBSJsoIKNycACcpDTNPpuXXWlclT3PHHXEwN8dkSQ9JVdO4E8v6Nr/E7qVcR8mwnby5kJu1I+OM
LPLeiED+n7gYW1JvycFcNUbV/MTLK6d60VNLXgfdJarhcY1gdAcsHO4DwJT/DhO75GbSg75MPzsT
JvKU5fEM5+ZwCrFhnibtsebuyENC17AuO02b48ihqfNxJ08zAVSLltReDy5F4jaPm8WUo+1WNg5f
11CVz03a5n33qS5K0IUEKVY1DkMF3POCIzmLx5bfv/ZWGL5PmuTD+Qk3Ve2BlzTYpDYJf75VbbAV
GcjEhRccudzmopqUVnfUU6g8Hm3FVj9CghQfnHfXyWe+ZnwSs89T53vaDYstL8Pt0L/iH1YbO6NG
U9Ijf7nuKWFY4gC1O6olxOzR7wBDkYh/PB8Sz2zT3WinBMr51+7Q796TzGwo+T+omP79hYGJCm28
L026miXBg5yDT0Z7Oh6D93bsGjaDmBNNN6zX9Y8OXYF/fOtLx+PEbyNSVYxBiiw70dKaq8iDJ6F+
PAZx774rD5Ut5+jPcQt7kpaE+o0uU1MYv+Q0iJJvXlf3YCy7Bbv6NVIgnSxiaIzWYhYF4LJxtnaD
Rgwn6BF+tLcSQqMqnD9v5bReKgNxQqxJHG1qsz8Sd4GrU/Cxs9K3KvU3A01K3HrVlBT17/4FRao9
dqRgZ9GMB+OJ0kuMNDdRqNHxKI113UeGmy0hQ/fGkvnBf9iGPZKsXsU32YO6tN75UGly2dZKenKX
bXifUT8aDpnFvjOHBs6aKXviFGm8nb8B9r0PivkL2gJGeriLM22f6woQnEZyS9qKQXpNqIDo3P7U
xKWx3EIvP91glq0ZhIzntM6y+17YWiMjg/8uZdODrBa0uA0gIMAFbqRj5cMhLj1PiWHHDPth/tys
2qVAKlWKnrdmihx0JTVUUWx7C7PNpkGpiD7g1U4VK0S3fWC0EvVvPd8zgy4kAGrzz8bgYRy2O2/r
CnwtPTLr4WDrd+R5hjLSEx5WmRlmvQN6b9hbzkHTO5ZZL1yyz7srI0sltlL18+a0uEKNcH6Q/hIE
HtRhylOy2p/ICrUpnhH4MBLFxs96fg7zU2pux5pnD7+tXr+Y5a0kBYVvZulsB1fVDMticblabT/Y
/sC91wUmLbk0pQhympq7nMH7XPJI9npYAAD/19ikGz69zMtrUmWceWf+SAmZo7Y64MvSpdsYgRGk
YHpNJbuYpSjJ52xR7GAk5nOnadbya/XNFI9+99WxCvIHPGO0S0H7Eb+F6L7agUQiYYHmuPMZu9C7
HcHm1zJmasznBSuKoumGTgsHFO3pf4FjFgxx/Be4C6ZvjFddeCpKps6bUlVetxe+l/4hePPV6cD9
GlKRaT60z9EJtOmgyZyY8khlgYdnX5ReGcwRZaaR9jy1z/j1YGexxR8Ap0jNtkUst9f/gmlCuqbc
E206tUFNQ5zX4QTfjKydpk/boVD4iB7lr5CoZeLynvDIKBSo+LaCOa10qPNyUsyRaNW54EnIHDc4
kb44FfR1R9qzIK50Rr1LvCf+K1VjFZnL4PbnMnZa9pzE2gGPmKIQ6lsEKyl69ZkwpVWLgu6iVnsz
PEKWxruNb7zqvVTXALyj4cQooX4bhH55K3kw1kuoU4Y9ttzZc8/yeVuQKAwD6LLl2P1b8a/qG7m9
gei0AGM+17wcCGBu1dAYSohTpZYsTTERLg5RyQH41rO5vKjn/q+/aLOjNJEOf5Em2M+vGaej3Ixz
g4/ux0XOvN7ckwEHrg0vfdr1X+eZZC16tP4SIQ7/HoUXhZUqWa9MeNtTqRel9NlQSRsLgpAGLHdM
fv6SDZ3lq+M221FXk07ThPv6pude5hyz9fzFSUVHcU87hmAj7QW6hA4P1FTOc7rPWrCv6QafS/T8
9fOyCGyhRO4kKSN+YrvnPYyX/1Fik57JHHVI+DoZwj3t8TfyyeUgKy+faVT3yszD2r3G/kdcBWgW
Akr6MbeW5HJJBlIG8kK9SyEqoPrs5KqRYlupZTbNJu3KFlKUCzkxM0sdWZ50G/T6GvBvyHHVIVCT
wkTSfIucR2fkCbh32iM15kVulviVD3SagRoGR0VZ3kn8RAspp3j66M53Tl35cCX49RiP/eIdTqYg
ladK9wkEfClljizI7FtihIpwfnyBFQQelGLUBpBpOt8zLHEo587OyB83D3Wd2NoJE3qmCkXXU8SD
UcZ/vlsAn1ZdJmn5QFN3srJ/byi7TFlwy2KTfOhAH77nwXUhT0jLlXil6izMxoQr/iJwRVDFsr6R
xFk+98E6SfH8pAfw9G1NCAgeEnRo8UuradG/aR5l890emnTlWYwPAxFiWIRYbwFBmhnP1ljg/RdF
gLPDpt5Tnm3ObuGZ5fl+Lbq0ymqHhOskj1WIaUrA25bsCPUoMC4qyd5vE5B8ShEBpcty7YhUq63W
lbB0KIiiGm3YCVbSjg9zde+aplsuNM/uUbc19CsoJGO7oZ3G/aKK2ZWBdnkaZFJ5HEHX9hyHnB4M
05/L7QL3Gse8wRiuKee3RoXxq8ewixWq1aD8tyWruMWSeN4xP8uvbDI7MGeyU0KgHn/JPvxy3M1C
gxUP1gAONdct0gx7Mlu4N+bXwv7ncT3NwHcZM3nL5C1wtkmQvYiwqUZQYDFfASTWyEje/TZyCJ4a
lNIVO7BlPM5nIb6r8TgCgX4eQGpIA2cJliERZP/vuq7txDDDrPO/LyCstnYZ7zTLlRka2mT/+Q9S
CVtyDYxe48QKPrWqKCUobKQ7yfe5jEBBvgzbYw5HBvAcAjI/NdhSkrED8HHV4I+QpQVYVKwmCe82
JCIZa0PWiO1O4v3f1nJNMJ45eus3aeLSu7ktQzRNLHPHfhADqreiNHRjrGugB5hxd72TbmDtDuBJ
zm8gkOz4Hhm5xPdWCfB5wxOWe8bpx596Jj3/bVyhcC0imOwIbSn42iIm/tw5kud5ZguGYWcUlQp2
eXlXBYGwIOpaxVEW4EL2mIlpqA6PK0OQl+DfN8i+esIKO1VVqfJD/3jgBp20q4yg0tdDEeuqvMsi
R26ZBr19ewcfwGDd40ht1WXu0qixRqL/d8McgMihy0DTfRURwU6JzekqscoKhP/dL3sGhDbfB1jB
WhrGpXu2LUcPTkjN10IyXPsdfXJ4bs36HK6xy2EdVwkvVJ1EuaiX2dR/lvhIMELA07nIsiR7y67L
VxupMF+Z1q7Nz/rIEU2aKbXES/a8CCkeNhyv+kZ4K6rRzbQtnSvVcVyHOZXvQOvDYN6gEvuhiXA8
pYwk4qSQAoQWUgT40IZdS1/uyVQ5T0mb8i6mJpktzJtWTyY4fdiBiqa76srJpR/mEre5Jq7TxMb4
a2uiPkdVOErgAGWlYV4CQMIS/SvOTUBr7KWM+FtWoO9wVizyBosxE0RhloIbuSsSrMM3E25ECQnU
GZqbMhjmrGfb6KOU1Ojt38vKwC29E8tXgcf7oxqeAx2fJaQRcECn6rgnEXSi8MP2+3P/0PjIrH0Y
ZfiHWVg9s72PKruWTFcNiTm0JcDP9KuPAuWqAek0stXI1oo5PPT7tQnNnv1tahG/jNSDkd1vOXub
Q4KADFJ8juucdRr7DyO/8oxeu5n0uiUwei7+M7DF1jiFriwpF3u12qKpbuhe9O3+XFEz5Gg8AQPi
chns8ha3JFKU75nZj7CW4lP/ZnuODPSDyuws+u83+i9e+IpHkkoJv9um43PfBUpZ1TmeB9p4N/7u
jPThgjLvLqTzkoNQ1DgzBHxL9t9IVZQ5OaHcZZTQlwZWWcNogmGVhwJeH46H9CiQG4okK+Sz8gj+
cj7TmetczPMeK/u079WZjdNmnzTRb5XUo9uWK8cHOlffoLYfcvNaG6GkXQCCpR4nEgYxsC5QSjXG
H+/YTsg5AHeKJF1mOZyVnx4txn/1DAjy1omGi3l1av1pKR10NvUD7M8i74lgEckmPhIZKdPNSRZR
D4HxF4UhCtQl6v5BIkrH8pw2/DZlb5W1YjmyQ3HeZewxnBrZ5LwULvSjve904tEs6u+5uzw7ouZ3
H4tqpfj4/saTy9t5cuLc9uvQTRzfMKbhgXvSvQd6qDCdVGDhJCZtKzmI5aWBmbjyq+8EQq2SLZIp
Qmao/psp9Ul0pUuWxVYap+aze4+uvtbnwt/rGtqNyFv77BCFy5qgMJdPWWIZXRcNWLV+AQ+eSCdU
vIyN0qZPO4cBmH0z2YRw2gu1SAXSiOMZ6KbxUkt1VQ0kJiST3fHKAybnbFBx+OmWpF332ArxA6dv
tchVsxQ+LtYDbHD7f7EyMlBusnkbGIhxqRXURVmuIoXSRHf0kVLr7lfZX+aaEUu3VGX/Ia2DYf0l
gryqiDRmQiD4BwTeppoW+A0J6iA0NNXUTimhBrws2lyxGB/mk0/S/9fNSPssEJDnSUQZSvoly0p8
xjtB3lncehpzeGMG1/Gwk9DNrupxAcWb1US68kAbLTAXWiEuer5TkADlNQm842t2Y8jAD6L7g0BB
uN7taAOOsyxn7BdSALc90yJqmCP6Kt7GzPC0BnGTHlgV6kL9fF4ve9EbWG3GDS2Wb+zeAE/UW3N/
4e2inZQ7GuhoNf03vQ0wqiD4pJ9ISN7Te1/g1ViHg0503l0zMWtfrvXyQyncwXiGV8fpVRGKt4WG
uWvJ6MasD6Dbh20HqQSVYkG/S3eTg6vHA/FGWR3iQnrbNBMH0u7EZQVEVIXeKJ5P1ZpQ/jzYUjSV
0FHqLt3cOCAlnewXL2XMkk7FvZ0N3YzlBIaMuxeY9H9LumpUVX38qmyLd5qOmSvYdi/5EWEAE58I
RMEAqB0Cj1Idp+70RyS8GwJbY7iVXnno/ZFKQ8bNnMaCPNf52/466aFOBBEov5VAls6qIRhK55Ip
89OghXHI4TNvwRtsCxrXUxkWJ7omB0la0xz+ufyrVSwvTel9ir7ULiDLgBHlYNisTIHF729rIAZy
+CJx2BRw4QuRIhJZgyYPbhSh+35n/muMKiJJOaeVmGWotdqKDA5A+Iyb+XOtaHaIRwcM9zYASaeK
q5uQ/NkalX/jVXwyBpt2PT1eRS8j456Efh74Als01LiyNxtzJDQJeTXD9dyKYLGjXQtGAGW8o0yJ
VCIqADVY1YhjPBjO4G/+kKKA1MpMtaAa34G2kWM5e1PFhWC+bdHtAZLyydyPwabjLMXc6i+3usqs
f1JqSkYksiz1NkNFm0DXDuoModj4ZpP6XyV/Bv0gkBRKySnVOtzqbwxfOLJAkuiTWOI4OSC3vIkw
nw5a4BCOeWl2NO3Xgj0A5hfASZMADicuD5PQvT2wi95vUgtPxV1VWKtE/OD3iYHBkqRAALZibYkK
JJh9lSdrHSHZ3u5RXJWWgpr8p//pF0y3RrALhjRaPIbgpYMc4PJVPrZBcXYT4t+vZaJurtdeA44K
t8JYtGfZYxKY5Y2n8avWB6TJ+TvCU/dFFEc5aFWgT0PYbIz0yohp9shAjMQH8uIapc1rJ2FbLrud
KEIGYYfdMzsi9wwHtwcZzzAk53g6D0wqAyM79HrY2sU18zBUGQ5NEJV8ayK87OdfHdnwueg67mS0
Ua6GsHfXk2/169ivRY8DOND/05AtuuwJaHd+NeIRIQXlGir74suOpKrGLAwGwpdVOzdYOalLGqFt
OgDViqTa5AGJTov8Y0f29U0SlKRhfwZGa0a8ujRH7ngniIZOsZt1Obf0Q8zDgNnDguCw6LyGYPAC
Mr7SQxLP0dBlH+2/AXKHmmJqpruO6EmN5okFsmW/7IdkxXCv2hLWLMU1s3Oai6z4b1riz3ZZevsR
rqRkijRA+c8vrSItdwPAgcJ36CEZjuyN8uFE2b6B4x20iuRekPEbf94gdzS8cn/9pKwKkNqqwFU5
3fxMiZjFtsbWBJmegc8WQ+SwPHmBoCX51qynvO9iGnQmMb4EOq029pdj1BoShRCmfQA3NwWKTgBv
khbibicSns0deL1lVyZt5zMl1XN5/bo+afyGZP4AoM3nJF/ljL/3+A50rbYXiYqRP038o9FCX4ow
0d9I0m409K3MTSlXd+mdE1kRORu9o55MvmsWG4x8kaK/i1xtbPRWcHw5z4/L+MkDTD0vwfgQOG5w
gl1HkhpcJOEQBYZ/7e+CDmYFVopUqaFS5NcD1QUXoo06tYW2KSh5IiMfOOdsMUFjYxWjB7AnqI2f
v+p5x5RJgPZFKGfP3C6EH3hTsiQ6a6DljdrjJhsCcgVuLo9AzyN+LdYZr9gIJQqGrTm9FMP5Tcwm
yy2lm6VwGOZA0QNtm9owwobveETnCJ31KJ2uSipnQQiwTDWutZIeRruWteaCK5quchQTVVN72kWj
QxuFp9LA2805X0lwIPIu9RrWNbptpYbZKYiFPNaqv6RD847a194Fj4N98uPEzmTYxDTONpkDffWr
VVvHctzu7XMnvIWyek8FBSS7qOvxm0RUJYCxDRlPYdGgU3OQpBTNw0QuN82G9YaBOtmQvVS+NJJk
5RDaMhY+IVpjnBdwpYSN6B0HjC6g/XmEBm8SrFXMPQrPGveIc5WLHyCwaUkrFr0ZrhW9O3pdd4q9
ESOA1DNysNgGcvfKXkKgxJdx7dELV8e6CJ9jCuDTC72zXoxesCDDKYbuM6kSM3txbD7qJsOHQlei
HgiuNi40aUtvgMxoJpfYt533GADa8vsgsTicGTOFqF+CoXjPq96ep+hLMOBq91270hCO7ZXuEtNQ
REH1gH4bn4yh0BqAhjCoW9+wVeschHtFCqoNe6U3rrJ1wwvNxoagWZrLqAJz8gUxD0SGFUmH0jSl
NVJ/O2AVS1IofofQjPiMvgZn61nAjz/fNlx2HVinLhc6ssiJywyZOp4Z1xzE+AFbJ72+1PTfJRBM
h7mDMNrbj+l9IE4g/bdXfzofeUXckxEpbhKFg/FiWeUUCHEVHb7ftn5br8NRTBvzwRLhHfrSV8P8
UPNC90J5jmsqRZPHhzUq7uGVoz0NI4wBQgkbjw5EIy/ns82THzYW2TJpO3nxmy06liWU1eTP0HuX
R5KvTwIZ5r4JvyjkSHXMiI2wKPNwDvYQGZH9E/QcmqShCONRnZUxEoujA6thVqByqU6KjasiP+NM
/TZ9ZOzsyvYACCYCr2C33rMFU6c/mcFaStdRYi5SMrknHzUJuYOqMNYohC0PCTEpo9vPLt+Dedua
acDgu7bm7JLFIPt8wApgM467VzymrX7WWoVjqTJP2ygBQtmYpyv5YFNuBaaJYZuz7t48QhOQwKSD
8z04iIZU7hwatUmQIBfxHuaNFBy8VwmIGh67FwLQ8Vq9Vr3ykCa884pQrFXY2scOYv57t8ywB0ps
MBxoPqaiyE3o2d57+DYzUKpgvt1NW9eSBqBzOcvMs7eJYzA/2kY3nTBHuwmSwAeUK1ux0l0VaRgw
oEBp860Bps3dRGucQcfAEbonGXAnAdI9A3nJpsEVGG+OU7xYy4IEkAsvfYSUpJb0W14ZA+OH//DP
1fIRKOxHz4/oTyMLpQ2FTeGZJK5Kshbs58UH4f5Wyi1O+A2hAXDqZgB1o9raZf48ZEiyrt7OpKBQ
wQmimOQZggX0avGgtgfL/Cl2/gpcc49doWfd4AxnsLF9G1WY/QmOXfFUxZg7gdh7V9pWL7pa6JEO
niLLq1OuLC2s3exWMai/pEh9irA3DS86FI6K7jgse9iaOPFBtxtHh2OsU6DLHEiNFiG3yLPzFGIL
UKRONH1WwYLtAlt2dFr1DXQsrXPVOz0NkPlZpDhDTAcnSdsqvaRYsHC1erFhWV+Wc8wWHoxg3Tl3
xOELJqIpBH+Us6PVAPZfNEXBfkUl/INOO1K6PjdbJCyHjpEaPUguHuKLuvhqBNinVLNvIVlMl8A0
XreiH1A1j/14WKzJEbx/csB3XrZ89hhTNv0e5XvpP5uaLooMXPorRS5fsBq2NUddTy8ndABzyo2t
hK5TQCZK1vBh746EVDGypOcC74ZvUMvLzNpoRBV7l90aTY1E+9N4q+2ip5L1ElBY4E2dB1MkeNS9
pLYKI3wLgrPX+6aOj9p50YN3/lMDFk/JD8FCcGfBFPO4MIt+cLj5fvgwH5xEcHVcEk++oMa0Lrrf
Epfn+KL0Ci0KBx0er2lmY8Qcyl8oh+1iPOh32Dz5ahDgaloG02rIKzyhpCvh1LBW0gK28KVQJIYC
fvLcDsZlpTpCrHIcawsuHKixbdLYH4mheoFSXcTla3REn8rpEpvNAxxvi8cZIakDUCqGKaSvTxV3
O98yLg4JTZ6QrHx3xFDLYtHfUKlJvPYrkEcrdKE6lg+basn2415NReO++1en8H8aQ/T3SR6IXnQm
ZG4Hmll3VcFR1m/EGGIfWc7MmJR17M7oFlE5X5usjEVv8UQmQB8sntXyXWzLzFoxl0S7u4YiXVz8
BIKxAsbdl1Zti8qKOHWQRwe7hF8saUC+UOYhztyFc7PQ8FEg9LNmlQl0rUIv2CeQn+j0HaDzPrZQ
0dH+tq+M9a9kUfdUICyAYzud5TgQdFYFYLK1Qost6bxbvyE56anYcr3OQF4kLkqdHLyoy0mufak4
4Bw2ZgCCOvjWkThh1nI6QngmLHCSMLSBbjRP5+OU9cpRUzMmBZKo1j9eyw/ZFKJz2UuUOAzPpYbd
updwEXc/BWaqAxDWaTwYIPd0m9d58NqP9DULduDjJ+pmXOYVYpprt+RLUkzewlfEDDHcxHQFv8K9
uIIskc6XQtN5ukghvq1bF8q3dAF5qX6EfeJrzNb/dAjyC7T64IyKBGPj6lgwZCihTtpJbxkZqpRL
Cp0WaZ5tjqWnmMP/wrvVZNKlqm6EVr4KKzHzFZvoWFq643rbt2uWe1Oj8iMh0hLJXVtlk69B8wCW
/EuRCUROVf2LzOQSOGnhBG7Lgs+Xp0zE/NNPUp/TxbDCerBJ67AnGdTPI/WdftLkM1CQMF9/jsl2
sYoR0goYcMbNQanILev96wGtGSZH+O1h/XnUiGD2p4eoEMwEKSFkI0mD5Si+0jbwwZS3dBf/8nDy
cFaVXSExW5+V2ixc0yjNRIop5wo3avaXd+bXZQqqzU73Xi/hKGoGc9AH4NBAoyWmnFUu/rtmwVXl
496Csqs7AQHzwpRUpsFqAj+UVaPGMLI9YEgZ6PKAYZ2L0Q43wzvBypj0WRR2TQ2azrACHdfWUsPq
Ki1k4qErK/nYhvZ3v26NKugd73f+hW/gryNeF6hEA8sHIHfNrlISDZqnQr4dmTA1a3EwBFGQFVS0
ws9YD+6+UTGT+LPN6QBC8zcESzLzd8mJ6zPc2q2A09UV431/tDoZzKnXr9FCe8IG3GY+YUK6pvP9
CdJiAuLoTiLH2xocJmmKQvwZ7JIPanBZr2DW9p/P3mHCALgHrXDPQNUowtsPlWAc9XQiY9Zcas5/
JiREqj1bmfhjXYkge0UfRxJlY4vst+xYOMzd2IyL1sbulSQfMPOGx4vjq57GIxRGaNeGSS4198iU
8N0zjlVRBxPDivFIiLg1ZjnQBHF3GIMsQsNEQI4r4YxWnoz+eVoE2AAuj4BEFbjm7orSqmgyQktm
AYVREFz8yVI1WKsqkBEzOJEtaen0W1F/0DL53lCx5ulB6v7Y6uBjbz9xZMCbgoDHKkBEeBc0V5Is
sD96tdfcMmzQ2s4wTxbrnrAURRCOzkiH/W2Cb3OEb7a1JTJkidUKFY7XEgKQPhb0RHcIpLvpIoWT
g7v1Rmq/iTRlO7uo2fdXjCaoTDvfe7Yqm9pcscxqJioRyA+0Ph/+GGyTOJj/4A2eUaPo20tPr41/
veHo/LRNADp0/ObxCGJqsCcJ0An7hrsRX011v07xQpNkf7hJQK9SgKjgTMJ5tfXjaiGyg1i5Pa6G
UEGcMZNIAh1/mgMlEUYKVChTyjySbXwnTFm+Ol3AQHdt4vOjObnrjO5Ww25GIrpgiUm+/iBhuCgC
0Rwdi46W4zsy8w7CUHAp+wQjKbWnUYjf/zZ+QWB2ptmCRz5Q7ZvD1WwQS/Ba/Y5mGsngeiZa4bDr
GwirYETXZYnChgd8qE0npacA4yHxcOJg8+/8NTEnLpVPBlNJSxSkqlXUcaIv/3LMMB2ibSxOXrt8
EgAjOUOJ7YdQ1DTfKe7i+5k8QrFUf7rSsUb7zrvVneB8OeoELCwjA3tWpS7XlAxp8doeEEkdnx1w
JgfYMEac+cZr0B48J32nU0EF7DkH/r5r5Vl/SxQ3ou7UuRakgDXoHghydcLz7aau4CMnovHOlYl+
bFt/G/jUrZYKnxs+ENtjddaVN/yWOg5zYX9orcR2nVkckihQSv6GpQioC77D7yF7YwjhsJWhwKZZ
g87fvkaToZk9IjwZT30ibZmU90zgFltYDMZeNn6ecb9m9OSV9U41S1rQBQi7Q1EwO+k8Gf9f2jiO
U3m06SnNb0TfS0jTpGqpjPH/JhHOPY/s/fNfxjmqH3Wr2e1xnMxl4J6/Qh8Zehrga1/Vn49TbgSl
zjSWJcU8nll7L7pk/muYQ+vQqYcaRBGh5sJO5/JNKUIjWoy+4zwWKGHni4Ud6NB82tV6rjEHeXjD
I+tbj8Ey05EmpxS6sBWK5Hwi0/yiXxysWu857ZRkzX3ufO17+viOnAOE4OOm4Duu7QD/CXctTwhr
h691Z8S2xS6jzM9cOpd/8J1mKn+WX+hIFNTs8jZwKjl4osVI9xSwajhBNzSVQK/+WXUvKXOYeWxi
ckdPJKSbJWfHj3gJ9Pom6cFOxf9VS8qsNth1M7dUgdOtZ/tTa68do60hWdzMnI282RcZgQ3cJS4L
UH98KL5TVi0Sl/2FK23JubFJ2YA0K269UyXd0RbDm/qsyTk8Am8XF0M7YB09FERsieOA8XrEteaZ
egNr3I/3jKMvGP7aWqjifuezeilw04vz2xfE3a3Qyp5uYeOd1y9y/EVvZvVex2/AVC92RKWfkqJq
7y39Hi8/j0L/xE22jQQgKRkinFiPeLdBhPmerxEBWoq1dGR5O3EN+DK1zRmr0K65f0eWdsbLLNtU
NzPn4UWGBeWf5kRO50uCJkTMDHFwD5nfwQFTHw5Pwgy92+z0qwQ9SH6TYXiSFm5k9NnaPtxOS2mA
NcFS2C2VoVPtVX/2SgPeZS2FylS0jrEBZ5dC1i9EqvPHo9o4kZ/P4K6iO3cC7TTNaL+FQ8Ky/vRU
qQ3wNsQNUn4Y/Sai+VEN7X/WcYpx7IMa4RCZ5wQY7jMMsuelNM0q2KFFQOabJH8D6GJt8yCdGX23
MFx1PhI53CMyxgHbJNVNyUdKCv8e+Ee4gKrO5fzwPU5EQ9Od8eYTtEA/PNCfay0gvtKhi96RM1+d
PE8HsxvyCNja4wNOQyBndrfCvs6o+cSiAW5e0oDop9p+3wJHfkl094zAiaQCm8br/8Sw8AXM+nvx
XLKH5SOqkkiICgTe8qv1ptoHrT0w7UOgCNhYN3xUl2qOHXpGjgHKyIHL3IRuV4OojMWkUfUA0roI
SpT2pvodEKzEDE/J3PnOW/5O57THbDO/wgl44dcWI8g9mAvVlGp7U5Wmgv+xgc6NCO7FstP5ZIuF
6CA0dV2JwwN4c/hZ0ZjIzopnA+VE8rSnVzmXYhAvO0xMxq+oDRQvFgjXCG5ZYN/TSQ6uS8pPiZXy
ME1fCNU6TkV7xtku8QurCELVY+AYhtohG/72KauehlNF8r6Z8XXEi4S+DvWzOGb82yYB7aDzc8xD
6iIPq5Yc/tJjNOWYTqeY37q3WuIwaxNl6W4LBCw8PQYKovEgweh2qiv2533VgoLStHy8WA12b+Wg
qK+D3XM713+oKg4d+dHhx8tkcw0uaDyKR/3uGfguz1/2BkzFqCkYOduxFkaE2GPqzYUUR26cqBCw
ZdCsf8DyHs7imx3TimuvbBDOzj4hUHjGi+SWf+aKGvb9taSDmbdSZex6ah8jXLoEezLm24UaDDhX
VZcIn0iKniJsT7yA6Ag2lg+7ixCKeDCY9GBzl4i8t6RylcOGhap95sV51D1Dc33XI8hGf4tr/m7r
Wj1Z/oSeM3WlU6psmJgJUPIXr07r0YmPpjiCDiZltj8qNrWeDtYLerGfxUyu92lYDPw2UvRSAQOb
kWQvS9c+hULFZTKh3MjVyfs5SojEC4HBpz/eidjU9bYOUx/JPgzKKmqngvAI32bAVgr8aG3zOrwZ
C4YLvZ18CchsIu1+v4MtbPjGL+lhQqA79nqej7re5McESDvSbSM2peRI+zbwpSNPPhZ3ypCRgqet
m/BG8tWYvItKxrfq0uuDuLtODYM4Bq8mBvSClEZdcLVVJQhU9tOdOdTdZAc8NBY1xy8W7xsG3JKb
YGfJvaPIBxuU33tOh6uBGQTt9coeTY68spW600jtZBy74HUYR85p9LVoKYacbnOFfOzvbHvFh7e3
DslGalawQnm6saFEBM1XJWJjIVz2dZNORBI5OFLGLee1foVVBWClmCpvbUmIbheIyON4vM59a7Hc
JfbXucAlc3RjLMSu9d0XxPa5uBNGKyr0rlMc8qYrb0vR56KfjMCsTzqEQvqn4OkuvoYYu9nfg93n
6kaZTjqhHvXg9mKzfBkceXlVAzgkiM5XppRV2ZGxDm/huMCMBtGKggDGsuiwWWA1q3KZ+rIdXU5W
eRFK9sfqpbkecHgawH0zH4kfcYzCDlFSGXL1yu6xfrMESf5yvdYknSNzY6P9heI9zwlVbOKaNl4u
4EtlqIDugqhc0C3YLMJQiQSOwL09qXwSidIVHydousLXXPAZxHkUlEKPZxrjID6XD2AmDK5FL/Oi
g6qR3pqD/rW9TKcCklubpti9iL61pjg01pcB7zFLWJg3UwxYI2wBKGTPnw5yt4sd9DF3KxxR5ujz
E4vjG9FUSulBxE/NoEcbEewP7k3SS6x9pJVxLwLbeFsg3jVZvLttCJZYsHXeNlclJUtnvwXIQEEy
zD9TtiPHowkyxNx9UNff+Q23rkp5+mMv+mxAoNSv7HYGzUcjXlJaSscQAb5KOmrDJC+83ZeklsGx
PWV0Y44o5ExfFYu4UI9d6uL51MV/0NjVhOyD6X/8apvTzKTpPCvtErvnwhp16s/+ILGHyjm2HKsl
CPfEJVMjLxXQVNv3pBaL08tya/eO4X/tHry7ckwxzgnm8pT+BP6fRCD0yhfa0QxUaP6ODqqqD9sQ
1DupgaJzkVoP1LkzbExQDc8dnan7W6tAlwJAVgLW21pKxO5LMj9ML1EauHhZjbZuLsIoPrU6APSV
xaRI4PMpQs33rMsTQoWy3G8YbfV0bG15AU93jueGXoKvV8yrbWkncJDAPdER5M5uuUE3UT9eOPvs
HLmyW+Ebue2rvn9RmZpx4m7HTPNz/tu/uEtSRVbBO0B68dPlTEs3k7OSrXUWHjLv5e4kqjnw0Muj
F18H90NVBrafQ9zD0hDs1jgWqXKGLJgm89KeIhenNHb8yW0vA7+Mns1ZsIvJjTQGaUqk12xnUNok
S8eXTJf328aZ1dy4nepgmOoERiqgNn67GJSqqNjG/hl9zt4ykevYTkLbNMVxSThNDTa37HvQMDtP
x7emnxRAYl4lIMWXfZvH2/Mc8Xr/7PoCXqOCJj1wGRULjL6ivCXO9Ab59fHyoo/mj9yrzGUfmCF2
kCiN3ihMsIx710PeYBdNkrhKadW8PskMUuduOyy1zysTtNB8vP//+tQ3zZ5+5pH7GvBHpb6hhJA3
L8cgL7xj6182hizUAwyWDeEhpGa6X6O58DMvruqajvJ+/wbRQZUgGqzBUr6IuN7frbvysWoPJXuJ
qjey+NbgxyW1YYx7MqsImt/DgMW6jf2olltDZcH5ITs3FrTU3iXB7wBxN/NunHNtwgrTB8C644hb
DvlkQCbFI3+ITR0ath3u5h2qj1RxeOydTCdX9XwGDk4ZVrH2zhKhdbewK+NKyFoQ3FlbqFennTXD
WJv9tsZBjweej1J7hRlJRp7zei1mSRNbTHGRGaEcgWRMdeL6e9d9s6mYn3PAAgXrjLW8F+dktO0h
B0Atet3cv8hv3S60AuzDp4seW9uLsYTIgKGSwQ/mX6P1FxpbbvwE7x+ok97rDlqvSFfs773+JRoR
qkB88l92O6be8ZXmHY1tbFwbCl63L61GTaqMPYaieTL8tR6ITvDG5M2wta4ge2IES6TbAFcI7pFi
p8TtLbsGeuJ6a2uQCN0UZ02M/hWHfR1IfO4f65HA0ymq3jGf7GH7ZFQb+7Y9SkLk18iQ3xL6iF1u
8GkfNAJYIsttGsQko/jS2ms3vmMDg52XrZOnZlgKSmImgS71SyBVT1hALbnuBRsq3vzHQ8tKdRrN
ftaiZc1et2i9Zqat564QPW3r0beWVXkW9FAEdps8XFnnDSi18N4WnpX5DvI51XDE05P9UX5vXhTe
+NN/ISj2XGr+8UEL5uDHWHTh7XS5Km7kCOWqsVjsIp8mCWeNFdJW1uIIWVYKQO/ciqVjjPu5AhCj
D7yQ88Ws+n0xgdfSCozvna/6gRCaX/VqDgti4Z+GFYpQM52wfZo8Jq0THuYwY5pVxz25oAFdz+BR
xaQA8KJ26cbFbOHLU5X5HX1HUMfFdTkz/rQcIGvfFm4Z9CC1+lNWF0rcn40iqGAlLCWp9UdaW/FT
gd0PqQD3JSFU2EtI1kesjFb5+Mbsru8w6700UBI2rz6RMYcbBPssQk2fVFoPtBrgj+XMUqPohlBL
IR8j6yWwXWd+ploekN5fc+sgyEL6vAVHSzppmsH8WOHRBBf4pMsDguByo0jeuq9fVcZaz9sdSsbj
CVbxq4x+wJAExX1ZSoGiE+hAJIBpkoCKt30IiJ5WyThENf0YIJzjG0RezBGYUXY+r0vF0a1AUWpD
rlvOZBj9+AYe0kMFLbTBtuXZ0Ik5w4EnRzQqMQyBiGSdqCQwqjdUDD2APwx1qg4tR8QYP9uCQ546
gsEynlzdlF+Z+TPouyxn50mO4sgcj0JSIFV838Zv4/O8MobRRjXOXcIR8eYRVg4ad2MGnuX91zoT
6vzbniQUUP2XpR/FbqJv8mG1AfNEXHgf5DqZ2FnEoGZvnjDs2Cldq+VoGhXNonJfutAFYBkvsPkV
7jm1AVFkZ7zK91q/p7qUxNr4kKmYFL728pekK+ndIw91X194hmGlSy6g46ht7qTAtR8mcHaXxcze
j3n797KurVvU6U4ApvsSdGdVXZBTE0EIc4AFmnPrxIKNsIVvKFSxhEOZlWfu9Ix4NeNBMCPNl7mS
D/MDvroMbuApGXLfdGl4fObEKPjntdLVuZUms12UZZ4hvRkFs0Liw2Eqfwa4GZ55ZuFPAVk3CK+s
sHPjvZkXlVnlLOtcwy7YRJfJ1VRztrugwLV8Zkp3NKJSxMyj6SfR0jIe+kqNs7E88PRjeuna3LdK
4C31XWG8wFN4T4iXFwpAg+l7eRiEEyC4fL2NLrF1I5n1Ng0HFSqdTDnrNXSp8so5RiKoGa5I3mOq
kHt/4l0eG0urYgNiojqEWIEQAomPeAMFz1K3nDyiNm/aQQX8/7BtXygqkInWE47SS9gwcWAKNVIA
mUg/oVJV3IpzXy1ElES2fKhEHhI3PvPtAR79sdgys9xS28XAvzncnhRMDtVUHQriEf//pmF0P2Db
N6wJ66z1gx8oOwJzrbjBpHm4ITpWX5BhRGFdjN6yrPpCxt7tFtsOma4zsA6q2sks/jGAy411TwqM
ODGEphTviIwixpUCuJUOM+nCg66M/jYaaeCH06EZoJVVPKtj0B9b+LJXO7lXapr0RTpn67JxTM06
btJQZJ+p4SYP2Z8nyQeqzWpBcN40L1vmt86qUXwNPmQMFQWVFSd3BN+m/hC0LNOrYFEHQVJ2oWQQ
8KdxhuD3Y1v+mY4+8T4UTQabMMPVZglXq6t2uv1XKPcNv40iB+NPicouROLVuVc1RFrzUMCxYl6H
qb+rrmcj1HtcUrPYA+sPh0IVEHt7Rgvxk4x6CXREGo7pWp9Q00aItzOe2RlgBGOkukuHw3fbNpQF
F2+y3T2P7cDxhrclnQ9xUniQGtYIalzmjwyV/7IAHomwVHI2KdEUD2J5RHC/d6YWAH9lqCP1uzhw
GxJu9RpJvPiCpGTjGupraDWhd7FGrdqDqZUPo+gPP49iJ2pNc+6BWzQ4WOEp+Tui2vuCGi6xu03U
V2y5wVq4HBhtpAcCCqK8Ojyr8wb0LpoD1Y3uRy04V0R8tSYl/IpPL/nSRIIGwpj/som1iRx/rQDS
XcBb6cIyYS+NhJgx1RI+/viaAavkEX5bOVp7gL64YgZ0dfSwdX21BKRJQ3+25Ix9lrCTGyXfFkwV
0a6DW3HpHzyqjgVFaFYMYdsKUg914KNa9nSgTDrG6dgKrPa4Ro78aL/zan2fphnOdDD3/J/pVxNh
Cw1QSlpFV0GojgeqyAHd9w3xU899cDKMbFDOSbwpLqCLq0gKrkp4KJGrXdta2GbQduz2o+Yf6m1H
TOQKBQh8n+osXDKzpN7ENCXi+ZoQa1d4IfBpbT+mDnUDN31w4bU6xQ/LIGGXR5Jbu5oQHRWof/Ew
FMIzGrppzRxt3rw3ri71M11Z+w/gfE1PKqAJq5UGw0VhJzHDVGk188aZr+KlxLCb7tx5/E69aUQg
IWESJBOqf/QboRYzPE81HXxwal3bsqJEFz2XB0U8fRn1lTQngevCva39jcmWXt2jtKUtQjmZBGBB
Ele0Nj+DCCytElUBp/5sOtv4zU2dL7WYvf49/Udf8ulKa2Zrjdw50p9fuZLbCqH4oY/tNoY1jXQj
kCgQOD4JniQ7yu78gOGpNgBzF3QhnJ1Lcqrs6QN25vm1z1Ol5qvXxQ+cS/6AUuNmqzYYY+xhJcK/
n3dNf5XdoX4RHp35URpeDH4LNZBsMJeGnqR/UxZUswMjb/rT3Rl3sZ67qMqBmfLy1QjabCGhgDh+
73odvH8zrytHEGPRePHBnq9Kj0twRiM0eMf2VK2n89zUXBki+uWErTGJ0pkW+Lzfj91pl9ffEosV
4AirAVEWW50SDgjwn/hJ2VOnm51vLBPsMA03WiADpaTs3dJb8yKW82aTiI/uaXh75GQ2fbql2R4f
InE3fxwtAIwYXprOltRTZxeag7nhCAp6axp3XovEZfYENF0FtyyNpIdPNeOQY5OHt2jo3BdUcFp3
RZUXTKgH6dNyj1jv5s/Wq14jit/0Y0V7rodFDrBAA1yNhPjseX/mcVYHJqyrc0++ExIVTHNkiJ3k
k6CgVV425hnwCvkPVdttKbk67CnRsRhGIkuecXpI/VbjMAX0s6e4FukqaOvBVCPWIdJClwGmA71P
zNl9h+ELQcDjlFjGZ/O2uezbuNu8VdgxteSlH0lNuys5OIBZtwMoZ2a/qWtuhw2sjFvPREXCKSW0
P8Ptr3RBcObwV706dyl3uVy67xPAVzGteY87v8w/oG56Ta6mkIli2G23iHPdtIOaXFtm5AXem6jp
6WoJvQpjbR4MxDCxbQTjY7Pnks/oLln85bWNPw1SHa8+0oHSV6hjM1U7SHgSCg78XvVFxsNBGhl6
iBjKGIaeNf2QwEFyzaeB1vKI+NIX8X291GM7TC3Z3sW13W+qeUUfvmG7vkihckGTlDmokDe6+gAq
eZurLKSaMPu46a+6CHOipGYz0Ccxc91F5GZF9vTrhBt4goLw5J1JJu699hkVzTftfgIL0reMTvnQ
4zsXtL7sg6ig2FaaOgaPXb5c9/VTj2wt3uc72DtsElD18mka6Wb0CFZE2vh/en3QeSHkzAGuGJw2
/0dS06LYdi7wSbwSDiI+povpABJRA/Ipq03lFPyxXJRc+iHiu3cTyXQcRgS+/OmWzWt6v6rMaPDK
uO/mTYHjXcA7BZkxzSMJSlxBaIOniAqJHEBgF1QQjGhZFnZ9CaCjMkiS357TuECvG5I0A95yXerJ
KOrY2rCjtaZpViV0wPEatx6cO1fdmwVZF/inIFP8yNrP+inR1V0d9zB/1y0s2XAOAvkaUoczRB/R
JJ20b3SoKjgx9o1WysIN6prBucws0rzj5VYZQUW+BzaMlYScKrg7fXQsAuaXXmMJgXVsLhwDYayn
F8NhP0RPGxcvpbEr5tw4cGJsIq8+nKrXjFp80s9MmdU5P2tyXxwvBCrQ+HMhlOsBrCDXz8KgKyHN
XNb0vlcwPLnj/zCgVrqfExo+RhtJL83GGqFAHfJrcf3yUOZ9slHgqQoT5WeZR6NM/1dpgYRNFV/A
x1Yzwxn8WVeBL2XcWw3w9M+ov6b+VEzVIq08qERurz2434KtNefAkhI2hFZFuu532yISdvFAceZB
iFIQ1lUQw5ZYe1KZo/ysiMBpRW0N9wHIJ3f1JoK65RRbbOl663/NbmfwLLaVixOgrzGY4VkcKPdy
84031IUnGVShOPjOOwiZNrBmhidkwzEd7/zF1mQNgsMZMhTq7meGgTzyuJdJGCr6YUYFd/YxXhc8
gtCybZHUMB+H6VDYH1yqwsygNhw1P9d/XfZJUj/HrEEfluuEsUFamM9uOF9yCbnmweMGCwRHCZXz
ltJmi6W2X9lsgyiYdpYw2SF5o8EstX1LxWXCb4866ucxpbVpVy1FtcLHaJrI8nvcNRG+yAPcfIQa
mCEe1xcSidbr2gzzrUl/W2bTj51T5833Gupyf/mVpb7a26BUxeNOXIxaavwlwNq5Kxez/kgsNVw8
DiZGBWn+5o0dDmZqZM+jVuhgV7nJibf3xWpo5D2RGTsuGI6XugZo6DqD8SMAUohXQlPBsqoyReUp
6QcEvW7g7Jp69o0kucKKgcbSXF3m9TmnCqYyXRcaul5cVZnaULNkP5KecjZ0sCfd8o+d+H5Qt95P
jCYarNZshCzb/HXhLJxRAZEsiXgeC79M7d9QjlTOuf/zAc9da9rhE8vWZdJgYNSn2/3RCzeIqJFc
8Xu5JSqEthFTPAJ6DWHs6MCsfXi/9MmiNLM5iWuNsxI1LcZYd3VxqXtDqxStMcbXcIowpjSuDC7o
sHe0utxbpbGe2mnnFZguFY1QHvULfVYtniBL4x+rsL6auzwhA8MVGZwexbmwJ6zXuVpYTFISqbNe
zaodHAEykBhDo76wLzhl8FtVDpc0vboubbTyIUvrq6KlzVUVhfeSeHbKA3YkiHh4ZgwtUf8NhRhC
I35JdSMINwCtEZiiPPzNpdlWBSsEgNLBG68JPasRTxLZokMKKKmjdPD0mKH1xlmiYW/mwhL2V2lQ
dGCzLvruXkyQwnnBByrj3iKIJc7rwcSgTD0HS2PP5u4E+0MTgi9NPBBOCPFo8i7UXxi3QbmYSMsY
RVUY/W/B9TX/ANrBcB7UHKq7FQOdAirGFMqbsy63v/TW8p3hB2n14HI+j70PCFUEugievk054i1h
u2sHt9dPxn7wRcjOErCaVyBTqIVnQepTNR+gYJRhJ4CaUleH20pnpudGA92T4b4xXJa+sevyBP1K
L8zcgkZEO72b7n+n70nLl7/DSPvJtjQ8G56aVo78npDZw6cGCS5Q+p3iy7ayKZrYuK2MpdyLecay
bPboL/5K0P6sGrRiAy8qo+u544DLkLbFyaSMz72PI3HaWHoVROuPJaKZiC7q0u2lzx3tjHxtGlZK
2REeAGR+X18Ktdu5LrPUTVm8FUzePmCU0UT4gI76H/LXWXSe++hhyH/2AbGk2iGtCJEXJHFeLXyG
hTkAEIxnzFhBcFqFntN+Ge4LgK+skY1o2oFwBWeA910iU2ZoVkXjFHXyl72DRQkIjiowiujjg91b
adK1MgixOnSfU/vLHRM8yv85GmT6NAhOHgBoYw4cRRgtl/H7OlaKilrJw+No7H3aVj/VIuUhWIlR
HCk8YXhbnqinuoe7WTsuRQM0s/tsloYhKh21y00P0Ftoa38RK/I1FGqmwcpWmcsIlfSVLDs4kC8A
kZrnrcIn4pxqwRHUr9Bsm9Xpiyf8vA4lw0Nz3vJVjn0ZNn6nV3vJY/6/7FthMIT6GeR8mj8YQGeS
py92thGpmmzV2NLsAEuRDI03lZ/a+xWe/vn8OS2gSlCDIYZr+hLa8iKD3EJFP9Bp2r7WlK7iP9m3
qOJ0QB5UneRCudo+F8IJVRraI5qLwV3K61uubV2m93oyZaGW1hEpvNUKmD3+vsZ5bJsbkObKwzY/
jj2EA6YVuoWnEnwRPFOaBD0Ixs33K9naHsnraDLS0TDAiemBTQjRl/DK9hYEgqPjOuurLzoU67U0
SK9DSQ1BHPQh0uG91Cg6Rxr/p4q8YnBbMWFO1BZgnnAnAvv4/ShPhPbNUm74HlXk631L+hf6rN35
kDJmn29ddVj1UkTvh+ajVTI7eR+rgfZn2qx+Kl3whyhoqyjUQfFx5cKm1XfAxJrGw4pt5otCLfBI
nGgPdDZanvml8rMdR3cxjkhpBoXY/dKXrO+2RYmp1Vz7WfDnNX2whkgKHmnLa4FK2G7algtnyiIX
VMrM9WiS0YA/EPPYGHuxyr78jpnuSEXi2Hrmy1/8DliU+h79dm8CNyaQzwVxZ5Jui4NuMffEnWs/
oZ2aILiEmJ54c0MpsFN73fHoVuhg7WYQ92bRR6vFLwIAigbYNeIBfiHeJMrf2IVYdhM3vcS0V++I
979to27djcNiJLuyE+IlPOwlc2jB2Hu1cgFrdSAMAFI9SkfjRQ0hOkqSevKT9QIvQOYI6e+dgWfH
M8i+GbWU6VvIrJsYy1CpiMX1xurp6cpCJNZh9j7iiPjCCzhDDBlgqT+P0RpbJZLxi9oaAmzB+igN
PNF/sg5+718NmsMbGz16wxctvp6BrO+5UuwdNQ+aIS3Wede6DYlmaqq5FnZsbJAE+z8HtAzJOVDn
OrWSWK53OqsEzW0+tgpNl3glOcHvAfS0PUXNqFRy8ijg9eyYueQi4QQ4NbypyRv4TlXyJFSCCHS3
UqpAxKIzSv+8CfsIHei68wX283pQXokeeMLtEtG3xAqcvDLXW34BAC2kzNLCLfYxNHAqJkzB3a8R
WWsoJ1tFZz5Gcq1t7WbqKZa9s1IFZHYabYvk9GbovphVXkzSMtKYV1j9U0P4a2kTz9hKke3FHUBI
/7g5GvgBqwruj1Pg9OBalYvpZ1SSkYTdoqhQV0APqNq4OzKvmPws57hLzyJTGw6VR2i1mnx0z5h+
c2JIjDXS/SvLguYocssglOBwAWSOhzXwu1eDMZca0J+Eu+pCam1Rx8QlWoAPjU3ShARBlRu25ltY
F8opCPaMlXz62icMzZDlLUfjpfzCT0NNVOmvl15oaQFAE3kOIssdtiIh9S8YQ1bEna8Lzax9f7Zv
hI2yo24e8LAI+TIQz/6M1lCO69yu8+u7OHU1lHdvznzHo7S1CwSjZHH7rCQmNierluZB4VjfUzw3
hiKKrVpvzfhINdE9RdgV+Pw+aod7h8qTuSdch/paaSoFnNP67w9VoBOuicMEsYMs4L51HmLX2D3U
LcSmgvtcetJVhd4gBId/oyvYQslcve9iod63Tm987L6NcjXDfTpj1Z9K1sZRgkYVGqLQipfS0H1f
XtLMJWPzd43Z07HLsERmbi9qF9Z7unsNfqj3ojYe5yyR47ZvGfZNo+Ogh8X3/cGGZvcI2kd5Pza/
VuGNdcZ3F1SW0W2s9ySP925iS1Dz00aw4gZhkVDG8WdtVBn18mJH3oIrLXDueOGRGuIE3UTN2kmh
XMc8lH/p1nQ9HNir82LR1UqRzH64kiytyNqM74jWmKAHB8fU99OVf+tEqnvXqPUl13UfMizbhgkj
Vx2GCQPx7APh+4YpPPxpbdCwHFJQi8Jq6qNB34Grzr0Lt2Wmk1bxvQ4CrkELGNGKrbfPdDsp9DQc
M5kCenisd3LrZhkluO562XzHNAebZfSWXCYi0+JDFciQzhGXZoIDIOpBw/x1NopeKEdcudkutY8n
2jjxUtsSNNLgoNoxnZ7kn5NJ6cY19/RDtmyCouB4+xulmGXj9KB2ETqSWFy9zGG+KfL1g/mBVYR7
m9YBVc7dBCL+UMOq15nfkhxlMS37WnvVav5IUw+cP164KOLBm8N/Fslq2O91TFBCZlZ1pJXTg2bG
YEnYUDJ3Rn1NjzJcVOT5FvxBMmKOGK+xcIQYkRQGOj5dvmrD18+jjSQuMHtGijVu0YHHGotJ0FSd
1dKOrqvhpvnV/LWx8hu7R2XJ8etomEmk6mI4ihAMJwF4r5Agc1yJ1G9YByYFb40sTYLoJYUZv+Ci
qgBQTivIRH2k995vgvpnkPgvaS8sONL5ZLBP0w2tikXduIw2wtxBSddh3jE8nJ6t9o05BAINqEyv
h6N4g+qdixes4yvATTjH4sylpLfO8RGEiZuSutcNzKHdmCnV8nb+ahxdv76JBElUZdMC0RkHquSi
2dBw8nBDhy4eHKACW1IY+edEE3mxdDUIyWkr3mNXhQN7vxa/hDUQzkh6+4Kw51cMWDS0TTMcc4Rl
6LSR9r9qh8eXjglFVVTgcJW9YrAod6OokqcVtXpTEc+n2tZxAo8Lfp5sOsGk3ZYThehxh3xA0GES
wSThrEZxW85nXZ6qxLlHODryl7LCXeEd7Eo83KQ8y8gh1eDdQKg4Je6wv8oiDMqYUngLTdnQJJ1M
dbJpvcV1Gzf3is28b6aTZ8+IIdTG8CRT9At7ZsG/YzfY2j9Hc+IJjn6ztOk5gdHPZeFB30/cyduH
IOk55GD/94IJcpJjO3lGPNzzMQSjZYPI7fAvs9c2YqMjcix6+E9Dt0VOHaIcK/QVskhhWsE3aDIc
ny6qcF3zAIca5ASffhoRTkboJmJ5/Y5FTQfy3NTBvVjD3uMrmogZukzg9zXd/A1oz57qrJsHh5C4
j/3I/jN3DZJ78Vwj1Lhkv8NkKMKmxKt22PeKeuC+qBjFsRyPNXXFwYxExhS7wqvFB5+NKdQoKhlS
/wirCpONwAyDjq03dZrTyujfLru2xnX1fltv/nX94Qcg6BA8d42R8TPGQLkYWN/S8Fm+tY/Mi88R
QEblAngZCzOuxv11VsMbwnL9YszAWdx7WjZch86eD4/FnZMw1XFBaBoZ5IsyxWSTn9aVsEYgXXLq
bIxQ5AowH1zmZKQgG1sI65E9nagz7BLEB7bGgyL3Ggt9oo5QoZVLLEh3zApr/5ffnANvtJKszVFe
Zx+I1AvPUopivYCTnly1tFBd0CdRiEdhvN5fGSoalR0wEIWe0TWX3nNmO/csIFGm9fEsSyb6al/Q
Mx8t8f9bS3fktaWzyiuvTnMwfA5V1QSjnjjbuDxpmY18E38ExeMZho2JILMD0L2KxX43TmJbCjzC
aGuc4fMfT6GxetbeKd6qqGitpzY7AzraVONzuf0WeVUTV63Qn2K8CovTFVx8+ZlVvM0kHUFHCglk
9IAsNw11wr5W++wwdbxJmsReB1xV8to6LmdhoOeR/BlsGOkVsMbNbOvShuXuceNqJHVH5+/Bb7er
uvMbJJkQb1GwJMrtTq+I5ogw/yJsXXLjxkFie15bXxRzI/wbUp/eYlLa2OY50x0drJdjatssH+0l
n3UEPf6pQRKUhrfqna+6fsEh8djgcHrWRcl72FgOzY+l0ULiMdAek7yi5K0jp88rsr1Lns+JneZL
0ZmVTk2rDl82FavKAuqZBFqvHaEi2wLoBBeSY9/wQewpaoeBXlMH7ZpPaK1jckNvXLzLW5lS+VC8
2Wz8eqswIRGq1iLEHqzbuhumW3zAbAmpqcx+vCeVhdyr4YQIINyCNR2PnoGhipmViajKFqzjNU53
d4FFyI2lPxb+7qviMFUDRZipLiUoeCUohReyZgZxP/9Ir5sXvnN8Pd8vL/tP0ov7+dK9y0LORcT8
80fAErRBN3qDfZjhyYv5Yp0c2T9PWWhklRRLmlO8MiFlbaCpWe5Nl/PmdydAetE4UGqnQXr5T6mk
D6vw4JIXL3sgMp3c/OT7EIwusKQw75A+kzOXBbFLEFmU+8uznixdjgbxj2M+P4PaCD9LbHiiYJwq
v5Sw6MhEM7QFGIOVSzFzQaTRJW5hH5om0GMphl+3i7fvy4nkM632T7JSVCOT2C/cbqWDr/ShLNzJ
24gmdOuCwIc5vSME43xMiM2O8/DCwYUQw+hI1Trsn1ORhvBiuiyeTPgYA9JLdryiEFOVZA8sgJi5
YdqfDKz19zibj8pGMx4FiCIIig7+grEYSK/SXIlYTHFufklGY9fUz0SBwX/npmWD6CB5dWPRfNQT
nl358POCfTADXTNy8wFBSXFkvjEsBUJWU9UBJamLFgmTS5rcoklH+9tlMrnw6B86FaOA6jhbMezQ
euvlt56YA3Pom5Y7C3ZAcxkff2UNOFEqJMxMssjSm9k+//CWJvuYpI0DkwSwGPYpGFEtZ1w38yeH
8fCnU1QS2jOJnS9w3tbh5KlSdWEa16wFEqhzx/nMK8CZJ/kDDXUVNgEgI3jqREN6pIuspfV9nMEU
nP+Pn++Wlf5PDNQafrIoEayU4cKGJAyeCgzsokAQ2KBhD9nUsqcCNmju3wYWI8K+Frz2gcX+6RD2
eqcL52k2iVuxTz0qTEHRS2ymLB4mKBlPCaJOF62feKLoICmdGPD8Wgn/BauUf2zNC8Gu2dD0Y6bL
5Ex96pU+7+yoCj7wNAosxP3LjbjkjYG6JzbVtC6vxatCHwgZ/uj0Z+AdNX8GzxzuiMlf/Lk7HfWG
drb5FaAjF60Rl5AaI3rE0C3zn8D/jqsdj25Zmum6OuA3AQuLr/Sz0TjFLPaR9X255rX2bmxsmyJ0
lVAJYcQSMlTDg5dv6MVx6oisjhOO6kBoHkbnJXBggKesyIPVW412OG6Fk87Ceeen06D2gA8gylms
Awl/Q/s0r0EDPAda2HtvRpU+JSsD3X3euYWUKV8fwihibbl0NYjcHb2FspcWgzaCj2zcwzqhVwTi
e6Kd5uUZvKNulWB7GwYQl/BLX3kSYLUyYOucBbS8EowU3NCM4NBlgGWvzxJrsEfLOZ5DU3VLPU2Z
gL6Q7WFKpTTeIbJr9HURv2cVO8zwMiiXofvwzezFYKYRP+BmVBM6lrIiTByDsuCqGXUT5JSWMXpo
lcHwe0nEPKx2HhwUkYAKZ8deqcc6GrgOjc9IgxXAXzrErKfvyTNtzlXXM6ZxUPD8EHeAPsFAoObi
+PxXuD0h3/IirE/NN+sK+DGt3VzFoCcvHP3qG0PbEUPZOiVkStteCTbPHwDNDhy+M5xiFL/6moPc
0EKor8cKBuFG6eLXZKIBWsooZeEJzfULsZ2qyHVDQzj69nE4GqSF6i3J329Ug3aI/JBCY0oVPLpR
EbRoXMQOkyoTjG11gogVnXK3nOXCEbaq75dxYAWSPqb0T36A69kRobvolGm/YIMQ4SQ1ihNZqTb5
F4W06BJm+xGco5Bo3biu8ScA9YGLg0fDXWfxQvKeyVJ1kd2n+5jjdWAmvAB7MgZbMPiJKg0bdhcB
t6rfFWuQNEg3Nx4QQgY3n/dGyAt+pGfv+BWt1THYy/zezjeqJKaK03lMvxpEdqWM/rnlJfgu8gjH
UT5fMWSJOW2oCJ/jD/Jh759eDpK0odHEq1uxdZSjI6bIrJHw57nLTwN7lpUACNX8B/XTo9IW+6Xy
Nrpk4YvWEJKXAfWXf8KbIiEDgO/7ZN4KJ5kYoZ5A/V6WN6xQVOn+JeWWAwb65pNud64IdxaWCJ7g
Mqru7+x2yDSwXmjQoW0+HD2evWCUOLbwNlWeCP5cmOsrPU4pJ6FQN91x0K7el/W/qSt+3546PLLI
/H+CzaZ7XL7YQV3x8hIFFV06sI+37eFQBX4cc3KL+uwFAibNxTut1PmVdN4nf0Xi/IzMskcb5+Ry
Fc6/cnGUC4Bcj1BFv8dbrjV/IVdDd4vQqQ3pt2Swd8Q7SOqnCvrDaiZNQz1Sj6+0+lB9vmfK7OBp
C4aIIYim9B+AfkbWplGdPMdZJD9XNWcmda/yXE/UdPhWfY+IOeWVuSbHFdQ+VxPQAN7NnhEmMJWw
Zc/rsjLlz+CUQQR5F2aaKjxVxjJSWwVC8s9V1UKaPnQZtce+FbfcrMdPyNPjJ7V6e7z58qNpH31F
/6tXtnHdCyCQPXV1gjI/Y/uuENOVeGA0dX+FEkZuqWkSeGMjQTauiJBCKO2u8U1AQHu6FiiTqjvb
qiKS8xsWnL+teDE3foA+8sSB8rgoMm4Hw1lsmNCi1XDr4+4lK+8gwWPpztMYeRdx6QVZNShBp+59
QmWKjKzpwN6/9gvrBJgruokOqunVcUNi82J4st348yC2ZiPjwp1OrFcxaolXMkyX0gXRGQz25K4a
oBPhEO554x4S6pI7Q7YCdJvTW+p4521st1hrWQucwOhYLwjkyFWH22eflxSfdkP2NYb0vncU1WJM
s4VRcjT2wimGU41DbdD2Zzodi55/MqEZgQslf9OyIsrQ+xZnEBr4F0QDKGd/juujl3CsLadSfuAP
P3t0/s8svakXjFSjVO9yTr+ppcC7W4sBId8N+qFwig3XjFNOgEHMNQEnXAEspeFRNGGMoizvVa9k
qoFsgoubNiy6sf+OU2IY6B1kBLwzNIGJnOlKxLCYJTLThHnznEvq/Bbojx9ahsl2Doi+kr2UwfS1
mIQbGVqIso3q9LYo6wQNDLzCD4QrLDETSJkVeJehlcOs3WzffIhDQHE6taDOgcR7IxYChUOnYZEX
XioJIq6TZZ52V3gr3XB/5XwUlg34vH8hfq0g2t6IXVEGmhUCYxOa/h2rh6ni1aRDpLUwBGrgKdkc
o8lkxe4mUhmCD8d2aL5lqzqGwusTYbDihhm/i/Sl080GbFp8QIk035Kmbmb5BdPHV+yn1bq9DSR7
TttNzXXdVgnRAUVISW5QmKBtsF6l5lU5U8N9qj03FpslPyfKZxyZKkluA8vC7Z+tc3B/OkQK9wrM
albRJkm87alhjJwgJ12oh5s2gEJw8Yr+eUCAnCOCpA7dUEKB/iliCBU1DFU8kCM2RGaJFsDevJhE
JpPpF9Fu+gg3lVM+B/Flw1BXDXg6Wf4PnCOTcfjUdvw4HlRtYLPxdx2B/CjWI7lTbLjAq6AAwhlE
Zz5Rc9j/F7e9Muj5oQL9NKhD9Sa7maoGSnmbVrkiLlCaZt7SEJm5+iSvXxSKSsiXlfLmcHbx+s0F
foKkOBEyvxOQBkARDKqvl3QrDS6bOpcxGfVZC61BZ1nfh3xbbwPjZer9D33zROxi8VuIYYKDcXx3
wCGnxFZEsgWs2keH41iOw4YvDLdBMi9mqtfIOVOLtTyrDazVCD+SNSyXPsshN8hJWBHbxjwd3GuL
3i/EnSNLSb+wGvyErd2LK+ENP72SaltxWrKrgqRFkit1VMKC6zJ32PzE9VrsFF4W83lQ4hnEwi7N
nBTLRnqrFZ9+vjTLtVA/0SFM2SRCbv1Rl3MOWgelvyGmQAS0AHrmtU5S1sWIILtCY3hQA2IYWpZj
rgi1mjCLh+WfHiyHUOi4a+BJRrPItG9QrYJbWei48iv80ReBE/xJpxuevNsqMwXKMM5U773GTy8G
6Ejl6qgUb5EWN2IrSs1oroRarcdQn0RWz/IgmzwTkmPDylUEfANNzSumMC7mdx+WmTY/8XiqXNLw
3zkUsQGwoBcPzqmA8CUxe8NnCBL/469RzEkVIA4k6tqsQTeU5bKB7aWxrg3nkJ5vFZq9fcBBiMuV
go69HyQE0A1GlVYy85dxkmi/yaDwhRXk3b+UtQEnMxKstNV8WScbT84FgD0IqWSH5f/dXSZawSmA
F4zq1aSETvij9FsdaK0MU2Un4whRW4dkD1XACk4gb3jqwjVdwhHlArciGB9z2PXElROXpGueaOIh
S0llpEASZT70Y+0mYgwVyww72s2UofMlHlYz3JWwZnSKmST2AkzIpO3VH/Kdkx68XV+eOe8dUeyA
8hdnDD+ESXHK5ur3J03BSM6ib2bsBw5c+Lxg/T1S3lSXWvAMFB+IzwrWGnm1+uiOiCTcr8+jIjsm
YsFkPoKVIdY6vKEEPTey9MaAneR1tCdg4f31Y2OIS3rEPk1c7JwBB+44F/WIakWMPZwBZdtmV4je
O1o03VnHayLoDxXnebb9k0gCF6D+NVrkFoLr62DiztX1BzAc7iWm0+huqfCjZHA23HLVHizsb9Of
dy4F2PjWwxHQD9msad8qiBRYb0FFtH/3RfKS1cIGEVByPh4B1uy8zOt4dYw7CI9on6+qH5FOJgF5
WfyUAd602wt3SzuULc2Od4gNZL5t42557ulQf4CfHvjAQIe6CgWvag84j4vPKJUAMCwHZgRT3ouK
bPjWzCnqzXBXzWMTKiQV7+9JIFpbwiDWM+n1NXHc82+4qhx6aH/lGXG62zFrS1u3huivc+FNH7Ys
42VGTJBw67cPzJPQ3pflyg6oPErxr5N8ua0irTjHJ9ZdFRvFx7uokk8QePeswL/0OGtr3guChWxL
uSaw4mEaR4IHeS5mpmpHHd7N6Lim6ZkPRNFmA1O8yA0eRxjbJKEz5T2kGPxqmFzV1AN312VAF1GT
ihbewUeorlL8ISDURxlSQTRY2rWIynLy6f9SGp0gvhAhu99+Qjon0qfihb/TnbaBN4YA4Ce/r5ct
7GuEW7pSH37ILUBLf+KsgSxMav2zkQCL9wQk5wzXx2pX9OQOY8FNkVVEfVYBOHw9hfj4eDLvkjF+
Extblb35cNfsCR9qU/dw+Qry06PKdD7YCfUniMMwXf0WGZiann4AcV0vB0HKwhubVVTGF6ziC8m6
uAYuhH0FvAyZ8j49641z3+mT8KdA6DWFEdghPTIoHX1A39T1QpjMmFWVP6YXhfvhHznZ/Mgs9dfd
9uBMoNRWK3bANe7a6/WZBfbaGdf2IwHdz1wQUfUCli1YlmVqMM+rsjcUjLHKpWXMTpDcrdhQWTIL
lteB5Jj5c2Y5d5yOnT8SdQPpOr7wwgzob8hc5C8amnJo+BM0wkUHaGUqQ+0fJ3SmOYwr2LIGKbmx
RlOm01WfzLQogNQITN+tgtylAz9+GbFTbfOOOxWy7m1r3dsLoZ4im1LpC4X1MujDNGyk3uqY4ain
CwaOXk8SCTBWr/YyQgcIvZpZxko5t5KlyW9i+9lNbFXUHrEguxiFSygJ23aIR/ZKfIm5LXofvZSe
0UlutOYZ1kibec/LICUxe9/OoVqtSZ2u8cEQ5CugVIvEFUFdQ3JKBMuo4Ohzw3J7PCA6ARQGDEWO
GoPljbtKfeHGe1F81a5BL1y5uE86dcZtbdYx6SREWmHb1WspV+IM0BjOLBF8BBmWuj33SLWkXbEz
2rC3YPO3OkSwpisdOWy4BsX0nTqrQulvAmI0pM4xqzqcYpVX0CXuxoc7Pn5cbQ7bMidQdKE5fmM+
DK9xsQLd504Bmg1Ah7EFgZmKrJeJfn6bkpbcnEW+GVIQfrw92Q7uW2+vfXX4RTp1REnbk+2C/SWd
pBX0rr0MUylNApml64/FkJkrfi169eTbqrLuDfL9oUQV4EeGgV2B0H2EuBlk5wPMmcYXjktF/4r1
gFhgQ/KZQaSolpcefs3y+LcnBlaD1Oyl6XuhO+Xp1/GZiw1nx7noSR9SZeh4ljmPUzdlHP7gzWMq
oXSeLWXcHgDyLypCoShl1kv7JHfwo+x3GSc1MEnuMb3YozeUA5IMY+cGQmIGppjfcB5HRBTuWD0E
xR8byyJELwRw9aJfphmTj1eXFetgHNr2JR85KLAal+v+EfCIgNf09uyE0skqODu6l1R+gMG7CDxj
eDrambkm1XRyZ+aZdreKKKf7L+s2xeVm594nflnn+kd4c7wk76TZB5uxKLp1DGc1YSdfqd0pJwaN
Jqvy+68bUQ7WlC/Riq0jYsfDHFhjV1RoHwTolfxY3Wk51Ai8PR25awn23u3pZXiLELl/dKY5VdlN
GQ7ibyGXnutKeK+KrbUZdeC0FlpqECru5VmurKZQTFEuTHqcDqfXqcAjmSGHRUAam/pqudduGfhn
jK9BxQcsp+RheAybRYeyZpD6gE7cfXHUxMo4UW3RUYIHaxnwf9+gpWV7Y2JImPYI+l+eINNkbRGv
dIr1D1Is2YfGaPhkQjwHCsk6n4Z40QVFKmAo94Dt0oy/G0Z+vL1X/m5Z0ktIfGVTSPH593ei6H8X
d9P8HDtvpq7rub6BD3Ib0LeNEmf5oKBMhy1xUr+sWnMlaxoui9OuYM0zvakKUAkCUdLkH6OCLlCP
tzJO4sQb+mMX5Va/gi257ETTNd8vZ7EJH43owQdKEOkw/Xp6Nc/RU9u0+zC4fVgn9tfbnvJTs9pK
A1OaATzlz0WRzhHEB3ZiOUCLt2z/1ve8Lkw46+P4nMI9XALXGFHX2wucUtXWFAk4XNSDxPn30QEU
Tysp3GotZ3uAo1EIFNxWELt9pjA5hlE6lt3EFes3xFMhoGIO1n/4PwccGTlbAkMB5m3Rj514+mss
72c3jRDqSjgK116rKvG97SU6EMU6TNXDUF0/zDJ61yKXHsJfKPcMS4miOXd2FN9yvCNM5LL00A4+
xsL31X0t0yuy4ma43CKfJWiErdNMx6Wnc5R795+iQkDiL7uphJPaTdq86YxKP99QQCKLvMtnHE4J
ES/p1Lmdg+76xNNLYCtY9oYsztMViJHShH6pdUqkWHPOFAghG5VB4vIWwqLaRY6BQXpdS1FvOJIW
Io7h/YdlfVbyjxQI6Z4IgtsqXowEVSqZli5rJQQozQROXjpf5Pub4QyiBNcpWn4N1NtRC5DANoMW
h0Vc3EhzBi0Gk6nAgSva3P/unSJDZ6Nt584PX/j5TV5zT6dkOeLiZVF7nfmGcskVaqh4vvZ4YGnl
ESeXJVYV89grb4mSjApHGDRWEp32VYbQehVXKczDClMlQ17m8gXXS6tSMJglxO4jliRRAbYgTNBD
UtwCZBrDNNySDvHsuUHSEPxn7Dzdljob/Aao3QIm9L9RLAej2pUasWwxJGNIjw8TnYIrtwxzqciv
i0A3Mywd6zT3rI4GIh7G3NfGbvsKlASL5bvxRBD/CXZcWxj6+/IdDXL250982GZTcGC5UWfF+IBp
cpY28bRUprQBK/u8v8DNqdA+62VtuPGgY/I+az/te7H6RUHrAHzis/u6QF3+nMYKFW9mBO9x/oE9
rGbxuCGtetRRItZOhwvmGd1VGJDWakpRyq5DCbf4wlm5ICd3qB4wBHYah9rTECTnQTXfkvo0cW/u
E3XiElsBWk6/02bgM3uzgzxe0nNQW8wFvH1pr88AL/L8eKW7bGUpex5i/lHysjc3qO0HHrvV0RE1
jTyzrtS3IKB2Z6yTA6oNZfdfNIUudxhsfs5cgRgpmCux7mzJhe3YKJulnG3F1AiIzx2Y/neHaf/v
6otCa8USWdvi+iOAs68NoE9iG+zxaUCMgLbiaP6Rq900eMgL6P0nQYiWtU9ILZ0Tq9Tq5BDHm+db
HLgK/auyQWTn/G69UvFyVU8AwNyvheOWjP8AkhCdQJXa4giSwf+vNJoi9XhlghJ3G48J06/tgEJZ
YdHnleuljJElVrlAI2T23OwZHvIXhdYKrDgOMNVyMM2oyw1lIN0r212ffx0xoTEIGU3Ox3ohu4i+
8ZzK1FhRNNyGcLvowgHUvPsHPie67MVVZG8kdhJATjYzE4Wg4V0z3yISNaoiC4/QPcekWZXZ2OXa
oM3e7i48PQbV3bqC8gWsp1fxUGs8hvBOEwWxjcitSywlODSnEdfX0DLz7M4I5msDRuvL291UXhMk
mFZYbn38poZPENysoMKaaub1v9I7ZL2qVoGv4kR+CCVzECQ1eHQlsYRMosLfQQccPxsDlbKIHX/O
+XyJqo8cI85sYBTIVSXSUIPygWKdx73qeMEfwjGA95jKIikknAmtKOzmRBmRfT4r0bNgz74k1/5h
rbpdgWLeYtCFz2a5JqPytdP5P+XnFzLrB9ULRnJwt0G+7zSS3n9I4pmQikAkuBq+DPj0M32E4TQJ
1fEDJfrZfsCLFAmxE+A4XyjzVPblJZocsVVnbyT4VSlLCs1PnP5K/VMcJ02a0UUuQIMwYmEBwQfs
U4qIW0wckoBw/XowuytG/KpwrzOd11d41haTjgt3HD7bxcB9roMjI7glmWjw6bhBGyjYMlWyaEAH
4A/bTfdF3T5/Y5Vskl/eZyqtc764+GIJV1ahTheBK5UnWv6XOLr3VniM6P6/5WHUnVHPoYO9orVe
gshTN2N55Rf24amQ3wDazn/V02jJm88duJHkduyAY9xxSPnNATi9AepFzwUa8hapPBLELLBf+RQj
QPrHfNgtJIwozU8RAwpEosWmeiEOcPReK+YIIqx7UMjek0sXUzj5xcbzR06pnjqaYS9znRbt6Vd+
j3ZI0WnygKxJUQH3JEDcAT9EZkhV3OESgH7ZfzLZ2ZiPrD3abmleSG+CvEUy5pj6Hn1dynvV+SVg
+Ipw6npjZPETzFlCBGbdOKTD0wsITiD/sk3sK2GdLgXQ4dFC/CTzn9O7KkJqCPSIhd08jIaayn/P
gWWP048Pem7T/lCA0YC2qbKLRMQ9AHcxK+4jUbS1KDs4oflZUjyv7yNCp9JBtL5qTQjlfCw09vxH
3OA1Jr/P/yfgasre8u4z7RBKhvs1Nd1qnoL5h8LfibvF0mPaIUUoyxt3fBYJukDeNq1mdkPLk9Cp
qcO/f71CDbis6NddEEV1C99+0uB6yb+OgnUc9ls7R/U8NvGVE6J1ydoufRPvbbwKaH7iXAoKvxr9
rMSixe/vpaasb/SqEzAR0WwPZSXGWuKIEeTWdAqeGaGKSWSHVx4jf0GgAMAi3ifXqeWcWJO8tObW
Gb+v/tbgNLeISXJ25NxUQovMrTFa4fGMXkwUuwdzM1uJa+qohhfXIVmjpgG7YMw05YAb02Lw252O
I/2dP3TvMlJ3opmk+HQc1qTjwZ//1WrqB02YMnMAb97KlJ/yYjuN7V3o79FlGmZXWJO7mTVJoKR5
mVzG5iFNy6Vra97RcScHAZvyPMytm3SoknA661L4PM0ajCH8Fps1VL49C9+M0fBZNxUMk+v3EBnh
hy6+7vomFCIMglu3Gd05EBUBu8VWFu/2TXWoOJ3m3z1Clraqb6Gl22HNdsq8dC7tcxNVJ7kQWhbp
xIkMnLah+5B+hhH7Uy+LtE8/8dVC6spzd/l7M1rZB2QeumkPCzdYhEc+ZAqYedPZrJ7nYh7QFjOP
8H3Tzt5VkwNfoDeqyL/32e04+PVXLLf+UKrcKEoWl3nmsyxE8dbHnZpnIPhg7WfELljVHtE6PshL
RCm0SsPePg6DsHF0uxZ15GfXWLPzhil5Vodxd5+Io1406BPU8OeUR7sR8Q8AspA+V4PtC24euLOl
U6jtX1Dp5/TugUhYVocJecwYf/aUzDjBJMi3EuqXMCiEHLif8lRultg5eNUgWPyCGCckHkKRlp/p
ofMcQE3jTEVoEhDCujtcnhd/DzbMsGQ4vGuVBj3joVhjSXYvjjJ7tGB3KbXhqUOkhJrjNqbiQjzS
G3W25MAGWSC78MVHm88ExAoNRXXVkztY+1E9Q+tdKT7CFmGmTk/HCSws0K1Mua6YLcuBdJOCM/cR
I5eYy9jrfrf7TB2jOZo8tzz4pCI7KQ7X4WVyDq/JFEv9r1cJ9gZTUVn2tQQQ9pt8cUgYckqN2Rqn
0o09TZP68VBpeH7843efhhSNPqu0en9sh9TPOxP8njeOZP1gFbFjW4i7izuOj4NN56l2TTCqA4M0
3VMn5KY/G28/tCvQqBsqAxJicW40X5yK9+gbVigj48MEy8N7gpiXVUcSrUNL1BriyB0vB4Yboj1v
0xE//oamUWK346st6zCHE1oJrLQ5Jj5Xt3V8K+jqcPChQkk2krPjUrXKwIXL5fZHaePCjt0Pw6M9
b9dygL9dlpfmFO3IYnHX9fhcpal7aozhfld7cIO1GCrXZiI/MHhAY5mJUppHPWhYBq0/uEkRhIUO
hLKuNO/ldnevQyqFVRmGdbSdiz1BcGBBjNgblCX1D5VyUqS2AabW+WptnXtCEUfv52+0dzj4BlBC
+S30rOTX2whO43jcLxicSTRsSH9PqweRCjOzNVlwdVsu5Ldqax8M4mgHmvEDe4yuhvLMt4PG7RUU
Ldi9weoemsDM1VjVsb24MOfrEL0Ll+rOzEWULm81MbHQVQSEZf0tSRIDo7neemIDvFRoqS8ruwQ4
sK9Y55jEusMgy4au8tdaSOsuImqnXZLMUoRIGfsWvrxjiYkbREZkQDg9PZcaxczXHox2+iklnVU5
1pqZY1UpDk7MFST73bRcwjyQh+BnKW9XQ6yZAs438rDx/CqfxGHjS4AVhF1FlhdKZonfrOA02fud
P4Hn/7FsknygSDxpfZx7CcmR2hhwOGVPiy+H9l8NxPWnhkWuDY0OBqqZf5ACtxGKtj7yrNkUIniB
SDbobwr75LHcM8I88pmLJaRl98uJPFc2hoO3bozsntKOrUDO9xKIqRsJX0Oml/3upWqtPH4DHuJM
Lgj6xHlqGqDzfSNGTgFIVh/6Lt7DwCpUEYHs8gnPw3AA5Mxj/gokQ0eMa4YfkYurbztCS130BkdR
+wIFXb+XPlztlMw2iwppr9hFiProZTBgeB7n0WhmSCyeM6wnfP52+iGafByX0sbgdBtrkrtjoj54
539S5NoEVJ6YfcsblyjS07araxnR/bnJgAL2pLEs0jCt7Pk0s73azK0Ba5+uSm0jdL9MVFyhSqc0
zTO5ETX4ArwJiAHHDY3I3e/VVW8TSQHGh3L7agNejiwubREQYfoLlfhWdMhLgp+NwqqjQSuOzFlY
D6b0muqZaUeZFLybAD8Equvy+nqXxNbwzB2JL1nqHQj6s5KAY2tUPaWbEOlkyZLp62cusDt8VPlq
xBIftLmQYuBlp/6XhxZcRldNLrR/qMfahDgj3lMWbRVBnN6lK/t0CxEmibj2ToY0x5gYHRom+4T/
wj1Z+lEY4uTBA3DPT1asHtJs2xwrZIVW5bjk2LMYnoSAMnW6GFXsPPPJvI9M5vpUZOjKc/uX3YOS
m4ayOs/b4PsYKHPQtt6+PhSmwP1ltyFbsm5PEEg8BICjz3vwTTXzwqEOZG9tiDu4LYT2fs7i/kDu
E+U7f4b7P+S5JnM6Fh6i8sq4Xa4nwBovgw9tzSgMcFK2e/i0GsBDfdJLVmEO62HgWRsYVRxm+2jA
/ecf8HxIsgLj4CNgyYRallaiHbw7q7pTpNxwBUo06WLlQjh2zMAx+vJiNknk70P26QutoWdSv1ZR
7ZGPkg0rsTi1gKNlkT8D4gMgpaGszS2Lw1S41ebITk5ZHmM/4LldS1GdoefsLzJKetaf1gCL3qjB
u5CSod91MyquglCGxVFjeyu3H3auiy2wc15D560szVw9B77ljA4xILYPUeo+X1fQrEq11CyYTENX
Xx1C/9r8/LWAibYTHOHEIsPeKsdF4ZOEoo/Z1DddoV8dvC0li7Ts73yv47C5Q4JyR6LoZ+uhKXGY
6eKqUBD4kx8AdoVHN6ADFRStzFEXoSXi4A9qyS/Q1MMhD9xLaWApmU5On7e67WLKs6izQmkC9QvV
3PTatJzhGpxnWzqK4CpltDRGD/RHf/+9337omN8EK/NOO2BA/Zbp5h831/Qh02SDeDKe1ahZSXfr
7i+QGtfYsW4x5jS4y6b7unwPp5Sr1NYAYZ6WH6/sESz28Y72K+fZ3sLhh5Z4kyH6K+mZT9KLedcA
Tco+gHfKoeIKf8d7L0J/v6VDbFfiFZLJ8LfTiU0rA97iKlzZNrV8IXhydkv3hElwZAaTNWDCWmeE
nHUsOOexDYKA838CMidQpXtEmZNXTDy/zCYbcLPcONMFrv+yJlbp3V9DjaPN9OHQlQ4DMSKVrbr1
qLUmvDUxvCb4YJ/0pGztknXPuUPpy+NxTUB7DwN+ZnDQ08YA7+h6wcZqBI7Kzv5Bnh6jtvgRDVKG
GEA1bYVQhckX19AYgy9TSffLsxfj1ZmM2UpCjpiMxjG7vFRgHTOeLf8mhwnvZ79Bn+aQY5VSy75e
BKMwNiFK3AfjKluee74RlkCNZ2o1qZMv2AWkyFEebQVjbZJQJBqiSYRfI6hsP7GjlslRn2Wpdwml
SApn8+JO79y4soGOzjiMNz7atCqDW2PQpgkdyKcps2qkCWG2cGlhksrCAvQOe4QiVKu9qrTEK0CH
X3GGyFJgDOPltqcAJwj5tqc73e9Bvd/3zCNkBfOoVOoZ+KgID4uNmytlC7sXEY/EPsDzIhf+Px82
7VN5OYV/Xkxc1b6TbKhwp8wXhPHcj2CskMrn5QRIUkOQR7WTH01ROHBglrwurhgE/fBoOxivROIN
Z6s7nojko1KBsb4KPTwge0qauMzBdS6XPuxx9of8F/PMGHtGTws2cDTSU//BFF10Xw9ZjyKx2771
G5eu9qvvalLZRcXwSK7BQFF0limYVuzbrYps7MuKjRlTN9xkKgnjgtMol9RN2Fh0N2Ec1UHf66Gw
KGqa+fzNtKUDv7kX+wNlB72yg+mb3PFqH+B6EligxYOye/QtiX2bQHIqV5oRmC9HNfJMClXgOebd
//loFe5xUYhXnZmrlgOsoNu4S+02cfcyn/jKQxv6wn43tnfOp3/Xjt0cj+bTTpqOe+VuNtIN+fkc
XWddvKH1LAWZEFvgmdvuzw1UnywW4F6EoN3eLMNbrT7f5Q0BIhBvLTjKDvX7wh+l144fptUdxbXY
mcEyGSUp4shu63EUh7mNZT+RCZo5ft/p+2oMXCtQPwmiufBEvt/jB9fcSe6w6hVjKaTm20GK0jpT
LCAs6iTR33arvvVjBxrlc1OD6lJ4YlGh+60avAOAWc39XmM8Nk0ICajyNFIuemXAXvpjJETtIXhu
6WGcxUMzzSa2yJ9GXR2wsZR9ctD5dELnqVtXiLfI7WQ8U6jtrGKQtsusjZDTY1UAmowzZttpdiVw
8eVRgtWm1uFUxiq9Tys+EuXGdVjOq+saAJ0yZZcVV+3alggB8xPzQzIHQyhh7wi7HQ6dxcBNwJ85
u/sdu6gPqW6DsHmmQgptLO0kFEvck2bfq9vu0t5oEgbDD9iyOX6NCF8dJloMnycMDOv2vi3sRJvc
S1D1d/YukAPL8xR2YNYDwesa32f4iwmpy6KrrlAKAxrMPErolbf5A5le5HOoe7Rq7xMTr/nPkBt3
umQ3x0Ux49nxP2CPpm4K5RNa3TsW+k6czXK0dMWS+KWqFMhzvvupQRWTpUFeztB+irUMJPHOpJFT
VFRnqCclafV3BxfCSqcDh7luOK9uyPyJ2slVpSRQPYU0X7zTVlucgI77qf9j40IfykwN59U8eUs7
IfRW3z5A7i1Wt+naSEHhxdch1YTIHX7NwqkNZLR44maMbkJdCF7uJ+RSeiZguNmV9AuluVDTZ+aw
0wzMIA1eJomDCS81DJ5n9kc0d7eQu6B3aKAXbWm3brYjxkpgsi5CbsdwvpFjgOCK/3G1Um6Q27nR
tHpBGcbuCfrOLu4aipOk8ZiuKRXi7QQzOk5pn6lusBvLirfKqw5b0i9fXQ4CnOAmnfTNulXhPxPk
tAv/6vBysu2WpjDt5fUc1Nhg3feVg4PuEWBcOnBqTt42xCj4b9H1VxcNyC/twMJHkVtV+q8LD3Xx
PDrZ4wri2hNX2wQByyymSShBVweKgwAK4SJyOxpR1ouOPNnrzKjF4st7m7+NTTXw9JndMm2Q/6mr
yqh32e7N0by8IDj5eD1tW8hVuyfRa+09qulFuY38HhEKg5o0Tv6DK4po/8tzqau+EOOK5XFDmldq
Oep6+PZLbS6b4/NE4GNpa5/8pAiqns/ZYOaN4iFeEKLuugb2OqJSumjneS6BI8pp228vxQTtT7AQ
zzxmpEvQxIKFAxoKji4YHWeUT01pZHx6Io2bY5Uf0Q7Kh2VgIAitNx9SGxebR4GsUzcMna3L8NoF
LFeCSRnkDlWJOkUh+fjvZGK6Lm8FHoE/H7/FnhBtW0eGnSwNMqNIlzAniKhQVtz3LOV2u8eZ8xPH
sBMAXlbSmd+qFBHJjn+/eqRO28rNUyv4V4FWemj3P0K3tF3CoMhpJ50yK79jgtctgOznC+WNb3PC
K+cq/UhzZ2m5yDZKOx04Qca42rXecMMiM4F/mbLhTIH8oFY9p6bAabgle5/Fe31fWMBXGmWsRL8M
mK9hHXGmRnz9hshsfyvjnTPT4DiwfEW/W9KhFSE+f2/bZ6ovuiJjNKdsfx9mogs4/06pWfZzt3Aw
fSn1n1bucQ2OVrffmd0KISLkzJWc8ZiVkX1U6tWVKghmuG/7RK2tGi4tZGL13UOe851Zww8pjxTB
9Wi69HKiv53caaFKfH+QNjZAH5tuEjs5Uk8BcwAUhSdPpEqXhcHIgXefHcuHq3bcMe8WOtobl86U
YKnWwvsrWhW8Zog3OUPaIlQ4hJMnfc0Q07QFHLmK7klr+WGykop2Ayh6rQ+qnptUxr0HVTt/+kkA
h3Q+WZ+LaRgpZdDEb9ckCSmSn/M/DCcTGMXaLAxsncYBKpP7ow4kwy2zx8RsiQ7VrKBUqEEHLjBH
dRKOnx7o5CGIMuGGgT8Zz+m68xJd5Fte4lASsixKcOkneIBUuSzNDL7JtC71IFE9AXrEiu3es2dq
jUr9TAsqpeArEVZ4T6IXZrOUQlm2iC89eK8t2znsbEcv+3Ew3zNVR68LLtneTCGy+nuuav3QnNMP
wJmwRPMLaI/xV3fzVxq8NauurRQuZPzvWrW8+byZsPfxlfGEocYdIpFqsyCKrUzEhjfjGfEHrKzr
8mhC3J26TV1ELHgkvIOsbjLEvFHWMKcL06R/R5ZMqrMyrE5teax7wXp2XPfTT47AqdUcwkjVkY7Y
FOV/lXWS/R0yEx7O454Q3/fPOMvbvgen0RkoZ5/iYbeohPoLHgP6w7hsZSCjSEvADvF3uI4SSkYl
UCj38Ry2ntaLhC2B3o2P6TFLGbVDQIYr9tgPnv85QopkYTfR3NktVZxMMfOlLHTGPHlv/EE8rESM
BtoZWMu7T1iRWcla2GjyaKlcf88Q2vSf72kL6RPYcn/kidVfbeMkT7VOMtENRexupU2bdB6Lm7yf
9NZi+x6pAFm1+U8hd2PmVQyc2jGSQYsDUB0UJdgU+H0oZ+WdH2/rLgVElO8vlBOCe3LCRvmWt2Kz
8+VjOcMs4c6BE4r/GQqEXLd1HWsEcEDUDtldldmRc3x6HvgwY1bzRyl1vrbcGocz7ab1OG674gw5
0SS6K29GSWJqcqZR1pb/XMEC36aPfJVYsZDnOuX5JnYRBJs48uxDts1JVYyOuhWJgnBLWzb0yJdO
IpH16nDXbInSJiJecgitX3fh6i7xlzDIrAI2syy8FPftvnYbCTqhucL2Oi1m1Tm/CxasEWveUP2t
SODWXLAmSwbWuVJv8F8vUd/1LvrbIPLkzbPWGQ2+0n4gKJ8+fvK1ATd9enQ0TrarOldE0+FocrIj
axrU9HN2KoRAKnJsut9UiZDNaHrEYFrc4LF0UZIWCzVpVZoeRQ1bHZ4zBJTB5q4/DB9HGfoafPMu
KyGl/sO1sfGIvw2PpTh6+clfR+xTT0BIzdB4WJlRhkEJjOFj9DnLYPvwxdSgTzNdGsx7GxNNCDUt
8zPQSusAqLm+H63KOVKHGz+LOOzajXDofweNynyE8cfnBGth8sncvH/I/OF+ObTByl6LivHTM7uR
0QdDQaqULBqf6Fg6Hv0cSfKMIDn9HfpORg2r6/m/f1EU4+4oYU6bc+izVcyLFqGHDCwXyJJ9B/qh
/hzFxy+OTg3YHIE9xfc0b5ZmpPNoJmUC+0t6t0xXHsb/lE843okIrhEbVs7coXrEGNhoW17OQ3/I
T8HPQwlDvWcs0t2Ctj/RkV0j3+2V6snp6XBLTgL0gC+B7Jndr7U6McaHK8GPscyM51njy3sVlRdn
lvT/9xJqR8F+mh591uPTIH45c9hWo1pYC1+DuJ19sWbluLr1Tzhr7x4kXOgAS/R6thvP3M4G+626
dFa7tuJuA+yFMo2jvHdF2AXLbpR3dPefxI7Bkwyi7MtsCjHkz+fMcVizdBjm9V3pK1mwbiOzvr/j
by7sPsGsKRNFdUM730QPf2jb+iTsLbo22SHVb6qMGRaPEuTdujMZpumeY55wgKA4EIbiA76+Jik1
YgbaA4PZOtRRDK5NbZv4sRDbWDV6oErOeWTSRS/jS9JRNxz/rICGl5e+6dsfDKhi38iGbSsBTZtU
LqBARzBMdZTf3eaXqSiClGcycDf2YDxE4Z9bwH0jOP1oo6sLNiyqqAml3p5vZu7JC9On5/N+833I
rFLRKq9pRotTOUhcKhWVxyvlNasoWq6EXW7Q3hWv5AVSZhOvrKCOcybe3/fbktIOmD85e9rh0bxy
ABT5ix+bTUqEa/oKwoFrqT9J6YbDX7UepzRb+qSv3ZJJiOpXkKo+du1wuRM3EU4mkXhbuWTIYDyI
6Vg0fhOYNiZBihi8MVpWUo0kyKz+TMTAwuwZ+Z2Mb5OgJfPpWq2H+8NS6qvxESs2wOsELtWq8x2z
tRPJt6yC8EF26ZLjTCW2vU+xOTsf4gUZt1+I4LbuYDtlIeFdm20T7w4kmfzzO1iYY0W2geSkVbZv
4IKEfXS+QGcXUXlWqAQ3ETTwunC0gva0Bs83cCTspa2e3OtdhNezsUjq6F2uS0zMRexWlBgybhXS
C8YrVJa0X25FKcfSu9qtdWadpSjZulu+OEyLh3zAXFJ/EmyL+DGXBaiaHYJnPL57BrdC4TAuK7UR
mLB0dMeFj2246oAc1gbip55RqJWSRNvBlBbdmG2mTMSdfXGPK1pZ4qeRpMM6+FFKunBrh1XBt6zK
XTQQtz927KbtZeU1xu+wjgn+ejfAUuT5ebkFVxGdCK9nDPiyHKdR2lNKG+7wBtfDseLS4BpbWmzX
Qsep8L1E2urYuo9aA+d3FZOprGKmZVs2gFdblrg5JOQXvW17RLoUH9Fq/5SlfIxZ2TppyE30MQN7
uDxun959ZspqCpqKO1+uqB2tx6Bm+gvx+yElre7GfKjBfnZTQkguFqI071v+m9N//bCiTTtll6cV
Gwd1PPm33HRALOS/FnIZwJS9VY4q/+uU4pcmm8UTouN+iQMmGdqg05mRvg0CD6IppJgXqPf2GLQv
Qyc/g8Ql/931QJTd1HpcegArk2N+w83YeZFoQ0o5bTQ7klFZvrG06M48wvgsQnGgdpCchtre6HFQ
rcSShCKtfFG/LPoNTZiL/+ZZFbjL90WTmkWFCJe16bVojeKGVsxBFka8SCcT4TRAqqO58sWDzm9E
YTptnlosEw34YVnaeNIqqYG+NoILhzjQE0flC8rWu+EYk/gjCzwhmlvezMRcDLi/c6B255VdsCLB
hsUSqYo2eXrlnYRIm06UbY0bEaWgSbcyx+a5vK7ZUt4uxapedpOGAeDPij1L/5jrt/o8susTt/3y
ZmsOTvloiRs46l5/vIz5SBc/gVQnZ5ktDUIEsxlt++113tY9XfNF074J06Itt6a51982cXzyAWXY
PVw5rMXsvdnmoO7w6rmjevmAYKKagyf4GuLroJvy4RtsmlHIAJfc0i6RdOlRUrlzQ5wEH7iWe4q2
QTUpzzC/46sczADih0X7U/2y48MhAh/UHpailGlnLr/nsXVAx+2zXvwwTtgASfkf10X9QcsU2M6G
l/4BULs5r0oqJ5QI8R11lR0z6GahWhBEKEV0ZkFQcgFf1FSWPwF9pgYfXvvsYYAhh4Bi61STkEr0
JCufMYa2kNMy2GLf1rRhrT6S6Tpjw5l2kMMNjIaPQM5to95JXvWA3Ub9KBin2AjT39qU35xbyOiP
7ib6Z5MQQ7kc8euVZ6GtlR6gK7b/ietr6d2aZdvloiceaKQze2H1KV0YeCGmxe44DkkVEcHzFOnu
Kn2o87jIjcv/+CW+NcHQqqjuyy+wAop+oXk2Rq0bIYPpLnZKO8s0PiSFOi3ULeGMMMUZRTQLHKZn
+Fa6NbOqbZmMF5g0pgugTBFvJbiPGg4m1+cpEprj78hPBDQgN41wdeuabP8kwzWXjkdRva1b7W8G
YMKvgcktOJd0H5ioy3JRZOzRiLizfQFPVjwGOsHqx0QmBnSLisXYf4vt6Z0E32QGG3+mjAeI3d2y
Yt+p2S1PvyMrbhlFKISv6ZUY47p3hgyGtb82kS/wjV8LP49KWw3n0uR8MLBUKLUTKFDbpzQF2g1J
onH+uykMTK2eAvzB8RCzqA5hj9jrAAElsJ3H2qDPHoAwjqmzfpBPpPma+CU5TlQKONWZB5UJHlja
lD6DY9OMzRCVa1bT3eTeotPWd8k7+awhrkIopqqvpnnsoL6kX4Vkh6pbe7rHPDaOKWmDzx1gMAn6
QK38yI5gJ7mJfQ3RrAbO8TGiH7roZ7oUXhKXca3znVPpSHVqfvkwRqye2zq2TFPCY6NaUXysmzIp
V2NlEH6q5/gFw/Rt7ArKL6erc0Omfs/gu/nWq0j87VBcUYzRsfKMqC9jvJErcOPTWwHzy78K+6/K
qDwYFXd7J2ayYReT9NnM6wK4FRBffrmAdplP8vnKvvHi7Px6/9CyCZZmr7kgcsEtiVWB4ddvxzr5
F1uSza1IV2CVqPP8ieLhPWQmpbcZ5956YXt7Tfq0z13DhVxym2iAfQM4wUx42VoW+qRdgSa/OFut
A49kFdfcsXjVLgYH1G8r/RMlSUQ4Wd6Lr5czhzfnPEulnUE6Zbe24nYTyaHe8zUjbKqGpHTkGOWp
8zKMuxtjI5iL/4kZ2f7toQlCrmobLJlokKinAtX5q/AJnXKt4XCyTCOGUsGGU8D37sjg1svWPOs6
R8qNW8uZ0r45Jxc3oMqmgu/KL6ghjTSc7YypbEbvjdAjWrD1hIrLN5AUJt5H46vepJO19wXydnwX
EgidxRRNnF1qzomPUEmpnDW/UfEUAQn/X5xuL8at/MrVK/ZeBuTOClNxEOe3JHZAtlLVicPqQQcq
Udih5/MlXoOz07TJuoB2v2bA4/wBIBAQOedKvXaq9F4eENqw1xp2ExiF1/US2r8Ui1CeJmj19VBp
MFZADJaKH5q4TXoaDltkEGCkFirpXL+EMsK3nGkr4Kc1wF/OO+58C/8b3/2t/0OnlOuvgRgTKYZm
tmjR27hXpOsaWUfkeTn2YgmbcoSkdHxSX1nW/lDYrmDVzEJEsgiA72qbYawrC4XsH7MhOyxLc8yp
9qjR4xeb3dzwzjM1xsMHi62e57XMCRpjUljw5Lm+LLzwXU9xGlgJ66YxJnTZIj2yI6RHOHuVH95/
VFk+E5jyjXlFCImA54lq2Rgl5iOiKgdRS9/d5RRSIKxIr9A3b+YsfQa/Naarkza1+QZehGJagdfU
QZEtMB/vr8NUtG/CVbsb577SS52vFE3SvIlkgyK4nIP/wFYOI6Wi85aaoVjrCngi8XTzJM0jmA+/
JerLPz8oOADLMNu17gYiR4SoicqC+Y/DaSmz+2rveuxchz9pcvl5sEoC2we5S/Qc3EnOfdmGqzZ9
ZiE8KqpXsyyHpP2OThM2BdVE0lga/uSy/b0ng/NEVXE6SP60ZNZS0iilTU1qv1pPrgZPRFTpPcKc
pukrqKdsPvpn4Ijh/y/v8bv/XF3N0RVcNHrt7Gr66nxtVkkqIMfOBGuKMkPBcktCHxOt7/16ZEJX
z3gdFZS+bK1QZ0hSBiQLEmjgg7dq6HOMnsCQDR4+nEw9kI+1TdWWHYZ74IyLEcNzjoFEIBmcpKz8
tZIO3OMRfHJdioY0V9vMArYvCofe7KrpCz8OMEHJhFqrsKlTtLEGHScDndl+7gWVuExaQdl4Cobb
xmT2hjdk3gjW5mA0mjEdmPyyKZ9Gxm42DMaGijFWVSkaFN+9/dxoYGZ2aSKL5z/Mhi5LZmHZEEvv
OEZvUnMW/Yxrw89y9zfc5XOehV6RusdRqQRfiYITWcjYSWjIbgZoXIribe/7nQn3dePFo7D6hlg+
uqN4V4ThxUL3t66eM2euIxB/GD+lo2JmVoclVuznnZQ+axIsNDqtoBvf0W8ft3pTVdqQ6K0Jw8t2
LHfLo3SwSiXyY/1iRkyOF7aAx7Ps1R+J9COfl6P194UwJjN05vgdUvkX5YeMZ0qW2hhZJ22qiT5E
RGk6hkAILFqcwEaCdvacLS6VAZfaOeBvl5kgv/droxQZgHVJ1sOhgef5bQ7AeMGajEgrcepEwJdH
BqpBmJPDqCKcuhchcxrnwMnQpbl5bUfvfDU5XF2qRT8aQCiiqO+YlnSiCpXu4+mQBipIGkiDPFHt
eUxbo8YAt8/Fr/gpugiwEFgTqlNb11mYkmocOXRxpWuYaVYAP/6ofs0nSPCjukkSIXdZK68ZDBpQ
vD5YF124wXkZBaCyOFxzkuSAyM79VRPFIIK8hwIAcyiV4r4fi0ND2y5fbiZg8Hwe1hTN2jXL+Frt
3indt5jUIxOFyUanWVtt7rleFWuUbCV6c+RXqlxtp1rfkDzTO4NIW3oCgQnCDZ6eoxU+Rz0o14uz
vfQg3eDgEmPu39t6mwJhTwd4p96z9dJobYZXT/yTFnHYf/BR6mr4NdOfrFtomFSCzCQl5NdP9zK6
XqgKaMFylUBNIhRvcHVicI2M0PpNeMDpouYMCgG+CytWJ73+XfjbRpnLFQG0GE2VAxR85iF2Em/1
8SkaDQdxxdsCWAOBIvfBGdF8klRSZ7SXVwLR006iFEoHARzELbdYjjBqDBBOMlq4czML4uydrxws
a/S7EZLblrubNf+TAtTPHeU4I3F7tJZbM9Ktfc3MA/FMTtiGlpvCheoyTwPC/UOBoF3Rmk+R2nJo
6CtQWNSI/LnlW2admGtgkjiU/PvVlz2CZVrD4Ob8VvycREzDcIBfDPWmk7AT/Mc0H/hsUSW7AX0o
VduB27uDjmO+Dcaqx+9GLa1N5OQYUub6BMe7uajVxOkF12jqwPR6dY48J1xTBPhq6PvOx6/XlwlW
usbUWY94SZLsJgJj7PkAc5sbmHlzVFjAgcivDP8pDwZTQ9Elr4V4jVYdRXwPDNNXon7OYcyc/+mc
eLXYh6deYXmo9akJ/w4bqMlnnnLXuFZTsHC6zcTOInDloZonNygrJe3Cpqi9CCRIX78OpbB0pMxu
YbpMyN2YwkvgCfPNmc18qvy3ncpjY/lEgK6fVJKR4iciJO4hEjEBj6rIKnPWG4Sn1m85g55kaPiG
S7Lt6qerzSwFq4FJth7HfiorFTnzO4/RF+E+2wgTXZZTDiIlbGKPN2gY5V5EDwDcFX06DEbM2NqP
KirmppAwUp8X76wrrcW6KuRdgsRQjv7cyPnggiGkZMzvJwmkfZ59CSwOwRbpdFlDScrDqm/nkrRl
xpVY0dhk0pR81sSCMfDLvTA+6CYIu4LHuwyEphakF8qL+Iy8TY9C2VMoUysd9oWsYzw0+VJMAHCA
4D5q4q7sgRcdMpvRGGT1X6k71gyuavh3DxEDj56N4rKullLzTwX9srqeTwCuwRU7du7KTXdqY4GE
cbQ337j/SQmvvV5OzLF0J/IqwaKFC+6s4+HPTBPXo6mJPHyIAzW0N1t2XQAXAueueti/T2O0gCeY
k31Jla5TtXf7AAFO3SW0hv5I19uPEDbNJwn/cd33/Dtn16hC7HekM+tYI2xGhxWCMuMJorxhQFG2
xs3D05WabNqd9XmuganJt1gLdrhDZkQbWa+3N1tfqv8cxNCKaYLA39ySORXvBk/XZCdOocNSI5LG
t42Kah7YFxQzTE+wzID0E6CkNUcSWbCWxog/aeNeE3WX8iQEcG7teb9R07vfrM1wYSj2Kf3hucpJ
7A+xk0q0CsiWrxTghYSdyvMsJJc0IpeojtRDdzlEQ0UzP8qO3cZsI3eUmNxfcEUwfte8T7b+KaSd
7fFnZw7uxHZ/NI93BBEM9GJ7wHZkBSF4dMjAMFScjWYaBJLXMYNHH9oChoU3NgX1IqFn3bRTlnWV
IWLOZ430MApWKnLWfVQbTQ9gXYTmCrVAaQjp6vWBujme2J2AJn9CS3Yo8cyBKW9HkwRex1GA4IaX
3UKVl1wkqKVB85AfQi3XqWOPYai3fSFP6n2dTuWGY4zhQLRWID/YQ5Vygb/HYT/KXE8Ucahswyy1
yfBsiIk4xClybgU80Wdd2cQnj0u8d2WHjypGCQ09hObPWGuXINmP8iRMU8A1pKKCDBxsE5GKsKF3
TG0o3lJZ4PKIfzXdthW4J0I25/CCXby6qIbGyEbO60wyVIjW3zAzfEb+ScKhWMbw7hmICScNZPjc
wJ/GYjIiBwiIc1hpzY4u1kOPefx7eWkXzESFv/pmA/nqoTlSWC/qzieFKlvK2tkf6nlWk+dag0Z1
boQPzDoX5kEsRQul2WvUiIjLssm3XkzbFn/WW6sSRqDnLs2nolxWpIBFQMwuqzHLVz+ngkiR7Rf3
YUq6uZQJmBCT5GUkp2Y9/8m5uctdiLRmfuzvB+9S59va8FazyrOiTqZc4vy4Ch2OACfsHZ9UPX9M
6rsvxMbFcg4eUyxMh0M+jPgdj0+G9aqP3KpvZUCOUuC3JLDbE2xEK1FMXWK4WqS9Zwhy+h/8uuqV
s0gLeqmXqNdzBXb4sLb4wHDBjwRPKkbRCZGcoHyPVdowLr6xvAanY5+ubsKAsjKtpkThP9AEbIkF
jomla0ht+I+7mY2Y9BHina/6wU64OzoVoFqlU8vTSkrM5JVJgelqecSExY9iWavkE1anlZiMNSlf
cq049T7Q03XPR0gwV1+cJ/eWic8RIRfsbtLVsJvRoaosxcMFtdyIabI7/17wUvNC2IfVPr+2aRWP
5jto2tzP2RxxEBFYWGTueEcxxuC5hhSsm8v2ApX4iS6nnmrJWO138oNx5EURmFgptplJZp4jEhi9
s/iAYi7RIcHekXh939EqsQXvYydnOwZr5QzsMry3VqYDysJs6foccxKxPSN21pVqdKnsq5Gra2Du
vgWNDPLKR0aOZOCxdwTvZEAd9gzXSxjOZ5M/IUL52LPSRpZcMDGFJoEN7/YIw8N/3Mm8+R60Y/rN
O/1ThWmrXVeNguzpAIIkNZ+AOZHPoDxFf5GFu2X1PrqBJxbPvC0qVtN7PoFCFHtzZLhBprxiiSX1
3uzwkTmdNi+RZdWNAJoa+Kx7sboZqrf2OvPH279o9rn2Mlk+j+O2uheI9UA8GEJaT6KgZZ6h4xc2
Dnq3LNbv1Y+yb64QpV0NCpd1oQo8cxHMRE8N/n/ii5Or+ZJyMSOGXEAOz6PhuX8jAUyyg2g28+L1
zhDDuow7gquUGJfqWE9t3irR8F9QvpcUxGTmdZb5Umu2mIUC9FunBZ6egrZW1QVW8pT06MDodJHQ
+HuCwCnFA9tMW+MxUPh2H+z4ATIWzlPmZvgKQd38f+uMUNjRrTJzVx/7YHSPjtKajzIlvIhZU3jE
Ya9X7kfN15RwMYkoPu+e5cE4kro20RTKqleGJ3KVoeENZpyjyPgBrxQ2aVhv7Jngk0XAjNXwxjw2
ZqLVdxyMEMYhjaeyio+BjqWiYSOPS9lM0B882aKnFFTBZ3+B8TYQ21YyKUCRFN/QbMS0R+rC/l6g
rvyosUj0wI8Gd4KC8Dxw5GvMSKrnt2eRjotKsY8AbFmvS1MN6BdSPANfIfPfx0RKCf4pRSfuFuQS
M9t++fscjeUZZOZtf5kqZkV6bNWwWusR7EdMdL8F6d0e0B08S0OzCqoLQ/7ZniVriwbT/bJMkab9
iUAUNCmBQ+3MnKNKCbzA87RmrpI4B3C2hBuBvDqgvNlZtWw8WgRQ6kMxfUanLgFMi+f4wlDf2zWv
RblHzbMsUht2SUkk6XhxPzTOxkalbtyT4Eyrss+nL0CT8Eu3SAyzUgibHqX3xe0s7dqcF7BiBi7S
AjWMg3RfM4P6vlhZFHawM6kmPfEMDRKxINH0DHBFSKiOE1du5X5Wdoj5NM3q4/uTNJypAazvEJxC
p/svL5whwwouFgkzj7wDgb1PG/iI2e7mK/zK5v6fymoJEaSVK4jLv69bm9X6SGFw/b1Y0rs/QG71
sCYFy3fEBr28fTVqKsexy9Jvti2pwGQrk81QBuBTaI5HlydJUi6LghrP6d0rzmTovLms5TxMbJod
eFtG+emjAxPwSNFSDutlPFT0OLbMrdHOYICPakC1CWKB2aLrdQ9OORV2aOUfDNlUQMFeLy0bVhYR
NPPCoBnsHlA4fgRK8ehFjww4UFYt/GW8XtvJagAYzw2lACMVe1VOhv3+VmNKWb+/9Gf66djgLI4I
2Q67EI8jCWqsp7UNLnOcOGa+aUGADlCo65e9EEpiqtU0kwE04ApiO5f/TxtofnimK6p43OyQZ8Yq
/WdL0odYpJ5R509BFCmEnHnFB4uHZc3ME+vQO/xPQog28+2i6aAPjN4bR5yDaJsXAUgQ3J+1Vp2L
91lr0neQT2MIz7k+e0TsU1g2cClKNy8sk0J4Mx0r0PmMvY5ZJ+8DFnF4dRhjbXNbALjTRi5RAduR
+GQlCmKq3NInNQwZhmQPotNOubLZnkRUiJj+l8y1GzNFaY8RQ9JxLWH9WyehUicxNHJRpRlmX9kA
U73r3WZrTMHrHcP9tkHF32qZ11qKokj53EIXa8zCT+oNSpViA8cQXLd3XwTPbA+AQBQVuaeZwvMC
f4sow7bUHAYQWsmV875ZqqMzIZ/yz99ZY90xWaSSrX/MZdVIk6JYgLyrPmtxxS1vKSIZTCVxPvvz
0g/my55ucWzsJntmp0hyW2FbpBjoztd6qiiYnvFjLn5aWLg8sXS7xEJLAwzj+XieLT1K/OmOOty4
u9Rl4ko2kGtgPKM6MGBL6VvzmmZtlAiVKSglVBEBvMhT8Pqb5FH0Narq/+0QiaQzgfvGfZzKRola
DkmqzP/d2Ug27bvxABMPUjVpJGas1qKPjmiNJQpgWArxodsbe7p9ntpS7IrKl+qTtT0SWiQHs9HP
utbL4wTH/blEyval9rIxQiNq9U1sUAZftKue83lXZYkYhJtm9cMztvnfTpou39OSyocYYrIO38Lc
GEjztCJQBpwldVQRpYQqlTxls6OTeicCCDqBvqXVulLvMDpXKim+WEh/oEmzfaU16dyXgSHPbU5E
bIbjf62ZdIgPbr+WLroaDAOufwpRzJaGLbteY4s1on8xA5pz9fMwerNcpLdeGIWQyFvI/Xr+k5gT
E/Ta1h8Pxda8P5ADh44o1cacn7LQFPEqiN/UC63AuYTbr+4nu2r6k7B8iWALm+tqcGoWF9UEuOsH
11keMAOcsRj/Zj2mDS3L+iLiSCp4tJaTrA2eSYay7sw4DQbqGv3AodgvVErMSrzhgcQd+1ParCdy
nPtmn9xszGNKXhsYFM6BKoVEs6sCB/M2LLopxdDl5a1Fojgci8NQgacq4gSj5gtn1eiulm81CUqa
pxU5zrA54qjSi6Hw8YzNia0Jh7M6xibgiT/rIuC6SQmxgaP4LV8OT0KdZGeixiZ8aUpr3JDH94IN
wf9aaIbA+dAW59U8jaWbklPWZwlJLQ3JmzN5zkLtTBGCj9I85I9lztBdXP3CbDaQ6/OFsPlByrtk
5WhvTydoILiM5PKcXZA5b+fy5kUwYqGYKT6oCa2ARzLixKMj6yOYhI9TDtiw871zr74+oW+avKPa
Bzms9xZVEZSoComZWH6O37OCH7HjbxLCUcSvbpvHTTuAkT8ffVHsOPn3REMltjGAyrvtYIvnTMfV
o0Ry2dJRMqr3U1Ck44U2FnxZ5B4o1LVOU064jlmvxOPZMYp3LA7a4jx8HlYSaC79NKs9B9AA4ta1
Cw5MSzn9l0HZ7I7Jeocx2c7Aw09OaUPzV7Ml+MaPsNb/SgwkvRBP0hJxK6EkW4IvMJ0gYuxm+rOE
5FqH+vcbPe7HjXT0+O9gTdOjp0Ljm7yoOQnylAxjDNl+f8PIJ5/UsWJcj6n5NiNcrNI3bx5Tjdu9
epswQuHREQqGHxfFaI/2b1aNqDCQGPcePD1KrnQj9dp8xMjSqbmT0K6T2m+BddQpUBzbp6fpWdz3
ru250e9hSLdq/vAoQXvYsxNnaQ+s7K+mszG9cuU2q3nqjE4eNLBnx6Wx1CyrDXb8ImjxGz6iBCcz
61lpBbzvnKSA3x8TxjI8zzmrB1/ipzd4aikwv/PK0DcFhLC8peT6UGatMeY754MCzS6Zh8mguyUO
hfYx4tPbi53BrBWfx0Kw2ghkh49zrrGCXF9hvCqtYJtuQ9xMYm8F5ydgzvfwUwywLOpk9Mwh+1cj
LIzQbnnUzs6/z6rRfS5F8d9bOQMl0Bx6ctnTn+yyGDyD+zRsizNZrkGLAr9Zrz0y6JFfsRah4KN7
/jjTdralEarYgSjBVpdri04CoCO38XXuVQ7FL6guJGCCQVVoyobyoyLLmH1OEpau+IKk4l3AJrPj
wE78kPAAlToT+dTltbnTIRquh7pFP4hfPwgpZnfRZlWM5WnAmxwL0k9yX+oRkbJCPiac3AdQnVHB
tNVh8U7H+n6w31/i7CtNoFo/FCglJuXTXDCRwuy8cEnLFxEiep081VgiUBWrJK/udcxG1Ty0Pbe6
PjjbLU9OMTW18JSomWNmjbmJej4UlUPjM3+NtjIN9RihokZJcWZPPW9gUtFZvQDVNst7I6BKtG5v
Ta4uP7dUhGd3hS7XECjj374CxLzYvs49vAzrbD3UAZFimO59XPDnr8hxwMSeO8SUTiyNjG8XCquT
vS7zzFknXh9Pa2qcZofZaoqzsrTUGWcKcD4bNG539ZlHUpCJ/Yf1iE+HmvC9C1g2I8rJzN/YdVJr
1HXi95gfG5mpCQateJTYweXyI7jpBgRJgwB831uLs4U47ZfN/a2dVXjxTCvOiyZH7MxngLQ8l9L5
EVKXC74QbeAZXd/KNn0ZryXCLBb09pjkJQAmeYMTMqw0oHThfRmzHsDi9pnQGuU6rHPVVbwjVKx4
z/YbDncYdnu2PU7SueWFeioqJ+y3WKvAJz5xoR+U7xUS4cu1K+a6zN/mKMWUiWwPmkIjWO6D+MnF
7sT7D3qYcONkwDYxCsnnYSKgd3KXIwffMqg0EaYCSr10pfZkPkpRiVlhI1+xCXpBNmGK3ni/uMOk
S31TFtnRPEG0HHIJ6CDbjk0hARj81G6EXyZUM18Y3iztF83GDQ2ghYNlp+TedOhM1ZV4yBAgjUbU
Qp9YPywat7PLbYKhA9VymgUIe8jb3RkuvJAY6PZ+xOOrn6UzDEAsftwsHJu7+j8kMZJnK/1wzg3i
Cd3olGHM+C9hMZcmR7FxsnOowhd/JFfkgm7gXpqfQzjq4q85LhrJWFft/NrTdA1ZWit75sx/twqO
gdqML8LV7jPgHxgynku7POrtC0OYyxpfd4bXQtswDiRW2Bk/fNxDAx399aGLWOohy3In8oU+bm7E
RKklA5XoScuWwZJYiqEIvjPK6gRKiuiAPgq3q76lOhcFY0h3W0TDMZrPZopYcKkUehx5xWlJtEYH
Ce+2skTihRPlHQXYAR6jI9Sp1A1pO/ufRxc2hFC+9053iDMTknyL90AqmJOpeKTtRuQS1tBVBZq/
pP7AZ0F8u/NRLpf6z/GLKR9MctiXqVLyL8c9cK5G+oCUV38eu/LAxk4XajZ7bMexX2BVoQSg+Kle
Mk6yUNdKt9J3mVjho8eLn1Vb/hd7KustWPTPNDYzDhIMOkt4fcMu4u3VsLRwD6EyOZBBgBgkSW6R
uN/dDqffNamyFyIPXKi8Q7YLN11NlOqrdnP/xA5bIhQvJwuZgFapzWRi0WWpVe+FUouolH5NMUuG
nFIlJp2r+GlxJUeb3fgJUGY+JQ69kp553geDkly1FI4JgFuVAERG+yWH1LwXWGM46mJnTkC2NBJE
SnHHS2PdkZXBc2gOt5RHdjI4HHRhuhSy8AVVs8bvVwZTFV7Me5d6xLnjEIY4oJwhczWVTtxSMUCL
L8oly3sIkcdwV1l5tR1CmT4QwW2Bu/ThO/+9ivpIM6JCIrTdW6dswUv1jnKERiTb5uXbGtxJFRRn
anzgu7ZVhHldulwpiPkm2kAR0/WWSERoRh5G3XRyqwCCfV9GUrRSU0qOkF4mKzL2kHYjibYQwIN7
WOXI964K5bBp0bZUQpl0amNkwqphmRlypa8eMJAVRiSm/D9OWFTuJpotaiReNyuL8A9Z3gPLvbvs
r2QZ943MHXVwL02JkRT8RTEw/89i/jpudy2A/t3bIdl/+N+p//wG/KWBvUUaPyq4Q3ZGDnHND2EB
w36ye+zc/YScIFbBix5HIlVMIJn2bmpE7J9EU01l4pZy6DdFdq2FTbmr89egcNYCq5UoR8AdYa+U
q7YMzDWs1JhOnoWE4Yd+UHwdEZBD/9agbnfPAB6TCFZjQ92TGwJciPx/FTEzKidUoJpbAgBvGhYg
eIqQhNfu3P1r8URJqF637QctEucvX7smWN8JzP7/9MKSHQawO/5QDkztvjwt0SQcs1yCEZ+NaBWj
SB5CN3320otwZZh/q5EcMq1FeKsM2bLEeNwmp7rHQ/IgE2qEHA7dBUwdV6chpTA8zFrjF+Oes8sc
kjsBqokj8D+j3LOzZHwDqiDNU0YFFvlToLR3EQ2buYDNQEkRF4lG42gzy65aHWsUsU3gTHiE2hbj
E+dnkQJgaph+6wy2ruAnkAP9wbtdxQx7cUuE2xeuj8CWv2JHZg2GNk7ak9T/r3pIukJ6TSkXepjV
eZmIdFEcuE8mNbGlG5jbPydmWb7KlrvOSJXArpTTU3B5ZyaOF6RRJ5gflXvIyCeE85mRQGbkCtrZ
6/tDD4bGTKDzKN58Y29XhYqNlpUvbnE1XSeqc8vCwAOV1vS29dSijWjFaQbk94bALcWoRQpwmPSV
tLyiUGWgP+BIyK+YRRnbIlCs5iy3ndMO4BjRQ56/6xAEl1Ec0+JPAiND3xv//sf4R1yx4Pef75iK
L4MAifR138IsWwFmLSlqGpsBobQFka6lpM7Gk/gmy4r3ztGLNzVZbVS0qP17vI00r85iKOJKJlYR
d4LqROL/pKEE+QVNQtfLLnljqUZOLgGv+bbcOvfval3jfZabSCjM8/z4blaWxjg64SjDA+6N6u/G
FWAb/lThkzEvZlnSSoKCGd40EweNJvrukSeQeobRQL5fxpZmhho2rG+fTZRQddTAw2AV48PoQm4g
OGZLU/EDGIY12g024v9dOFpUHTeBm0m7RdLzNcd8NnuGpe+K2LLm0WOIUN5R4MWf1vwfYArwy/4e
2aNs06pYZJ8cbXTnFWEURSEU4yXj8n5syySRsEthb4KFy8UNZ7qp9As9Qj1uH3RwuA30Pdd33gjn
CWe0UKW39vmFX2iBqJDrZYQPINrRHySSOXIGR2eflR4Vu6vaRnaF7NHa5VFlC3m4aanJViQGSBd+
8gLu4djnSC3r/Z0y76j8GacemxyAsGYe8rDhJix9FmUSBQ7GFw/CmewIBRJ4N0Cmsrqi/S9xNx7d
YLm4RH70scHvByH+aOk9FdIvkOpaoykTLx5tbleASawC/2/sm8PqwXF0znB4Hi+d3C2Gf8Xz13Z2
uJJ70iAuKmT0Mt0LfXyOpDIHzRm7P+qI7L1noY3zVSr7QBawEUAJRa+FNlhE/7f4H14blKed9Rx4
JuE4szgOkCK7ENMFU9t0k0hgtB5zjuAWJ9eVS2Qwnau3lnoN6HnvJ6VjRg/8IpfkM/XOgjjHhmGw
w117QhdylBUImnfIobIG1qeAUVnaYVO2/wmTpSZt9VvfID7LsfUXGG5/aJoLkCyrbmbL6uY936Yh
+PIZuXNM4PcOp3ezkcQJMvvNxmbXl2K68+6tFSyJsG1y5mJkwTzCx7fZbiwLcubTeOnrI/UPtnDg
uxPDdhC375os7deF7qM95HVthYgk/M1Wt0XPi+n0ui7/+fzc9faNzHzSfFpEwdO6EbYNGk5Tx27c
+AiI92ggCtHBWqcPexH3hPthkyzXtH38nWC0hnIaAskVS15ervQ28TkwH+Qms7AKbFTfcpmGSxqV
AFoTRfXTgnVX2EGRAS48q5smjXgL/hWjdD2L0MhQ2LbqvmRxNATp5ZoLswe02WgA3V+BxTP/fZvs
i/euxOQz/CR715MBfFZFIK5wEPpXB1y6vYEho6RvB7RQWDm08OzBBBRDDqTzayhdVVOcUejypOVO
h5UdLN0mB7803JYPuzF/zk2xQpzVfee4AXYpAi/af0Ibmt1we4ZG765+mlqcx2ZOomoP3rz/u8ys
qCWzh38/3C/+Bq079wRIn2+ykIy1hnzfwoovlPzS1u8SdajJ8LYGBB2WlBwd9atlQBYfzT7UOBdo
bT7WJm0uTdvbwBqeQJDvPwratC2qQJYEzAivNf9ZSjUiT+VZcwJQC33MHypaTYdaQx+dyH/NRvnu
YO1/fjHwKSfM8Zde7YuzKO3pXyNpWvdC5XcY/5GeWbtAKDlmkBN7YIfEm7nHW/UvmNKDNMNik2YN
UvflrE88Q+e0VVXtFysKv0XmVO284kCiFsOgxx80OajU9YgpG0TmVn5rsK75bnh96Ioer71yxMud
tkPVTad7flCfkEqa0VQzi17UEiL50Q0le9IrOZgKpb1RGeaRHCJK10pUzWrrEffGXVexrwydm8KL
HuTMt681wHHGxUar8KsL5WpXrmG9271QqCSzlyGYkJxGWFbv7ZXjTKaevkwQmRD9M71z0GjqI+pk
r906aABT6662TLU7dBiXYNMWX676Foi2fsBBnEFqOnkGtZJglYAP33jNPjon8B+/wfupYT0wyi+A
Ut+Wral4wNG6dbBO059/tWJPTm5aUO666Zu8OocCoPUoBeV4UEYgO25XZpX9VodG21mklJqW74Yl
FVl1Qm+hlvK6b6gcu9skFOftmEWkJDbcYyTwDHYuVPpQ8UToIQkywRH9f0m79tttepr9CLb8deBX
n5M89AiKrefKCjkJcddlyAplgr39rG3cMmR2l7H4mgVF2EpEBmTEyvzZIm/qVKVTdfElCx/kbq48
0uM20tOx88nrCyvRLdfGFGfqlZx4OQIIQcL9Za7H6XSiQT08k+/qVDIBSz+FTQMBEWLqDAzeuCCD
6Fby+O5kSdwQ2Rd9WguWf1RreDUr8ci/lzJmpEax4SuihRisRTsZiXFnIrwjRn7ugKbG5wdhbvQT
zPh9CmSy2fYh4f3RkiN3ujjeOJ4da2tA8VKhfT0i7kU07GrQuR1S/Wns8OiS+NY7lIzN/oNyTnz3
2g07PBsCZxasp6xCJKb6NdIwNtBh0I0bfYOro1wslp/ccEvh8Tvaqf73SP1HI4NmwtT0m8cAvx7C
5jWny7PVa1Brkgx2ZyKmeQhp5VNtCnaxSA/8EtY1G37tAYHb9f/HQvNxQ+HF0sWzMhHeciINsFGK
M7AhxQABZ/8UVkowrRh1jmGgnneTQvQTt/3y3zWOu0r94i5vpxRRAI4QNPcTDMEsWhp21QLN1jnB
ek/J3ASwNZEMV+hc9DO3P8EKcDwGY3Cu0l1+ZWQcM6BSgu6orUrrXnP+uGv7wLYeS6qd6jUI1jWZ
g5CGGRmcrEDfXUzjRRNtLOYq2l8IscEXQFPB//cQPrY6vUvcWFW0SG9cR1Hv62HkI/VJ/26Pr6oh
3cuND4IISq12Frnj7yMf+wHHziMAyWXUHDTM6ion3+0jLn/tnczOD5wP11gWm1a0GkYXwzycq6DA
5kGIyyP+IISfBsTpWWoSWalvPNv7mmFBLLdi+T4/MMLK7XGwvLSIOCGK9rpptVOqSCMCylM9Diq2
/632sGh9fXpgCncM4WJ/o5IkG2+lYf9yCnn3TnZhAK9/TJ1lP5auHdgWROgiXE8yaLCMHfsi65Ao
4FqJNSW6RIEAiqJGoZTV3Qvzi1lzHP121GBwsAbecz5xKOVBRXSdW2+5+2UjBGRql5dYZaNs0IDF
SljMLGz1xylPHHo4E8NYEvXiXigjAiNI6RjhiC6Oyaaimhn8KUr3ZVmTgUFm0G5bXDt05WlfXMmh
iS0X2zDTO1kRE0QStuZIdTtLvbI8jeo4xdKDcL1ql8/F4IgNPmciASw5sH1+Pi09tjKFD9SVb3zt
hDhEpyZlzsWcBs4GRN5kVpjsofxuraUWb5kcbzX7V2Emr14OPjOzmVkp4XdaxqHROW/cavp4bn5/
B0mEJRlUu9DFsd6MLPgy7SmzPJOGx2MMf5kY0vaD/j8WNDQrDVeudlOSBXAT3XBQgQnmX2p7QLnU
B2pJGTYImtM8eOkfxavLrYNx8uaIN0q9FuYlTDzoKcQZYAVh4Osap/9F+x2Oi8zvlGaPr+rBI3it
bUVGmiqG7OVvdX9MxBIB8PR1NfKKu3l19Qbryk9eo18wyo62iWlk3DK96ANU1dBp37Gp0csszaq4
nrB3vj3OZIeMxVrv/1gRlkGaDJQxLEH+NPCpwJKY2UrGosz1nBESeW0i4paRpyjTils+huFEEOil
bAihDLy2F/JvBWSJWH8IbI03cINsaNjnkAfWyHK5sNHBypDq0RZ8stSoLoTA1FIluW/wDOTBkrZ4
qYIs9OqfrCWXkY8eIb/tsrn53WFvDMG4ZgY6wFtbsqPnM900VckKE0VM7SZOm/65QF2o0i4d2rUp
JpezsOGJbngV22tgUfMrIAVFHxUtZooeLVIXZU2M8rB+oNfn6LSGddDriHXGhdPGIzBlzucIHYC2
dTq5kRHGzpRGVGA2+60TQyCCABxHBZ5knaT40PORg7WlYR66uG18rg8vFAbWvYDy79I/FhvjFaHv
dAFUsuEpDKv3y4IV2sBA+FGofAYnfqO1IUMTr8MSqm7CqdoLHebuoahubG8URmtySli/Ws3E9OTf
0Zhfwx+UcSP14TZEdNhQq/vrrNDREdTW1pw5+bUMxh9o/W1CqyoxF1A86x1W1xS5canP2/UGZzxa
qiOiaKwcov3gVwH9TSuyXQSGpJFkQTH0bdC53Laci+1To0n9rYPcPSXVG9w/ldhgrgJhZ42mBEcC
+9ItcVALMfM3kKXRLOaleBjqhFv7xVKbWBYrHkgLjV3yusCCtDsEcSDs1NfCGq/3mp8MIMTeJcp0
LPAhzUgtMTLdTtw7HF2RQc8qsiZBQMbrg2ujNqyD4OHhZn2VpPMyHUXeMcfShggNK9IiIIC+DMlu
feGleoDCiOCsm8GbO6XGIBRBtLFpdLYEl05pIzI/kdMrbhouAmrkfXh6YNpofoVNH+feJ6BLxFiK
iKuOxW7+q3GkbDSN3HzEg68Iwuhfnqg49dgq6Qb3hiI5L1u0bPMf2idfan1gVNpPpzzOX7eVAzk/
h1ONqXSstrap+7wAvG5Kf5x3Z1NULYuQLw4+lnmHceVNGHxvhpbfhFF0CNj7CubNvB2VsnLz0z9D
CTNxmAvrJZ6jXmC4WmvQXfU+Vzpg39WQGuxK+Cr7YxlJHXd/lDWWxTF8Kwylhq9su/QdUPV2Ntpc
L17kIL0GX1XSeQueZCDlnXhsW78ThhC2PhZupXtraK59CgjE2LrglCJcfqp65+JaQnxkiKW7jNI+
ha2AaB3rSWjXeq50NYH9ToJILurcxg/lw9X/5EjxfG6Py4Aqxkn85TYgP18wg+Fuvlc5yIN6j5gg
yvTc1an7mSK2nWczn9p79fLVsvcjxef4kFRVBAI5NzNi5aEH90q5AwGVr2cBsD3+X+wrTy46DU3K
TQxaAabInWG4TALiJqQ+Qzttq++9CBEDSCU9t1xaApd3AlrsKVicS4QQfrLs21K96JAvQNR8hppN
rjhyubxgo0g9cfTX8X3dyETJL/bPyJQJn5n1jjwSYWm8+VvLJSR5CvrVNCXmUf/GqU6B3kxvZrkF
RUP4nhAcxboxGgsIg7l80gGsqF2U1Z+gnhPkFD7z+tbU9nHfFiFMQ5ywl4u6W/ELiz/hGvTqPoLS
bzYtsnkQgYUhlzzTjN5HKpmrR1De+d43WR1CzGy3GhiH4CLencnje8HZCDDa6KYqeYMRKEPDntLE
aTdk4Q5isxw87GLePuRZM1Yst0X6zgIh6MAznRJZiaf0ovGNpSvmMI88v2fD993140LtWhyHF0G6
lNB+PiOhEcLbJbw8z09aBmIevRD1XPVfqYetxcuFlo/LNk4GmQG2IleMBG7b0AYqnQZNKupn3reT
o9Ayjy2vL4Ax62wTBUdDo2TK0ABrnsjRS36BS7ScrTClx0DuXVSoshY1ANH8qbZgd7I1cvPzenA/
vi1G98eKVAEHnkyra9ER69NhahGm/xnh0/WpT8D+iCiYbHggF2T4vb6xojiJA4Ce2jXxrTr8u4o7
7/EONJ3CbXEgtqf8WYNJlBd3+PSECjsyt+P5ZIXQSeLXXD3cepdANUTiTmI+nhM+B81q6Fl9rCl4
dfRM+NCjuXIM4unaYPcRaXFQvdN5ac66uVtsY7K+YFxBeefMvdVRcR3W2VbuaWKfomnV59wgc+e5
k0ZLflUuLM2dftwR31Jxo86rcBz00dQikMfA9q/kJWa9QHJfCh0PhyHV/HXBCoLBSCgRlF2/kQne
XKrGrFaqeWAwelGXuPAHVRAkHYla0REsB+FvFVQhtEXS4cykxjcPBvoKpZ68iHEZGKxcypgNyfVx
nBji839/tOmcUsjCH15ZOC32Vy9yR070tWd6Se4EAgODRqeBsnIlir2hxGEmBL2fUw4uaieddQLP
OcZD/ctg38wBKgFCJCmVNn6ua9X4Q1DdFYGcbgNWm+sAKbONqMCnz3cM3wrxYDlhU48efB/pDS2L
lLnJ+IsV/CADgt/3MdA6KcO63U4B1QTD8wBOGJOL1IWI8XrXRsUBCoOwF/ImwaPW5scXSAdCY341
S2ifJVPn7Euej0hWLI8chc92MnP2V9VE23bH/5GC3jrv0xejMJ9jJNaWy7JK1yRa/pQ24emGLsbN
vZQNPKBcY3YUS8/HMlRuLv3b/e9ttIfidYlF9HVQh16jkdYSc9m9WanNb0tv/c/5+cDnAOKIbR6h
QytUKzBUGxB8zlEkCRaMpywfpuRHKZvtvVCAdTjyMnjgjjVeTLuL0l++sc1bgh7tJ3e5kfPi6t1L
YI5Msy0N7KVvUWAtDU/BJtahCVTNF8MsTOTJUZXPqR+LXxF1LpzwgCyLgR9luUa0WtVa0gD4Z8LU
6J4P5tkLOR46I0e+dPULpydgCobt1zy2/ra1Hh5XaUngQyz4Hezp+H2FgLrrM2Ksv6+1U2ZIE8M9
s4xNlKocAbnvIVdgMsicIonAphc7Jre5x8UySbY6xb3RYrii4oFMS2JXbUstjkqhAsTJcKf89ZJM
9adVdejFielNL5BXrW4pik9PPaUJah+9/pnrDqGTA6TGTX9WKBbnBhwHRM/ecfvKxh+p/9xqWZfQ
eii/TJSBI3qKdrnaigtZChEsrgIBCcRbiHhRjFFKtrMF6RxD6ZYUG2OEFznxx0WrA1ouJL237tBe
yh4AY43gUMsefLunvPsSgFzoycheOSh+tbbJxnpGQo0R6atzgfWxMuyweBBARd6tWQtg9S+T9JYd
7kO+0+//irTKqYSEeMRqcjGd00s0Cq1uYBUT8KC0SLv1105542+X/UxPbcOWEtDtqEkIyM18Umxk
WGuGpPqzejHSOgiZtGamrkwmrXf07CNUhtEvMhtkEH1ymyhzXYEJwt/3QVxLnQ5XcMSYFi/vItWo
/rORRyON3EJmdv5p95Mklixl/P8af2idON0dw9R7xUS5+YC9/FA3eh8E5fEI6hHSLPcrOJN671hS
2uZqXBTmKRwwr/BUO5bHgWAkfkn8G5AD0k3ZxWxs+fTA6x74eQV7fpiGuYFfUZ8EAARazlOFQqSI
rZr7wp3oihORSGtJ3AtEsLehcu+A64uF94+s2cfwVglNSpO7Ig//70odPymrfBG63X2UEPiNT7IF
91Ew2v414BrJzf75VuzchulOk+rMj3dtsC2Gxo1A4LQqAVLjV34ksc6cCRjWJrBoHFC2pBlhCe4m
tZVmFLsNQnATKZgInNMjTqdkFzweI8avlaGC+FSwJQMp8iiCgxgEm0ETXqGmJg9P4o6ZQBVBxwPV
GdYHDZldNyVI2iL2kHm9M8tBXQmHM4bmM07oRVU32KJdJ71GKbLLlIM65SZr7ls3ddy0BkRzxNMY
unZ2uSTGmihkJzZMdhdchzogaVvv/9gPh2gah2NMI7OuIlgX7OvZ3nULUMdeSUdPYhYwfPR5L2e9
CQsHLbm8p6VG8GzUB+NVLNMJjMUgOy6Uyj0gTY5G41gmsP+nzHTn5UWR/K5SSQRbb8CGuvqxUkZK
5OGrHOuH6hTDkEWKtXLdTjD3+ssHuQqeOUbwxKmgBll0EtTLU+py9qkSseqM6n/dSdCYwuhXTYgB
MoCuVdfkQo9EXADOzJzh7hlbwOyhScOhLufGSL9ytTlSxzjTEFaANrUpQQdg6P8+Va2NbeulvG5q
lUG8MNjHf+Nci/Yn4nf6g1BsdU/Nb//uzgPujgBPfYrwcXL/NREZ2Y+X4EcDeqGrh/g6mDdEX2pt
TkcP6xgh8viEkdy+In+Ar78H+xfF7oE70feSM2+9hdU6NZCCjCrNnsyjm+KAVd1PsGEbs8v7mj4E
zFy3ffso9imHrjXbGA68y+xy0zrg6A8xQwBYh9JL03XxPhr4r6/jUtAugDpGPz+/VEUEKDxYaapE
rHxLxwYwfYJfpY6uYLdX3Z+VbtDb0n5aeeX6ZC3DD0rfZmmgA3Gai6Ns7Yqjk+05a5xRD+2b0tg6
+lrJ3qOBFujI66dT6YAb9HWchGZrWDRwIH58KyQ+hbRUPX/45fEjRbMpi5YlO9dk7uzUD+TT7YUZ
l2dhtIAc2d37g6KfhaEQkXRgmNVcFqN4LcyEtee9Q62enE/vf2aHCgPmURPJ1so0jhdOibc0AWVj
IXBYhA+1A4tHknUyR5+S8l164TW7TpzKfvJQmb1+iDQO+l81uN3e5vyhnaJJVsZsNbRrBxFfzMK9
DlnmtC38wu+NGxGBti92yryZaCUVB3mUn4rlO33H3hwFvfPsjwBN1ygKIow4dXwpKKZwYqSjnYFF
8GACIkXnnnZC36jCWWnlAi0Di1P8rORAjTK35Wx1MX17XYU48tKXXCawFBIbQQAdA5NzJM44ilwx
2QaDME9HuNvzwZSbn0LaNFqY0H155sEa4A1t74QGFkbGesI1ZkF/s5MWowaRPWOJ4iuNKEW75oQ7
6BeV9N+cNEpF1p1Z1dU1M2Sxl1oEBODqLurJwd5T8QNVen8uw6xtsh7ZBFuNkwVf2OvWVE59WNn+
VWqDTR5ECNsdaXw1/2pe5tAzQHWlKvhUqwcpYz1vwCQfTtN4mEmDmh9NARrYdus3oLAtT461O1ti
tze4Did+ilp2U7+ct59HZBcvF4kIxHlJOG5oUL9+XPShkpMpJQ8KL/gBVy7vCGQv0jlkaGrqIs+r
m8+4JzDcZrSuivWGbFi9+XPTHnVyJ7eGzqVorb6HXZOuJhKflZteK4Wqd7BYU8uo5QHahWAHmC4V
zPT0+h01iH+23kt0ZjhvcgBPdn3+O2ULdx3dA3h7k5n45GENfQHxoWmrTXHFH5oumNNMFMJaGmnZ
mYtbKvbyNiBNuk8sfXcnKMVTo2Nf6B/wYQDFNRBL4WMipzd8PnXfpjwsvWy1Fm+sybZJnbaFwjC9
4qpm1Zfd9spruwA4t9ETMzYCS4g2rkDP2KUNVy5yXUeUMqBTinyij/Vr8RNbZ3GZNeRAVEhpp8tZ
uiK5/6DoNuvBuqAHAaMbVhrpzL5UWr0W7Wk5BD/yAz743OVlJR0TFvw1mqkAOSaZN0B2BYFHh6j9
CXTLLMpHZzNESHSybixoXpEU4BGoaUD0WZ+y8NChnhGcFMexHyeO578JasYApGX92NtGhuX/tu8g
3loS4y4udKTgeFocbXiofAHZGobzdeK1jv7dG0IVUi/a8Qx8ayw68VTQunD5oJjegcMfzAptmbCx
r36dPQsQhITD7xoN1TaOyVhOkLiBCicltSVdJm8nzW1GzLpVZ163FpNIBydtBR5mTVT4GAKhHQ7G
nX2ag15el5dFJ+nBot0+hvDE4ITyyfWHzPyHE9cU/K8ayXTfKlzyogPQW7DY2exnJOf5s3nk2tqZ
n9JwAsY17k976b8PNlWFfRvOXyWWZZ6DJHCkPo9mDfDU2k8sA6ChleTDjjGwSxVsp7CMXaBh0UQ7
FhjMJ7KBE2m4ovvmfawMQHnJ66HnVBMMD3598uhJHVS/60uKDYlCD6WDLmbix5HEispLvXYwkyvb
wv14ENRfpW1Ft4DL+Gx5cL8wOXObwx0g0JW04VJi3w+Q2CmfSFb8S09Yq00cKFBPPeoArd1CoTkx
Vu4VA6uyBEU7HemUF9fMrfWAQ1mgyUMPg4nWJx/f42Dr+5HM65eapO+yFCnHO67d/F3RuKqdklnL
yySAi19St1kbR2IqYXl9/aUQuwt5x99byU+ct7YHqGgtf6unjtO1y+yyKPaDxFehN96kyU9VCxXA
WDqZPZuISnF7tjbiWXesc+mFlH/p0hik1c+Clt8S3BcdIQ74rfeZAyoG2Xqk4vAlOqsOWJPngAm7
TI+Ip7HAjOvTHPffq+d/P6DLC84pvPzjphCfMjoMmlLO+/ePFaVJbos7y/Pcuz8L8fF1jeSqvZsP
vx2zQl2nY6AowWfTWW3qAKfR3jv4BkQVZy3fO/nzHdwrSFaLk3XKpgLPGYPYcm2Bug7LsmywJEPu
9XDZMKl0yHeMK+HUVx7tYyh/vSkNp5mv1ohvR2yJ3yTH2N8C8mtjX0qIV4z8pvW7pK/90WDd7P81
MW8ty7go8B0Ou/Q1q5c7QHF+BrZ9ItG51iWVMzquvTAzzwuYvgS9H92HjdSza50xNMQC2A34d7ic
lJcU3K0fOCs7Jo/WY5qARnQnrFvCuj5uXGWK0551fZanA1iHT3wKKanfCeMP5BwJlbQsS39ld16q
iB44OoTmu01bssIRHRaqchA4d9q7WDsdDU1ssF7cMrNLsk1+zVSZQkEUm/mcqbhrFfX68N8l9qUe
m3fnZALtzJPR96QqsDp0qF0JERnUbucNKjxu2jqqazwRzwgqLWjzsfLdT3b2qFXXEsfMi8MMgbdP
6AdJNWbwVm3KrFFp+P5ydGSvzBVmyseuMROQTbbqXB0DQGnV/NF1UJKm6AbolFG1sbnsKqaao4mI
grPgFzPCA+FSkhL4+aPzcic5zr/msfSCIdY64KAIhouCurRSx7bf2zTL25GV9itio00e5N1zDpEc
mK3A8Ys8BMLhdG9yStyjMxrp82LPmkUpSoAE/cxXQcy4tb+f7qJ9xrFK5fLR6aiVRG3V3Qvr72Uz
06KxwDwk45lnV0yrGATpAO6LE/2D+f7e5oOCnMG5lfYik+A5YwghFZuOYZFTwLeL7XVn2yEavtry
TH4z5mRyyaoaup7Fqvzrf6QHOUzJnNYun5hjyo/B+0XNbPRB6tvUWNNxVCUQq/U6/gjFNjMf6yeC
+2aBh4RsFNunmN7m6YJg0rRrI/wKOYCpqCaojqSLmTnJul0I9bX4FBcI3CVkFlRk8dGJSHAcOiQo
gJ3kWRDTaW2q6f3EvBcxoFGZP97EfG8FVWM2qHpgd/K19Fvi1wIXNQ0inksK688k7lO7xjOfVChX
SZgDAMlZBEiA9MuoWHGZUkQJkpDhoS32W5kcXawir26e6cwOScTqhru+rtELILkh7SrzScdHWftD
G4lS8MxfsiCyBvXAGYu7dxFH3xWbeCRB9oeNCmPl28tPquuPbWX4iC15Q1Pz3IDlAOxu6StMhhv2
gmmQXAevZD7YjJnDjaLc4rjyDD/STzgI/z/WbGQ6dziXDBB4zB/G8hIGVMvp7N/THozVqTE30eLi
SSr6WSmmTHlkYJKsM7dl7Q65Ijc5/Y9VqTIvaxpG+a50Cn1Qjgqy1Kwa+VFLfOdpOtNWU+zvpFWu
c4dZBWnWrvu6HZUpcHBvHShMtjnQCyHywQzMu3YyVi8QUWq4GJoOig0BeGzG9VV3mxNEH6KmY58o
j2QXVv/WWdsVbEuFtuEC4D0GfItcQBZEOvFCuynj4F+ugJgmdhqGlmjXfh8Tu1kpTbODRDCnHduh
Ungt9ZC+Lc2CNqoz9Lea1O20mjYZnKTLepzjbd9JxSQLaSyv0WSDL6BVAZbB/0GFshk3Ekrzhv7z
VwRvFocDK5Wih95AiGY6h6Hb9/6g0+CKD5GQMF15MkAZoKI8vp6nF4fxadURNblYBL0GnlnFLpHI
OnaQYrfopaS5Ms5YP2BH3adcamu2xGNf0sf4UW5p7E7719RwnMoGawEgif6/67kdRvt02wP/OSQm
rM8mcZyiaw5LEFMPLBaLaHaSCeDgVgtV8kY19x5qqWKqHXXPm9GU92Ip3j0rMLA/cu706ZKNeYQY
RmYeNfkMr1Qby+Oi/6CoseEwUXAJnugVzNqkkAP8NG0iyFH0WT9PQ9s502kxWgT4zr0sJ7VdalVT
6TkCb3AoBzN9GTQ9CekCnrZgod2BOGoa4p97bgvwyw3p04CX+blnQBGRUV1lYTeHYJjNZ95iMfeW
nap0lmI0nNwzhDqgIVuoWkzqjqY9JL5CBkn0JxpZQ4r9ihCNmLgzIJOP0Gl8u+xzCgzrBXhMKNy8
N3JmMSqf4KOb5xyKbOZU6VuXfhuUov8H1Mk/7ADEPGYzTroylh+J8z3UpnmUszmLsPgYbk+A1Q2J
1joBrMki+azxUtCUdKGCi4/zSHp5umAUF7BDNt6dKYIKOKF/tyjKi3h75kGCtAp1nnQeNFfbhYRu
Qvcro+F78B7RLZmTzxZXpb5dg9zUSGUkO4GsVaL2L0eQkW4rXggQG9TpppRjRlNxsy4dAccSxk7b
QKsNDySsOuRXirbIXh7yXkplNWxLiYLqaE8dUhNubc5MzCWtkSkClV/IiEC83WQ40MBXszTK8s2C
e+K3Hul+vM1VBAxb3NXU29Ol1hZcTkW46/ccoLMBfyKU9oIscQmxkLRKyHeTx2pMFokaQAt7s//9
EG9uFImR2p82L1I4HOgYhBwMsundOSwG4Q8SItrNaS+XSBs1Uf7jDpoKhltrm4kp4GGQcB1PjMoi
33WFSq50DjMGUGLbd6Z2FkxgA8oijOynx12nMWkWH6yQKgAbDNQ6Q5D828FJHJ1pWnev83SbBINa
HmPi/xsEBuchP2A6K9b809afOKe1MHlfzzAMNW4EMKQYabFENyqrjhkm3JVTS9Sbbqm98BglERcQ
13d+bkBG5qOM8UqcYW6wYcAnSfJzfwzg9B0xZMTuI2C0kwL7BTl3gEkXb6gwQoTG7S/BcEYdZTpk
e+MwzQKPun7u/EHU1woZ7IZOYtr6X2BSoRWtCA9goUmhxIdRq7rzjVSA3Drdh0vTUQdnNOxG61PU
va624rOx6Tqm1zaWJY4+9Iu1BmFuwWMBJ01se+C3bLlbDRzyjOPkb0xxmPC+lTVIipoTqvxu6s6m
qbYkNnDQP3rnPjE2imOWtHF0dEQ11fVVbBELnTzGXroOrAAzGS7j7hcqYl+qNz55ILT8jAkGJixH
ThLchJMm6Ib7n+nNH9oOdpfJL+IFfMaSnhlTo53KXcpS29VgUPU2mojnjsMbbNPhmVi41+FEkpXv
8gmg7psnFAYrxx4sJjCJO1qnirEwahx/rfXRfzwhjrN1ArdmSPs98mM0kCao6KVpRkApbdke6Dt+
59rOu3tiA89pRwRnUkmYg97CJFwPPfrzO+lx/izNf0FXH1UoJIuDsCvw9MxmZ9Nb54Nd49+u6aMd
OPY/+6bjlmcdkiFNJiPURNgN9B9GuugyHSIr/oyliLGPFvn6NT9WQka6fTF/RA+XRZez9jqafEJj
6JE3lx/BiVpaH1hqThxBnGHVIYXC5bKig+a7Kc1tOsH7SkZ5719ZKdsdYHBPmWA5DJ+ZpgvKQ35I
rRce1m553gjEkwoJV+/Bp633SDX4oHt3r+02TZ6pL2rmzrUVXQRdwufUgpd7v0wnVj91c2/JmO3D
gczfGWU4tTHE9dJBcXofsiwrqIsb0DRBZlaJtC31Rqvltp5U6eDbMyprFA6w4++WiZyP7pS1podM
i3Bih8gxbRWUB6696CpWWcL/33LEZVfLA41TG18DeVLjVikWY1i2pZlku8wGam+WTU2aoHCKt5i4
llNvf0AYlVlKDkI11V4EItSyNkQFDtyANGCi3TO/EB1dR1RYFsM+Sx6SiT8t3NGFGS4Da3Q/bOwG
z7vekw55xyyH+ZW4g4kn6q3udOEpCD/hR4tPPrRRXhpL6FItitdgIEVYHxCeutFhA7GvHc5oaiUZ
PG+VhHrsS3eRSX8cOoXb9fzhIQ9KIrM5jmwjV64H9dsbydqVmkpLE+2kDRDVgnI8Yn32gSKfX6xQ
hFd9CVMxPZfnogAtvrtMYKe+VA9/zltuRcJ3DkLloLroAYJ2XGszVCO4zOyxiTnUc+OWLjTQEtHD
zTbDFlCHscYBSpIF0+5AROkqTvs+53bk42gRI0R/m5SP3JShedo9weyV54d9vWqQxhVT9mwWLra3
M/Fbxxh8GMBbrDIMqNtX/YNEOaEtUiGr2VT+YWRvFotDSlBhUKtQyM6Qvr6ElCpJy7cRLL0yTKsa
Pboq5BJZz2U3L1IHjpwXbFQisT9n1pTK2qnEjY6wBXL1ozWKFFUhO9u4kqczPBgQ7Aolth1rPVQV
WxbgLZOglY/hFl6DBNeq289Y2Tnvt/p1SG1NopRbrXYwtzznqOGcg4PYz36Til5EqrKbmfPAICCW
SZyM4SuummfO/YeoZqaI8kX+7UUyFatsZkLCaYIVYTLqMkKRWRZXaYgYjfrJeF7OTFO2MOWDhXdM
qv/aZkTG8TqUMHiS+myZBH5LeDk8FztfThuLP8zAou/FebDIYV25Dzs3QT5t8FY0zrG5GNxqGGpu
EG/uGA49Mp09XX+gAEM7Rg/0tlmKx81pg7dSW4an/L6ZUgk8bXX1FS4xjddLfDtRlSreYSNZBo/e
zoMoeR08k9CrLKKw7uq+VDBVwXUtk0x3sIh4lOI/lcc7bckJ+JarDCR9e+kMPHuIy0+npiuXygMk
PPO9cLlP7X73BH3iKeNVSPlRwk1IDTYgDl7AOhA4safRekxjcqnVX9GjeH5UZpbDqKSNmMCvrscm
aNqfJvjPBNsRyRLmKLkMWB9IQTmbJMNzTcLGN2VnBX11HrH0o3xSD6QYfCco+8+4z982Hzcz/gSK
2AqADqYAEBEiyIUa8jBY0tBC1xQehifvpM0UDdUmSaoQdH+1bYzjGww2yBMXNsJeTWAV1lj1+Rq4
NL9ESdExPN0W1/Dal8p07Y/D6G7mbo2ASk7Vv2adQ69fm9KmePgpVBuzQ1IB9QLaN84PL9/V3CDI
MdVanvmpwQ+PBlwKdBw26WnQztXYq+8AghhTnvupvuDgXvHUzu0RkOiDssHL1jwNvNhkWnGiqWey
JShEl6XWsayHWyNnppimKfGnvtz+LOAVTejlXRI3epyKNx1L4/KZ5zCbKfyn/00E6cYLAAjIaE/1
P2ohRlbzc0sRaLY+uKVl0SgHr+al1amOZqSvR8XbEv+BURd1O3CpTmOrdTECZ+USYRZsgQaBnnxY
0pP4jR28/MBwckTA9bMJ+/jaOHEPxu639/JRWgrL6vDplm7qVpu5CbMpBOMyfv9Q8LR4dy/vusLl
ndZPGpI0YQ/Z4pchKf0OfLxD6Hp7AirEcaXw0sKhxC69fM0xfkHrMCUJYA0PltwNadYevt0oLxmQ
Vh78DiAshxPACePRjWjOVtfHTJk6mv5GaGdOmcyxTxU9P+4gDS+gKhir9A2tDi9o0g/woo/QYtkX
GfBtI1/05bG6lp2Bu+Z179XhUOT3xKzqY6P8d7hTtWEzShbjmTK1ScT2y097NUPn6LuidKv7n8SZ
9zOhbkrCfmBr1rH66XYHOGNzy8q8HsD+vjakh65YQPwd2IhudtkWbV0uSOU+Ego2Ozc1Iv1/MCgQ
+/X0o7FeEDiTlyRs4HjkhaP/YxZ9fBl8CusQbVbdefLmG5sLL/bFpqwoKKzlpJHvje4rTC/oGkYu
NkFpKuLH5ZSiY4xna6wxgfTKDvf9qnWwVjf1GyEzLeNCN3HZKhgYE1Sa877kd9IRegQj+h4E3d6R
di4FMJodn7cSloM9ogpqBHfP0qz9db+zh2OwdPoC/qxouiszFn1AoaZJfGEF/99cbKrNnviXdl4L
BIfW2xk38oYgmiaEct7noydMQYgvK2ko1yzlOMUtQXjUHoy72vJ0Fb9PZJpHh0st1rhB3gTkfAhI
og5Fu+a3jj4QojiNs1mvrvPpJuwU9CgGORjc3THU7O7TlVQvK8/UwkHEVlygSyF7xeFqRgho/P98
Ez9MCh4n20T9LDbD3qQYrW1boDYA6QghNBfS2uO/UuYOszARFF6y4Z7lSM6Y7GdZCHfqinC4EDD3
N97NkUTxM0ziBpUpqgIab38hMVj1muJit6c1gzeXUxXPmJZz+YO7XCHtYGc/rcGeW9FBuGJDVaNN
iTcujnOnk1c5VS7gsTP6iOhETtEkOAhfHnDw3Ln2lnzb3hpU+rWAWC9bDdWBtxVS8jQrvuGn0ylh
R4X926T3WPV4Tw/4Z9pQsrsYFCSZbdh0MRp2s1fmAqI3XVFW+cPoGjyaq/aUAFjM6TKSugva+w8J
q5uZ0YDTQ3j989ROyKpvnWr6WaR2pk9pNQ56SCFUJXkVtIefJYA8c6+29HBF6zxRWphluSCGPNOS
l3S9+EqFvnKgJ+lMbO+NS764W+H1PByouJRlHjobMGBsBkczLzab0L8SaA60LTjzxtq4hTgL5Ezs
ssjfevmK8MPmsAg4rTyuvGwa1ucKwapPj+sX+TfTsy5pzGFmWA++OoI9+cG4TUSMnrKsFwUFwjJi
v9MPneh7KzN6xOFLT4jB45S4SXadvkfuCrp16QHYVglPG1lDJdbTohBlmRx7pbQ9LvLaGrcpdK4C
CU9ZVezxTJyj0LWDMYnUoW7foWTmrZ1XQdkb+qLMXnLuYh/elBc0QGuBD4BxSWguOX5Vaj3xGLKa
0Hn9phYaO9//8HJCqzFCq+FXwKvn3Ou6uUGIMga/ctapqWMHAJCkNHOnNzSSh3XAudLwDbib/r0l
uRqarzx1hax17ElQM1A5ibnTWKC7isa6I5lI8nsTdjVIMYBXKJ5xejku8ZsVPs+Bp/amhfVInC1C
r6xPK1geBkkoicIpFYKjpR/KICobiGHTmjlko1BcbuG/m/YZZLFywnwXZS5FhSJf1EYL3PA0lJNY
Mas9hMf9D5brh/kX6PSM7q7IE5pdPCHB4QkJizhdJrIYafXLzCUPHrNYFcz4GfkmLzM85xvKGgTV
/+NxfGmJyo9qd/fvafnSTJi+9d0anJVYfjEII+PaBrOasRsFdpWqDIVC7SVMKC0Vjfb6aV0FpaDi
e6fnydz0hVO4uAuZF72NJA+BtOmlo0ciobF1eUFY7JJ4zowNGV0pwGSNTucLEcBCu5kImzXTV5Ih
w7cRK0/FA4l5R2QNCmwiqglD+xgab8mPzTkH1iF5I5T9wGKuBv8KupPvupH3DMKSmW1t2VuUrC56
VIWjXY8cusDz5iz3Q5N91su2eAPC11gsMUNLC9Tr96MNPRTjEfAy65ToTTDh/N4uNLOy8iyXwy7i
wwAz9zv+VXQkEuqHSoDRFmqgfXtGB6+Rhv2ZL3V5G0ADzCLyLv8t1NwP3fBTeuO8jiypY2TUboNJ
s4+zPmc6ujs7e9G8yqtB/kjgC9mos4/JrthO3E0QgrenBSyCd6FGNJqgEGXxRrZuyZFVfjdygjZ7
Wi6YX1Wb57wG2+lrFQ8RSXbcXCKeG3PbdYwwKn7eP2tTzx8QP5bDsDpbVW2cDBeglN23kf2TDblE
/gWnXXFHELMLGiXj3blA2zjwzyjcqprhIowbq5jW6E1Q601v2aaWhKJbQXYwGxpaccHeIFCj1wOF
d70GZPVUpn7duVk+UIwCTuzLqavJpMAxmZ5t2r321RV7nmhnDw2sv1PKVd9mdZxne5ggBooPhwpH
1IhpJehw21PesVCyPFXUyPxwLQbp/eMHztG2Gw/vzujgp2Dmx8uMepuSkwFOm4hBBTiiJFv2CcyR
b+YA0L6UXyy6PaWDJ8eed4tDqNA8cnJ4Bfc7GJVDILAs2kwuK03dXC3Dx4AfW836OIbHdpb+ixb9
OJdY+GrVaI4VTRSMqblpyxcgv5dvh++GtvbkK+tfJ4tRKv9Do9EiJrAD4x/vo9XehyxbtAimqgxQ
tiLrubFkrO1RZ05jHtz/1BEE4AbaKi9RHUjKheGcTdPyndf9vT5XiXvgh94ZyKmRZHNq0gL4ovFf
4ZDSzrDGx3FdeLRzQ72M0CQ0SFZA0PacPfjrcX8axx8YjCNdu+O8iJifml6UuzNwT8kJSLA10PzJ
dhBMLoTWu12VjKdTYnCXY3Owqiy/5Cm++W2lWSpQpkEuO9kwmtML+oH3QM1DE8qjTOtCCkkvVTgv
4pa2AWkw7QCNIFh8DhsYcLhwL8dkVkCqkmomrOAoUN/Ux0lHxZuIAMVtGyGQ+WsKLRl3eHP/Cbot
hDjTd00W6lBvjdBjupk6pNExbzM3aAdKaUPor2e0xFOkjQekZ188Ygm/vyIoDa82xZ+MGDDkxWVE
F7r89RIYCNS143AEstozZFtX0cU8IQH0SIDmd3dtbAWXx6N+VFME56ILDXhFugCa4D5bktEF3raw
lBnc1hseZbxjWRayxzeug5EMcnLo+RCdJBV2M+00EUJuGEw5kt4/T6bgGsbBc8HfWAu0Wi50kfPb
WsMgSbiUyOWNW0COAvyngJfwrAZUsnpszUhUqNwBDZrnfDc4bxYVya1onpGFIunvsCF20sKKR6ll
2WOJoy4QfnEO93aJ1Kr40n2pdqm1nWBp/x1VCCtuKtxeHXXblPo5xWLOQCDO9hOQDHFsJnokOVrz
JJGSjvQ6ippBKnJIdI4IegQ9tlL8MawfgtL5DZNEPDKew3ncAoUhrRA87dHk8JvG9pezxchh1ABy
SGy/PvIpnq/mWInhUf0o+PR6gsZicvBppr+N+XOPg9Aorz/0n6Ud7OiGaJbRRUgMCvPuF7feRfFR
ANkntIS4RufQg2qEojJTuTkJfFiB0leAvduUUTzzMTVPJiVerFu5uSRRQTHl94wCbCb2Trtr7bAI
ghRTREwfB/70eLq1V2zkchC0YFhV++uxCHL2JUmG18UNDhPIeCQirm3O3IWqjEccN3uX739FmZLF
6OYH2JClatxYRFiEru5yveTEeDEZLd98TodEQyo2/8s8CettruwMO+acv1gtFtvJr6wdz0S+FgWv
Umo9KETKxBX41ZP03+vjHwFDp7k8ycrQ2Zc9qPsHR+6tf82kSO0oWCGAsQzvKE2puzeD20iLWaon
YT+EHoVDEPK2VAR9+o9MmSfd14zkFCpQueFdvhshCBWtkFzjlEJUds46LAL6gGAb/5uRsLCBFNIE
lFHxeXR277GP/jsdf03rik5ToOh3jhAMS+yBdS2nFQ2i7ztA3+5GfiJkHZ2bvh1qQcs82FSPZDgv
iW85A2/zVT06V8N7cQcwBgEawCBt1N/pwZ+rK4udhDfZLu+L2QJWi8/j9uekgR5yy5LujJkal3st
0ZkVX5u0VH5buY3CTSIj+xTHuhZHjrkzpvqiyQuXG3Ottvwlf31qOaXow3Y9GR6KMSWkZoxZhcHT
SeIlsre9CaUljv5o6n+cBSijvCiwBGcHhsDXlpZm7v1yh0Km9PPCFK+axSQOF4aUHe8+bxSAlxFm
b7ug/NwBYOwqnuWSM6iXlw7UL/wxwvU87B0r9NEdQV0NFsfn8WyaviyUK/QkT8Pxr2jnCgTxzm2/
1q4ldhyUba8rf7IkZfvdPHluWQ7zqQqPblkxQUMr63QESr39hNRpQsb/xcSHfow5uqKU0LXVPF5T
828Xx3Ox2J3ux4XVMUy/aVPBaCdm6iaBscN9snWYG4TlX5YLcov0GgmmA33ZK/Lbae7ktNHReyTm
iSiWKUtt4tqcXBrAzojIuBTEIddiTJFLVVA3f05SvaC58k2SgBBvtBQmOcfwMJYchHrkuGneZo0r
n1ADZLSlLC70TRQn77uodYDVEez1L7pikd6Kb0B44U66c6zLfzzWuw71XykdjAn0QJy5SCwzalIZ
SiAwLDOfm1T5QQ9XY7OzAszpw2EtDMmeIWuhby8cv/I3qa5Qf8ftHHtkv1se+WYteTWt8+5W9Add
cHm09qikDdO/x/OSAPRQjf8IjKXGt4BCYxmORxt23zlGGpVs68sKMBb121i8ZJy0mOS5uE8Oeh0J
xY70SzTOFzS5uRIlVhy5rhQJINV8oFg7WuJ5l3WIjmdWRmCnO70tlI97DzC+mCp3NO6b9zU6dAWZ
PVCEDz9Zdjp+pVmhlVAOrMYvtAQVQnEhjxmoaLa5ZMWhjjtU+Wtnq+IaBAGAXLlcRP0WAPhLF5FA
V7DOlSvc8z6ByjUOAnmxwXh1/vFGLoOo0EK/a+TBVFBDnn05pZey5Otq5JmxbP6WGg5MofuDXEE8
ljT0Xl7aKo+RG3H55Dc9/4g23wQN7cmGVgoZV95Y0nzk9WEJ70WWIriPjDlTr6KJdeQEU+uaxgaH
P2ejHgqqawAcpVBd+0/XL24LmmtO7cvhKPdgR8l/Sxekzj9x4di4WXQEKeCvf+tTZOeatHMpLXsM
CpKN51BvwK5ENxjOEu9Qo1sG5K4be7j4zZeZhFiIQR22YB3mTURoHDI/Rs3bQbM/E3m42qhk2Wlt
9oDn650qFzMWfpRD0mTUBISmyOFONkVuiDDN65W/+FDl/RbRfilFrIhIYcKpvUXWwU8dy8fvgZJ1
vQTd2Kkua4wnUkeklwJfoXZHpUvQB1D85FhqwS7IoIQMf7asDj4VJyADdsVtq2WHAjisDlztLiKA
zy8qAsoVuMAAQeja86uPXF3J8CFz+vKb46HcaVgI6YgFsX298SOU8k9IrYxIUPhsFW7wXdrOqoUu
NoIEuHyxZ1lmgDUGJkA2i1VketoY1ADiWN/Q9BxdJ9qlXi7z2KuPrmc/PMAqPD2IXqhEzy5PWO/1
xX+NAp0+Gqws/Qo4OOwu2ipdsXWP01HkebsHmLmF+svxbvSdF26gMoXOJzEGxkkUh6kBTAOuZYKl
PH8seSKbfeGR0xKfH1Ae2T/VPuPoa7CVIq5Et+UKhN+zt2eFfFALeqJ/26opE2EQYhLInVXwen9v
kDgWgp3zksZO7JUD0T4SHBIT1+/4mPvN9gYCRY2Ma4Y+9PRjxbHbG+v2olWE9sK7/Y5gEahpNJD6
Ls56ST0o5xnDCWPnFdn9SXYAcGzN4eR5Un0ZIhiX88j4TfWI/hvNs5Mv98cAOODzyDh8Hyeire7u
3lMDWvc4Dxbh4bIy+af56y551MA2hNeijgA5DD2khDQnEMHoQqXNmdf55EebWvWa7GMZzF21lk6w
4XcSXyAgqxQnlqvnKdKfNVyfVE4TaHDriJkatf8ZP42dg3legnqECnyb2T0xcCwZ4NVDiqhQX7Cf
vFdSNfnpWkRnBFkH5Gxa21zWLNup6Z9eOeQhtvWX5T9012gflmm4bvLGs9noS24EfujBcTlt8C0C
MSPDrNvnHTyV3vR9eDlgCP3CebME5k73tw0MkYC03hT2PPE8O1z65rIUyqYutudNU9VmhK9MSyYz
/nGPiYU/4vlzwSMv5Y0RkABq5PkS72O1doMf7VB+dthWzFDhFBDrPbFA4m1eNSleNE5MdzyYKcUe
f01XtpUQSsbFu2vHt5FkyzHRv2bd5yX2e40JjUeoJb6EFMOo2WH/c/QQAjbMEG66jyvw6ps+SD4w
FzYF/bgMuXMRPpzgNoU1H8YI1gmsZWbgfsj76UeTMqXNWkGhaoj3QojUxNp7BrlXeSgOAdjUXxAZ
VOpoHRrGB5cLOn7dA9NR+zbqJOViDekTXY+I7mKk5MwUw33R2G+SNffU+LwAtGPPtWBbcpWr13KJ
usyYTCJJ/2IaVJeAh/DesXfK2n3i7GxqvjfUOhvQyqIY7FNYgdXz28vjQyS5FGR+NVGpSU8/bfJQ
zzzBluTdIyYetaUmwO32iu5BdYD5G6WyhpX7dlc+cl+QtTbxGfPlvwCfiX24TZ5/PZu6ooTmRT2w
Yaqgv/Qic4jSpuSi6lzfyxobfxL10oe/Vr9wVXRctbmDgDO5vbgxiCWYwHwDOrVf9ZfnxNkIlaYN
8idLsayGR+VX82ETDTZQJdvovcP7GXumq037PgoSo57UmVL4+OUEqOy4IZDNxED0Oe2Qp6XPy0gd
rko01AnmPzuDfN5YWJyRVzByp5tqf34kIU+AfI4PLklC0XE96d/4koKrWE8jsvzIsI3HAzCh5XAa
TStZzHkxejDUDJFL2yBUm256e9YT9obrL1mz72MSyZGRmXgU/e4Uxt/0sCgKhdkDK9AvrYfhOCCB
K3oE6tet9jbzIJZ1SATzvEj9gPdedYSCIJH0VTaFOQsbiJBtP9pZ68vrJS93SUBS7DsLIc6zOQ1p
7J6CPJr/RLW5h/erX9D79R2LuCl4k/FTZfa6k2Z4y6U/QR2JAX/a5ryOp/EzXUgZns81aoLl48TT
/7UXeazFDeCGfJcDHCXjn3qx1TyNmp3uT61A5CAMkEOZZLQ0wyAWSMa9bmvmwyX6gu9xrcSxqQfx
ttrx2cyEMXVeSSOljFE0NMQQwm5PGkgLG/QmqRULbmkxSVuAfF9n1Lc7Ejth4ovh0HyNPexZk1w7
Np3xzUkq8aABMqOnhA7d6gmB5wnGP3S6dZFigaySOvjt5X9v2vDSxYJ4H3Rqt7atlVt2Uvz2GRYp
C+uWWV8dBAcosdciRiGHOm1HxdhEYCMWgRfdt5tSLrtGnzmF67DROGrPGmVIVu2M/QFb2nt/TqQ5
LT/nNpbC2KGaxME9eCnirBjgzl7snTEtmzMl5QO7CzI+VH85AJw3g/XyO5prm8GnRz+Tuz2U9t7q
kwv664zPd2zgFeFiNcqDZPXz2aWx+IQQFv9sDh/SsuMQkZzmZTHvCPiY9nDOU3iRVbtI1X6cHZZc
FAQAnwPLuio2q1ob+swuOGXanf7ajbU4ETOLMt9tP+7qO60vkewg8znpLjjR+coqe9P9LkUbgFUx
1umHLJlyzu3j3qCvEfA76ciuFfopJEf6yw+guPxyfM+xbrODjEGOG+hGngLCx0pWAFKJiZYyMJvP
HSD9mrvwhmfxcyFrlysSp9rG4Tzozyog5DY7uJ0ZO9O0wzGih47WtJEoOd82Uk2qwwafvNd7HqU9
hlxnkB//pPjdSvOywH7EOuKaqwnHZq/r8y63GPYHg5bF8g59wQHqyDHn4vRCX46xmpBzPvBNm+Bg
tbJLvWByr4C4ZSz97UCK+EAL7+LzYJ9yQBPtxv8NxClsYXxGgQ9/YF/zyFbOurprOucnL56i2WGz
V9pV1vRwdxfWv41BO8cDsKnAitP72YszrO1MEDI65rhEHt2Nm9iuk/ws/v/ETTYakHeiqJWhcOWo
b82VDbjrKc+7Hzco8QDGlzKMJFFrI4amC5jXKzA8reQT6lJqBSItaj/m3XCFEFpvXPu3yM3pi9H5
ZepIGHdScK3NUjA/jgv/bNyNRm8UxquXSZmT3ILgQDeqQ9cZBXyh8svRGQJX/Hf9NAOTa34ZJjZU
l0/7rXnvnp0qCxzuuiZXFxQ27U2Z8LKG3HYJLS1jAxe/viWhaM1lZyq3GRhbVzkBybJDXF5B5tRk
U2jonBT5oabLQ2BdX500kB72tyYldXJlDEgKPixEWRoKGMW5mZXuksXRjmb2Xp/DYhq58ASTekQX
VjXm/t/9DXrJMWKdEVzqO4EThfN/wjqj7yYn1snMuyM10o+m3tlxABI1Z/0jsKBsX5zzjX+zQZWZ
1aG3kRcim8+JUcjJ3CybnuhaS5D/eVm+yjt5cD52Wz8ok7e1Z0W63ECyud9OlpsN0iHT4pVVjYia
BgST6ebc/qTSSI7RyCI+jM9eQEeP6jhOPBdv/5EsID9I6scKtzH0Cw5IGzw+tAPBTXunE9PTCfD7
eGyEygzNRMrmigNApsRlg7Pjet+X7ffF1GpkIQD9UdM7pAtoH5+WNZ6UmtphG/qn3MJrU/1dHPkq
1NUTuUuhcjDu5GMSVhi3xfXPHS1lc0Sk6OoP5SP4x6N3eUe13Q5DrxGEJyRolbTdhLU5kEfXOvr3
CfneixL+q3/zn74sqnqzBjY+I5zybEgHNLe4d586EhOe7anzsxAaRNJ6VU7T/kWtauhL9JCkyzh0
1zuKuU++JVobtNu+Q/dYd2RP/jquNSQTIS53s9mJnvkAcZENDJLHQWCAqCKKZgMA/6m5iqJyUJE7
dPaVBUvfrGZiPHbUJgRNx5QGON2gsTAk7/02zFFpEKdI98ekFKr5PGU2zHaS0XVsbFD1pOiwXSW5
b0x9sNpmfj1eWSh2jvodTs4OK09vf+VlMyNN4nvfTr5j+k4Km2MiSWAo6AElHU9xaNJa8KuMMnVG
it3ek/6FpSAOeBlUB3hoU860MRrd2dbe+Rq3UQeHvnjAd63XJfkibCi63iTAET7Rp+/NknyixUXk
3HMTfsgK89uLXm6QYh/UYBlWvHF0X34IrmgnqO+WleG3YPtQ8ohSItpe01L1o9S2O0WkcxGzV4LR
hc9BtLqBdklTzYGqGe26gc3NU4+4e3QquqV5TGcIs4Vp0MpU95bwQnXGbvcC+CrNt3G9dWs3NsJG
lUmpqXKfoaIQtYAxCx4gQz7IdIRTaJ1c/aMXrFcHNITXGS2I4O2k7E4jvZzMk7gK1NfwiZGHsMpB
B7ZYQEde2XQnImkoJBaibZtKRC+IlFN5QqX7uk23h95DUV9J94rG+zBEk6WZQyv/nWSyoKWx9KAs
ToPWvgva6f5R+VqMiW579CbWD4IVXN6YpRstoCHo7nKPI4O9tGZb2W9kL2O1EfzAGbYow+HzpyQn
XeByTGfBIGsYChogJuVt4L46Su+pJ0WVgnkJ6ZrCKvngZTHN2C0d8WUpi0izUxQIJ65MwRacwdqI
HRqbuE/lIgCRlz+Wi8EHi1jGEd+9m+HQtlF3MMF6rLTn1amtyMab3utWz7Aoo72tGdd038UsLbeK
RNSfSbbW2FEu2aoAnDrXP4Y/i1Mipbpz5YYL5gcd860ZEQ9tjOfXiyQ2gXyBqSyg/9ixeqcflLTO
O0WnZso7CryZ2M6rH+lwDumX9pJxZ06wNCZ4Csr8PESXIU6STd/k2AOZiuDxyd0eYUfqfmwsldXw
NDcZIh2rs5/BmRKHJWUanvrH5Kn+l+owN8hh8Ulb0l4v7+3GZxN+jWfG3ACG8hClP1H2WdkH8P5Q
wYkrl7DFMRE98fA4nv3OOo2f6eKj3D4Ov8y3+j6VwrfILp8m+nZ7/MguTGYc2i0712X0yxOG7nMZ
AWXhuIVltzn4O6aLOz/jbJkjFG2gtMMU23AeNhIx0CLPt4TNicTWdhS7ViaVawVMsNJCJhc0jnVj
9vyzy+lx3UZHl3jxbEr3zPqHWQO0q6D/VhX2G1xrin4Lf+AGcgPN4r2VO8aeHyuJ8ng5vPWqeL6R
xUVdPolJOkdQlT2HFOJif2p8EJG61ACB7hUwsSPKKAdo4YPGAczKewqAk4I0zGVO15mzLYlLYV5E
PwTlBoBnIPljETWaDV/JPTcepBpDz24BX+dlEBpN/05UAJ3Tz3dEf73+7i1hZQI4WXyZA+2/wrvc
c2e/bCpNiGoRBNs95ih+YocpGzKchBW67avNqXzr9SprlMBeTVHnmXoBcHDaQ0JNbN79VPwDv4Y5
6bkL+/KBZs2+cPX5IUpmyV5d8Pd/NfyRdtrVOy91Fd5vTLyGjWLHthLDU096YYgPalBh5CqM4HEF
T2/3pNgGngmYNF2guEKInZQ0/MxqwT3G0T+JRK83sZAAE7VM9THz87IJMRqMIniyvowKwlI0DfMI
F0jlj07PKRcZeUGcYlnKekgWb1icozlD3qfKFfFf8sEvtgNXtj809qnxhr/oL/B9hsivo3o0feQC
MzVGuN4NVqJ6ls43VFv5dNYVlMFmi8L6JX1SC8HgDpV+lqS1peU36oFnfBGJn9UN6gcG8165+QlG
FZK/NZCfegfCfzf7Yi2Md0CXPn3eY+VbBaL81B6BtHQAoPeHFjo2fT+A5oNJZ/oUv9jc32VyDNHb
mBH7JJWkOyrxqZFbegR1jkrx4lBC0z/axmjCzuNOSevT6bMd07uNCtMYavxL5mwBJW7/8LqGPxoi
EIj3/nmww25pzOMKTB3umad1HHTLe5gHevI2fREHzwinlIm9PszEqXoxC50KVb4d0d5V4OzqbDl4
jlhHOsLgssysDvXNKGrb9rYmE49i0amDvDdaMpzHZQtINgTFBR59YSdPZd38UdNRpcis9IcKYPXq
Ps0JdOSnHKWuQF4/yaO7U5r+8VCUdMe438zRh955CZYWRj/K9OrYhIhCo6pM2rmOhCkcdQrRZ5+o
KYl+hQFyQTaw9IAmlQ9YDkD66uw9UTrddmEWQFmlYnN2axbtzIYOtT37UNYDGS8coCdEECGUzYTd
XzDKT8PBSZGO/v/AB7CV2ntVHo8q8dqW9SlDYNJRkjUiS+45ziUhbV2NSQs4K7qAKqb+nl+T0Oag
9RjezRICxS1lIIuTE1RckjQnYsetLnZjgLoryMH1Hel0R13XrL8+0ubYYbj3ZV3h5qQRRJmOHdP9
aKvydid7eEOZRnsSMbeVzuzfi4xtjVMf6fBFs4o5xbuLI4EZNFktm2hGoHq35VZKWIgeWWYqk411
n3u5PAK4sOrFE2Pq8uX9OgjZhCcNeWz8IwTl2+UxqVrghO+K+gJucFvlT7p3/T+B/HC3fzi3a+qU
q0OdxbamcQrQmFaLUpDWBPug6WoOqgHUI2rDq3v/3ZpuMhkz9RprfpUnniC2goket8G/cSy8recg
C9tBwSc9GAOvzD4FpZo0nuJSK5yvUYKU7FwxLpRVbrh6EcUsBVwctnU3oeG+lLxLMH0Xsk8rhNVe
i0/lY2ccUOp/zC1KsH3uOM736zfuq5QuYj9V/Uep0Uu9NFhrqnx0lgK8YRx8Rg4eLI4hgREF+G2S
QsxYcrSQDIsVE1mhi2rCOMKdZvplp+pMZQr7jIAMlK2IZgnaoJzqqscvkzOihZ2r+wFzhFfAdC3N
Ys9jaa5ChUbh01kwvnJpL0DdZnbnVngweB0fha6Q/diU8jeWb6tP78ODDq7Rokxf73X3GC8UKI7o
aNMl+X3OZJJdEwLGUIY+1SbH6n4K8CfiHx9dGwqKl7BTXU0VUDrLItbpftVjkGprC6ZEbIaQMfs4
NB8YrpnmmhDnyFpyUm8ZfNUDnwmLLLmLM8L4HzDJhG/LbJpNL2nykg8FEgrWknMMGeL90SrXh1hE
PUeONj2xUiafV34oqBvjfBKUghoxN9sxllu9gP1FN5zUSc8nZqEngFgSXDvgc1H27HJV/CQ5SNJt
OjXambTJDLwBh053GXfGJLOpJ1mXQR/b/KLgvJb3vudkp2i9/+aO+EiMWmMK0tqpVLZRTUxe0qKh
9YmsvVT7N2t/wyozxGpkU1bkGnhCuvRCRto7XbbNjxmLU20AKncS1eeFZOZOHszW+uZduxRmK8tj
WgZQTYhxJ1Ntil2uqsJpHnx7a6U8lMNId4FRzsk6t1zGsa5uyAifWTJcTLFb2TRXmdgKKBrZ2FvL
fkeLOD9QqoIWzu4KKv2AV7LypuIxSboePOMI8tlDTvsZhY6tUXJCaNbRlrtcGYIyerDs5WfIUEn6
C94eE/v/I+sW5HD/Qr/DBiED+2aDRuAxwZjYauZr0SXUSgmPXkNR76qEZB7vsy1vVShELTZe5Fd1
OezgVV37rSo/Tb6seFDupZJDj5wtn3Kgj3+oKuVtSWvWYURxmNj9QkhnY24Nlqs3STMaChXK9RIg
FN6nSzMXXmaEYLaT39T2pwjQTVfk4cWcocLNNAsCACJDZyCGrw/rJXhxkvTmTFjx/uGRUlEanOv6
DJZueeWzagoGGDAx7ZRHU6dVHYdiqfjJAE9qMn0brMWu7lot4KciP42+cFjPKqqdHTq4R2ktyQBO
vBY4CwhypOG+eIQmzr0a3q8cQdomwI8hOgmSBU4rPgVfatQjrRgkbUwDzBlZs1YSX07u5Gc5PnGP
QMq0cKM7CXdEob66dGTIsDYNzQZrgf1ci5Qr5Gt+w8hxpfk2soToWDB44iPmCzDvMSojP0cAFMYR
xfoSY3u7J2uqhvr2LgHoZFs22NHXnvnekjy5bwX1FQFWxV3csG6lQFEj0v+fqQG+m9OI6VUbmHf1
V5Q/fz3Rv4TTQUd9uO0dv32/Q7kbp5MbwikJOOIxxG1D0/TL2N44UZ/qU7ZSbvPJ24LTdIoKtdrK
l6ebKd+njtakgHTh9HhdHBPDPP90h49oNqb9B0im/7Y59g1y14GkpPuT4SwPkM4EmUzf2IgLlnDL
Pb25A7RxdTZIM0j6Bc69EP4pBfUUMv5468BiQP+0qfSHVGLwjyz8VSxitiNOltzUYYkIg9KzlTkm
GDrvk0jP7WKqAD7L1Xwy62t1t5P5jelG+kjPSK3drSGUgH8J8n93ttl+r7yxDXePF2+JliNdEwTz
cuknN+UhOuQUaksmdhazv5mDTXcORML/7RHf9xp1XgLWYrtzuveDqWDEf0Os9O9UIm8fLGllSlpM
3EkNIPed9ivs9ZCMmI/QpV/LC6T1sg8L9K8aiE+E5kVOc1ZCEHykEjhu/LU6E7H0AKIUEXHwr3he
o2PEBH6u8wG2XXPM+EE1baoMPCtMEU4Psb4NRZsiJoCIVRRM5wwnLOl5NhJz8Eut2r3hPlMOOaVe
AC8zaRRbyxvTZRnHqmzQ01wKzDcpngQa9oJ2oSstWnJW31Nxss+pTWmMziShPGp6IzbNzPHHO1YI
7t6xm6sKTV+IUIe8Ltthz6Oo5RjzOIEP45LUhoDGc83A5yYj9YgBojjez59I2fiu0ZYBERFS0Jvq
XOQoggLxDwQTuHsHhGGmB1U7g2EMUTsv+ZLJr8SVtylMV8xrGsthNyZA9bYGGdHfIK7bTdTVLLxr
MfzzIUix2j8jRLw9dUWNh0buJ/myLndI0Iuq7NjYWaT+wBwfJveHBqrJWzYl2UM+GNTViOfI1mqx
QRFY90VV/mnfeFaJ7c9W+T9ub8Rxxq2uFTeUgg4CIsp/GHS6oPFbmMXaw/mXTnIM3rlbbNf4a+Dc
09xOFqQ/zjTh/uQluUvJk//8el2kX3GlLi7KJFRKQJ91EvkDNo5Ld8tPx43UYsxvhQRXYi2vgDs4
3pUFCWywLrvNKEdddPRLomnSd4m3RenE23C8oiNmrspR7Al8NJ25I040jA/drMxJTqgL/mNLhwcZ
7jH2oNgbM5YSZ91TQvYpx696qSEtx89r6Ul09V1Kz8vkgUIiXtZ78M2dAbCLhkUKQR4nnx1PunY/
0EswcTXPoVK6u+PtjXnJERyAcwYZZKrEFIcug8jOQbadUJoTHEIEcf12lQcPcq4a/HqfyCEsfPSj
SDyRQgq1X+Cs/R72hNeG5+wA38HJxMqPYo0pPLiSsSWoJRNylHzGdvIiDqwKlZGcfSYh+3DrCX7k
OwOJd8qh3aL+3QaSv9cfOKrJxm5Ph47QQNBLliYCPSmk+MXlv0PpCxe61L/6jOouxW8766QOHaUv
3Jt6V3wdUAaOzzvAIXL60GOEOnwuwffWN36jt9MNxT4Bdiv99Cd3JmZ5+jbk1XkWIpYNMXC+T5fG
ZypudhbMyGuWHQUm8qXKpFfYHMLAyfBVFhib+R/sIsO2B13A8f2FQ9PJtmjaYqEIn3PZA8Q3eH8N
2/ua1/7MaesviU3d6IvjxqQ9bMUHSx/gJ58UFKwxN9AhAp01cjIUSeKD+/CgpSnZZVyEPIgZIWtj
lxWUQDEdk7LNozHDaXXoGfGjtNwiGtmI7Q94oausMV0rvMukE38++AAICfPpbcxkdfaMh91U2Jx8
snoeX2HVjDTvj+TMFyMgC7vvaklKRRqaK1LiydFUsoYDNf9cQFHT9ajaEn0pQ9nSvnFC1gr4CgXT
EcqwKKSh2m6TLNYBGXFEaCTqKfoAZJgacuOd/a7AZvr+ABs5DkL0xIxpCutc1fG1TL8qQQ6/QhGm
wvbR/Dw5fpi1yTNMW+0e1pJ7IC33gP9k4/X4RQUFQ2TaVqEe1P3Oyz9Jba8fHjBd7MFa2XhOCuap
BQZcGjxke5NkfqU1LEgMEHoXZU3nQ+N+zeoCTYCHW/y+KP+FYEG6lEmAGEqjMAiTj5MmRT7h2pFp
BsJS6JoUxNA2wWNnBmTXc2M1+rhcUjc/njRQPvZ7vgfZVN9qwUm4CEQ0qg9Zos6N3Qv70s6mXPoE
OPsRfIhl27+QhIeykM1C+6NjhXxT7TjeBBWvP7S9xgV18UVtORMbUP1GNr+2Fx6PK2Ii0mMcxtHj
jMIOxMvaYqYcPlP3Gcm1qJ+dEL5nmMODcIcK3r8wYv4lhW4Aq9e+w5JPutEuTC5yPcU2YcD1yfNh
9T9saIfb66hKknJI3VQ2yABoxTxKleQb2z7Gy05Yl1QNiI34td6k/1OzxxeYlAdVYpJklGpTvogp
XTNXjzZ8KPRtIr4lGhz/8KLThHRleVpqPQP5bWytoNlk8TBb27TwfHEXp6XQtQ/tzi+pWRgGRYXc
Z2y/5F4bVx0oM/cfGhPW3y9b+iy2B4F4CeDRr8A+Pa1o87QwVvezDUILNBsSliMfkrd4p6ZIxET9
NWjqUlE4r0HHxuyDbQzeRaAei4xR3SKriDCGScc2PyDRuNRMEe4l9J5QpNmd5/VQL8UZfh0rBSg4
grM+j2j0nZYIcX+da8jP9P8Ue0BDFu7rHVvoN320zhyxhhNDLKE8smIhTd/xOHoHQFIlvOO3deTH
GNCJ+xTrtM4+oRY9r21+PVT+lWYJB1I2GgYM/BTxYfVTym2VATAdV8odrMyKJ2HIcCnCVdsGLg2v
xj6t8+NMSm+5joHaJZdG92qwZQnPJDCMYOOt+yg0RipJEz8qPhy4GJHQ+Qemy3WUGiIl1ytIp+o8
HO7djoihaEboV5TApdwJBPNZRs+4Fvu1zitJSNGWyiflkT2/cf84J1eDWYhL/L43mkGU6OgHJeln
SRsaPIvjZq7sP61Xzlaa3zYxy1tkgOS7XJCRjx1US9XN/Bgafu5L6RxzuYfnogdIRUuQGKs5Tho+
oU/IrqjcyjgSANBUQIplpJ+T/udXby+p+d8eQGMEnKZcKSYRBQhUpDFXBZfgeLmkir+ggqiBqh11
ouHiQ3ZzLHpErOjIhXy2it26IkROqYPoUYR/P01OLtK9DKfI5vfDxuR/iTUCu/Ovcsu/6WAusr+G
FStlFLHeJMPTr4VZXjArI7bqBDCdHtAT8oX+XS397HuWL365UfVq+XriLdBeyX1OPIW1Xg7Vobm9
aDJMNsrATNC1/YLYStjrjkNgnpDkp/baPVXNEy1683xI0kQBs7D9lWBvAOro5kyS/AU5PNNent1D
/sqTIUzEqOjuLAvN57goVMvHHaQ6pH5G7C8qxRl4ObFoTHLipEDTBRuat7vdAZlZwxEs5AgTfem7
e/fQHlIu8R6TcI1URibjXwXhybYtMCJyw8h5Z1Bacnbyn958aPFkVJeyPBsYQL9M9ny/qw0p/Cx3
ywPGAjoLVF4SbnEMKm3x4EMQgnBeMJXBCvghd+YJUSBkf7Dtwd3vcO2jlP7FgEwvZUakeXjtK+f1
gBwAAjhZGD2mh9U5hIfInkNkUff6BvFMYohBq2tTYgyhyx1G5+oYuwwBw+1Aa07Z2TAg89AS6o3m
Nt4tX9y9nZQ5xaWnhHC60N9MzIIEdPW3LyY/QePFXXPemvkCUQJYRgYe+gcjy7ANvz3ZTI3FUeD5
WUYzqDSW347ePkVanZssGIiF1hmUzLZk6etC/6DC0yBwKpf0jyDn6/8JO/7LZPSR4iTkKO/VdkyY
3S/89fg+Wz+HTyJhAS+9KB9H2AV6CBHrKxv2Ct19yW98iIFtE9PtHH4qY0uMeE0SCG9S41Eh8qZg
53FaUtROo75bdQsyLARNHCJO8/VuSZuDN1eZhJd9/uN+PFWXuORVz6obID+FxWwKfMSxThrFaMYz
ggpq0caPXHwOVTYghhXrKOFMIEW+ZZCtoLeQDQN12hqymG3B+9xG7JGSLl05ujR9tCEE12n7ddWh
XMh5mSM92WbWSNclGxWU94mX/ef7yAQfr/D/8IpQNq1nS7vbdkPF49F3kPrUdJmY/P/xnNHrdFaE
RJ1uDhO6ZrrvI8dvWwGLFK6BcMJRpTXHg3b+z0rZQ8yqM1RhZ5EwXwQ8wPe22pcnm5+gpwMgEtc4
FitfP5PT1bibqGUVVKhvyefZnlu0m0mwWo6i+sb9QcDFxkQJbrLelCLLluWz62tymlwu6geCqakx
+Zh5WqkAyrgpqFOb7gkfG48pDYKfS31xWYRMqEL3nncUO68nazlj9PwMntlw10V+K+A/UOljv1cT
i4IebxLX30QG51VSWqqFn0YgPQPd0VJbPwp8gQMv7Ak0auMUp9+DG/wHwZlsI96JyAGfcmyDwPuD
NXY5r/isnrzq6kNUYI+tYD1oZRoomBoB4wnuu/zF9mpGw50iS5CB5cV1SNryyCBh84fRkg1xLXMe
nDHOZtRCOLcRKEZw37DnYgUITrFsOTs8Bv6QOhCNGCuE/NwrNn1wmjkLvTgFeQg2sMO1x9djIe0m
qyCpN3u70owHCM8uVUusZGR+bET2jPELv/EXPf+J038YjWeAfze3VTCYA3L4SQEwGlV0J9o7i7fZ
Uza8QaJLlCMxrdOZmUIsY7GDzL/0Pc1yvtrec8ocBSYuo7ekSK9lLOhWLGtuKPi+8Zd9G0OkEkhk
vRU5uYwOILjtYohtBpjKCGhGkABD7gLX+iFtKK5Pb2IUWCPLdry4bRI+rQDng1biuvNNO16dom2d
C3aztnl7LDx7KDynVmn6rIEIJ9g188LDR6R3jVwHgNQcR5N6Iqoeg3ZnIVmiuTjE640gEFWXC3+V
BMgp7RDrLdBcCFLgao5j1sZFq8tqPwvI4Uzds8RPeRRMx9POgZTbj7M0Zgv6WPkYgcxEMA1/lmMu
/wPlzqHTA1gIbeTYds2lxNUEvRIBywlaqd4UqHIE0eiERb2l+0KDaDk94R6ON3sJfuQD+92gABPk
XNsx/1QExzby+gTUeJC9n5cycUzj5gdHF1ZrtG/3iJKp+5WzpYUw7jjGJG3cmsfZBWUovWxdVg2V
sOBCCy1mKoMD5BenBEseA2+F0JWat33mKuwY9TGOTYuws876vEt2VnGFNWeB8engxQbYkjWAZyth
1f2qwuetUNAAw4AC7C+vuUNqn1SvQqdY6fgDsUlcBsU8uuVmuQ79C9OIrE2/It1R0UrTgdUNqOHS
kJTG2JaLm3w8eMimpAl6cdckKe2VvMPTtmRXbsXtNi0sjbp5AozAd9q2cIVzaJLfhMB+xIjyaZr3
oKAoN3ACVfatud7nhtKBH7KopAZyuWqMBLeeVJjqDuZj2WiOypgpa/qcWAhkfXyOjr6I8lh12YM5
MMvgFrVCOjEe6Iqs0SLTsEiPSydZygM76OlEv3FWwjZ9NTmbukT8gkeCBI57RU9qOSJJN6up5t6s
d9Sh2cM0qzRRQ5/AhNqnviTeRlUtcgRXQlkQApFIKqd7foPJmg3GN2D61QnwLqfy4g0307a5FAuh
1XqrGLbeoukL5tdnwmaitXG/X7bNtEAp3MTFZXzXlHkbn2pS6nwjqZqktn0TL403GwOyzQOiVZuf
C/zSXWLEQFWuMy9AoM2eVqTi1Bc0zjIrP657UCz2LnmiqD9310Ff2t5jQ/gXRIS9fncGFFeExGFt
WwUd61l42K0+ClAwEwY8cMbm0jCiuBH4zkeMJ5usdGD+07dB7V7Vw3M/nm5aqqt19rZhtX+XUPkr
h1QiAso+lDz3SwbucnGT/nwpktHtMXirndbPhjLtN88XzQVFByT39CaDQ3TxktLCJ+qqq3epqZf9
OVgzobQSkn+kTC0xsGmHO1s+mEn1/lSymyh7ynObTcZYx7Qqta3yJgvl+fWfWdtktziiRiJh/Kjo
kWoQoJI604vUsnnSCJ8TzpEZsiLm9NMFODk8O0LeFPbfI0Z+E7IUKwOkwt3kqYSwnHl5I25do2PK
kdB2xqkNwvjW0Isc1IuvJUA4r8RNrdfshm3KJZz/BHvhNhJSbST86H9pW0xgEeTOYBt3VYSknae7
2OdFyLx1oD8SDVAf4WUkWGPjbIyg7sdr9H3itv833YfjCwAec37NPoPDwvDUhQL8Uhjul7oFG8ij
QMQDpjvE0bEygYWYG2JJOEePqthYxSPejbI3gLuQdflaoauwodr53VAZIUM6sAF3R02aRxpulyfJ
z48zmDl4k9ZSGo/aWIMo5LpOKLBF1sXfwRZoZ9mJ+pKrqWfF9j6hvlUU6NZFU9Qer+hDsskm2oNZ
LtIq0cP+M/llVqM4HziVUkDq70EXWRDUVtql2zuLueDNZqABGrHo77dbrLkK4efa2RW/yjHolKha
ypzNeOCmVJDMa5HpL+SVlcIiYTNbN9gcLoZqsyj+BfDd/q3/cPiGLmgjQIxUmUShEGlYNG4G12TM
+e8dCgCjTzKT7cFhpHAIqTes2zwCCO3Ew3LZlQerquhnuyBAF8C4Kq+9Bccro/xjAv3/C2D1HJZg
d+TYSTP7Bgi+SjK9MkBWmLAQVXimR3L+6s7H0bFsoXlsIerzx9lQtSg/miRg4g3NVQZ0HdYWxLLW
wv2+TY9Ouz0OffnUQkBa/mE7GAT3XGejpHUUJMR8fAQEnL2cqbZzesrFBBOJyPFM1lFc0xlIyXvC
dNm6jF8sM0+JE7cOT6Opaxc3kCLY4OVu72KrB6PDFRro622UHSTSHfxB70wx7yF2EuGZn+8kYt5p
dI1b5vN142ywNlFmMPZVsjnaycOJ8Vjm2VVWkDCoNxW60hJ87VSKskl/SX7xE0vfDL/2bSi++gKf
tzkoELbuaBHGCUgo+qSXqyJKlWyo0+jgWi9GkSBuHOe6OWLcChIw3b6N9nE7UqLg+nXmUtxw3x4o
/hYzaRcHuk1+P1KQIjlnMNz+Ogb0NckO1CLDTuwLeGPL6/fM/b7XCIIgI4d6nhNmmVPR8aeUQhNP
WZWQ2krTNSkiw+WnKc7mrkHo41FPo1UeXyxmOucbf/kJWk5/OoP8oc9hJmAgm4Aibq6YFNEeh5sO
UWfzsz+XfRTh+cLHmeKBqMueZeIeFjHiyrjif1GcBp1FiE/0bN0mRwO39RdY+O0IgFQXFb8yBX1Q
h7dv/zBpDqSJkb5veEYEHgHdEWhCh22ZuyCu+rHLkv9tiXrFTxwG1YrxdAqXekkbMuMBx3myz/4z
LFNk/OLEUgx5FqU0ESStq8tlG8aO2eg0RWL9vQyDtGkzdG5b2Y8w/m9nm5Cz40UuZmTqLzoe0kDk
vs9AxUmip0jeg3csgeNRFO0uuhTmmw2ywVlKhyv9h/p2KHNHaxvoZtiMQyBJQqnHDh8ktdrCy7Bp
zwMBXHhHWPItlCVtGmKlOrwniUI1q0bGAymcS3B6HOABMiwUpAXh496Xsfyc211Tdv/pLVP5U0jr
84jMfrFhz7DRvcyNNbOQr24nTWg51n4hJPozMX5cWPMG7ZHBqwDGFPA1BTAkSu0+rVj/pqULpqvk
+L45+gAdvKfwx5u4U+DvGmrFEI68QyrIllIJvITZyb793S14kfd+wDwfv00v/pGTeXtQ9kz79TNl
HVmsvkZPPrGkBaloDHKwW8ZT8RyPJy/DVzqwSw2Q265C6EN7c6zO6sH6wtm1oHTCplRAKrzBTfNu
TmwtE3+k+NzQM8jJm/81dKPnpgk4etizLK0Fw8IdQLacdMF1gJ+SSTn3QNsPrP9K2ER3CmqvVh14
/4mIoW4e/eoJIIYIiJqejzhxiMCh9yHIju3YHqfWijL/nsAhG3KRwxdE047u8MZbueR5xeWyNMnW
MeOec09gPR78HBiDhMGPpYpJrSMkdMdooKC71wWw1MHmXwPwvl1+srmg0frzuZ/whMD4reBPiq7d
GSX+V/LfwE9n+Gud/6otz6ZFqzxzmtowlS5L8P+y+Pep3+P5tbCNF79vOvNr+Fv9eQGwD6qeLWGI
YeP464WAQmSP8jxlAi87Frz4NTot/GwNA0ydQm5qupobU6ZMIHZujMZjzSdHWvgVt3lEddeWm5oZ
Zjm1FBXakUOAwN/WF9sTVtYs5QOEBI0KRC26jhXdq2d4lbVrvKmz3LGpursDa/tHN96tj1+L1681
vMypk6CPaV7L0D8sqXwi29JTbkb0yZOTPAsQ4M6mwmSWkw4HPhvHbZQx4FgHk50LSuLO9VFwoC3j
sqAxd2mxJk2zoxSH50drWTCsaXDL1pw4nBEatkMo/1nsIxew7O0hlnVtI1NfKT7X6ICd1Gc93mQc
rGbGtPFSAVTyNiK60s1jghHCg2++X5kX+yYpxgN5rLjd/7NvDBC0WKsu2CuwxhTHQyBYHQdI3x+t
ngu4HvuIu+i0hQuXBmE2BK9b8CEPLrc2qx+y2/GBiTNQ5FjKEJWFcVQ9hzClAkkN6TFucZ9RjgmT
YGYZ2KnqmOu7V7dBuf3ehQV0wUU3SgE4mYPyfYLYOLuz+hx2U0bL0Ar/mHemvRA/zH06BCHZS4ua
qyjO9QonUH7wtiIdOYu1iBDuIji3OLByT8by2KSPENr42BuFjSDObCgbWgNDC96GyAE9exmWSDvv
1c9+QXdybr2qskkhSKMEGfnPa+CN2/57RBqpoaQqixeSIYFljIcmePOj/m2xvM57IX4YKX+GOLfW
oyJnRoFvYCCJqKJBJa6pqX5RWK3NWs3iq6SmZYwe1zg+QG4fMOMncZ58wpu4TrY8jmzy7pYI6I5B
RRlMNRkaRjNWlsJ05nF5ZCdIEVG3k9iCNuApZfu/FmTTRQ6u8M6EJranxPk3XUvlzkfm+iItP1Qm
76vav4612DdFOKkUT1pAZU9SaUjc0omXc/GY0a5vQW3g+wx2E2VFy4o0pK20kpHZSTJ2caSeCU2S
n+PHzQHAqQObHsFKCIL5P6KVqXZuPEm0LvBkGZ7XhS/A6XjyZiQoLcOfK3Z9DpM8yt4rRdJaTwtk
6u5+eCYteWt250ZOzvRMwKtJlLuUJLpmVTzh8ZblN8MTZoZaapvDpRxXBAW5jkmSVPhcWepNqise
9dB89Ttx9RmIT5Vgjuyac5xoNIvUMK1IGWwGRWKYxs2cP86CGvujU3kKacKtxd2SYgCeMVQBRfAX
YcuJ0uGekJvUryprKEKHomif3zi1+6bx8rx+u6mslqO8xJUGxEoRtUGMphMzo0qQ2dY15uIS4Hm1
0TpEwF36XXhCzFX2kFVkwcFbpfdurl5e1mVsd/nCWLsHFtB44a/J6a3FDeWkg9onewNEYtSrpau8
0jkeb3A9Q1BTeoxqgJWmrB13abnsRrQvn3xMvkGDJ9FUUXjkHVH9RCIsr3gC+ILWubbgyifGM89I
EKq/8qTAecxeIt8afJR0EZcW7CFXgg5UUWgazb9jCnb047dn6PGsyCi3nvfAmykoNFZIoIuaC+Cq
7WWR09eVYXrC4nFYw/fxF1RYMRXASxBF7UH1K3yGRgAOFjCBxqksJoGnacb4ZTItDAvW3QGh9qd6
SNbAmUH+IOvp/MDRRgG3PaXEINiAgz1obclq//yG/EOEfOOnwmZPaasixUKiIcrkOyItx2K+M9eg
o9LvaQc8LFrPYY7GgAN38Ced5YH8K7JzRbVLSuGKuH6am1B7st7czSwwrB6eSTahxfxJkDilUT/w
5ML/mw5quhOkoG1LMsgl4TWe/Jv59ymrin31vDMrRtLCTQBLc/TYxOTQgTB7ccrbKoJdp5JLjTqe
UXsZ/3J/6hBlu5igzS+QdT2KGsvingDkzWKrL3t1bza/13miSRLxYN6ueLz036u96UW98WUPdL4F
i5LH2g7arTGD/Bn5VBX9jLO1lgg2SRNpZQCwdXDXqOwHp7MIGr9ioWKdenTRph+X3SGUh7YWudxV
tfBwy917cWPujnRWuSfWFCvTkyt1Sa7ja1MDG0CzEj5rAXY2VP/VZe9YvV83xsy/MbAgVYoweAE2
6acN2YjEQF0X1ZiuRpDCyXqmA0xUYgALGGg3oapLzStMJ1OBSmRRljz6X+2kKpZ+6vRXmPhZMmZe
gZEeQwV2dCp3qatd/8u7FbNXmMQy2Jj+8BEZO/X8LYEx2NS5InVUiEJ0MsNveLFIcaIvH3/pBlSy
KU3uRs0W+n473Ry0Q07BbWnavw/mVxN7OH14wwJtkTFFwZ6QM71PJHyQOtP+RHS20pBlIjVoIsue
v9Jhz5vgUjZVNFPyui2hkaOXBku/nysFZU7Y7U7Zo4kP0xrC+c1NNOwqsyKZ22D7ab4Cpu2+MTiI
uhzevo26A3A7IVNiaL+mE8akD2jTou1dFzDGbJoFnCimmuCTf/dOZwf4DnQeaK1n9BHZrZStBZPf
XzbZFPCQA+2HwRS4AC9yPAPlrnjaw8gj8Y+6oP0qYlkQMD9gwDzF/E/w8NhziBbYnoXbB+jZP3RC
wMk8Nu+so9y5pAlLIIKjChI8zKchjPS3PnFDOa1EtHCjBJ55MplfhvRW0HAFEQ+6LPEEr+LYnlXN
mfbPnMHGEEKdY9Cb6rkkCeIZ8JbM+MMAeo38R5ioCa9/QUjvmbAkSofIAnUGpPXoAQmF7XkiJoL5
KY+RNaT1bGkyFz8viUD0wa43aRrvb9wvkrY780kIah0cZDy9sKFXNdTaFs/KQVubqGELgglRFqF7
TuywUygf7/zqvJZ5SaTyie90x8ZEvr9hCKo4DPIKmUsfHIuXko4KSAg0cCsXKhLVxM9ZfTO9gOj8
1awwmzNMs0V8mHXAL75+ZURchwjI0XFwPQWy7KPBWEXlxhp4k68SW8WPeUwqer+X2s3omqcyLpmv
G0HwJUnpLDLcfaz71nskXUYukyRfUebV0kxNvyBG/nwq3jgVKbV4Q250aycLSW5XILNOiRVXiNr/
eiSVQb/XEpSYL8cQWXgtcjLlFAn0aB73dO/hgforppD5UGNqnF10nVGrURYgvhO4XqtCgVHh+B+3
1CAash1gvNAnSIWWGJMvoeuxf96drOvgHfMct5OUfStXHHK7X5gPFMGqbvjJmjufo80btIiZgQB8
317TS2SPYZCd06mXChVs9X8BJ8Av3p2KiM1mEGaPclMP/vFER3386vr8voe/+hQo/mwIFhS3PPNv
Q1tHMD9Rl3fOYUmB5WJnpbA1kJkgDopKVyr4KsNYD1pnd3Luh6seHdTGStWQnz/oA+OXtHpV0yKV
hebNW8oQX+7bp8FwvZ7Ky6mYyz024G139PRc/NPplHfmXMipPm65HxyCmB7BmWSbEVFYhQeEM4Ts
T1ES67yL4eUFobUga6ReDNuBXL/21QeQAnv+eNUK4srZRU3+exX01ZY0q0FGphjpx3c+2KFP8+LW
QhMf6e5sRBwc6jDFHYME9ATlQf9A8Nk3jycAMq5oztPhfsX2qyDAKJM+R1ubx0nnqTXh+4i4rIr6
SE7iUoIz6/Isb+fpvQWU/NryxjvoFTNN1dlAZW3kap+U4utsRpojGd1X2HuTvXgwifll+m294dN4
T7G2gyu7YVsNLSeqfQYNw1FpUcHdQz/6et0Lzb0Z6Fe90ZN5aDW6vjygfiCEM9vmPQWN5N9d+JHn
zyga4uQNYPLNEnSANDHRk04C1r/VvdTzJOQTF3ZKvFf3kJ76kldBruIctw1VrQQoHMkCHhDTpdY2
q77pASftQ0KND+KFdk1LK4A8YchNspAYYaKCCrxQnH5lHzFSc8yxlzkq+HwGiusCVyrmpnJRrg37
c0UAZDYjMyM8kjEljKsAsqmnLuXuvi5ohAQVUE9zUqSzPCGaUfdDFuZPVGOAmpws2R06V4Uvm2ta
uImHiBgcKspRxJ156J6vHWYyBw14oFxlyrzCYlqPFdUmJnC1OJDZBIHA+ygechZbx+4xnTwK+sWY
tVeZwOpFh1ZjjGi+xw0EoZXtlqaHhidX1sgNNtKNV7FTG8E1zkvSdkO0sG5fGVx3d7Jmh7ykSnr7
31A2xmHkFUeNd7oVrVrfDz4VjTu2C3O0vYgsk2vPjYPsxIVIh5nrjvlbtQIdiWJyP0ZxfTqDUHSk
Rf8AnxUSFpcq97oHDUDlyLfleF+9a1QKdqKq9/Qxe1XpnUr1zhpf/lbzpol5O0bFCo6+M83EjqNB
de3rX7+NuiuhjpnXn3BtUWDbzDdnOOP6y7SNz9AYIRVfrZnWpWV62BpBWrh3Si72TI8s0Qrkl1Dc
13lwQ+aUVkGqJ2CjMY+V2+xnNA0rO2D1j5gQ+Q1d0RvPf/KGNbP7/lWRF2IkpYQtEkGiI9uU82I1
SXrKDS43LvOkd7UBD8kTJToa1IAad18tpfH+K5FprZZ5WngH/vA1fcuIWpEJDnxmWjgj5z7Spu1o
wM8zzncqu3Jt6xSqTD+bAhr+xx3GZDtZnsJEfCECXv2gQAL+iEs14849hSB/+pu58hLRAOHHuoMB
qUZvaQ0/CkLOBsiSdNbuTcaIQm926NY+rtG63a0EIb3WqLUgRxNhtbSoIuo96QEtFp57gkmkyFJG
eWkty+bc4BzAr+Jz1aPrRDk1E1WRIZ9zjBHT+fqEvc8KA91de4HxWUQFdyK7pyXa4+dbYE1qOcWG
fbhE7dtuWQPr8N8atudyPj3bClBjTnUi1ME45Mmluh3+lpMbqqyvJUbaPt7vhUt7faPkgMd3BHNT
WL+PtDeR99X20WcI81iD06aFae7ccgj8I4hiI56+h//Jb+7UMgBeGjtGmif/fTsQ/mK1pzB/XD5B
5/ms8IE1K6foeweAZJ0AhRWmwDqECyM49KA2jQPTpceUvUvCbItLcmu2iDHSWaHppcsEqOBBMfys
ETzyYQeEOlHRQwFUBqZqn+9JsyTab66V7H1ZrLdJJQmjgJTJCUn4QSKoLLGX/ZhOcQjmuN2z9RQo
esHoEzO7pvtYKvBc9vqC4FapK/pvbXI0awZbsCdf5LlhWKqTJLV3ZaC7RhTwkVW2PbeQQMU3y9lZ
Fk34SEkXJzgNqO0GdxsNPw5OdY/St8I3JvX8feg9eQGFYi98/gA0g312juo4W2B40/YQa3TiRsW9
Rv+5G3GM1y+6oHGNm2PeofNkHBMye5zgcZS4qFoKN94b+Zt8ub7DZz6kGvzFTqGXDHVmtADRlZQK
zSFB0XyNH60xOogHFi1j35zIsacRBHuwRxptUsp2wxp1eLUmPQNBw3ig3QCYy4VdtKo+npz6B2j1
PVkB9aSw2eoF8u3n+HLnL9swHkWU2ijPZeFrRbwHVFzSN03KHil4zcmNyBijsbRgJpJ+ToG5zFJc
vscjoU+irXJ/Q3y2ESuVEOQsN7KCcDHtmDoy7ck3ekveYxf53NfyhtBomcZzyn9kednVVIoLQ/XL
vVz7RL4o41mkL0rYQcpE20mCbnzytSCjrWO73DHYDAlU4yfXHb5COnwTw9U3vqQJcMmLuWlNueZk
af82KYyeb6V5sSLL9871iUXQo+D8d15bADRUYZp4QFHHJ9sBVoNNqIOM0NGx0oARt1M4AKgnWKBi
IgT+3bkgp2c3tQXPlOEzf7YXNIiR1V77ee/7sWHBd4KWedPurBlWoZUbYtIQ3HXAUW7BuDXcrYxv
MDiDgiTe5+e1uayEYgop/Xvs51KW2N9qePJ1pZLHOMDO2op6Z+x2aoUgH/JnvAWP72QLqW+JE64w
j2QKmL7N7/rGtLSV+XSmq8Ns2tZ0/w3vN45iQtTCGOPB0i3IMjiIjmIcl4JS3C8rBREaVW8dNYcD
JdNB6jeCQvdvYmh6+5aS/mtgOSyk6r4x/TScIb/di7m67xnIibW5G610hXXRNJcQ8p86f2zPiCSw
Kmp8Z5fQNrbcUGbN2OOaD1p19yXfk0hpZyQXCnKyFOa8zZq/Cc4n8EZvoY1jDiEnli29tD18JbEt
n0/ETXPAuy6vs4gAM9eL0g/pwX1l1clYDIVvfwkYaGI4yOZbq3CFrHLV0mRR13B8XYrmF2PrwyeG
vX6uSa7bmWcG3Q2L5RDtzQOhSFUoKW+v1IEAS5Ef5byfcryvBkpkctG5vj/P4ZXg/Yr3LHmpTmPD
H1Sm86vqJwMZUJNYx7LJD1tR38MnE0Us8rjHomXEbjrCF33tJCWGRngedYIZo6pHurs1/2gtT7Z8
lif0+eWFRgfckCB25+YmwEBPEALhZet0tXKEkBdTfsEO8eTeO/NSk6qAVHVO3iDi/xreWi7T1NNs
23zO1MBspYizUR6rUis5O4/APpc6gspIKSYYZ9xXT9AFLwrzXDoy8aYo7kzFzdIH/qVUyo0HTjIP
BClyE5Cd3vl8nMAs9Z5upht1vUWO+dxZGUsptsSxQc2HABUO9wrC97WqTZ0RZZoc9L9trP6ZTPpq
0NIB9VOAdnkDW2uuFCR06u9IMq360ApbdwAjTxlbAjVPdXWl6JyrT5KpmhxtJs99yblwXxid/qh7
jNyUxLtr6zezlHcCCy/N730MiDPEgb8bSTmQ6vQ1VH2qroxBC76B6PWsUnI4pxDCTKTEH4PYih0P
RWJ9A9f25iLHQW2vZ8oXJqHGuCZ24cX48+60s1IrKE8ISqljtYV99qeEut6pBOwa0Rw0/Z2EScmY
HE4CAXvL/dy8LgrydmnGmfXR6MK6tycISR3WJwHa3Gxi/3gQFZ461pGMy7Be4LRjrTioVdvr6c5K
8elQnQ00MUJB2tFaQDEU5kMR64g+GnMpUzS1H1NkohQQSHMcGtC2eCNz8oZVXXSqbSZuUVsby1ZV
RhiArMu+lpyCUPbOwxPvGg6VfOJDsut41JYLc45gy+Bscc2Y8ngxq8kX1YSXoClAihyGpKsdXZDW
n9z6Fo1GcN6lFZ+dbhpnoRfJHaqjpIhJcKMLL0IfPx6M7Z5kOvYv8SlzpNRXUq08Mfr6Dgqte3zN
ECaO2JCl8mhlkj7T7YdoAytBrMtkwkfTY6RUske3t+u/1c8jEZwO1V6fmi0hudvuyJC1eiHnF9at
Fc+jje8Puxpu35IjYbD6qfW7K+hXtXe0uC16ky5mSThfxA/QH0qLGuKzpnz+h+L97QrCfAoNIsrg
Vp12xUWKL0MLJNyzhq4NPorrGhKKAuQHOBZQP6p6fklm+scZrvOsqkjhBx285TXnj1mlNYBTuh6t
02XKYjjFgtNfgcylqkVyeJekDB1mnmDSKLNoUPQRhDx4lVaz42O77Z0duiXTiF9gUAdVtY01rL0d
KfBRB/U3HHpUyJ9EH0HtZH+HdOWup9XsoegO7JLWiMqrEi10mYEOXziVZtYasnlxC6tGNzLTCbut
ceLLcb8HrL4kEYsF4QCyWF0NZo2aHbjv40uKQKC+T6pd1TRluoPKN5in1cPFdSQqcTaK9thMBvgz
38CtOSbxJkYEpnwQt2/SzS6s6zAcWw+Y/GC7EPaJKxZ0UN9h3WE0Zz0nzTxjqdO9u3CGIzyieSgk
dAhDFjkgYj5nIvTR2eq6fk5LSsov6LsLvlCiqJVyR0o8NwVTPooWtkCy9uvSlw3qY/XrrcvqMlMH
MUIJ+6BQYO1a7JQsl6MXW5iu7FAIGAhomHDMkII8JfIvwcrWf+aF1ER9IFdphblSutpJ4wKA1zFG
RmuYHZ6Vee+7bb4naNgqrMTgl1eX5AJNZLLywvZDCA7Ut6BmTxhY99+gExDr5qSsQWjl6syUwLqh
x6+H4lR9vySd5mdkDLMNRZRrDgIf/I8rT+LmyHg5F5xmR9BTaaJp27oQyZ25lI70ZvWOA0AI4eJ0
moXIFcBMC5nhIY5v62Z/r5TGliLL3y/HmLoVCn/pVocO9iPbOo+WETwPAe4kq4uElDVxHQOBUFYi
n4Q1T9wgdYQ3szyWtfhETM4lJ8T8h6CJeVZ8Hh5cWb22YOC7z4dgDW/F+fUCtVpgveuiNyCtS8kB
ZTD56sC2XmAw9arPwwTjagFeBayDNEOi961dSlfSTwpBKEbyfbn8DRG7kaSjsMbehJCIfwURfFvl
BKrDo4uiNoSNLsUW7GYXRiTFgfPJKeIisZgPeP2E4y3aIr+irLEGz7IaAVfODQoVOPGfhzk1YHuN
6o0m5dt+fzbLS57T348nZ5Tpkfv1AGI55IG0w1XWXEynj6lB3bcfQnuIfMjmN2TbWbuXeCrnknuO
KNuKSBIUGPDcFslssqKvSAvQwbuDVvDOYIeoov/KvJ3DMxWGQy+8xDCIiG7ObfCxEFzRWUTdkiTf
1is1tiNs5j6ND+FlVBgjfbkOfuJeWJjisAYxGSLAyc2E/3E2md79i12bt2KVQfYz297BcdVrZIkX
n9aJvgs3IQfuDVkagBDtGEgnvvC1ujrd5kuJPAhGb6pTmE0jJEZpjYgq60ADDgSDLFqJfIiusXP9
SCLkjA8ZtT3hrQO6DUuj6ieLG7nRt2+dGhYgDGaaDV8Nkp6urTgQkjyrRA8QPHgPK7sX5vfy4m0u
UCN20SU9zOAddpXBLclkDsiS7pXTz06s3mnuI4AN6iTYOmWdTsl/aSFcy1fDnDH2kIG1E++YzvTY
im9X+QkZ9nZW21FtNX4d9TEA1w4P3F7YMOB4JmigwqbOg39VOSEQ/SnXi22Ue5j+FugMZLLL5RCY
vYr6Qxx1X7M5WzWfogG0ajBI3Me/Zrr4j1ukudfe7rzmsQIV0MHDNL9h5T7GWYG3rNIDRMbJuHS7
afwIe7Taj2osE7y/9chxPVPF+7c/KVnyIsiO6bTLQF+egvKIgyHpfzM7YoPIIfvLvwKqPCCoHpWZ
IBRmV7JeyLTXVNzmOlzUU6pPBiPArlE5vvwT5m4W6NG9RxON1bw9MrZNYecAt7l23JsJ2JTqndQc
uHD9udcETxyANfILLfe2KpNBs54B8WA8ADhbMzpwkNxkAuFUNk95KGtFsDrv3V8r3ZFovMABbiGU
smBeb77E8CO1LmcdqW6M3Np9ACNGe5JIYFnITWDwNP+MukwOBl8j1zYuxIyaH7hJMLgsbKPrg5E8
Jnfp7Toga4g8Svsuuvh9Y4MjDEqcpyNwk2YblqBkgDmFk1u8rET5ZEvIxmtRTrZkGI0oaAioYesg
xL3bEwe9GoNFxphk3CUIY3iOOPTXfx/lgwCIM/1Qw1krrPu/zqsl2BZv9JAkrWC8gYVpiLAbBgql
O6ssb3RSswN6w+6FLsTj0cu1kB7two22GjKD2z/fUKdyq5u5JueprZAbNG615aSuCwJfQ9wyVSDB
zxlxlRIdKEeQk7Xg4JAj9n2a7CdYjnf/ARXOaZyBtXA10+5rwS7oirtr0yvKIBkr/KvYNIgVt2Rz
1Z1Ktd3hZUOWVk0ZiD/MPG82EZClnTzEk9mfGDGV1RYAPDZ48htQo0jrbyOdvfuYt6ABMHX9/pvf
jv3uFsB6aVx1j8dQhULqEL8YJE+B1CdDC/YsKyDAT3MNtN4KtjzYoqDgb5kg8mcGzJFxVeGEhG8O
4bzUSD3i2w69yc1FYywLm6/cODayyplBIdfGMyQJHRGjc0u6j2EcsNsZyXFGTtsT5Ejv2yfTAGUE
147ltPTXejUlIMEtjQH1X2/V/lcl6WuS6PWYboE/l4jXC542VGAmyFnmQJuVSnXjkEO8DlQoCQPH
ZiWcjAcNE+u5Z1HbCY89dCNrf4YKlPWJQNYtGEDeuTa9eDzbwHWV6eozB+s1NmHXC1LKRShqtviV
7jNG4goXiOXhD9jabt1NDWzl+P3MIjxV0jzncK0EBt0IRv7xUbiNKMldawTrLq6SOV+kjLRmQcYu
9Yhz9khQa+kXMHXQsW+o+bn/Qz5wC+53DNWYiMbi219nkv05Sci/1d/EdLX3Q0RkgZx2dlmxq2T7
gVOkb5D9KOniG+riGQiqWVjAGc/tmL0jnVfSHOmJIM/RGIv599xGOIbhW7LwlxOSQlZkOCBQsKmB
eG8iQo647vdIowfTFK8EAEigMkwWLtG8VkJfuOPvJMXcmxXx8+MnIoKy/Q0QMY8CXRIQlvKTMCkW
tTlVzDLC30D7QTgl/TW0urVt4L9nqPqCceD2YK1q47TVgqhH3Or7yfhXWHZ8gpNO8Pw7dce55aHN
qGWi2TOrVYMdH7Is1SD7GtB5s4EivmIz2l115TCAh0We/cUjRudzVJdDcPButDsD4Uy28PGPfLKc
oZ+SiiNod3Ls8Lztlvz4+XtQVedTYVPF2Cvoca6cr0v1AonzTet3BQoXPVkGnPjO0Mytg85UFojk
r9gBus8wSOaxYK7x5So9t6G++sG7Mp3H3mViddHYmSP7b7/9r0cCGr4GVpvLbjZIBHYRHer1d+aj
spet/tqC7vYxKgbGnHAcOu82ZZyh7/Ms0mTcb/HOrucnKPE5F9uxewSIQINen32NprWEOlDzp+JL
65Pz+3zen89OeCel/o58pNLUiM+/A5XzB+1l+tOAjYsaLB0mJKnZ6IqLICoehBpHpRSvpiyBqAw5
LMmtC+TuT6uH1S4ZqG6zmGFN9y1wI39BqmWLbh8iN+CUkZ0kM3kxsbmtSngRM8VypUfwKQ6FFStl
WXf/i2MtcUgFuNA4WD0al/fD9KBxeCLpvLifs6FYGmaHf0D59UyuQSt2PYNMgJA5FupNDy43fYLS
FmgtXjFt1R9BOyww9EZChEbukpGVUjvxvFmOjkTWSyL98Hy0se6bCNicGO4Aoc2sIjl+UHDKt7hk
LzaKmTwCatbPn3xj8d0cKzrs8WWMUcwrmPiOcXRvomiQVbbu4IE0SLFYgOE9cXBQVQdm/0NuNbje
2nYjHlvNpV1flEenVFDd5rD4VzjRS+NYBFS/IN8RCDaUf6KTgUEMxtXey3EBblNkt9M2TtT31OiZ
JZKJXuYlLigGF9BTSLWDfPTicWirYbrpUZJ016I6ZRfMn9nhTkv7LLjXcFUjWTbMwQqjB3unCeFA
OU+Pi+RUaxEkqoJWmWhH/hfQK2cvW/nGYZgsFN6I6k9MmpOETKtT5PR8ngyulvzGIVyPXXkZiT1i
Wvp8pFdYZsFltUQ2K6XVkM+yyOWd8yhWU8lmzc6MR7/z8Un8WYtAf1L473kwfQZgvwRqTqNiNAXb
EkiK9A3/jlhTyUXH98k7QiSoqaMaeXO1fJgQMLtfdhRO5Hrmw+kXbYHyIi6uHr6EgBM1is3sS/vl
YmoGWI0AX9f+EiWS0kaSkC32pddwH5TASGAB7G+skNID1rjkLwrAJ9etbPuu6k5VJZmJT9AisjaU
z3Z74PrFeNXRTq1mRljuaJmiOMiJhxTgsCbJOA6FuMovvQRsNMCql5IyFHlrtGr3yaNrBNQg9j+f
wCdz9Qqw7gcrNZ4YHhuqLiCAx7Tr2Z+beCp6WC4vvF02nFpWSsS+rdflrf2/PCndFJ0MtC8P/FMQ
2ngRdhtnqljZVB4lH3IMnefqixuIkCzhPBYH3qPLuY+3CQV+BvB64bZ5nHmrYGJJIoLCdRNtV2cS
9WjjS8Xbv9YWfbP/HYzSFGNpKQVX7pBHjwVNiomae73mhwVcp2WSb/EbP9tUyQaYhD9bqcsiJih/
Ec+lYwx+OmnLvdqxAiQW1oNM/tANqAvdq6ddtL2IaENsSmSJPMh9GLkmMqO+1fI9xpsyi/4eYgCg
wLWYswno8ve8pJ6HX6Fs1xSHO676otCQsywd6pEgr8CL1pQCmiaCJsIKWMyN8bWYLbN1pSFqve+f
9mhIWZyJNMnl1oTfdD39TbBsPqegTpO+HqE5KnwIomNUeZbc1BojDRStx2B6gTmCcntyXvwi1mP6
16puDBTfIq3+gc3qzhZno6XQ5O9wItP+ogUXWue09jX3QyqFnl2xgJViNEzOuJ5QmLDM1p+2h/rh
H3pCXRtO31Cr69GsQLxM0QPhie9brJS7cglMsnck57sl9ALi1zcFjgWNvTbaPH/eMZkUj+Z4cfG2
VTzTyTSFcziyzA3WhiyHUNarudxSUCFRF+xa7G87jPBhj9zUD4456HG5IaZ+1s+kgxByJTbDz1K6
5OZoCHajOeaaJnOhd6Tz473XFnj/espLcXcl2MkNBv0Dulwz0qjGMi0UrjDD25TcNa8YHQSAvHx1
bMHL+xAz+tLuVYrFoL3fyzzggBIyuN4abEvHNn7cULRiC8Q8pZRGO9GQZGClIDsFH18YE1FRIanZ
0je4Gp8ctrbp+wCzP5735FplsHwzF7t2wmOzpuhHgpkAzhhfcuH5M4Ma43cpFAiS+Qe8RsTOs8cE
c3OZyyxzKiYDe2d5nHWtI5eAu5lhQt6qqiHfr+70GbcW59/FisMpa5TttCR3Drmyi/FGT2XOM8Jm
YOG/DlSGI+h1t3e9VF0nwVlxvnjZpfvFCF5FL8P5GSfvmCFIznz0glS20HkjOoJfS3X+hHv3hXhX
N3beXW9tQ3wF6WRlYzyK2CqDBSIFtOa978bYPHlkK2RroKFkynEOpYFKGLvYOtkG1nMZLzE+v5Pr
Vh2wT7KHkhIiP8fJU0VjJa7AkOUFEh+BDjOCyfABLVyQkBZPUYvnNeczwJfGYQWy0VKLVF7/JC2h
JY2FMlzbZyaE3/aMAjohaisRBxjdBZtIXXjF5DiVh+AL0I+8UBsPGawGWMSP3LBy12opHap84vI5
OoZ9mbgj3kFpNzYILUim+4bQTgMDYAVjcsFY3/vaedQqC8tgddCHCnW0v7HYWZEB0mi6NBEowpIW
03VF2TtNVhKwVNzGUlWWM5HVHosj9CCl76EHzBRmT/sY8XBj0s6P4cStzoFoRnRNMNk7LXDRn4r+
SxPIpN0xZb619OGrhkGhqcOqmC8PRbcI8xejpk/uVJjiRexw1NETBkj8DvVGa2mJJj2cWalqRTK8
3w0qurwabZ6tIL8fll0ZIRkcY5hEHnUmJX4P4Gx03mawf8cg1rST2cMv1etXap4lAW76VvUzvtpZ
lcrPT+mNWp8P9pe3qEvtn4fYrkfdvo/+j3+8aTH86OgnyUG8Tw2d4WAi/OsQkARTD5yKz1Ml90fv
jCwK39UoAWi4Ny8AkpioS7NrQchw4KB9pKPSue3ryT7G6lRCbdD/B41rImt4VuCXxia4V5xWhpOO
7iWD7IUHrG7U+gSHgC0SdUqYCz3QbM9kSt4Qgp/qcZbkNf4sgiDsymlN3eT3ZZNtpfzSZDo/1gNu
NidwWmxJmkCGtbQgrHhhFyQ3hV5IirzBNJ5VSGwPzTcN4wFe8J3q83wPtN5eV+ehlb3MyXr5/6dm
rvBxtU+Nj4feLMSb3jo8IIByTW2BCDu9OVxpe3mwH6L9kzxuKrZNHfd6SX/Z53ry6/okgHErm9BR
wb0DFRvLAiZQqVc6C8Wlk2F0xkEuxu7EVn9QzYxo5ZkJl6CVQWS069v6G7Ny7HenkC7rvYH3TZt7
CdbJ9at+/r2jEBJVufdumbkTps4t5IL9EGSit8WzNjZZH32aDqo5CRq/NBk1AKRNl1KwGnOW4w4a
7pw5bY1kRrU/0RkON0rDIdfCQ1CGzyNR5Giskb2UhvVIWPgt9DjwseOX5N3M14Zs5ixHaKrRuyCe
QU4kOOMAS9A+LgFSy3W2Myc9JrkhqUfrHnw9UWENIxFDJ0ULsdz4TJpY4HFMhjlDD8dz7fklhk9s
L59OoXvRl/A4kD+eSVJ0ODLjcTWaSlqZ/puBW7ZmYy1MGJlQuASdxKtXYkxu34TKMQcVJbcC5kuw
vfvvt7Q/KAPs7Ql/TWdQBfDhtoHCV4npCBDgFciamETB3uJ2G/PQcFTNnHrQaHF4JkGbV7hDYj59
58NwW2H5ZaPiq4lBf96YM8J0kduS8xfSonqAtzHL5LktV97jVklx6IWHMZJni8Jseq3EyVcRR+90
00zU2zptGb0e2xply7VnB+ZuCZ6sIazcOWaPe8YIDR4wznOwZtyZZGdZeJO3O8z21FDwfillvzBy
lMAGNAwsKE/A7Rv/Pg5EJme9H+s4r1yBw0YVovDujw+QOVtcZbhq/6FkACX5szFycP+ORtNyeUn5
xgJSkKiKU8LqidgwVnz46uOmrEIqL4VlYK5XTHJbevjIos6/6x3KeRDT/OQCnFnfC6ftZeonXQPO
dmn/m+VfLliDceXVawvehtHsOcADVkFI8I8U3s7MiGPIjp8Fiq02Aa88bPvXgoCJdCqIKjdW9huv
O0Mh9jaSyh4mKVodm37KaoDV9TNBCidpFRMWrcNp9mZUD1cgrlAc1euA4WKLmgZEBD93+nAZJkYq
zIjbU40CvZVzA8j1ofoB/0GruJEtChKJ7L+9PA0wI7xM0dH1tnUqiegDGgSTqx+DhxbQISoLcvV2
cJB6AivVp6uMtYUy2wQHLrTctNQ8r7Ednc4zeFCJV/BbP7/yfI2wKterYbKoY34GhcNSSkJUrgBf
Rcts2bE6jo5nJV8V00yNJvnJKyiVEfX6RzxCQDi2452F8nLJMJ0/2WqfxpeKaIMPlGaKY5Yaisuu
wz4YMKC7hg/a66WeRuWWnfUvZW2NCb0bxUZKQBQXnoCN0T5l2Rt7NJOf+KeL2GHf9Xpeq/2yfBsF
+EyblNQkSoKfeLUMfmZbhVCQvHDU4og5ouIEqe3RCvsTQhczJFqYq5GtAXzQstBxKDvvj3YhVMtG
cV1M+GfNQPoKaJy3WexchOFs6GR7Jhh5Lhb5mK1xjh844tGROhuJVjyjRicUlSUABozL0Lw/4NlM
BC3NwbcqtaeQ47Y1AO3+9343pBepvM1XMfYS3IaklQBHLyUz1GDlSekSj8DnDOA23DXUbFL5H3z4
6Wor2Cp6QA2kyo1ft8x4V0jwCgdx/VIDAyEK76fLiSKz2z/i1C/Fh/lKoNpg5U4DRcteoWNPHibD
D0xzGw8CbEqLfgzrNiolJsMekLnADYdo7alC6W+f891iiVnu3IEOi6bYEdwTkjFFselML5nVX/r7
tOULAUPv+a8Hk5TDEL2QcFDU4/2BfDZ1JaipUg3vt6iEIxfk+TLmoyGMBVRpTgL2VLF8BSi9MBce
iT7gkbQ0mKHCefB0CKHpItFWrd+Lj9SSOkRNEOHHnXDTl6PulK2v1kfpYp/CfJN0oq4tB4emo73d
gA7a2jCUjuBfD4Ox9WRv613OhOqqmQuKeh7o48Rc/2Q6n2t/Bxz62gaTgoRSTMD8HoVrDkkTNnPo
GWK+AHujqMHG0QkjivMclFV+XV4misyW/3XMUdJQdQa5D1EzPgnFxt9/splvWN2nBZjsZI4p/xxp
h1qEJzlhlsO88k1JHebT5j6DaZPjxfGprvSi2BkNasM/5VZ6B7KwYaRh16id4jHFIt6Dl9U2XxZ7
/fY20WjCzrq+/3lalsWnHcHMLlQmZi2F/ZTtsh2pU9paPijrGSmXz4z4x+D3WN/+OG3Ou/9a1g5j
sF0SRIY1ljWzCKlYywCT7LzpYli4EcmY1eiodxvHQbHG/F3C302+/hsyMpNHbA0gDLYKxuTn8d/c
L4VzuDqN5ghpoANm8i6bUwvW02NlyHCn/byyyeOrDREbj7K+Frk9u1lnY2tR1piUjmkIvXuDbItQ
S2SHo7o6wYeh1aPTLtMubaC3T5rekg/4pTZ6+4vdx3GVbtZkoR7CV2LheaX06n/ikDA4jNEBD2uw
SnG8pHwm0X6FeakSfxK5sFb5hXagvG4VDon+X/uZHTRaaJfXoPUcL7BJMzSB5dNE0qVozb8e+GHk
LBf4KNshI7EXqRlk50FHiDpYgpt5zeiwebE9riytTHoBoChHzFcgR0auCRiwLYWl1GwLIOVvrbuS
M5bEW/l9RoVz6wwrnYAUPgIJpm/gpqOkIcnHpi4pwfMOkTujJru/FKFWqu0YvlVJxLTifnOHifUN
KBfHZ0HloZsfjTatZExEy+Wt98BPAv/w1dbCwAz2WT6rP55+5BJL+QxcKYkYRmtR7yl2vlNWaiJ9
riFT2GYe24pfg1vRiHLxJwdP7CVqObNZdZmc44vsO6hNXONOhdLR8+yLhkYLhNm6tyMqQSRkcrmy
sknC2qC4+LcUX3KBRzCNbkOIJm/2Mb6EmUQsLSsDNbXJJNZC31KN2MwQPwjkzSh4aHKZQeOOLQDK
vEj8GBm+VwCc01JkVLsXWCENtg/yRF9fITM5s1vVlHsnHWb2ml0QdxNDN/qLKdrB/dhQfcwcDWS6
SY2Ugo99zAT2gTcDONxnhtklhEZEerFPSPF0xTCYxL3MBh8YS6AW2tCsxCffaJFgFtcMx66xSpRa
L1xdR93YB/idRVvjyqbrJfLtLbONRiggT22OP0We5Cjv2//nhG255PGV86b9tTDAGK5GazL5z2AQ
c4MXvLe481IP8gbZt0CSliOAvA+FDJ1Q1mTPJz9PN+hTReE7zRhbgx+GWqjT6Kx1G+VU2lhjRV2W
BmV9mWNvhSNM2iT15JaOnRx5LPh8AuwDheqPSeFTUv5oaByAp3a7CM+FC2ERERfaIfQxZvSP2WmF
/JI7hdvqtIHqeRDEtk8V7y/aPc/varv4aH3gnJamkOVCd6nVbBQb9mUsx5WoUJNzrxUlkaA3E0cV
mW2+dPR5szH0vt14W7g7IGn6d2HZIZN38CG5FMyTJpYjoWvV/uUsWjIIYxlBT2eg2KvQeX53rdDR
ZY2P2HgNBRQkTj4RdDfGzFynjXThb0BSRjYicZKordbMjUNErs2alaO//CgGtBKSxoJ/FR1i/4Ud
tLu4Y/ZWOvyFk1b2C4kuV6sD7CsbLZSxiZcGknMcVv9XSs14TotDN1w3ouk6TVj/XjM5nUDwVFIa
uxgNHifRVqusMpGKszrRsh77ZP+3ubDXa3/ka7w4E6CLCvUq36bC14riMSl5YrdSWpXri7tGufsB
y8ZPVDcCnSvJeSJl6xPjfKw8P0fKT9ydXgreraBVaUoRDekI+yXy0iHPeUiwmbYgL3+TiqCW9sBN
1jFSMy4mJ+DLj+SrkXJ4wyRljdgHShQPyQ9gcG2/59+aEvTCaRv6i0wjjUsdjLRKChCdo8neEz5W
OVu3ix5CTAu60+9fK8O1Su7JJr7lJ6ILt9IGbp65eiIlJJD3kppuqiFpFAZz3zwXv4AnXv0+Xn7e
MVLgIyO7KevAoAfMzQULsdv6Jg8gw0isI7jmdn+BGqIon3f/vC7Uf5NswPoTzI5dE8A9LnvTBN21
LgfauPLGPBzYToDEP11fS+asOMrThkeRSNSmuVCOPVSR/LtLM0om3NSs2gvgN667O6wmRGjvXr0Q
Z0u3ODonINEnVxgD5rrfhYNX82L7et4fjTm6XD0fq1/8c7VW43HrL5ipE1q0cg/tP2fxs8ng0rmf
rGa6JH29kPgcXLDtP5t8JzNIXOyxqaPVDT+0/+c+CtseemnGyOYBsLxzKdCcVbHAUNyGneuwiB6l
TMfsZzOOmdSwP6q645VYcVcuL6gbBHAPjZDM4XcD8WWTxxw/80UV/0ckHNcN/oqfw17Nud16YxSy
5fUy4Y5s6A6NnoYyQv7nzeGEhXb98LNxUXBcA9wYc2e1fkZtONpRZuJXg/QYH0/TAEtUR8MzeZfp
r6KVjd9GX/3HQDDP8BHQS/hCZBoEwW8aQpMAP446Y/27IIcG2Ml3w0N0Gx5xMmlmio1LH8tuCq0E
ZkGhSB9v/bHf4k6ESgQVi80YN3jYLjeHZzqe6SiDT1bxbVEaBJaEnUa89ojdf1bjd5+AuXlEJfFq
gStWB5/Opr2FcSSsABGNEeEjgZShyJcaMzyS3YgpYEIhxsmpm7fTo+vbmoS9JzfsoTe+kd7VivYl
eBOwtUbTn7uvf/KH1m9ZPtnJjRCo5iq4EjvMZbpyqkhTGZ30TCI5eRlsjHw2Y3zCmTY2+yCngmoD
r06+lXHiXw09sf10pMGn8c76keyePU/qp5YEcyimmSWaVmxhLNnIcZw1WOERaLpEyFpXIxsyRFOm
m/G9cI99sRNlcipB2EzvtqzkEK/8LSO+we3pcP+LDBuPQ0N/Xj4+4x3JhpLrfDA7c8851v3bDC2A
KetEZhazaL3q+OJZo7EgOZuQVQMSrwosuZcI/KAo0TRloublrtEGvFno15oV5ecYfSKaIkDFW/JJ
F5iognAVBSmR8RDMrtGO7r1nK8M2qO3UMrV60mxugCjR1SbmnrBvI0TfrtCJEJWaDGZWoyEwZmcd
K5bq/TmEQDu2HRYkrisEa1SSnK/akOXDMdbTT0Hahb1N7zn6hMaKHS6XtrfxtxjL3xuk6JpeZxKn
NhYcQweBS8NOw96z89mxMJu3OXivMFOKAZeRNDx88DwHmlKtQGXWCxALC04rOa5q9jkQjbiZzSbP
ByOEPeFIlzCpy0xUrG70IsKSdu3z2Q+G92Z3ALEFcr7kmMVENupEp+dsSedJNX18WZwUT7CuPXjU
2ZIlLN4b+Y/JapC/yQ6zg/7hnyFM/2KlRSjGD1wieD2Y92GUtYkZmECnmL1nAiQLO9Gnz3TyYvCC
Hov76TpLxB8TiymbAyM97iyixzJnhZAuFxr/8lBYdxtg5Z6maRCYlfsCFLx+/3ayDTnH4j30ILI6
9CRPdwKVUlhFSo7XXIbPPqbl2UZNI4Psz02aqpgjFqkXKfBdvIbhncZVn5HWIu7nHV/9Jf4UeKbf
R/Ozkjiqw+Q2ijaZ1KHieB8YmjshH4Vfk9Fbz8A801uo3wSAXPEUCBuMI8ucJ+TA6xXBMGPA3M+B
1L8BZSUTFLhT2Yuzs6QMWFKypUgt0iCtVIMkV+QZk+q69z+SRXITdBf9FCS/t4bOMaxHU3r3+m5c
lsAaFD+8Btn9UMgLeP+VkCt9evCPGTIDJzi+VvfCFiBtqnu6BuUJPaF4CPpvE/zzSe2GK8GSe/Ii
enXGVip5JD9rXmlnTqa/J+vu6apBmx+NmnjS6iTVhg0lXGNlPh4SH/yMyqH+1PcYMenpkL2D9dwz
pgzqQ/QCw2fRR1G1hWU2uOy1noMEsKZmheUlgTFVzIo/U9LuFR96/PRo08usDvd5PbdkbkZrnga5
qJbeT5GovwU9SchAbjORgc4Hld7dntVJFqdAvY7zOG4vFvsI8XokqiMrFCy2JtL0vQBVpXm8/RLh
E+0WwsPuAKR0ujWlg2TD2nZRt2ymMGaWTf1HweJpnJDha8Cmf768Mk8C60p55YEkD9D9kuTDysWX
P2qShLXWi8HaMcGE4YYD8+gAFsif65vD3fFjEp9Fd5/tVm0V3hsUZ1oDi7dnzrZGRht8y+zM6MZV
e2f45nFx9Clr2vbnZ4REkf0eMx2HRuust/ll+sPyNv9cVz/AH8YTgIWmUWdnQIZRyxiTj+IzZGbY
ezQ5IjzgFK22/ndTXBEIaWsZtH/4CqrJ7NUtlERmTnmI/R3cA+33RYsNpWc+EIsZMZowgrth1V5l
YCA6s2DZ3hzxeUN2c6b4AIwn09lv4reHXMWmjZm7Ee+G2CyD2PZzdsMcfkmJcNQnDPvvUvC0z8fk
o9y/GbKNbh7CnfEOE9Wwxdz+U8IuayMKmveqagcWFEf4uzuFJJ1iOeOWSHJs++BSPAx0lK4ichuK
8NQN3asmhk8/q09qGY3DRBw713DMcYWoXoJukrfrdZACkbhu9sxboonDnfdrtDiHVf6lz+Fl9lO9
WbJRBcCOzaAcPrN161KjtH+p3DbwYYBd1op8Z/XW7kD6X0pZAEky5QtwwIxyx71SG+sGVmm/9Bd0
rLdtBRWgvKtIyJ9jJDWqZsbdC+o3tAPudR4zAgGbs5YYECaABcHJC6ZDgA1iTTXsd29Csx1HpaiG
44Aj0OTukC8wcH67IaBj2X7gBaWUroxPz7/n/m+R+4RLYUcYKrp8IHM/KiygJH9+QGDoQhaRNk6y
ZrmBMpFfH1OJWR/FSSIiexX3MyYI02YVCDLUzKP8IKuAUomJ1pFcnMlku1W53i1rvYpG6YRwHNwE
t3xoT4BEui6IXZJzDH//3YxjSGUyIAc2R10r/WvuIKhlYgHk7lxuBcVYOyFKv9rhGtqA1hyx458u
vx2oouqyIUo5UZS2A2DWQq+MsVmHTRCQF2IFdgbLbRTtEfl4pC2jM+okTjOkSxo2aSCPgeYZih30
wjz2+/2cQImgr+zx9LqRw9CvFkDsh9mKcftfzHMzTmlbZtpyQSlHCHaiZxf01zFJQcheSJdCcK6X
1zUWx9hKJzxlsVZ/W+Md2yg2MdaPTc2hU2FBE8iZrcee6FnH8vP7EOam0BS8TUwM/y7rjqqTSGxf
jKC0oa1eYX5RJfaAh2dFW3IyNDtVeEhOFeuv92WwsbNuQyLTiDrzyMfLR0dG9h+P0Slt+XMaYWOT
oZusZiBCexqLxGhNzcdE6oy2/m99s7CvGG7aBoov7pzBwkGPz7fXJry0MvLT8eJc0xnFB9zJji12
elwwmJy+yoF30MCgGLKzysCHsO/NVdCRdIegZDNoELrIiWnPtYTISQjNHtQM1lOQpdue71XoEwDN
O6WnddooyWDv9zm7r1Q1mazvys+vZ6l2msHQ/0bB7aYsj1DVA5xms8o+OHLWXINOGfMlWGH06e3R
IGKWi61OHt0VR0hKPHyPjExhWdYqCkXPAhm/osCNBULrWmLiYdcKPlcJXA4Nki6zVlerJGJt706Q
rt1Ta7Na7z8nkAmZV35wzuqKwV/sdDgTv3hHzFNkO0/vunJCqXyIfYO2Y+AVujr4iSA00J6UfEUI
mAQaSXDe6VlNeLnied8CrllH86W9sxZooMviqIkt/sNAMH8FaRU/pUpuVzH1Kis0QIY8uQwo7pD0
KpHp3fHl6Rz1U496eGhWw7yH2HZ7vKV2xwtnGyROo+zAuN3t6Spq+uScCdrClSrDx3bDjIo/U79y
BrWAR6mz0LsfMVImjCZdxH96z/6/ZUJParvAadGJdwjw2d/7hLZHnv+4RixleWD01/ZSruI1A+nX
gK3bPtFtvEtveoAV8g7Idy7U/1u+uOj/gDXpeLMw2y2La1bQUwwKMCsbisxyBCR70AyhTRXlnnGo
eGfSYcT+XiyJEpsvNnYMPF/njYPpZu79ET+E6His0DAoCE6nH8NVkseT3kQOWjposHlX7h4+vH2c
tT8OX0EkufLe+wrNzChjfECSUlhRU72rsG87MW6Ea8eKVqJvN4FB5rRzY8MvAVknI5ICAInLGcCN
gDRGDPouPfNYFTWKSyIsXHtbVEOWxQAdDVwmqjdv7Rl1yIFWWOMULkU+gVa2nRA5XOKvU5ZMpaZR
VCH+eSWYqh/zNmMNd/FkbNHww5uELuZ+oF1HKnKBUGGV1DZLJptHMibjf8PzfPEygokiU69yIMIj
1QiXzTpfKeOEssF0388stcYQGKdEN7j6klDUva/wMZdljpLXM7SNphe/tV5Zxpaj86mc3UHtpaIt
BSQwB6N18CK4pzlw7Op4PYsvRmdU6PYEAfufM/nG8dFPOshkXWb73qvcR32a7ZDicBx4Pogw42Zq
f/oHB3CBrV14ZXW+gLAslNVHXLOl6xj5vxqmvSPK7lVbPjijUVN7Tje+/E67kWf+YBiXi3/jUZNt
YvAow0uNpccX6pDafTj4PRhxD52r+N5TIWfcyBrJ4twvjfrLOXkLZzzZmjOQcMqR97Qi9fLxdGwR
3X6unW3AfNYk0RkPZZ6t1vSdf2Nw/k3mjZOfqkk24XLSX4TcLHDEEIpdiyLe1mo7A//Crj2i+p+E
zPycGwcFqCFlS8QELCNVxFRZTttvEdjg9cS2yYXbQg0f8CEBr3kJYmkhpBo2mXtwgjN9NwN+iONz
PvNYc2M8iDVQvZqTBCw2C2/2knQFOlim7HsECMHsdOc2sGJj1+hrqI2JSuGb0Lj2kZH3wdGqRIwW
1LeFeDFB0trxoDxKqfcj8uSwNiN7thkKP1ZTJ3L1STYgaSsSYl1AGFLR97nYPGQjWHLncqMxWkic
BM+iyQIwkNI0CYqGTWEjODBXYf0F1Dfo/MGGo26U/bm8Aot4rfDlN6srnT+u0bNhO8NFJN4k5SqB
10Yx8FMv/b/w3mOEdr7o24O3tyTwpaewqwbaT5TdZP9v5zncrAoAC0c04k+FhPio2s4E7e4zuDas
bb7pG+ORkdTitQvePqEtVl5nd8jcn98Ctxx+AKlYGy7F0TzhTsKahSXnt1y+Wsofh7vnhqhqLlbN
1xw2LHfqVmAoYRrtN3UevquMMFLzAtST8PHDyKDis9iU3nVWxHGQHOhVRLnxHwOIu5uHStjuYe4W
wjE5zvhbRgrtHKZFjQKbDubO7JNpmMxP4YOjFfb1VPOfQbTazZ2lKjYlh8zlWNQTQz2ZH/VG0EGa
BYNXdHNdyXHHndSNT99+7VSp5sQUXViMPHNvw9XjAAKlpggHxxWxetdBJYzNpHyFh9iBoS2cTX8O
8fcaazJRlO5ysYwL3SzAjwgcOUPsir5XkQI+Yc5OzBF0dvEoBc0AjLvgk1jfDwJY4PsO0cQrOA+q
lNEj8vN0uax1nu2Or3OsrN/nplsuCEDcGz7iZg+EUM06cU43kBlcuxKfs9oP/bZlD+odKyKzf4ke
AnyTNNUB9VdjnofpMNSh0LFv3r6jQQ8n/rtn9fECVmpr0Us6oBCk+oHSB2iUj4yxDExVT9e987ok
zIpWABu/Fukp47C9QGE4GTT9UokdVQr9i6uB0GXZkcC8NJEC44iBcVthGaHd5JIkqvWL2Zkr62lV
pJla6aylYD8At9gufdC2xaRMti2iCvnrrmdMchkFXgiyl9ZpAUXKzvjDhfH92+F+Vehu1gogkNC+
HfN9Zq1+mq7hOz9904uV3njVeqBM5vkSC6ZcHCfYphkkihca3RB7O/L8xiNvL7D1ia8SZvn84J+d
oHORewV8GE9XJbQNGooetJeSDMYpv9RnF36mdWNS3qd1qeRPyMXijD2WMKDG7tp66PMBnk2r/iFg
9JiAoK+1qsHRu8VUafXviaXPrAqrmmFy8mvRqGCoH/KWosMdMncJcRC33yt7X/KrN2rIpN0h/WjH
wfZoCiBw1CHl5cgjVpqi2okV34hvs7CA3zJkp6hZIjK1N29RMH2gltwXGB36VxZfOR0++cWFWn22
r2+YbA2tdjwj2HE1vZB3+MZRdwQdqMjeY4n30Svc4bT3m2EI8Ky4iL8691vPSEb9bCRL68LSm/fY
fCyJxX/Rb3XxKbDYD3EFmjRYhCYnobMN9MSFwcl2DYgDkIeZw96ovdt1FcVx9Tvg/MjwPX+NeosP
+0UYb2TzlkaVrv0vmdlicr0ShR/6SZ+2mXhrCQCFdky+vEkCSEnOGLDSieeSxAq/sSb+SxRtuNmO
wSF2mm9xfldquXvbji+0lS8UDQqgl3RF+u4ow1VQXYIuZSIjeGJyTKlhGXvX+bySrZo0V/hCmQMe
exvlU+UEPK/TuEDVZH0OOYkWMgQLJAw7vO5C9qIlKa7jtvS8uzI4yacyVMVNetE6EpdUL5h+KTuL
Wer2XIshnrYpVos8Z+1w2TvEipnwT2bmMr2WOo8OAZBk6Yfe34v/c3No7pwMKTaHyFcEsg5Khgd4
HIFlixSf0xTXT7+Bd/9Ba7OiytxK3Jtj0RfhrevRRAWyriNthD6kLM/e1wRzKDjBzQ0/ppAJWjF3
aGshr45hAJezehJD4/6AT8phEOQfV8fCN3vdx6rbbTBWQSvNSfpxCzjza7UHaI323llvvALnG5ac
jlE/1IS66udRtWq+D5fuiuqZnS3YGzxeNL1KCiRCdAPQF60NQ3UUPe2v9Cd18VKlG8rXsZQyz4kQ
dGd+ay7rJ3uwazmbgMzGCaWQq4hQZvVnt0sT5xRp+9iCiqIoHYGfNX9S6p9O2C6IfpYiB44cCM+J
JJTRQ16Qzx3prUnDUU3LWH43gD6NInkXFbuFhixdTEH70Chf7Q254cWn6JmYVZtSCvFKxFeMQR+N
bTKboDf4U6/5ouo2xmVIahtjdQZOl7XeEJg2gKJI7ECKeSxyYbFwtiigRkteRwzN2+cvTcVX2w3w
zMhCQn3St0yzeHlQkwhzw8FUWH/5ULfJqeaFtqBB59rFPNSnbdwy9c7wS6Rb/NLR/NatKHx9SYzj
JQUaO14fq9fRoprWoOtWWjI6nsDIRcMqKyWxtAGyGNDzpussh8yHb3bG6dUEZzCMGVyM4MYnhGz8
/3q7CLIHr6CeQLeHovkipQnFCKifdofJ53/hHo+0R9FHDhLCJvOzkWBZU6seuu8gSjdqUfe+kgBe
kHVsneuhXAJU3lfPwgqS9ZT546WOQHPgN7QGjyIetlQ1Kmv1WEnzJLpvvi3DL+rTcIchWdRjinot
Btx9uMdOohaMmBxXfRLNjmayJj5AD0qiYN0+5OtbS8Uyv72fe2caL7p+Ni5j2pe4mVR9MjewRmq6
0XVdMbFJvEdQ8MGv764X3UpXjCYTQ5NWmoq1cvHbBiEbZ3pjctpNokwMpH20k37JlWkTBGXR99/h
On+haI5pYDe/0Lc6+q+491OEMV1Eqfdwii7Pzi79DYjNWhnWpz9Kgg1FPtj42VYLm/EGe22J4clN
osLGvMzAPNTJLOK0BAQdH6PcNhwcIqQnapTM9rnDGHs9Nmrrr6me73ihNRW3coTrO8ytc0ZfIyyy
1XSllU7H69/djNIDbK24adEtWTsxmD3dDIjvktZxYAeSP06U4uVeA0pVJCj/IXZi1fwfvbw8cULd
gFV0ov6Igbojbqw8NGzNQTpUvJ49F/aRxpqLh9XtnEzhzKax/wxN84W7+wkZ8ePe7ysm5SaH8qjF
hf5HoFR+CqumfXW4YjsXJkpu9JpTb6Wl2BfIyrn2ZHxyzPkEvdYW09t6nz2guAQ4PJS3H8pJ5za3
CQoxgxYmjvFs1bt0lAV022w8eNFIoitXUlAY85m2HOUhlp+DQjRzyi5dzmAqU4s1AaofgMabGhG3
og6KBpL9/l+HEUd9jDPUPnQi1ZbZF8nrN5LUqZGCI4w+c07wxd+lGx/K1Tfel+mkStCppuEBmOWR
UrCICdUZaQ67C4/zo/6cmWbYlEpm3JBndOdTYGvttdPYmmDwjeqBCVSlZSXt29VJePEEVuYrtc8Z
0rNNjWNJdyt3eRiSuSXxx3oYujht8vfhOGjeI5gMIabq992xELGuetjD29GwiYn6Pi2ofT6lV++O
7yclo7C7ShZj2r9lXbCl/LnPEKFKYn5gSyeeI2hOC5WTQHBbTrndx4pbJonCB1IGnbmb2ZVL1BdH
mxDkpeKJ8uhe8tT+YlZdU2H9ijc2T6ilF2AtxL8pWyTlhNqzhnFPLeQ0sx6Ra0Oa200JDEJmd7HN
HlMv3zU6JYIt65DciJpeYPwZnP5cmYgX09jQM32XayZqQ1tREmEqnoyi/oEdNou9jAi0525RRP0x
JuQaKfkPaF99RGEK/69tw2jCGOuldqkFPTN0TkKQwZIsfBY0r4K2i/Q0KGyV2nwuZSGjp3eghtB2
OtBUNSybO9IJ/dBKss+n7aqpoznQb5Y3Kw5saHblLUGXyNfZ6PKhiFpPMFmGlWIb6xedoipcs7yd
uc2F6NNpe73aIzMPKYSEmPPVlj9E1MUp5DeyrjgfRdvRJmNjsixZAxtISUSbXzEtdJSK8J43cIft
iu4bVB4BEk7bmfU9J2cvClOYMnqlyuTe/RyeR/4fiq+ypQd9XXRsi60UBaJqBI3hdy0pIUrvt/LO
ciHXPNEFpPvStRAzPaJx4D52fGXuMUmZgmRhDOersgZYrj5910vmeiJh6yCoCfYpXt0osA2VQOHW
HKhP9oXniCQmbcS+0r7JneKdgLBuFHE7t4ByBJG5oNBOsIu6pzo7A8eVxjIKV6IMQVGDxhLGxKcm
21u/TgFUO3a6GLxqeYyioKrujkO1H7xVpFiGCkR1HEgCsbwzsQDi0Y72jHGaB43tg9xDGQqwF5G0
nBVAHHVzgdQD9liD4gJIn/LhHZlBVLSfyETgFM6HC1MZEfsl8ph3a6+ovP0wJdUDTzqZ7sDP1iRM
YgRiS8M6U13qfrOch+RP+koh7V4N7bZ3A6c9Ul+ziekrLyH8UszH+lAoGl8JA570BYQNrmSn8NCW
pgeJIY/d4mxpneTVkLAkGPaJ9WNF3eU00NZkcHB5twy/k8jmVKG3dZVDIt3hfpKbLrEGOOS8NxaB
rZDy5eMGxxYEajRHu4AAT/z9GR4bKGncYFzPcuH/auAta+2HqQVYAoZvrE3qAGnpRTVzc0npRXmx
VdKERq5PYkKzNqKi/kPePFNrlKPWUVJl/sHLJmvQJGYre4rhSoahkiSVE2OH2mlNwiMSc2M/L7Ku
2jp8VUqMyZVbQhQU+KHw897Lda+dOo/7Cm2/zkhraRBf2pmo/zklwijN2LlTPColVRV4ICC0bwf4
zfNCxcZpRVNjwzrlgSWbtBv7FA6CvW6qNzVXZ9liXRbELyti9Zo7pDO+F7vzptQ3fnlp8VQPMiok
3f5eUmI1lUKkmLVydCqbW1AdZtkYa4NwqRjdPPSM+fcC8YIOQW8tVHurReJPQTBY44bDRJEUoSh4
wnxV1hc4GaKH0SEz7px7JrjsWnw4tYymK9HaeakjUfnWPpRCIjjljxvePEO005y7DxkrHSE41ecR
qaHx4XxHl8dAUmRMhyk/gWQ+8w6ya6xNFl7OBkPCY6rn1RoBeBYBPWXkpswdMo/w7A8WyX9Olibj
QxriRl+HmWkxbakkZoq05XB/6F4lEf0ZHrdOpKG0BvQxhWierxTHy26a3C8oc16xJB+9aI2V6CjY
j/Ruv12f7Ddbc+ZI5Y6gMfNOxBuokldihvwnjUcM5xr5h8c9rU6iGvJQi1DyHo9De75q9E01bwPi
l5BNXOpeM+wvs2eJZ71mm0cyA9Kv6cfztrWjOKZbghl4fh8P2o19sQVnMA3U87ad9XOL6JT3RYAM
is6Sfk+OBDChl9u2tBPzsTm9JnwWIKbXZvmuIzKFoUkC1LyH1gAJZA4ZVl66rz/hA5XWJHGTMlY3
Osj+pqpJAmknWh82Ap7RP0RURapyHNfZtDGpb66rg4EJ72pKmZsGmoin5Vr2mLAXAPuoZtMXiBWi
YC/sqIamczPOzWrlsIb2cQ3W5Ctk1S9wF4B38LV774ON5UY2bnfUfB51MdnhzEDUypPZ26inJSf1
9eUvPdcGe7nj6SjwKZCc5M/Uhn/iiZbNulBqZMqXOY2lsJNTlmcC5lGXAYkHQ4Df/2DbutjkrmmA
RhuXU9iHtOxg++/T93/LNZQDHcO3Y8736HA2eiFnkf0KMw5GQI3TfNjVM99zJWfW7Z+mBRH3mkEG
cxc8jqFGkrRlcwPWgmvOrokTGCTu1+Ak8zx8sGTjCou1VMQ9rKzUQDeFW/mr8jnBtZ/IpW81XZNd
wPWdN5a5QNNzL98uFcQf5jXngISIY3imQvRB2VTNJ7aOUJR/GNQbZYsSaKx1Xt/F2UG9onF7Be+X
+s7/nF2iMBnuoX5Qfe2AvUx0qs3eGYFGCcxjS750JPPL0SDDmQ9jfkdTjR1FCAzmaty7DT+PWCOU
V3fjMbMstDaPPbNa1+eEKcpDAmwy2/9yJZiYZlqV3Hf51rEavUR7ixYaZl3c24i8FjSwTiPnVGpH
E5h0iksB9vpSMPtytex2+NLNd2F1rt4/Tu+IFZkIZptQA9CULzSNH+YAC3KLY2EICY6wWuW/HfSo
gYYPBdHokJ3Qq0KA2ROxmMQCaiOUycXH8ksNhvDomdMYz4KJiksPCBHU03cDpTsOI+RjpJpvEB+P
sHUGRngmXMybe/qev84Xbs+7IbdxO2vZGMPsmMSmskAWJ03eDjUOXKKKYGouH8skV/eCtPUT4aux
0eIlhrdo9tIO6uhSxEIwikS+XS0x1XWKbe4ScCyWbBsgez00E/zmO3PS/ExD6qp0rDcQwROM8+Z4
7NUlEsg0i5zdF54U3FP3+4lW/YGSdBFV6HQfbnzIgtly8dMcpopDzrXtn1CpcUuV9Mh3TXCp4yMh
rr7ldi3YdF8e6BvSu/7VLcSd5VUUmVaJqsgo6s+FruNvUbp0vATJ0PX/XtEl/dmj0ui1TXTL+MpZ
/jqseaT7jJ/g7f23a0alGkiELjK0iA6wACyhAMEwnkHEXNpDqs6ftMZOz4Tli23+6tpYgvvO7W5U
x4PFKHrgJTJ2YYXaNyiwPsgleJIdJHluan5Tbq/tKa86RYWZ2WbC9941K25Jx8Wp6xAmWD3cydn3
cpnsTpyTh3+R3OXiMWMh8+Amy0HAPLemUcZGvLZoJWzmFLGI08Chy3NLOkqg6PQPREdIGrdqPdU0
zh+QmencgT4siPigpnn5NBWeiIbsWi+mPK4ycibsLCtZE/si5Lb7QerryBQR+KhABPCk4jHR4L6A
BuGFDLZZ8Nx+/V8wcH3YsholH1Wp6ygU04lo0FgB4ucyiw93UDnfiMOFrKYQwfU93y9auH0xkPIG
WwIRRxmg6iX11x6wFWtRBMzXr9JR+8h+9+v7grlBGyausJXoq2pOCve32CxUpt2A4KbNfejC13g/
NQ7ByegutN1F331cKeFMx0zGUFMx+if/Fnw1K6g57cnIXlGuD2B9aQ2mCY0fLZieJb3LH4JYxMeb
+nPKV/GSrN2TByIZtugC7KP2p1Aq8tDy+jzwEyVt121xXPWTbAroNS4c4uJCwyd1Z9O+TXVuRcWk
SP81gOXSD8Nt6wAKCpsxWFxreakoLnQYMI6Wf5N/Om5HPk/8+T8xJKcyL5LI0C/yshKWe1vlwEfA
Lg+kv4xsFZSf2dnetxGGm9md2Ywz9Qi7K4RRsu0ixDBAOLkX5oySLpmikJ/crdsFtAY3qrmEmWcM
KDplxZLCTSQqZM9g7tZCQW+YuUiLIJPeYhpOBLXEFuiTiNukOvL0Tqc33LqRz3gG+ekArUyNX7oK
j660ZZVJHOHjnCtji8T4/WCQl+iIRqgoJb2o5FylHq7LJ9Pz4PmZVRF4UtuVMWbwOHMkjDa3lMo/
tuE5sFDvlFES/1Uh4sfXo7CSu1ZmDAvXOiINtpQ4AWovWOVFdkNo3RZ2HTsPbK3pYXFJTyt4GfAD
ef42L+2NRsgsCj0JHBYKiddRiFnddSjTGhYljhYyA+4uCdmHcT7JD/7J8rsCSxdcjLK0tjuv2IsI
HOQzixuHr2FW0hvPmL52tH/Qmid3keC2fSrflYfgfTjjqP7UVZFJtmrhNkdZwTNck0AUnyeb+p0q
IblNQvSGinz/Iye6qJV2Am/Z0ri0T+ywZ3h+vREz1Cg41LI4PNflxUNqAENBkfEeoLQP8Ewta5FG
q0ZniVltF2o2MGtCIfER45nfkYzxEdaGXbqlcPaj1LOsbRx7NtuzjrIcm7lvIjtMofkh176JQvFp
sbnR2Fh3ZxvKQ+uk+DUbFH4yeVHtpFb2qoPcLcPQj2mULaiR9CV8OK3KA4LP43Q080OlYSFy1iID
Iy3ByfU3LVq8pI23/HGxWbrJa7U6OwXtd969U3bGc4LsIBfmoejAifJgtXl9R1Bb37OuJlM6coeM
LVJsBt3hPU0liFFNSSY7dzl0h5KxjfauKrUdQTxAt/EeR2kIZcdLK1aFnhllc/sQaNjLvBhbyLL8
tAFswcxS3i859TvJ1HPC4CWExv9yWoXh5VPFfHqWw2VTeDd4529/8sMy6JJQ4gcRMoGVamYxjU/U
sllJQ4tiy1B9BXeBHA7X4zsi98n56WN2ftM3cqM352Bvt+Bo3aF+DZa9tESD8CG0NwWriG56L7rg
DZeYKesKk4tngtGCwJa89RWBZUh96baa0t/o5Z1vuhNnXgRDFAC25xKi35400dg6/PYMnB+twxyK
Dq1oXUA7GSZMjqs6gdmbqzJOTMMqFt/Gw78wy4lFGcaSd0GZ18L8edtPLiPhfslMT74gdkxaVOr0
s+Dc2PI1alOf+EjadaoWRoOsASvAzeDVZHaUnz/GmJTHfCSyisqkyYf1mmngxOuXTF3pai/IGylC
j6+SHHFZkngiV6yfn7pXn8KJtNF9TgL+2xLibBGPSS7PEMGl818Be2eMxJYWBmroCzC+C3+Jpxrn
zA0mgR9LpQl+/NCVHn6JKaD3iGErJpOzjbXWcX+zlwZBCjFfACMwnhcclx/TNW5dLJ9GnCMuAiGM
EqLO8S9K3e7PW6fsBuuAgLmxNdczsC2udjgKVhxMZoC+2AT2LFK1m0yE/TBWPZuEzrQ82YxWHx3+
POmL7igdmQhfSPrh4MUNxksUgjy6oYsqtnh2woCIBKgs5JWN9FI//aZTMKYXHYSWpp9csT3qMpcQ
ij/gpuRlnD9RX4ZDqjq1n6xvxOvdNt5jVFiIVPgmY/dvi8RR9235YLfF6czC97NLU3TAnXVn1cmc
kTVZLY8pIAwPYbFgja7l28FTu9+vYdr1om+VOf+XjHGPRidPEwng8gw/cbXYkjqG5XXHRLoCAKXe
Nb8L4LQ1QGGeWHhP9GGPdJtnBYUqZVVbnVulFPzh2nGia61nfQE3eWLIuG9WXtxlYdKeE9oTXCu/
ZBxM7o+l08fkcxfK44lRIy0CcPWjAYvkI0mPyb4+9PJpReQ/E15Zs2AqWiYeXPz862PxE+dBx/0Z
0iszKzRQdHI3dk+BPiW50bFE2bsHAeQz3tX7/kWFPIX9W6wS2yn2BcHII7K3We1y2k/0/P3VHY90
k5GkNanulcNiHl5YUiLw0FYZ5qBqRR6uBv5rD/CRWGOFuAsEBTj9PRPe0301UlR9DoZoiESVXN/3
+WwDF2DlKu3/kJM2THXJnv7uUVvjIjZWTE45XYZHv7zt7LdVemooQFTp581pGjtUOfdHboG51Q2u
1re72t2OSNMDocnaQDLLxhflmYVk6Imk+Ak5M42mVS46U/3E7dM1DCBzCl/02JwQngUEnt9vF3HG
+9NswC2w83gxQeyOzflW0n9gblmx57bGrjhNfDAdlykucGwXKSsrl6Qe/AlFFIiAFeFJ/KfSqvDS
YDPOLwoN3eYIP+fzDEMXptkDLt8gXZbirBr8acWCUJEFD53kiA9tr1PAwvoWL0aM0dy96pcY7mk3
J3jPtRO5jkN0D3B8Jpfp+nwk3bDVbYrkLUMtlQ6f+80TkGQLE0zER2v67tRHrxGVVAJt+G347RsF
ATuGQOqqI/T/GKfeU7LEcY8C7DhLZ3yGZX7L9Fz5mvhWk3sS0PVzlaFUL3nIWsiuIrJJ8UR5Wl9q
k4dmXIZzceJ2ITdXYOPmjVEA/X5PsloAKIoz7iogWzheYxtCwf7mSw2jc9WqIK7qDCf1IupFrJuQ
JvOb4c4gbkpjj19f8JP/Qwih2E/x+hJN4c01YBVGPND8M0C/0I4rLhYJm6YCHvvB+tTaBs0usJSg
ekytDuUyP0ICa0uJVDTUbkiL0gOrkzdJHuU8kPkCPIn6dbKsneR7kkeEMZZ0Wle4/v2vtCMYhRcu
JG95GrDaTeqjKUPHhG9/5EIIWyK+KkuSGZ4e9BQb6G2Gxa+AOHv3clbf4SEOVK4bCgATg3Fv1LAf
MFH6rwdpGr/rwB8cUOyRQoo1uBle3OHChNteUTQ/BwJCzCiWrou9fcFMV0Xnh7OSLfPOXavoGKPi
XjB92FJwhsKAhpH9LL3CJXSPXwNM/UZfeLwxS8sGYo3wbHtGRO3Z2JJnMoHnXs7BrKVe1sLsJuOJ
7Q5JiiUdtcEQQd0P+j6uOf9PNAAszRd6yDLx/kMvDgYqfbpmQaNO+SNbPlE8vNIed+sv6xsGV7gn
lVCdknofkR/AzWdilXNhXODwD4q5gKRjBub0dd3sLhho/xp71SDt3o/huJHn0aaif8la2VDMZqnP
+2Itt8HSl2SFoB7hcPRrihkkxWXdtq3DknscMd9dVwdRKFDgdR78PNGR41iQs1GWWHy0Rd9sJu6q
P7EhHcI9lpXTW5uiaqWRBqM+VAkBDWLnCs7NZ2Tjt4xK+6Ib8CTUqcAf1gmiA6gUgh0Qdltz4w7/
BIrLqNV5yuE50hqO/OZvCcLJq66xRREls2PYXxg8HO3DDgoEEhUYpqXWW6DAGBMKBTD4m9vA2Rm4
DQgarYqewGJdZTXo2v6/9Yg7kVnkGmww3BZcbqmWIwRmopI6c8RSYx2AMbqI6sMsjef2cZCdFxVX
VZVCLgWNcW9fA/ygUbvJ/M0/QJwYMYHIoepgJ3Mxzi9iXARoyHr7NWYPOx8fxwBwgLUepNIHTVf0
qNtDoSNoA2ChyZWsNQzzpkDzKwIqLOt+d2pQg7txn1ECujDN4xgFs8N080uQJnIIQPxe40oX3rX8
v/co77FlBhA2y97lTAyRLJQR0JPmt5Ikh5pEjW1L7CIXa90Okl5duKu+lQ6VfZ9/AH6vdj7zJP1S
cIZDqnNyfG0hn4A23YC/2slQOLg3CKc0SOkks8/yj6B06B/sGqtx8jIuoj8bIwuLxkNIY0vFNBCK
iWdsV7YVRQouTo0TKZg46N0DG7qf6j1/m8V6huwf9yaZMvAhnOeBgSDtgMPW1oFY+lwlUG/UwHDs
DRYiJLCy2s8LaYB+HSuGegRJrfrA4E24fka0r4DuOIXsPUm6HpZmcDgXtqe6pu4SHr19UvLoVHnT
VY654q+K8pvww1BB5G80NDgfUTYd68BOn1c/UNcNW9TV1sa66vQeoAM62jZlCRDpXAFB4idtK3Mg
zEzQe/gTnQPEZrUsS3fil+lJh7CoNqyex/awZtRYf3GpwL6poxpbnb3RwixjcfKRmVcmdeb6UW2M
vnGMWGpCCHjGQVGlso06prqtd7OpcvuJveFjuTv73DzxAAVO2j/xra+pENO9hIlU3f2ar0gLWM+2
S3ESp+Jwc3Y0khfRr7slt2W+yiFE+XfFZlJQ4nnBOIMGm7SNQBibFeSPfBwrKh0X2fhhRbhipMoV
q0m9SxHWBeTf+iTMTjUdqtht9Z3oLKQldo2yq/FnibqUgA2QkZ7Cv1xfz1aA6z1wM4Cg6VkeYoVQ
dHSZlZ279PNcD5M7zxd8ltNiO2a6RV54sgtQZVlwYR9Rb4/rX36q/AOCYL6hH/SD5NTcgTQiip9o
DN+4ZlzuqmPqcBzEgkcl/zCG78EetTWB0359z9XWtvU4j/Btuwpb5w51sskYSbkF7pc72nyGYoks
A8jXW+/vTELg/ZmZu32gcooHQXIGpBd9M6TxhlizzvnINlClt77L55LJII2USx7G3NAEg3ljG7Hn
erZIz0myb8xUHDomh5XGCDaJwtd1FYohnHCSV9oVc4x2nlOF0KejaNOJrfmxEvLhzEbXskPEKvji
rR7rJ/OfU5Np81ErnUagQgUzjgvipSKA/5ib3P2qAnRiWjw530gMdEv217j2plHpehBjKosnaF1x
PwmAUkgykLFl8CZSxdRbaJ7pFhQXjHq5HgXwUMSsmAzM9rkpoJoA/C7WL00cqIx9RpmsrSjXgZcd
vIcgwnmBdY53yu1FaaOtoZnIww6ZgiEfUvLdWe6g0hnzwgWIpsFFONAQ0KXeE37H2l6TcD/ekLnn
k+Wfy89tV53dDQmPiSkj35nvvFnT5jYZewEh+ID4GvVdIR8ZLVIVq4HwzSplKlTjkKAsrIK7hADG
8/xrTHVDtAdfFdI6KrdqS6A9z8BNAQFwmjzW73fOyGW3s7NicvZeeSFPHhSS27Q5BtBYfu0jF2Ge
jhHUeeWGtPA0It0vHQcJE4QAUSZQ52If+9SuBPfXg2zTqItkChOO6NVJ6DqBZPKyfWH2kUgUx1eL
v+hmGetUfZD5SMJVeaupHYY49Uwnlo+kkCZWDgjsBNh+lcxllO9qRHhGRSTUDOti7C1+lli3dwfl
76kC3uRFAqXhtZMMPPgXawtjLpKSZ4iopIihvd+yzoKh0dd+BHoOjophkHA6p2mzKvPVvv/KYBcV
aUhxFtMsFdO7QrXh92G91QaI3I4mOtsVa0yfLz7w4ahQfqJuvmFH60zVg6SGrmuvMmD2N+BOHcuv
G6Hqihmr0TE21QAWTosEuV8kpDAJTgmcHh9OkgRWYMPVCfiqsZUidJzjqyEtvQ/VTDvSa460PeN/
geoArprYmftN1xxwe0rKhhu/yL6UrSvQ62zUFuPTbzwmQ+AJhQTMVHk4KmPC+lxn9JylBr9MOlzS
Ved1mCg9xn4c9fZq45p56n/BFyL+w/54GpokDiRqp36Cd0WMPLc/08xgDaJ9lVGEgHk12rLhMAKm
gBHqXjI8oviW6eod7NfMqGLW245b1CTxi6ZNtUHZnSYu3xwHZ24s+qIV5Q5VNtTew6/puR9UAWNm
5xhrCSGA6MmfrlXlo55DaXSEaLwpSvQ1U2wlyaLscZJ3VjLvalcR8C+rGQQhDhRaYuLvNP5kh94f
/2ay7gxEXN8sE9tN36gdqrDYKi7NbJfWtAoAjfCWNkqDnxNNAbP+PNuRVYrC0wH/Uj+OayJFU3b/
Wx2ZmGc7WYV3i4WEd+j+XIUg9mxZpfN9KBXmYY28RBWbBX8n9jSvA7B73SAF7N95mO8i7uRfxAIi
zH5OU1SYVm/eAQGsObUiQy4SBcwMgVhXqbP3O0GPR8NfUNfnU/dJjmwN0aKxnqgK8pQx557MJExr
/5juPNNnevqZ8wJV0ydh57Sbe+oe6/zrVxy+VQo7Qy12ylz4O97cqO8Hh2rk9MwhxdUBmDngzCYJ
gzz7D83az5xFcO0sjFz9RyyMhvkdg8sJVf1RuDBwNOEkyz+BWgBjnesznDX69iPNxI+ELblKUFjU
3ipB1uZTLAFVdLhhnGXKrETxslYX0C/uJGyXLHHuO+k3JDdAm9M/FytwcWHaI1lCzlGkqg8N8ORl
Hbk61PFthZFOBchi1pcCq6uD2I0mbKWPbFU4nbIvM36guoc3h0s5MUSxoNVBSzSp0Y8/tkiYc01p
5CZm4MvE/ATXcbEkWjPjwYnhQpYXXhSHYozs1E4zK9URJ3SZP7VZBlVqX4GEhN+mxQQV1o0GETgU
NjvxBu9ijC9BwpPd1pXgQGZKOiDSCjefeO0f0VDqI56rlkPYqplWUDPfMEeAWjxU9/rVJ6qHa037
e7vl5zqgszYC8XzdNBg+ahHKMwdidlDA2pN5aqU6hey3B82cmDP4k4kfHsMYIav5XdO7MmMiEv3X
UZkVbdCDOC2yHQ1LydOj3TPZh+4fGm2ez7+Xn4N2ZWbDjy2zpwP30I6H43Q1ebBmIsrGWpzcTgiT
YVG3Oijuru+Mwp7OL1MfgzSzSGF8iemE7nlxSRqSkpKubpxOuIkw7C7wZCEe37dp/V71wBBKFJGU
fXbFdS26opiw5nzyntopJyYALrDTwPTtqY17Fkxn3X3vA9GpeeATTGlN4p9+y71WPvGEDzFoHREk
Hyrskic+sZu+RGnr8P/WK5s2fglgP8rdrCZNDXk4VMiq8HvSNyPnziVjBhiOE3kWYBFwd8iAyNpW
sx0qowAjUbPJsj0vJhttOoEiFXXH0LeOIUShW0ZfcWsCB8upSqs6p4YZpfYiQw4kHGGmnW4QwlIP
m3cRXBuROG9IF8wHZxYKNfOWHbHMnK/lW/v9MgkvMMqRjcjfLCwyBX7Az/OYrjpxszMqAWVCHv1j
u1E7HkctysFusZ1+ghotsDE7tAR26PsGt3mKtb3UZ+5JScwUBHODeY9NlPPbmPIYVMVymxFl/AoC
NbefRRJ8fdus1kAUiDbaEw2jmxaz9tyt7gT/N6B1NYjtDkalnboCZnHzs3/qs+ziH5Fuj8WZco1V
nNXxhaZvRFvx/NxlUE8XmqXlgSCQDfcDV1HkiPx+8MU/noJ2WXn9+jd2lq2SOIGL/pRrKeWFEKti
okKwdsxFSE9pIGf5ZF2/z6Bj2cZ6MXs0x9j/KnHAXDpeuxcUQLrYa3VJdoHlFRTtV1WiyVTG8h7C
w/PDP5qWt1fpA8Yf7vOrMvfe5qqSQGj2JC9Bv48o6y+aBCbvwxvkmbAdr6ITp0PokUfMdIdmw/ys
vJzc2s+uJ3SPhUjbe9uT0wRrJ9z9uJh7Qo1AbIDIyMOtS5WcMkLi6YFMAoWRcU4gQoxx33WaKtzY
hl+1RLtVtRtWt7jz9MIAURD6I6cWnrvKtq/eypp8FGcAKqpJ3SzvPVRQYNe0aln4YX+iTXoxgyhL
lDy/nuVfY0X81L5d0lAObPiiC0ZFqGH8+CQZFO0zxSljmQOcL+df9yz+kXHemniL/X5hvYnBN5vu
q+1uQ+LX+5uAldxZBNWjl072N9pXSECHlcf711HY7mkp9Y/1RhLWvcG59vSdhn9bzuldxRxG+Gcj
bWmQkO+Nh3yXUbBPbER0wVJ4wM527jDmfhKPXOJwWzoloitVOaPt9a2rIAuTInu5e9iTsOkIvbbd
veabMUYtIs2M6LUv3tWf8hBxPXUBdYjrk/FtcdUSstI0/pv0ibicr3kqi9T2j5LRAnJuk9Hr/PIC
CUKKHCrdBQg37WQLAoCSBDWW2riwyWxUn4gQz1a8W+VpgsbPxdaIW20v0VWMV8tHIQC2ypE8R7Rw
RjEFKY3+6MzSAMXM7K/288xN/4gIkWejK+mL0jVs9akzZW0puI1A4uH9PxJ3i43vQBJEFOSChl+Z
sNbNbYT8OLo3XVQICZaNDTebDOb72sEqOUeSvtScRRYrKA6XnOtfkYHREy6T7WM16bBLo/nNAtZ0
1e7ujcPfhgtT1AMF50oYWU49lAfR02Pfcel76gU8Ch5awiYetC94zKBhuZgJkSW6OQ/YwjzXm+u5
Yq+4X+JtbMS3b+RjNGDr30LLLjx5+V5mSX4fKiozvTKCYI8iiRrYWa1cMvhCBFg2qhSM7kVwtaek
+Ii/PJGafdzcFEDR4tn+J5svZxVE13KV5eOeIOXSHptj3A7f3h0lB9xaPurviReMnMQ75Pnu6MVv
4Jrgbg4ZLffuO4q4yuz0amsJ8Xng6NE7QET0RJLzmswqwpNrbApRZolBRLgKgSqKKW2jRPeK6kP8
U3RhmUc8DFb2bSFAzC1KLi4FO3Z9GPkEXw9bXrOFKLRiO7ToWTUIktCD6oy0oHv2pmQ408ljHH1b
uguzvF4riI1MoBiot3eXaubLK6nsgokhT8TuUga7pnwupEa7mlNxSeJJegL3PXYgbChH0TxJdyKm
fq3FG89b8nc0XBIyYBmJg8EL/+Bkl79bHeZC84GH+eMZ6OY9eoRUG3RI3mW3Q7Lz8gB3uKFJeK3h
HikcjNg17arg7GW/4QneWe3+gmnrerApebBdCz509nfFKQEjog4pKoF5qtMaoMhW4og8aCRYPHCd
DoYR4SXXh0EvHqgcgFL3tsvb6SUgbulq77As7Mp7wRcq2/73Dln9C9Kj9R0W9B9HPehzqAKf81+V
sDTrON01M4Adbi5PzS5LPE2AD8MOwGj6ZZa1355Yfr6ks18NBtalN3f5gR6LrSzAAR2wnvunh44w
CT8Q1wupRo1qdA8HbXT+9ZaYPLQ+LYnIiEGHStIKF4+uSckALJpCO/2mR8RqhGjQVKkYRB0ZujaM
LuyeSRECyXAro9Jv3p1Okg0GS0ZarGGctQqpiBBeCG05gGG4v0S8XWAxOPPOdvBKIeHAOurCFbqw
OQyc1KHA0NyR/JawTU5LLuDky0Q/Muphu7n7v1RBuBGfjeYfiU+1jGOEA+fy+S0F90AatwnV4PV+
e68vBJMgeZzs2DK/xSi0bLgjgRcUJpNLTN0JZsE9Os9dGW5qDALwwrIsZSU06/Pd7m0XlMMQZTpv
gt5op4ASOGjdOZ1GItQgts29u3h8RLJJtE7gdsIgkBKx5Fl8nSN8843EES38U77eC6XEu8dAUxeP
2/oMSy0GA43aTY7w9AwS/IwQjeSQxLhv/naQFIUVCitlrpKTEb1sfuZDqrFLdjsVCi4AZtn19V/x
kctBGlIy5Pkt7UV3GDzlsGpxU12LaG2/C5lAKz70/rF/7gcxNrmq1RIfE/FMAauw4ljoKbpgXwDQ
CReafbqm99ZehuPMJFbu61KzVxSpIVecStCMNfe6ZvP6MAZ+r53GuCc1XuXmZysjvVrhbsvZanlb
bB0sm4a201y9k5jYRRJyI8bxv4gi4cloa3xyPJC+vGvwo6oXxGShOCML/kYuaQ55J/r57ZKSwhGb
46I4LvdJvEaPiv47ml0K/ECau7XMFqxcIZWl6ZRXLRyD7Q6Uzugxq1THSgAsj4p8JRXI5SOcNzks
SjT0UBBVma4Sqo8zwTpMBQ6sUYjI1XZqIh/WaPEhg9mfBo06KKhcP9pOQObHkrskd4NZN4bm6HQq
wwn5y4RP9uY4pawjRECrUL66beAcD0++ocd52HeJyAspnApX91aKzsXJKVVwxrb4fYKnejTsYjvW
FQftPifMX4HTQX+PF+OunjUW61YsOSfsYzWR2+EoyjUhOsmTLRuMZ0v0hUd8/bFXnCT4QvYy9tRt
jJyDk6MfGRFcLzutC2HgX/skXs36qZsiKlhGtIXmqEt638wp/5LoRTx7KG1BG4g3a0QBFyRExI6o
tqn85+KyYUBos1dcBzLbKiIsA71Zo8hZPEdvEHBXsJjZ2VXoHvstkLXHS9qCl2uenJVFjwemriiy
JedRo7ZzT+tz5/ABcA3gD24RTqp4CVFWEHYaFEYZMYzHkkAH1AZU5WQtbMVUjNDPU9Q0UqfA61BU
/aspzju+eq9NW7M4KRvbgXg1zUIjbSBdws2JnNpOk7wN7tTmQqhCoQbmbXSOdQfrY6ixozbhuG8n
F1m2xqtbdKntiwcmLW+40bvd0zcNeSL+PCdQnEhRlnx06kcguruOPYWkyYdj88ViddP+amfMne60
4I5TqDTwPoakNGY6mU8cEBmkMMLSjmWKjbeqn3W3sbmCGQpqR9cDVqOYpQE3C5R+OYEA/7w/pkfZ
L1tkS6CV5dIGRHnN4X5jpu91XaDfJ4mOHOCu8EFdzQ1Aj28/934Qk3y4qUqSyXSmaMph+sGphwxH
jCwzRTF4Bzn5FA01v9M1qAEK6GwaGppTa4czsv35U56FsFHAJpqXx3q2ytiddsAis94zdEJI6kaL
wX70+3EdLB4I9Q5a2C5C7AOAK0DhhoAwOa9zh/HZZwGWZILdraNi7db290JjC7vmzz2Lrqgm70zO
KjfXcmW3nGFwrebq3xcSEP8s0E9hCm9SemibT5szPzHqU0adMCnKJrKCgPL9iXrrx7RHg6gGkFjF
xJ7N0uKnrDzPRYigX96zCECMBKADnqMZoFKOkFL65KhFvpMgQdDaygr9ZHBhfRtV0fYiXS7RiQjZ
ms8qMHdSuEUmo/PEfOC3DU12P5MedNOs6emT9X2eMlrWHj5ujzbssjXh2aPj76H6OCLk9Y5zQmeP
B/3ln2J66xtQiiKBqocXNDVZFb1Jmfi6NITdpIVopDGeSHzYFXhSmofdStw3wfmnyKPFfFw8UMIp
9EystL+loabomvievBTSe/gSb/eYcDhho79De6dX0jvxRRYQELjS9WBjNr3N/lry1fStlfIWwJ9n
SxSB49uMZPoOOofVyukCNVfm+mB9rl3+ohnB7HKrrKOZsfZz4agvR/zOK274xQuiN/5M7gPbxsTY
/mWAhJP/DGnEcczp205ox8/zUaQP0bu1mDBxeKKouQ0/7B27xIzv6b0ZL5eSlYqrTbWl1OvSl47z
BU4xoLGYao1CJoRliD525n0jhcn4L1PbZzf1ti7vfs6os+ZxDD4abIFPihTJjVtRtc2IGWM04JYQ
dU91IRCOApUQSu2FtXs5K7NkIsAO9Q1+ultG848HgtNDvwt09IFm4CwQ9WmN6uGv69w11Tw8h4gI
kAdbTLkFF8wFnS/mq7ydhuYon8nWSd5Ycc1pSBQPDnB78Z12LwKTgnCZNQtrKQ/4IvQMj0j7lXPQ
zaxplvIqirJKB6AUkxDvkBsn+ciIZMNy87C7osBpUwf+HgYJmH8gdzart0m5JcsliNT5UzIxg5ym
rHippnbPHEi2vqhD/VsES0t6lML+3Y3xTRSgLBDN9yHZHX6lfUYo7+cWMSUoipgasCzmXXZEJkAl
zIRASbcPoFUC1iYKim7iUx9L5Ut/DBtFF94oMXs8qboDpxNCIRtMMt7kLpltNrbOzOamlcUZEttf
eWnBny6p2o2PCK4T/STEId2xZfZBKa+/JChmCN9NrzNwe8m9jitWVNiGtrQLIqnULGGzfSnr58Oa
87dF2NsLH1dUKdkObWoQkGUqM8oKw7957cbApvexaLFsQM3QIy5dxtdWREHvT/RQeGummH4jt4YC
qIKMHj7rm6zO6aKscJc4GzgDSdSkgNGCr9s9UtQ3Y6Dx4NmAK90FLH1qosyOYoe/6Gosobn7H8DR
dM5XBG+eDemMIegeAKCUU1boYbzxh8jXgtNVgYHzHqlWheSqTYEQqjWuCDBYmTUnLyoWuKnjvFS/
uGB5CuyFbudwZYStNPf0XYPwWk+na76NjNY2JGJsbWc/hV9LucgxgTP4nqsNO0IyeG8Gr/AzI3Mj
EUcDOaQpN64A1ESzQPD5EA0VmwQnpj5U3vFRbr+8A4EmL5LXyBuv/X2WcHOSYP2zcrERjLtLsyvD
niaD1Pz0ySIVCU5xVGphg8vMLZHt9edhR+L2Pql2RO7Wj8Lkj7ZkkbB4DalId4+HQoVirXRG+z/I
m9LIsP8xqSkzOG6gNeBKu3iAEJbBFldBeV3PVktpP+z6L9lqYKBqa7wvWiw7n2ja93+Lo498dFAb
nbP0rCXzSjl4kBMVBixSObi0aaHopQmxlL4ZELEMqft2ezTeArncct53e9xJ2XyiTkrIV+XGlZkR
bhJ4ChkNrKfqLMrC2w0QrJspUdPLUDwaw8sY/4mntT2afa4D0k0qcb6jOYu3SD0oOZzU6DFs6Ks7
aPRTnKS816YZJjIqWZAWBNkt2jYYGL93CMGg/3ItXbQjUB2eeK7GNc8S1Pc9twf4+haKg0HWzpnI
3O/0MfIqOHs4tL+c1+SpMa10jozAFGyQ6aza8y7G6iQ97JMcdR28IYL2YNO9sq/iMp3p1Syy8C32
16NvX2UTyKy1fSEOi4HAaHGmJsOjU+czYL3b19X6C9S0AC5zeDqCqIktNQD0W4VaOJ+X2kKTLmj5
BFs6aoKK+8hxkiSELGrBJrUktRQJZVG+6rZhOnVprejMZfAYYjtGhABR0E5cAbkc+maRfBEHaV8R
GJvE/ZgvDI9ofBhCipymVpuUzxWLjdXFq65YSHd7W9Y8AK9GzgxNPBqL9+77az7DJ/rPpQpkvw+q
XcaI0hVH2ou7IZyVU2qJOQZLCQpBT++cYIxlzmpBbhKiONq3CG9RymWGc7Fg6R9pPhcgdbywn0/U
LBNWHOdJ20jSrKXGhSP+bqp8NAqYJ+xBvlFqt2Nd+MAdZPo63fgZmwdbYkAfHWbcfnxUDt/4RrZf
XetVDr0TwbbmUuDty7tLIljAepjgCdiK+gvUCog965DANftL3ydnV9dN7+LtHv3TlOxNY0/PC6iU
kZn/POzkX+nVgIvtWxKx0pyTy9zSi49xTLlXxz/lM/sOx2Gf3Smg37RiPusxqllTzaOCgckhjuEU
sw8fuzzdsWCDlXAulPzbO+ExxeTVcIyI2tTn3h0horvCheJJ3+dl7Gil8MGDB7Eu0cgx0BnWmSNr
mFwMEqsa2HeBnnsh20s1rAHuIffjKt4zfX0h2KyABXX+8J7OEfj5xtRdezHNASeKMT3133/pTGXU
ehQreiYMrthR6GnsArb92UTTzVuJkqMnKs71xaHX/vgjh4iTAoZfCZvBSclLFv6EDsjAGkPCM8Sj
tqmF9mqICmSwSmokMwEo6Iczzpab3TRVq5FTmUcSOn2+EgGxzIPbkgkAzK5SiohPxjNdVQJkhvx4
cP1IQqAx70HbJNmGHzNo51glUunvM+mnUeP0yCXODypCLwVMCiiNYAga/0r2r9Yw+07Uz5jDpxfD
8Dt7GHalhHDmT5Iy97TPVyeAaG9KTTE7jh7ocBGrp1GD3D203N9dIzBoQl0BfilOLEa7rGChee+C
38r7svL0qZfjsyB2bmLI3n5OHIWIJKZ8yi+9be1qgC+xghK+qamvKtib291yG0yWhOFxD9CZFns8
8FNwgRr6KPicWGFjdAUy8PS36pPAyrB4bQN0pHci7EUqD8fvVWh9bvMpp+m/PinCXoGBhPg0JN+C
MtqbgouDi5qrJ5JE7QXvWWoxMd43h9Ya0V1/hBhEl4Z1CARDAPeQ3KB0m6O/fvZcambRYMh2o2PG
yTbdwDXT5ahjg6F42oid2T6W0V8oVhHwVU/vQeUuV6H9dWoTWxATLPC3FYDpVz2B5sYr6xe4bHXa
12JvPdu3UQI4XEem5Xv4rpBOvYHlQjJ3pPQDKK4f3NLbx61TYIeJhuzKG4qjw+a9+b9YSTfxi/qD
CzEKt1m5jqUS7ByXmXwk9GWNDTqcFQvxwTfVCcrCjTNHOfdrI2JGf+WlVtLHvTg7CUTWbnJS0jv4
thEi//Jhbg+C6ZAgVONqr1EjcsVnUehBdHWJ1px0Tx3B2Zo7vfcc/b/hDc/rE+FTGu2pF7WdUr4I
lOOfoISntuSAGqMAAZnV3D3JpdGAWsrWLoeTlJ+5ScNn4KBEqUfojQ1B7I+xuF5pTAK4Ltrt+UZg
pvfbyONP0fxc4no6Ud59lhpxO6ogIz45Y7a0delNsYTVK7crJPneL5TYrYJo76hgsnV/PGy13lt6
ctH5uKwD1iVM5AVoN2BJVeVWfge1CpI/RZkOXzsvrjBvYzvP/RqhEKVYDOn5aXu6qAkDyVLB5tGD
FBoK/7rS/vkmhSAJQ82sfkJCwYLUxokK5oPXO+tGLsj2Z3p0Xv/8O0qeJrKEjtmhKRujeaFSJFn+
VL5kLmCf9Q0wG8/f+aH58JFO8dNmyc2Io3kQ1B/A9XSYy5kUF6k4IDXcqm/asnh4huudNblLxBRo
IPPG8uq5CeP8EqN0mwhd2V8NXRjB+FflnYD30alXJ13U53sIlGX2yYBDO8tR3WwBOz0Q78EMjBhL
sj6HxJot0b3M31ZsDYVJut4ZGYY+gsvJKlr5t18UsK3Da4MavkjuwFx6ewvTTV5b5khIKB0uQtCx
U0GaO4L2B7iuBWrgEhQxiU9UnlEPlWLgVHie0HQpyW7qkfrJC5kSmVJl5ggpwnQ29uomqQ4PBUbe
vJSdO9NejtBoLUHKFjM17Qiq24/4I8YxYhWmM2QsVDJIxaVg3+jxxH9A56UkHMzcF5mc1LhvmTD9
sxHgCLkBErbl8eleBC4yu2E5Vi/yXe0b9EIu3gUvstr1WV0AZa1QvwA5QD5Vq//r8PqW28r8lr/N
ATzn6BUvb1eBc3StAJiTKVJynHuHnMe2CKm7PCgGgWNXx0EHlb4nzurzv+5dLnSXFUO+m6/VINaY
keYUCw4mZnL6rsBbR0JNhCZYuq1Q1Or8dLTZCt8ux1DkgtBFtr2e4yPnn+7fqPncRsTMnggGg9ph
OMKAOevKNn+WREUPidaM1XTOL763b+P6PG8xfIUjulATT5LjDK5/jmKFw6cesUu7xJN3dQpUYykf
W4Xmx3/y+gi/jWqYkva9yWpDXFUt4on+RgIA7vQJgXCqZVWrvdjiQsKf8Ky/D/3WmRO5HDjK7LyJ
8Ltb51AZJcydeLaxzCGJqFkx1MOG5Q1wU3vV5S0X+ixMGq9M6jIX4a0g/8CNeZo2Jyiho4NaKF1E
e0odgNjaMifOKNNgUnDfJBcFvEcUs2eHaqOhF6s9nyfAqJ6O9xJIC27s9R0P8bmS59StaSVI13TZ
INBK9e0XLR/0oV0Jj3Ht5IZFixJsTaONBH0trmxxWNn4HCzqHfT+c1J4w66SAMYKXbwLU+eao/i2
AVRI6SGUw46E7c6oXpvhznPtNBzYwfLT7PnWk9WGEsACl7XOKTaURvpmo6nuDKPV4SE5DuX6HXk5
xQTyzMn9JISlfDc4Yg+rpWc95l3BfVXloj4RBRUV2bV1tMJDUvfCV+g6tOBrw2sj2B9P/0BmNlZx
im51bZp7dpmeJf04KZ4z3EzN0h0JmHexFC2hNmKWlVNCep/NPD1AS1R41kGWnftc3GIhPpepGYg4
mkHaKWxEmzzGGe9I8jNuDb5QZtEiiwEcRRM0m4Y4Ur/tBgt61VpPq4MVCNhYUPvB6DHcbGFFm2XK
y0/imLvx67yOZaOH5tij+u5dOqkEKNtc6N0ISFrFDHpSg9/YxOQDRGRcISw4oJq4bTNv88KrRJzI
4FAkM08CrMRblVM3STl5x7jEJoim2w4PhQAE1q+cXBPC7yYfYpUR6dGOIl5fuGbitP27TaLlwXiq
eSUQzWaNMFcbEeC7AdlzlMhvpJpn+DZjMu13rlrg3TRJKzExPhMKOUm/n16Brez+Y91p8HBAGG7v
5Ja9o1iCyYN9M8vontBGZW0/bB7WEmcvJwCr+34OJR+K58IWnoM/KWMKtFX54QSE186lUf9dYw9J
ukSVQwAqRg6TZ4ztPoADnh6XCLYm9lkBdwP3QiRzwd4adjw/ye9B3TGPxe/bmKzt1BRo6b7W3UPF
yTwL/srDBwFUeBCLabmtwp1vB1z5RKFQ1vSM8bAO8iRJ3+ZmZnO+fqffgioNIEGOGDIHbYhCPVSA
KMWFmcnbG8HsIuazx7oIbNnbZ2TI6CpxlAWss1MwC1ulGHzWlKvSz9X8UH4kbHOPaVUJhq5ilSxj
s6yqMvZaDI1hltVq2s18Ui7aJP65Q6Bhut7+eoOak/x9Gs22bDujh4n2h0cTvKlTJKXMhXU9spfL
itr4Qp3mUFzuM5tQVqnXENUKlSV0YGCW6nbNEW1X1NbYtmIomnVkpQR++1ucFdL1kX2ExqEbZUVh
r2rOJYSPU5vPkqfGF4hfsVJG/Kot2oA18Km3Ov4+xbzxsU4TExlRdpHMPbvQEFEIhQjeu5YnUZVG
9bB9aglD6W5RHLtNF6YDu8jhAyK/r4+haWUvCGsoYSWgUleGcy3SxblmK6CRpgisj1xozIhuAYL3
F8DTxixoeNKA+uARbQ2FjKDuHNjkbCc3ntI0TSrEoOHtIMiXN+nOge1w+6+FAnbafmQ9yNVHTmY1
FdlRTQ+cu4I7gig+7C5S35CNI7otpIjcM0X+5/r52K+ObtBtlG11lhCiaoP4UFfqmQOKiAurmAT5
TRF0Cs02GZnLGicTNIatHHw9+jqW6hoFp+zu0NY8eWEATqVAUIiI3V8vVKZcILlhNBNdxMwzpVRr
SGwIOMBd6HwL9drA1BU9b/MwDQUTi/nS0gBsCybcj7zVkWEfueXa6feI8vNLUvK5dyzqnsYtHQJA
9BjiN9xsz2YEBR38Eqc2zk3hDWfj9/sGeV7575EJtEh6MVDv5B7b9vU4WAOZxPiOXfW7xvVlpSgw
EJucZ65KcIcZutrBUWAT2DcQFFOvWI7gN7m9X9+E4ZPbne9t0GLoWw5eoOrM8x2za8EOAD0T1HCp
aYLrXCdz0mVzvUJ/Shb22Gmj3ePC5CxyDJ9G2nGGRf43WIS9ar6p5oIWm8H4eO56s+xRVPAtuY7N
cA2AiFbt/gYhsRbGfQbUDQ17qlQ2GYsxn6xDc8pcDvOen9cqDygT28nYeKu/5JwykSs8hY925YBV
dAHMcEjs7IV4V258XyS1Ri3Zs+KOwCjIqXwn73odc9fFfkVSSNh01Aci9LrGAcA3GGvQ1+OkFnge
OsZGEgNW3rjS6nklr21XEAgOlCjIEm7o0JOHZY9sa3pe/LhZSPJPWK7lKQco0Q5E3Tdcfcrmqxpz
ssoZZeSPgpWnNEzH96mAkkd0fnaIHUNG5RV7NDuWSFQI+q2EDgMtgjTgBZBmLXX2QlLkoBTOH5fR
jWpnDJ12jt66tNKu1pogGQjU0Ub37+Al+gzySVdwMr9NXFTFOhasWqx5GTyQVws+MG8p7wDyeyka
YutS8WbpBkEe3CMFgi7gVQJunSRlfz8r3vg4tC6bergt8meqbVtK6YkaQ6+fOWTVgdlcGRZVdTHC
pJp3MAg1sA96DxAbOSxpXxhpRlcGMTxL2H2Dg5EX9QpQjaVqxnE8M3Ilok/xQLxnHKc0JYiQOyOj
vrse9oLBWAHLht79STuVsLBJDhYizGJrEr18mn/FNDn5sbr+FMBsPO9x7DVN7Iwo3cBlnhZa5z0l
F8pDVXMTokAw/SGpmL2LaxmyJ2tg/neccty4ooACXaULzNFef8p1QX5yd4GV09UGYtQMy2WUmN8H
urQe2QJEtXTYGhtDog32kUCPW8zHu0aychB4CJrcgDu+yHbogKGS/Os5daSxPCs5S91tqcl7qczn
RRDtFd4ZLbKMqQHNiDDJQz0rJJX9Zk8wBApm0vLZ+z/vKTPWUBOacoXZ2bKCX4FxIY1epLxcatoL
SclsLttGUcgPdF7wsJWmPnG+fXzCmmeecrrUPfUp6p+XYhxibrRf+sT57ck82WoGMtQFCnxaeW8s
jBznO5PmqmmXeqTiyTfpkvzMv3ETxYnKD+pEvhZIFDMNcY1m22Ck+4WgKYtmzOglsI+tydhMDnjv
hi9JRtnY0s48QyExHoLYkS0kUFbPbDhYO+P2Q9WFqfKITz1WaUxX0nGOiK9YLFSnFqt5H/bssU4d
6zRhGobPhYFUom1a1dfKxm3EialKa0A99GczDZNccsgJqn2twWmfAL3AaU/XeEdeUd/gm3D+i0fE
XJ4MDkQrh6lDrQlDAdE+Pc6G46gvrLg+6Z5TeQqE3qyzvzSuLGC6awvwVlYjSsXZoFAMf8MjwYq9
pzomrUtNmMitqa2qalg20OTVXgRakCg0giUq04cZQL3CejB5lqhSbDW7X6UtuX1KxWjhLXuCiUKp
Y+V4OvP+y0C1tyipqSiYh0i+Mv2VTEYnP/mhaFNEhqjChIG9Lfvq0bd8q4C4fDF2NHJIX2n1j6TK
9suQLVSHfy1nI50g6TSDQ4bJcA0ekNiwUz07Io88MmqEG0jaBVSuHp46NCiyJgOw8AM0HphO5mtl
UIt/moAQk+oZIVKOHvDeAClp0I9wRh8wWlbr8P6X1Aqkg9btSpc1rSq590UhyFEEu0e9RpMfbHLN
q25MOyf0QmU+YT93aZar2DJB2nC1i2YEveEXwo80djc6YPfUqIs3J5pynK7CO3fUS1IGRwN3TH/j
1EOw9uMGCmXRUXh/Lmzk/XZppZ4a9B9SUJgRqHgWVrbeA+CG+xF+xvXDdetXOK+1dgHqX/qKls/1
J+To8adCnNXLStnmTrd38hsQe4g0xGp7Jtn3R9RK9o+Nwj9uQl/6u6Q2Ykmh42pjeyEfEr7jiufu
+uDzcY8WNCTci8d7mNTIGRYHYTGEt4qd4YnAVrpNLhNeVIshURsqM5NDfsxc5BuwcMJGrVrwkZIx
QYl8BkHffbTGMTBssn4cEmICFFTJXx/6iUkHOA2xwnzF73I8lf224EKVvrudGS1vy/XhmxeYE5V6
nSTGj37uVSXxt9OzCOEfQumbCOI4ZYim7pw4rTZOLyAZTv9cOffz9P1OGkw9smrz9o1y/wNXHAtS
4K7dW8S4raaZ6j/jxutAvZNTKxJjA5ea8pUXdeHfIy1eX18gWNJ0BNmEAumNWDE4GVrMFbZ6/NGU
l0w0uVj0erWa6qXXN9z/tOgP8qLjjry1RXGb8+CYIf37cVt47Y4PuF89FpUKTyfdgzV/uJExDpyN
P4RyFCVTRDiUKI/iwFzVtVtKcjJt46ujbGQBmN7euAEkY4dVAnD/enq9RVBWwKmRn07sF1q1BysP
rrm4R0QkU3Inm6xwo/5P2lsrfG+yslgFVq6SmRN8yFKV2fR+SjAL470PmkOrwEYN02ItnGcOiD0C
6yZJahhnZ5P6EiAe7GuDy3fhlBB2Aj5H/7Ahirm+CUYxOD+Nq+L083SMfs+w9b7vrKRqbqppmYUs
CM7VPXgQvAaL2/SeiaQTLZhIMUlAfuww8nwrCSRo/jOIzMduaO9ruImXcUwDDUMiwyFL4FZ85Zws
LETVEyiNSDQ44PKScreLMYXYQ89VoEeTg3kyAvRob9hqhTByQfAyyhQQI9bEsJmK66BZeK+U4nPf
hQTaGb2ziKwrgSduFSffRX9ikjjCPn8W5M41k/fGQXPzoH0TnF7z7fik8Mq8vuYlefUpqctdufBy
MB4ltAjFfUHcff2WdM8TBO+G4jN2RmNRrr2DB1RuR/bJbs4szCQwKCOcIsOo9KwMEdpon50cHSLz
gvDjasCod0cLPrrtPODNtw147ZESowE3nRjbDl2sqvDOJbeYLSByAZ0/CHo5CAWhaev983MVd+IA
+dHm/3xskIsC6WgKPvLq8JaatkNKnktc3XpHLoljQbm1qAO2MRq3sweVnvU8hT4P11R1O1X7/Q9j
zNb43sMLznlsVBgAhyYD2ZuVpAzdw1raPobblNErlbIu87C1AWJifBs6EoFPdiBGnaByxdL/A600
kAU6dL7RtNwp5rXWDAQVG1HKFat0OxfNWf/ERQ0TuBSRjhXf1mDuKkwbrM3E2sqwqURi9MRvuYZq
hEtRe1eOy+GsL7m4Rd4dAio5Ilj9G9wpZ3pjYUCptdPpizqiQN2g14cI4UIMIIUdMRcegmupcu4j
hwg/PG6SbPDNyjZ1WnL14OnVxVP0rK/ER/sUiSI8yEkVLHBJvVfOweA70eQY6xUy+4tjnZkj0zeX
R2GQfWuguLHqk83F47LCdAgKJUdfMdWBCIFM0l0RZZoZrYKCu5gatwDxfIDa+2zkLh6bx08y/l+h
vrbvAF5eyQ/vx2CoomfI3nibmaD/mHncsj6y/0JRfrx26XNTtiSlAuWmwTYd0H+mrBlF2hlFjjR4
TR0GIcbpSijuwr4fzcVbr5UPJ21aVbUOwQwK90ry+M5mFQzY3dP6cWKaJiVilYCF4nCe0SAh50tA
oHaqcBMRe/FqREVkydfoLOieD7pwOR3Y7TNAYku5uCn3dxG2SW8ZdNc1u0V0U2c/rtAmnu2p797P
D6++8LPfG4dkpAC2VV1vL+Is5kJ3ZokIkBoJEeSqFsMJGn2aUehW3rANgHscL+cg9cKfS2r5ruPg
WCPkstyqekNd7hlx9t042YExgrqltcrd8GAVMULvfEF4TgLnRY9pBmhpZYgztLHW6SrDNTYX+HVu
lAtqePkLyjIpdo/NXcmvC2bvZk5iWqWOEP1J1pbeDv51sAU2hgDPos19IbiC/o3Qs9teXltcPspy
ReE/v23mnO6ALOmlQYOs/CCyjeGN2hFz1+B05FlB/KKjEu5ZWs5R6q4b8l13CXqjvMP207hKqVRo
xDVLprE87oxDq+jBtoT2c1WktS3TfY9FRRma9beoTEnH9zehBXxb5AXq9k7RkprnXOg14Jg3mo+Q
Y8S5S0yq3cR/C4Yxit1eDf2t+Xj/fv/GbuVs7B9CVMVrPegsvCXBkhTgxbfyr2rWpNs8zm5NMPQU
4MFfDfVs1j8R9EyxuGxPMarv9VI3dzvUutNxqSSOIkRah188LsAhqDteaZ5KKF9LxAN5g8cYKI1X
qtB21fb0NdmWpdGe5JZ2JqGxHGR5tos2wLzv8U+Ds2zp4ZkN4d6mgm1sYOit0AbObK+q33XjwhZ1
qDpiDMvzOG8IqTyJTWfkTTxzOQkYoswuClvckn7J3neFNFu8kxHhqHDt6MG38q9s/J5fZH95P9ni
ebpTOw0ZWs7ycFnvXVoi7sBKaOrhTKaYd5YTmdgvyGM7ObSjdU6NH5hde0hXODB23guNDJEBjK24
OuY1PcoQEh/gY5iNIB6p743Uk9YY1WeRgJXbcu31QBuFUy/0EIdfg+/rlv/YAft7B74QdTLX9ZU9
dMrZMf4zrXH3eRN3HyaYDpkykAJo+ssVoUOa7xa1ywKIVESyVyL1MQaGiLGb6+vIuUENjp/k3FlD
0+S/CBaTjgSDliWtibEHTslrgyZbctiULJ87W4YB83VN0w8m72bSpvg8n5CJtqVbnyOrvkscEAi1
fkdHPB2Oxm+roVvm2G9SiVq8RJngv3/93W3j5WzNF5gRNWFZijR0vjCaSmu4lkB8l54yDsMhbFk1
XJRZnrYn2pbliuNQqLXztC4n7/ZJfMpt3uRiEY2nV22KZDnpJ7o8UKIm6vVdFKiqWDzL0a4zvPP3
fFB3PN5egwM2P3gQP8imhU61v4ucPjZbpvX+y7B1PFapUnl3TRf0MNouVAhQkzZ+l47YtLUvgv/f
J99JB3hc6WWDbTHxCnkXDaDvA7oF1XaUpoc6hROCqGAqywYq5xkJlP7GDlscwhOOVAvvkfFUzSlw
nYezrGx1LoRFrHA6psQlStoAYlRs+PxpZNZgDtmrE0vonwMhPF9URUapxn8urhZ1uY6cDsC6jpRT
3zK8ZnuHWNXOzc+wPeMB8YFP98LOiAvuzXDIeJLqA9fuhWBvr60cQbWvmVZbEI0neJrF1rvy9hz0
GOErXp0u3wjwvblnfKj5qENvc8+ZZTIOGo2BBRvLUwEgDESPc10FlJkh3rBTIJXQx+X6j0xA6foC
9kPljy9JJ2jR5Doj1ejp7bm5w+d5fCzVwsO4192m+ySqxpFu6ydfnzUb47W7ivikHYNLVkoteVyF
ZkAUO9g6wMtWeFy4ZeCOEyadERQTYP4cvh5MCvakOSLNYjj/7DY0mTdj11Z1gkaoMzmw2QjyQ6Py
Ob4B0z2kd8Uh8bFKJstKYlliOkgjSW0qQkbjwKr02mNwLKfNfrg+hyuDsSLGBGYneU3eEV2jn9dl
F9s10sXbvDUCvCpwroUc4X/mbnhVcS2yujNP7ugg++nLUwW/4dTl5RXMbgtc2kt67GFDR30V0j0t
yxn6C03semrVZKeSpEYil6oED/ehczBnNUoB6Cx9wyl/uW9jPaKpmgUK/2oKBaKeHjBfuCVA2vYy
aHo+oIu1jroA3OOTQ/ekwnO9PflJr9Vi+YjWtl5cUifaDBBsG++Dp56d+T+7PgyCAFLR06a1gsxG
vLq83MMxX5Ge8iYZ74/ytiVa6th5ixbNOo7Me2PL46ryCqml5FBjOQKiqBtdrmONe3sJDYrJiah6
YqccBuKCsxBbkOER+o4t4sMto8ej86sFpmy5MNP1uVNckHci8xp3AkkUFQmCfq5vOemMgv0k1wlQ
0XGlOivswBb+sa7nVJcCfzXk5o5tMuzrzB1PWiwPvt7qwP8v00DLsCs0M2Rh/DK9msYBI3vXtxfm
UyZmmKKPu5GHzIJRRj/jdeNdeRSv3qw2WRBWIrbaU/oEUm4YGQtM6iD8TbYDVaq6p3el3twoAGXU
Q4nknjd5bBs2/CAvtp2viokOx6YiYbBfJhL75ln1UEOtdQlgvMfTDX6K80drm0aH3Kj9Fa8Vqcc+
y5L3+Qqrenc38ZWwQz+jLUz+hKfi6ESL2slenc4Jm9E2VNgQnx037Rjr2bwvKm/2uz1I34+ayOZH
ML17OuGDeojuB/zteo6IS0okAczmVSj7jLzjkp+/xQmEENn5pxBQuqFBH97qq8zLXPM4QRO4ziND
dc9B//lmiJ9oa1SH0oJTOj57an8nPJVCmkeOLxpTpfgsx5RQXaLIWAFBC2R3Hqnlu90sFMPgmGfX
CeYjDvoDv5OeFaxrG7nWD0v0JMfH8wFB1XzUkE9yLsXP8wvzvISbfwWolAfwd8kiDDwTUG760DL4
eTv5dZyJbGAYjKdsl3xLLFJe4kq91YHNjVQWto3jS50ivTRzQs0xO9RMJKYmlyRAtWrA9hzkdQxX
cdaTOctHlpJdwqKuBmDMbLfbNNH/TTjgCcvoYkqN1QSmPnppp/OJcQQXApOety61sefrPGkTtrZP
ZV1vaV1Cs/YnjaaV6lsgnhMuaTDAo2QZS1VV5ootj23vz76/EBAQrGl//MANEc7hbmS4EYiBvD8c
WfhKr78mBC6DBYnWufrbNYWIsDQJj+PgXcHJqL8SInsGIsccivRjWVDLzoQ4xPMQar7rY21OuLr8
iWje1xuWTpzwMx8xOKuirs+dhU/qkg1CSIqeWcN9QgTKEXumCX6ir0kyStsElQnHGSCqmSXqGLTm
TtHVjTnSr0XgpWR3F3rpADiovUg/1dGiDqVKdVE8iK7693SdlhNFlkrxjyITAADC6VhQUO5/KZmK
0XCtx1tnvAXSDTLj4RGwFku6GswRmatzy0xzI6kLR+ZIPqV22E/xIBtw5KMH+0kEsHrtwPVFGwl0
BYUz8flkVwwhvUBDvCy9lB+sPcQGd/yi+sEDGsxYGWH047TrvVU3DGQNvpuPH8GN0EIotQFo5Yh8
gxzyW6EdbMESVR5nsGj6LIMNgIjeXBmzf2ByV0HyIblyIGVaUCqy4VYw5Y/OSfEqXolDxxo8TkU6
OUIwD6r1m3OrMMleOnVTmBD66jNnKRew4O/s3YeRAsozbV/kAZxjkUwsdMbAS7CMz8GXOu/Sixq8
cY3mAwr+vppBEIphoq2qpj923NaV8giSUh1V3E4sWtawj/zn9+5AdNCJNJ+iCLKVh8vSafPFGXmO
03zhLaEBejk/EDzXrEvb255Df+uFg1GZsiCmGjRTMW2fkpJRfrCH7i5H6nutQ0xeUtuRCQo1UL6i
mM1yXHoXexkl5HOUEzJ/QTREKYm7d/QwkUVOBWLC5RDTEERQxFpfdMRQSG+lcYLakG3nFYQWGsij
kEZZqwU8t2NKRZ5DQWALfWjHhYgK/bctBXCtI+JxClXVnPvBoKE3QwDZenRe3eqgSFVltFG85PmC
EzqE2fiPoUA6lteP6NMnP5Q7HBvJJrtbHaQLJzzTTF32r/e+7HcHP4eVrwAcXNbGtOxZJH4WRVvb
+NWnQtF3aujpHPFTNWQqEMhce1yeAHHHtTTrAQI3umCqsoXpicjEFENdrtYfkIBgfvZwyiWJAf5e
5bz9R0rb3R5OrLtxk9kVZFY9Pj6M4cLkAQ3pW+FhqTnNU5uSGNGhKaHkl6vpteIuBNUqWL5BPCqv
RmprpfhQEM/wjOCR7Dgxc7dmrr3y+PVAtYvrbmMu0BMMCsmHtRY6qKJVDhm+hQa4Pu575y4ISnR7
pVsiXgkm/i9BzrLgOGbdzPelNE3lWSv/AryMCFHl+Sj5H+ATrEtxtmlwqVhg1XDX1u6vPET2ZGnd
lzR5cFl41lAjEUB1Qhqowg+TZQKAmwrblEj9qq4hV2MkjN1bVQMvQTHDqboJHwYyvh9JOLuIjqoo
S3igVJcx85KXfKyKv2ivM6SOH43raFttL1lOzkUin+M62hO65kzD7Epbp/gidzPSlOWXPPjOuUgz
5QsIDXKx0bDN4BM9sHJL+InlvqpQ4jmJaPHuC3a36O0TD5DvyOh8lyWJapaas/BCDfdlm0pwKESU
/iheXwP76EvIHxKqPocNKb19q1c8vfGNOaalVIfuxhtCWJqcxT11+MKWjAy+GJjK2l/Y0vw32/yM
iRG1otP7V/uT7vPqJ6zGUB1D0hURjH6P7CqXgkLGrh1myo/y1x7CdnzCsHSm/EJGYsz1rlks7dcE
l1y8GyOdidJYYMnPGSErnrB7odWxuuxYSeGHowrIw14mpMt/b1fbImjuPKCLh+p9bmTX/6kc4nrU
+oZl7LXFnueQWxm3zpaa2KnhUn5MJIkRSWWC0hHIIj7HQ26n7bK7xKvoD+aobfiGsedLXlhfeSIm
XGv1tNcMNd7dTVw8LWe78lCWat8K3tk6/4TXeDgygOFU14AQlxS8zXHMHuX0k3jgnjx5nD1RhG9y
zz9iN2KvTCCfN0AqLVwOBLC75Q8aJvOPJrrygp+XDumTmrav+QJ4C6xbt8PYbTfe2XIuBlAZgowI
VOCkL9+IERyVzIJISTPXqRWOgBrJFJVUutPMgBS5CwW0sPZkKJTMoJWdZEFs/QVjVBlSPnvKrQMd
bFLI3HgVckGh24SdZ7xCGHBMD7uUPlgUDjnPdbcvmJXrBv10phdqDopqPPNt0mbhQg/mhzpi0k5T
ykyi9UhDGkw55X0/9DPan1vDpBFF/pBtOZ7clEAdrwzZ3KGSzjZMo/5GcO0nbvoPA89eR56rrfJ8
8yUfdwsSlcfU4KWcL0aJnyrQ2BLSQtLLaBsdorWFCqOpgALi/ohH/Amk8R1Ud0qyeojwIJi/8Rhn
fmW/oBGfiu++xOvaNU85KuAGgBNZGrPY/AJ0ctrI6FkV8VwLxBQHPhbYrW8hdNG2iO7jj/vbfV7m
G+H7++quh/NNRBWAH9z/Ek8i9O7XYtMqbpL8f9G3hJyUzhNNK6HvY9N52jp0ZCs88C+ZQnvQhWsG
U8U1H1wrquQMZ8ixHuh+m7Qy1eSDAu8lDUyBZbr3WHnH7KhxFNok1jBwB7mpaYnghGcSGg46vBgf
G0dkm4QYS4lkBqyN3mreja/9NG8zKVbcGzmISATMIG4ZWPitIm8EpKSBLQZqzMltK1qjnmXWCw/3
JK77CEwNO0LujWtwGCEOq6a17TtLfRmpN9LbawNTBGS1avrIjC1d2muQrgH4h3fW9kBf7Iyy3x0W
m8YSB6EuOsqWp8IGJWQ+hCaH8BhjAmxZEkDF3awv/BhZaT2LhBA15y17WWQHv1S2H8vaAQ0hTisP
FlEW0zaXouJsNnSE0lRSAezXUwkneTT7teeGs3JQFZIZVyVG30W0xglpSlr5/ohoX6UOSAkacL3X
VkpjfxNaBz9WObexRyR9o7I5SVzPylKDxMxjjtfLRh7We3G9bD+OM2f0JSdnD5lYRzkH6V5oxBG+
jozkjQcStvpI6sHmctWl9G4f1GGnwuvJ4Kmj6nWwZvYdXCVlJWQxjBX59brkFDVfXltrrqbxRiXx
BmY4RRwMHNeRLs4lqavtXe8c7oAV2mOCVGRVnA2gG9K2/EIb1zJDIbjP/YYoUxBMR349x+eOkJJJ
F8U8gAb/hWfrJJVDr4zx3MLU/LCdJsfSASATXCy3CspmMXdBQqPgm3Fkl2FHeiEFIE0mQFrcMufH
kzlYk8oC4/KIP4zAUFm7qEQm/nihUy0Cu+dQ6xRBsHhvmikr9DCvqIL+Ro5c83VjyBhWi9zBFGWl
hSmoDojAKY681YbTEdh1ypUmEXJ6IottipaxVChIp2iiHCQbTVGSYhwwNDji4LZ/A3/V2WVYu2iz
TAla7WfFSn09J5hUVhcHovBOM1AMy0I3z4i66Jma2eHuH99CtXtufu1D6X5UM1D5kkNWIK9rwCNM
XI6k7N+mo0u2lbWpnCLX3TvHpHzvCdJWi4yNKBNVuYLONC8o3ZWkKk5k7uT8zMfyxsvUvo9MFy4I
55cxudtBW02z5oPvrmT3qGk4odaq1xXqV2UaILOS67PI4LlarTb8hsspPJgrQk24uzH1HTtZp8jc
CMH+zLLYJ0fR3bFTQJg2YKyD/zKofoEPoBZ6oa171zebt0vJYsGfyQOTLfyI4oFaPGxsJ7rHdyBX
DLthiAsCauSzTZNirUFo1FgrnEAGv1wyNVpF+5A3jQ5wwLhlCfXXrt8e3oWJFQNMregTdmKeDgu0
VBNlAYp+MnBZTmf85eOvX4Q4X9FSDdyQccw3MFemzjsBz1B4tL34Bo+RSwRYj+JKEdcFHQLzKHGd
YqBeMfV40gGSXyz0OdV7N4iT/gQeA378kYO67ydnK733R4Qf3IRp6GhOqVhwyckBbiFq/9DuV8zS
z1weuWy4dOv8WLg3cnw4QWj2RWeEnj2QLs9ce+cuNobj8610XvZsg4s5xR1u2cnZWDFIXZSRLcQY
tiVSmkquRTLjIoZRkBshGSN0H7pzYLcc7H85+JlnvEV8Uw8JjwZeK73WWQWH5gVTRGqJbCXulzl1
FvZ0TXG2C0fb1n+CJuaWB/IODhXLlB3fEM4Of6CEqeHh16itGcAro3KNHStWh4/7qRu0Z8ngOz1Y
5SSflIfwRpUXg5rPbaiVMoM2RDRskdtyKLCPt74EZtKzFaiWCF7RNTnnuktdDpggFlvi2+Mkfjqb
Xb4w203c3rJn7VRp2XSwObkxRypD7bilF6V3SkOj7XQEuHMJZRGHZIXfzIhC4RIFg1gBH5rq9ZtQ
DhQzwaQKwlxaMm/uV2vVsw+C5oxT0rpvTzociCasRSuLTfhYbyRNkTwf1rOkq63Nsu6uzPP+LTXO
fbeF+Gh1scRpEgdNbQs0yDJ1kgWRLquh+LGemviSteRab+sSRYWqVB+0EkQSeLkARa5WaqPKDnFf
AIAHYrKKfJvxrgA5qNb3xl1Ezblre1Zocy5JP1HXlReJtE52v+Sciu+liT+1kWC8ie25G5mGTzZP
OV6lQo0X8BflOTBgqCTaGD2A88l/jWcwsxROGmPvhNsGJENI8lFoe7IPpE8Ply8+IVhoLIsKMTxa
Jz6j5ePynXIg91YOIBBNY2L4t23fAnKWi3omCKZqj2KixohAWnhwSYOjSETOYyQ1pH+p2Cv9B3Es
wB6JOjEqU1WRh5aNbR319V17uRyOkprIJOede5j0AGBtNONMjoah04RnTmOMpwoR+RBg9KlVW4wU
t8e8XjQrjsbPz7lwPk0pYQzPa4NiBjy1I3THHvcGiORZYMJs2rGDTl2yXKoM75Fv2zpKH2YvKdAI
rhCEJuFQWqbZV57c+/3zlKq2b3kA2PF4r1roEYFqNM3Smp9qjCLGujD7CaXzd3nAt5ezgLw9kA98
sjUyWpSm2tY0GWHC3jZllpPIYXQ72Bdp+T9dTNuwN28yAinOVQQ0lHul/mvB74ZoMGx2gyyAvFT4
dcQ6z2PpPj/+zljyJnPkIyvYpKrHZfgQdVUNtbNcxlJiVkYyHbnPVpPXK4ddjvXC2EpiobKadhRh
5OAn+Mm5B7SqW8hajM9ixUPhVqFWUnasZztwzg6VMIKnpP92YzRST4j1FrFe8EpF2Z3rYPyN5Ko3
+MBFNWJJlxnWeI1/lAypGaOItibL9dxG2vUHnO5OD5830ZhMbjp0e9nTJMAgjMFjMh7BK3iZ8GeO
RxePjzQGKytY2M7QArYzhyGqW/+dd3k5ZBViMuQZnJx4gKGYJ5g2Vqw8SwH8Id3gcyqA2O7LmVYE
XgNlqRR2SfKyNYU+plOklXY5bOMViLD1ZSbJU1px8o3n5V/Tc3967k18WEaA6r6hyp/3Muwk6gry
GERK8pq1RDQmHm9AB6sZQuZVl/1b6dNEYI4XCKEgXFFrHIRvhXLtp9ozeSSIQMNJBGcSCeejkbHi
45vulGT4hVRn1zo4EN7cGgqR9kviL8URZV1IBM03fpeNTCpPgdaO+1Wbu/CrqDcB31i+chR5+mmo
kPKEmz8wQ251c3fhwhGAcUD00eR5D68vpw+HL6eCVIUnMBkpx6+HoyCgtJGrZOykkFASfGwUeWjP
dn77HlB/RIZGuXLiXXyDjmOrzxlCeNH3tQgM+oBSsH13cSGBmNjfrZtNCPGAxJoXzlHHTKFOFIiU
n+LeFLYC5DW8q17eMBWmWfATjwfZMq9lVAmxpI8oSUT39PtivDAQ5eQMu/pAAjOp7XtWOlhzZAEy
hxOPJK3V3RxmIfxp44Uv8PWe4NRNIuWgoL+MnGfLNVb7OLR75jAo+xfEwlLTYKmoeIYa4+0AjT+y
QKMx7Rs+CagVdKve9Yjj1M93fm1S5Jq56jMyr/OBPm24tzatsH6Gx3hNj7qfy2qj0aPv/anJM4z8
kpMU5QhkEeif64JIFcYkrOHNYrh1MqJwhZL+LqgU+Yyeuxh/Q0hLN9/eP2bSn4cn3L1naEg41G6S
pJOxIRkCIxIOBcsmDzix3MjMtamYXBm+PwOnxJU5eIBkXTJ6RZjyuiXrBpV+YDECnZmduhnKJvYT
gfhsf2XyH61cYxmDzRtEopsQC5xjaIOhAyKwt0wnQkkRMFQ7UEb0ymBwOm5bi6zblzagk8L3Emcz
IWzjLLjqZh3OQJKGEcUhKSuUsKQN6YsfQqaWIkYHaRlqnieI1vxHQ+KahlIIdF3yy0uDkFCsBGta
98zDs5uzXG93gFw7XYWSVxBzWCkd9fTq7yzhfs8aF/BLD4V8BxFfDbCpVcF1bger9sJOhnTnGIbC
xiJBuYZV2zZpk6IQe1wzRmFHVkq4vv03vKhaGmNSrFFs4FrlIU0t1Wux5zWCehXPeyPPomhQ0bTn
UHsz68S8JOamVCZ7gyywt2RTky2cpYCItx+lxSHMNxC0hE9SC4aa0FU1bCU3eB4rqBzNhzbrSBr1
8PL1Q38LlK6QlnwIK3OHuiw1mqVTeYgoeZo3r0ftFfANb3O0OSXRfZmqXxmCFWgFVdKGMuuxnlLa
gQCW3aW3wMrCeMjH3YEMdmr6PkqBl+nfT2uu8dGC9pfC9LMxt8kU2JaWnOAb5sGs4+8rF5bqmmQ6
o+VJ3L5nlAo2Fd9husUn/1mID5LnYIhH6lTlt/Iu8LFxOrPMndClH7RfKnM0XzTMkVBDYbBuKbcN
zlktC2YKy1CCuyMB2tfpIz8lqeCe0DVolh3qFHzQ0/aq6dyIQQedX4SIOL3TUIP1qCH9K8j/UVLc
1pYUCuIqzRjxaj/3i7R0kV1NUoclO1nlCNfUbWpg4aAbVw3oBcMm/dGngbd7uPlK6Mv9/eJgPrmR
7jolEZJWdoDqQNYJuUg7p12ozBvC1DvKwzgxg90OBZjwwqlQ22IWRDV/vIbZM9xsEaVOLALNJ77a
muEz8mAy6tnX96EPVeyD4hKnS35SNEaNUzvhicRhE0Yfs+f3mS2C+EmipcbwTEotZ3YOZCX2lD3v
BnDKZkQs5pZVDFay3QpNUGzyRhycN1xjPOJ3KWEdj/xgEx4WWbzt9JGNt2wTKqzjs30zmsSLSd5B
Fy21CSuXSox6VzXpb2D2a7isOtLP5Wj5aZITxW/tElEFcUtszlNIsqbbisTGNbGjF4IKQu3Sqokg
HSrHkSyQRrKmGC0RFbfamwacOPQUy1BkBBv4wSWYtOEUbuzZyEvwgljZHDD6jjMFtjbzNPfyvSPm
FYo/zhmdBU7C5x8NDggHJ9XmFVxIlLbLGeG9AdGymLNZJFR+wZyD5gMy4uwUHiCsQbfEA4ILvn+S
Q9DbC85Rc5/IftmqJqV3T4Ym+ZI9+FxnsZsSLtMKc3jhzllqXAt3vypry1vFlzVem+B2bcv4cjYn
KJpTz5vM3i1t533KzjyaiIbJoacIgh2gNAI6W1P0BIePSnhWsW2Yh6JRX9rBk989gVJWAEUEVD2W
f4iTgZ/OuZUk+PwTkHLi/Qmn9SQbsg/nh0YG8KeCDdZkkx/a4R0uUh30JPjx4Rb9D9epWw83+KTr
3SJS1zmMLyjzNHEMDvbsDF+IqNK1x+r5gASsw5vFpbxvXi+JsbQqUyZxtTtkNmbty0CCJYCRK0U0
7MEHydMW0WnpbY/dI0P4a/HS8x8XIsF0bLgKrQ22qaJBmCPoHkG75t5ooE/AqVY58CS4rE5XhHcF
FlCnh3Lr3T+K+c7ljk6N2C/KlGYTdAyz+kO+cR22ahzITvGGDtVBQLH6mzM/25YcpfyJLOSuPfQ/
RCuOPKobHYFoQ8aR4dyaYNnKVftqZF5BFEzCcIS6zjm/FBzdiBXHr1VNVANRXxRHDQjiNTt2X+h1
Qb4DjG32kPTr6Am1wprrjgDzoLaLg5NKS8fORFZlShtM0Wn32cXlML+jQxmsAty68H4lV5rZtQaT
9XLQ3mcE4NNvk/SMLqK9M+Z4jzZPPzbdqLQgDYzMxMOTVPMMMh/z6yC/TIDCtE4Sz/ra8ByCNPko
gh5J6RMGE59Zeuj7+hn/2cv0IsB7c2PmyXEoNsyoxu9VcJrW/3TH9yTYXkytkmozAkErZonptHAK
FPfhfods3qoc4y/DA1dt4z7w6+fkg//m5uS9w5AZ5U1VaFN+cbxDhxi5IuimBr+DMxx0KT1ypfBw
WRtkmLSws5gNDCTYBCdCZmvsPYlRHjDFhXaeOwmWaWre7qCe0EhCgIpH3yAz5VUn4TqgTCrHLevi
GkMgC1ykv74HZdT6ojCmHKj9t+fpzTlngHBFj1C4tVtcxGxu2VKgBYa6bDCOwT7Izrc3oUPSlxgj
7/D7w9lK+1csBbo0RNT3wr29nJmKL6ctQf9xoLEDW0T51L2o6pHDtjhKd5DkOEl+Q3UtQ/1Qh944
z3rx6IbJ3Oyd7W4M7CQS6EcGAixvXoafJNtUy4osMcRZEOVUYYrftWn+EcG3ApugtWuF6B1cLnKt
7v4rrxpFqcNFBqHIOWaTXBaY3h58tbJiekb2UUNeuMe0ge2bq2Z1lKD+udYurSfi3aZ3aNo0JUwg
wObs8RkKq3Id8pB+8vJenZoP47yV4HLqvErDhPh8kP6rQKpsXKvPlRsZ9pM5eyLHJvEu2ICcKxyy
GgxZo/9gd2aGTyeXBAPArJLuAfiBhCNP36g6KBtvzEDXU9uREp5nHzf6BbDkmCBCtXxqKR7m8ZYs
gYP6V7MqQdppGZ9Lumqg2jyBaZo/YLCMx79lRrM6WG/yfkSW5BLr16z4A1rySzT19hgztT6wdDnj
evmFJaUwIdEMhhfDaX65IzQpz7C0M1Jb5llRNjHgfXMjtCFx9L+4hTpHC/A+ft9CkTeWkiDlXEhI
vsZI5vYD0KeWD6C82LUEOD+4QHDeGBb/5ymPQzHxpo7QSoZ7L7GxOLs7+Pwx3C/o2wyUMGMILHeN
6b24jOWfp8MZM+BQlhj1hOaIDSzo1Kasc/V+rdjjdVKN/ZMQNEdBY9GjMsDcqKOmJZSxtuZlnlP6
Ppi4avXfTkzxDyI7nwO8eDNabUPu1GgE+EvOS0UQhtLFFbsndroEed+98wFzBGFWDuErh26nx3OM
eJVofoWWEQTWfMB3uvJQxBbqNOBXzmyG4blNp9ywfqoIedMxtygbZfO753ajdTkNa4kadsOzAUlf
lTHyabjSjK92g6TBVR07EpD4P1ozT/7M1Ns4Mkl6w/wfi99Vb+7kNm9bdRFGUR4HN9+s5Dbm0dtp
0OytCONYqA791m5dU4sgMHLVUMKuwxk0zVrq9Mcg7t25H7vchHOJLAiyJktX/CuU781/+rWYQkK7
savBAN5YEnCg5Mrba/bb22XQMwqt6lg0edwUrIRpiAA22afR0lJr9ZI/Pu4t342UDjfRKrExQ9Az
/WxA0QLhoCEA+gASlMyP0SPdgiCEXxHZfqmB2EOLbgQvbIEWdKaqHuBpOOBRx/FJ7iqYGe7w+rWR
TxdbRnRAQic/XMSi7xspdyG+AJQIfMnM81IZk8Klw+GfBEGQ1wkN92rabglRbQFGj3Z4gAzp8PNH
T20jcKbh1QE93pK9LEQroxBFDtzD6ni7uOKMRUYsRU2OsOLAM4f8F4Ts/wmwjWP9LGzWGGkN7f5p
tPrtWEHWT/bWsL7fm4v3HsFf4K7fMWTyzZ4yPvVbq1BGeuhX1o+HWeNabf1WP5xJtWE4y8J6q8/d
MyoHzqdWpZP2Z+gcU/XITvDt3wAAOFeM20JxMVkG+6C390N5x9vA3hAyfhnOeH4EKuic69eRoGIN
4w4+DRC63xEw0fl1sYNs+cp8o8i/GMV8se/vWrwD9tYQ2sGx1xPOHakyY+jrIc1sylLc3lvboy7Y
CNK1LvVq6hi8s1EVngo3QzdHkN9G0G95/VyJB45YeM3BLJT2m0JqRr0r7lVI+CzZPh+TRhoGTUDM
ogr938xvP+Wud8FMyqDrnxbfz6V5m173hiYhcFAxFmED8dtlblu4Zdq/tvRwGdVWr7+JXIfNTk7q
jT+SWvP70v0THm6MLRdZzpfCvDA7FTZPv0wlT1E7L92Vnj9oqGGLHVDyPhKd6EuZ6OUCJdNDV9f8
L3ZUthc9w4Nwfpwti1Fr2yUhOHG4fy2/2nXSgf1tH9FsQ5MHbOuwag+1uOLFNhF51A8/q+nyQazY
EAS5HEyxDUaVefdIbSlZ/180pL0OeJI70XR8vxh7HYiGVsNLMRNqRVJcojTy6KsdqcntLtZU/95h
KsHqrNoleXB7Loc5mXmk7HV92pQlDuyg0vp29AAvWUsMik5wBPlKmNZ8ur/wDKHqcbcI1l/e57u4
yNqvxs9Bj3NMaA33EnhKDBS5V4NKi/TuJ+PQEjrLrvq2Ldj9hxsiesf3zdsKUUr9MPv+tp4o54JD
7CZy94YRZaC/qoKQC1rlRp7qF6LyCv0EyxVyzIxTdO6YMaRFhJYUkIoQOQpUKdGJLlpAe4f0mFOE
siplbvtwvbqAkmEr4CalZ2o4DAy7JnGGcKsxChnUJxcEHdLOiAV08paKp8R+S4nu2B2rOB6aVC07
x3zabCe9/z/AbtZqUEfq9bcgI09F/kXMJ1iLQJFbFCrvtaXQWYrjvnc2vba26Q9JzqQm4se+oDWT
ZD/FUp+ktefBd7srfDlq32YwE4Zj/Na099Nr5OUHD5Kc41kjIvKAHGIUMWx7CAYhZFGXioiJWtM5
cYsKW94fnBHFhgfHnyhYa+YVQfP45kArB/biAnyAHDf15h+9thFzzZutcaqkMYagJJ8ZfZBbMzA/
2mPA+j9bP073rDdcBOrfZxybZfr1ccB2/bLvH2yqI1zkSPo6tlQy8xP5S2/oR6N8b2kz+RVagYHZ
MMoBx+rLP7Lms3MBxxaDr3/d9aakn/uqA7Ui/9/IxeV9alZ4PPEGHmgjOfhJIR4snA/VAAmCgmKJ
a5A2f8vHz13k5ABrq0fEF9egVFaMod5uH2w3+kPVH4gwT/xsKjNEg3hqBqC0Wq/gQrh+bVv2si2J
BHZZeTkDsYxhik4BSQaWmJaSBMJ4C3bn3aKz/w7EeoG7zQMhLeS6i6pXXa9gvvR+NvgRHwvgc4KD
sfEaciOQrVFvKhrQL08x0NUh2VtYXpRvQc+F/aSWoiaez3/6udjC/eagYbcDoqXlpdxBP5ltHxZ1
eeiZ3wZ4h7iaKPaXmKRnXmQzCAR+x6495FybEaYvHGxrjg+EjG94CR0VZmsn3Ln2prjYxZ7yejqX
mIUwOih6wD/J88macvl6Ro6VAPTxxuAOzih9ROofwknC6wja+l3S8liUk9026lro4vTEnmDxsB77
P1ivw4aGG8jx0Zwf7oC6tXaMVTAWrWWFjN2GE9p0U/h5uI3KqJFS9Cvj4uhvgEZYgGA2FUI1ZzVd
ZFQsMpmGpQSDl2Yf5HEOfsmd5L58knxC8yarVmmsq5O7IZgkfpV/dp4mLyVSfI4q7PVOBmLfQ5AF
8QPenZ9a0+xh8yrgJM7sU9lQyNxaR2PSW//hLumd27yPo0tIWkDII+/RkIfHPncmzThiogdKJptU
no6dGkeVldKuA26Po84tPJQAophWaqhuqkbjUNvdMsXBN7DK8MB3XhxMssuoPbA4lirOSSXnGWKu
vzPLjoIGZJCd5YkzWw5H0SjuqRXtv/L4V2Tc9I4IdPZeoufzV72wOUfs4nvKvzkSU91TjDvKvXoV
s2RoGfWAK8Mc9+8FyKcqiarHw30QgnA1ueTxIBgPbMcAa2Z5Qlfch9jZMKaNpcuIp0JQ05Ax3ujD
UX3BDXaAC/B05uxPzcRs3NXtmpEV+8AkOV87zGKL4pIPPYiPj9Z9M5yLutKxAaVXdR8sYqKFRUCw
uTw5aurhGWLiBKTeSPJjvtargmAsArVBsdNj73jEMpbowHKvohgUnovdiu9otpFiRfTtDLZX9iSj
455UUuyodQBTjfJR9jBN0ohB027IJJ5rzmr6lk7pxQXmo05TDBdZ4oVS5Ais03Rxt2ScqP0DV3ZN
0TgJqFEdiWPO5gwsbPKssVl1sD/1M+APsHL3xguDmXdW6XglpqanD/tKqh9WQ5ZEoH2lkq6n2UWt
4hB6FUeV4gnwbZySEQfh9zTEs8xS6BzwvZHvVgY36+WZ5h/sELPZmv61ZqR5DVOsybY3MO9RFAsp
PE4rgUOqrbzWvijWOuEU+6Tuh1nXwU2fg53eAsklX4a6hYyCBQY7UxTm7c/fJ22y36rZSrSTgqHy
ca7OGE6jqyeA2AfSZmUlLL42DAaYOB6R0EaTfVJHBAqaudOtuymkCb4ukdhkFqG1sWtwxvQwihhh
VoMtuQQ46np38xZTMDV9O1RnMWghv3S7UgNokNd10EaG681hCu/faUMKelRZb14CNTFqwjefdVax
JmhPag0pcwdcChnseSpcGi+JQpMTDGYEa9RT61XkK5O2XBoyxemkHhVIbwFUOBuBAKkvuANm43qd
bBEg+jcRlBOwxpqDGSiIlxf5GH8aZvONAYaNvMCQ877vHz/pTQ7BcRBWRadHGcOFqn68AgNE1pCa
smIeNSJURNOsF2/mnc3FmM5luNRa8rAwb15GdEdBDyx1F5CZSODx3sr+UWRvSamIlzY49qx2p4Wb
tqiPRhuzHNwiq3qqN/FDFJaOEGL7RtzhPcjf6PaqB+/8C9qvulQ2AHy0D1LF8JWYKU1AF0phbKDq
rF+L2NTat+DIhArTsH2qGA+1AxgV8csjuA4F3ySbvadO7maIiARhCMjcIf8WMLu3jdVMgr21EnRD
rKumlZJbDdEPNdpfY4/RwNqZKgTGtWkmKBpV2FurVxAINx0FnhiHfRc9mb8fhWkXFbSe1OSkxDy5
g9P+Nr7yNchzXc2kgoY+Deet/oPLlYFtKuTYHpeOqCqLyDNOxW2wxy1El9I5mbK7rpl5DLRFuK4J
7Wvmj10NaHHQ+Z57+AXs8JcwsuKMQGhoaWc7Tax3twkzjriEAgc1X7HzHiUn0T99gJ25bJtasfAn
UuaPezP1aXR5JT981b51KWA6N+ZoSeMTYMNhrNbG2JSMztFZX6nRclQcCDsu3hfE3izNmGj1+HLb
7opjIuZdC9I9RL4pr740JLc0CYFj+x31R0vYZZN+mGAnDoLQTieWdRH04ZJ+OU8HTBfOf+qQtH/C
ehEeC3JooNay5YEpy4EQtHYsVE0pXzZDKND9XQEyFE92q+VD7swJGbdY0sf6FmtIuVVwg5fYFM7I
vIPJn7TFyT1uf4fvHAfR/ZUdhK58coGiAUIbGBcYEudkKVOvPinxlt5OqgOWFHNjzhdtI6qt+lg+
jKvb/bnnjgwRCoEwt/TdGoGhWxeBpGiFsuGTvc0QNbWLttHVXvR/54BQkREvgG6fPWkzSptzhHEe
KF8lvBAnxSCqAc7OPc/nnf6GXP5cOER0I1xDcgq+1XJxUMPmDdaAIB0NqXpowoGv0xOVK/AfMEYd
zFHJFjlB8LOtRJaD+iCLGBRZawnS15OxyQAfNmzO0cxO/81LDhCbeJeBuky57drCvtdT4EtPeQIh
F9FHyYyn5+H38sDqGzPsEaz2DAx/ldzce3ut3k6r0RRxaImFDnyFMTMS4FG7TII8w+yy8NFYTm3e
KcBiu9/XG+iIqgXyXlt5KC4ovHU2Sbz7XUb6vQLjKKjIUKZVgZuxv/8CjiPcGaTQXO3AZOLjZc6X
y16QJRdxSvYqDNIL/0JZjOq4rgtoHw56ThJKKmw13X0z66wWIW9qpwqrQ9tx0oj6Hl8OCdl6ZT1w
/JY5QdVncj//E4HqDOtNQRm6R8kseClQGSscsVh8wnxkfA2fKXmbsRa83slyeY2FySFW6ngOjs8O
0+zwKyxd6ZqNOlknwaQxN1e2Gz2TLnv4aUN1ua7NqTSM/DBfBc7jQfY2BKY8nXRJdppuf/HhvhoT
pOF9N+MsVWhd8vyw5JLeaKNLpwCuljSZARSNX7nimYP0AhaT309O4lgPbleiDGQqYX8395PsfGoJ
Prr3+kox8i4VTrQGAow4z3cIjfhDuXRbT9p/5RqeuL/vptZrT+faf5A+wa5ZWQ/NI7g+1h4zGq4i
Hto386dTkuYK1eXuLH0Qvmoo+kfiiuqw9A5F0R3J7LXoUR8+iGosBG/B5XKJ1WWMJVJWMXPoE4Qa
n4CskUPp6B+nvjBu9yj41okAXnspHEXP7tBzIE9OOdMqyPBWCzSbnCCVJxsUXrjBJXjvU1/jP3Zb
IrYBnpM6GuEfkZdoNgmOF8Yb4TsSqCWmy2G+hRF48RvTIZRXYyVLFOXt2zMgESoYg7SWJMpB+N1z
vdfru+3YQ+f2v64hh3UzZa9C4v6UAdWgy/p4OhCbvs3c076zmrk35e2z0MRNdf1TluFOsMEC4Ykc
k31P2V57bjJl8DeRmghvqpl7oqP7kANblNHoPUgCfuUFCp3O+Di4MfP99kURdI65IASscUNrO52e
eSU/8Sz+o3QEEqHc8lYmRy2KQQIYxxDo0VpQjW8abP6yw78+l5kNy+ANTN2Bh6iLUaWeTONXJeED
0JydJgxz89CTg8rmTpn7/lnM+9uCtbFYeyPxHCyhOQRI2xrIwHK9RnRgxLzRwkiz51+1Igi1zppU
1fSI1Y1XlIV3oSzG3+0Bavho7LDBTXaJEA6Q0V8ZTneVK1NGKKaxrgkxYzQYke8Ks92xq34Po9TF
O4aeOWV9gLmEudQAaOx4lKHuEEBK8YaUaqe5nuHQd4kw5xW8PS/ljicXjqYw+J80sNkw2FRudBTu
U8aDE7d9Ecx+4yvzlhTZG4xcF3pDx3ti/wc9sGnmw5ZIsWACTrSZzjQnyFCEb81OPF2rZc724mXX
vYqeSP/zo9IdHNy75e3E2W4qXWLckuoCTv4DycJA6ZYD7NAKOC4wTik0SAo9xl/gBgHLPXou2yK5
yjhbSKZF4jRbdMLGQc/NTs38NbYkJkT2X+vqQbea6ZQ4ZuG8zqTo26vZCR8Ed5Dazg2AXVez46r2
PPPhA5z71kgKuRV38k+2XjIiXNSvHj8heWtK0LsJRp5FoWVLXbLtDTDpIt5rXsDM9+uRgTJUD39M
9I1c48nZ7gy9CghC+rIHfCw6YUyuLCcXiKWCtgWQ+C9WeotTOqaIBnk6cXeCLcwcoEny9Vpocha1
5ATVarvpS8TMLDwoiWqXKFpmgIsLegilO8iVSgVRGeRuu7QKmXa2o5f3cePty0eaG+tW2SjMFJ7K
hFGthufGs80IPYhAmaatH3txQXO0dhitI7/fYNXqaLRSyRMY9+7D2MPQn2xoEUs6aK4vmzszPYFM
eXnRKh3hOPZPXqbCPvkOh17M9MuG3lWYdPaQ2SLWiedVCx5kJ4NILaNfvqgTSd83BIbs8R2rV0cf
7wi1MSpMwAt66qYCyerTFXDFnAuMFRTlXuQ/MzAdSNvDfXGpS9gE1OHSmDbNR7Y1Q3oHOMGEILXg
pFjnaLTS+znSi/zri7mn2izKwfqF7nxY5SroWTPK3+a45hTC1zyZp3a3G9LzXv0m6GAPL64dXU0p
uRMEWA0DO5ADSCS4LB6s+AmFWJbunor+ObeUGsMaClhycaAUUCqUR26D+wgpe5gW6ToYWNFaKe3t
z+/Ry8o5H+X067DOfuaPbrW+7Dd8r3B5+iaKajRONYk8r8A27++qe31e7cvBFNXqHQHilwAXJNBN
5XPObLClSbUZ1wA4Nqh7WXfXrIbUKTv6nXjUZMsUKQR+hhsWqk/aHSTnyv+yrsWnwz8++6QS88xo
ixkJN3jcF3fYo+A6FHMUbSEa3bA/31IuhfU/WXxKMqoo8ZyfCbWjIM9OV9O7eNYnxV7IBbcm7djG
3PNbsq3Id1GxrJ4s4EGAunr4Mu6Rs43GX/+D0J/fRFgiZAEV6W5CKrdLLzLANa1rRSBWMhpGF1F/
OR3HfbgUJpf2XXplKLMk2CkC5ejgDyczD5WAJGWd6PoPjmSdYrKUJMTaWRSc6ba1br1tgDwvdHz9
aqA1gx8N+vTOFrcJ/cPBStN3CubEMe2GaIM4ulv2Jkn5CvxDpAFKCOHUjdESE/XZkdXR3IIUOZXX
OWlFi2CWb7lRHW9/k/Ttio7LM7+9+ltLBOUYrmso5533+5wv4Z9V51ZIZ8I/3DtxxN9WUiimre9P
DYhirOxYy9E+ePNvWBsuSfTcguK7akuBjnJ+bYVHJwly+MlosZL2br4gL21GRyOeBekIPc4IJhct
Z6xxmlQnQt/ROzOdy269xtEQ5LtPdAuAsjLRqPWjCaHhTwIDEIOt4TO4sCO8PKAoiSmT608PUYkt
E8FIDUgRPRgcnoawnqMcI/iXZ08uyYbB2wpypF83IaOjCKiarBIEwjLR6YfJz69UL3wPkYr9T0hU
Poh4pDpTlyU6dTDHfJlXKCWAKyKBtK2KiBAjoxkmqQMi3OLAeGOzYVnclEdIdCU0S49A0VUWn3rB
BVV8HzunqjqtAehRV149w2i+U7PxK0Y1nZio1aVun0O5eEZDnjVRMAivOJpwX5leY2krUN5kI/xT
AHMzz12r0WgLG3mA5XkP5GqWAcuhLd9je96u/U9VF7REnMExgX4Zv1Vx/3CK+ZXXYMLCeuwO9Pyj
7lI114Ne69HzrMEYpCAPzHpr+vhzEgkvC6eE4x1rx4xxUP8AS0qvEXR/uvBlrooCNnVsJWosrbXm
l5FCEYDEGGZTzwYf70WJtlKY5Ry/cMpU20zpuCgf0DlzLDQHsyWrrD4ycGvovO+mXOsXfe2Wn+gB
IHVtiNgN6hQhUNUjVlU4trwkxRoFOEjJhVGKqMtp/Fe7gRory2QK+Qt0TfYguOciW5/DZEEZdm6N
AKmAbrM8xkFuqo2WrzMwddu0fNHa6bR5FSJjZSkiqHFV5L4FOtGYphrlBsXNIEQ+ljUtThFcEekk
zhYd+mpsmpvsKiV/i8l2NWp0UNRZbDp5sd1RByU0s/L2u58gRY8XJf/JyGF1zvSuBUy7Jx6um5EW
8PmeMcSISW/Y5lO25ib0umim9UQ6DEiYHk27pxR4OLvD+KXHiM9zp9yTn6L0wJlSnukur3jqMmxT
SfU9VoR4aARh01gf6vQXjUSF9WaxnYW7VwnjX6saH1m2RcCkClqeg6fsSrw+j1tqpJXpy28gbJwn
agdTWUIHQJ/I46/VR4Rdnrltj+gC4bMMUb89o7gEOZOYeko3sfpMW1nhWDvYH5Adf1Z23GlyVxIX
R3IfOYV+vWN1tpHUxjNq/nokLHxHPAFgmR6M12HEtnSGyvk/yBxXQlG5IoIiNhKNAEWBdPx7k9YG
E9EeopfaEImX4LOdjJxXkED/T0xGqEPaYPIO+8LDcUYMqdHo2QfAJGInfvtIL1yjkGOW2rH9eRby
0GlRx2K0wOGhFTev9DbJT/on4s1dka8c1k9k/HLOZC3ngE9Z2mlSgmeMfflcumE5BnGGWHQB5ohb
/70yGh5ZjLq7tDDu2HidoI4OdrwGMIWAUIFAMKhOwvBs1jgpXTDvOzAgUTkqrXjBsDHSjRqVw0kV
sWw4pL7lcFpAeMUmWzJmKIgRcsyBuQCYuHB/QaLeMvdYYnhbgKHxQgZvNU4z9nYNOKWgCisLd5zR
iWrPWr4XMbCuTieIY4XKKhOCh2qZUlBRWCmNzVdn+DVOuu4dldxt6S0CrGZ+biTX2r02Zc+rA7j8
QaOjmkUmhuItjqZJBzPdzeJOYDey7XWeUWwsNRiTOz5igGTfZhuaLSnwGLcTo6ImKff4MIz1XRRv
9GwmlI4fH79m0kSVBQsXGg9pXj6wmTO6hiqcmus+xRaeX7kxQzcYNOcW6yue3KcH0eqC6sShQ/qt
a2cxGtaokXpKbqV2ZYa6kzC47bpYacYde/RZA3IHQ0UNDKmbkJk61RSuhse5cak/HAwHBWPwSvqw
gZLdQ76yeoEH3D28gEGPTqeglaBtpjivscm9XQSS/arY6ZtCYjkvu0mvIBxTD0pDHKeWBDPsQWGP
vkvkCT2I3iYpb9F3Modp3QbPwO/kILXYYf/HEruW6STha/nwNW3e43X+gzaLyX2vidydbZfjY8Rn
kNVB1SGHiNOyHyQ9Uz56Su5w0CzuULWg/NCdkAK1sMNu0aZWQ3ve2lI12AV93rTITjmt2ZKHpXGF
NZezafgDCRgx1LdonyHtZpwzgMho3drAxBrjh8IYq+T9iLJr2a/37Oo8syU6SpkB+383VmTZZG8R
KpWz7T1x5TqDcBTkxAnwV+gMq7p7jsWwqWWEAy4ymQK8Sj4wFLagJp5eS/pv0PIVSJMZ9G1+ti7R
qb4rqt+GzL7AnZs7WEkw0dEIRj0cawlyZF4jGBJniY/IpUo0xIleD1TDpuKDbC9FhGR9Ki39vfRy
dVvki0wXaE11+iXAR2122uN/j++frZLR/D/aOrVcO2csk+U2IBBYEkxjMt04NwlgIEjq09CVyxuR
ZWPp0ZclTjcwyLyrV9Ri04jZEj0mQFX/2QqVXDmizJLyEZyWm88w0Wix1hs7X/Rs4JmVwdAHDbEP
Qrl1B7XlZ9eBwf3fCEZfNeXYB/d+MRBLYSkYF+6V7NQ6xQZdFVFv6HnjFHqQkC7ry5nrT7XP7H3/
DBWra9OJhHnNhj9aRdnIFIttAXkCd+hYYz3mV1+gZASAghpro6aoEnZaMI2sN1GUaWCp6j5ZEC6B
jazMIuAVZcBI0riJg9ZQ7WEwlOKlxkL6K+bUshD1RkMyUhb+HqNpM7l95o+T98A7mpHZOxTmaOqU
dV3ZGjZoFdVz2erppyP3BbNLw2O+Z9c4FIPqCKPNhe7eGCv8xD9dCVHT1T6S3NpKI9hDUMjcmLfD
bCx5sqKElEAmR5KWb824hP+ZaNlvp6rMCfxIGBzD+xjbJ3qyuesQCSBj7iewXKZB7qcxxbmC83Fd
PuYgkbrw/cLJvbdJ2mcKkrq3oso+qqaFa0KoENrG6+06f4jg1v9Ji6kGOhFpbyT5DgqMIkgFlf+E
dTyYZwyBzllXsbY51+FMld7B7BzKvLCExxXjy4nHRQ02u96joqiAvzH+BHC2Uz++gIZV4Dpmbln6
OgZo4l3Ho/u7cuOTbonqCNBJWUXOxsA9vGuPhRGu5pz0vEwdIw+LusWY8AUUHmhG70A+Mv9bzjHD
ylC14+2/i3MUflxjjvJpOIhcK2aehCN1F7iNjdYVYWu1Os3FMizeg5oSxbCQ+8imZ56zw8xZZqKW
15qN1Ft7He0F2kgZ7liTK25uYoPPJTp5gnv/64vlgvAQhhedZlVj0kVmuCJhRfJjvZHDxE49AZjM
4ilG3AWP5HTLbDP/B/poZpOzri69YhPJ/yEAX/kkTLXX3SCINeHFq2CanmwEAc7iKDd4zDNLEOan
rCDaiWB6EDYO5qjlwk4WpwlWipotHsNK665wjA/R3+E26WUnMvyRGD3vf41gqm+qgmbnNBDjUeId
xkNnS2WXLnOp3CwVrhL072d5ZEBfzarBP/CIFw5LLVZ3vCdJslwWlpD+x5MZDbejub1wR0nGIxli
VGAXX4QNqI4DFXbr2aJffIkpAnQXLXhHSGHAt4sl6Fuk03qZm+9dMc0b7HGm2SlXr6iZOcbxvFk9
9ouACEJ3NbTSwoPv2+9w/vmobUl1qELR3JElQ6pKjj1mMRj6hT+XqYA+blrNgzru5vEe7wRa6GgG
S41Fmj7lc/vTRGKjHuX56RSXNHH0o2CCfFEvnidd9XxQe9kuP2aCXsP/ZFezwf3BfLtBAeLse5LN
lwIpTN8xKhZA1w4FfF64HDSP/BUlpYQsKyZo8mT+qPjkaUWSJIQicStwkBVo+Z1YyV+ylCK2dLu5
HsgWT1s81x+jAauPByOKQHOpv2PQW3dIAP8C/aYBWzt3a83mAnmOECdv97wUvbQB8aiK2ZK6IB30
kEd/RPQPLqpngaMXRV1HEMHjwb7Kzkou9qQZeno2cysRYDH7zFFXSeaQCgoQqrsodGEVvKyYjlEO
HujwFm1AfLeP6Ty1bdYtNLDGMPOeBQvxSks2Py+Tknq4JMAFC9yZOmI1xnl9MBbrflMhHoY+XfCr
cnyK3VndMiWMsza43CQKr5aiSwZsohJuSr8xb+/6gVbWxtw9zini8cNmfFNCo3OfPR5Y+fz12CCV
osxzLEaPubjO0ubItSMhmRKFYF7V6dAwGMSW5GENtFI2mx7ESZ191Z5eMRbDHtFAsoCHRl86NuxK
7zeoZf1HLXfoM4MENRkFE4z+NxImAxa7yYDa6hwMc8HE+u2ZX/tjKomEwRJTFv0+txbSzWu3CsXB
CTY6bErf8lFVkvIsDL36NMuIjRKLY/TvuGMFiT/HYfEpkrfOgStlPC/GnLQYVuRZop4IW7TMpH68
ls7Z/zK8/egmS1McXG6tL3C6FkKLcUmFkzQIy1D4uZHxB79xImYvjDEim9kT4bVQ/Ikg0IwWvFOk
YDKOzugzrEXnTV+8WVG7nyoKVX+Jq3MoqcdL6RvBgPAbZ2WnZfqCRVHCpopAcz5uAM/YfZHzzYO4
NgcwgGej8QVNSOsQB2weiMMa/BXoCNRxnuwCfoxEECE6sdamIZmU1asWTCfynERZQZUgYLdjMM6F
4pKoSxevU6Wcqil8Vmjw+2WchadlmVSldV3ty5ElRRfmXDS0HY/6BRmdouZU7vqxveUSeJm14BiM
dzFVqUM7r2b48OgTKJnMuTeDfyOMYhVgOyO2kokNCCtnMmCHTwE3cMqMWFJAvNKyNHWHmXgPkJoP
ZHPbGsuW1JbjaAG2nvurKoptaJIn7FxD7wvBW2+WD2b3No+mzz5SMGgrrmGsysIXXCEcpXlM0s59
QSs0GjuWgYlstL3GVJn4o4B9ZMLQOxwhkSe+/vPxFOgxK1Qh8yry3lYBtlFHidEpB5PqEyNlSEpf
mNJFYXbBAFa0yhIljEOfNrdaH46mx7wa+QR8msRr6408x/B5djzrt7lyiNsF5rXyFUvcliFI3hTT
Vs5TlrLlFu5otqpL8bemUeTTGO5+8FUqUAgImZyFXPNRia0zL4JJPZJhA4C+ENutktEkjE4xcV/c
elwzE6M+rQl9R2GFqK6aVXcvtr+y1AXZaA820nLlwLS8bpCRHRJAs+EmyKcWPjvqxNQqErMmqjZW
W8WFpI/eoI2n6dE9/A2/HPIF/0ML5kdctBy0umOzityNgCCtoCKb6bCB1T4KTV9rw624ROYDCsu7
SEcRdzYkn3rRpHYL7ziOgrjLv9D8aXocsUY8ll5flwP8PtTjBoc4bEEsiMqFNmJSJAXF+EELx5sV
/rZJmUy4RGRUw4/D1j2Yxv5LqnDMJ9w1wWRS0rQrrBznxeg+Ds34aZ20APx8flym6klCqFIuQ0i8
acFS6ucXEeK7g8sunZbOPnZGcLD9OiNeIVq95/s3bi9+oRKF4VcqUktd0ACyE22qeiLgAmez/hYh
yXXXYaXjui4aobm9KFxPzIb/efdPMPx2kZjQWjQeBuGyBPBf/m1uWwAWw2aJOiC/Pb4MgBh6XGO4
KfDPK3DGtXYfLb1GiEYx0hIvrKxVeeYjOsmSfH8ogHE46sllrkHmy4DInjUzGby81zTd48W6C2Tj
Znw8sHFJtOA/xjH4I7L97Vos0hKhQFFKSAQOtqjtrclBd8BhZm75KwbdmMI6OcZiN9DZ42Br2Kjx
NGBMhdODcXzgUk9hImmkkxpBh1YFhZYn2CV5O/4oRj38+zVKPSqvaykiO4ta/k73wiNfvEvJmRuK
LQFugTx4zIgGVoazlLT/oFCGoTgdcor8h0rOPOER5RswQ9IdSCPbp1VAojrPzmwVdZhMJ/ZGd2i+
TvMRktI8Qk9DYrkTHMMr2P0Ba4U44GN7K96ag8QFr3U05EDlA1DvNAQGyVUtYCX1qeFAodmiJ5fk
d1d52HsXv6G9eMp2n7kajupE2sWsMI7zlHvYwOKTKZwCqUMMy3apvDxMkpArxnh1TBY3Ye0D1WKs
AAi57zC9beaUBWLRcom0rMpNSObxxfSKty0i0mcmMuq5qqE+hu/kT1yjcXa3HyMB9IkcLX4FXH2s
j8oaIdAE+hV0y3O/CBCAStVn0sUiAm3x7aaPB7d40ta77RCSTZm1D3KLO9h56iRqDjgXvz6Tlmyc
6jxYs4DxAZBnLOqEGaEinZPIjelA/FbjgHe1Mh0WQMUAmE/wsLTlM2w2tsLhc7J+ALLBz9u8LP9w
bueUpsp8WwJEe6B+7Y7q8USU+LYkssDZ9rB0I1vm2n7whQqY5VjjeIiLo5T5JKqmnm4CdvuxHWSM
+hXazD+lMj2sMe748Gmvcc0m2k95eOe9hPqoxshgU1dcfv7WlZhX131VG0217LptCLenjMi89waA
LEhFeXF8LONCBcEnWr8hKz8Ibf5Gu7DBNMwMNapFgJoj1MsSaXRKqfd9IhirKrs+eSEUYa+6/8SL
Fvgo6sDAQ6+Cta9tZ8LOVDA1729/Sh4KlRAnbLdzotUAaNVOcMDL0ko+ld+Ew6Sx3i0YN1QtGJDd
nJOfQL+RO3cIMQssuCWYRfiYlQkn3U9fdUcsTyDFSsdN232H3vs4fxFSgBKpandClpJQlBeh3azI
geDozUmt7Z9A0NOVZ3vQW1tmSgaZ/cmKtZ/aR7CFF1EOfQWU6TYwNcRzx6JqCklFUG6ZFL5WxuJW
oGmAXDyn5n1Dsux0odCC+gPD485dSwExL93oi1H7TFtPtBPLIeRFQ9My9GwTjx3UJN+tp76CX9LR
Nz+pdixp3wEyFesPGFNfwi/wW1K0Xck9cZJb1cHK0Z8wG4FFgRTDFd6qeEXOcnPewDhkA6IkQcvL
6EvM4mTbgd3q3NwYkWfPV7CN+86Jju9VAz41Jpb5mX9F5na681XRUcjb4E+PbnxUwxUITqh2jCV1
ozEOtviWVctE/EEqUArnUp8kYqE/lqJ8kT4fv79WNJEj/tpVryIBeOp0t9qaSv8p8avFhI/MBKHg
ymGDhd4jqJX4IiLjE7ZYyKKIggaqWn2jIRdeVjhDAaxDd4LJDgSJL6o5E934k97AStcuAiOr8QDA
FJMb0gxfJ1GV3zQFI3yaCUHZxIXlluPF2JvohG411jnMzyLf+zQloOfDQSxk2NIrg7KhwvQOlMhl
LZG6QfMrt3tfVBcpL/IHp+VvRuH7ro8ZQCpqWmfLWtLIfdGRyVYe9k+30egD7Bn8va+1Zi6LtZjn
xMz/WRIT/Cde6bOHZp5vYj1vyXOhgZdZe/qHUXy+6h7QOKQ4JzVgPnDU6zxKRJxw4jfeDXo6BJZ/
odeQiS45QJxNO2veH+jo1nsIAn+mItXabraqYPCIEF22AW+iU1Hq07snquKLSbGAAAgaEVztfeWh
I0Yw7BIKs74JfbHwV6fM8wV5VDHrNQwMWMhMH6+03Hd7eV6uO5g0VQ5yQES0YmDpq+fOj3mogjcK
wt7TicxtVhkFvvSn9RPNM2OhIHdlnko91ICkOVPR4O8YOfQ5mg9loMdC3CGRzcx0vPx0J8ufP4SU
UBMrjH6Y2H/IYBCZ7mBtrsHQCSSwwRyXfiN56LAnZwwNjGdcYUMKkGzrfY/BxTZOy6kOTC1LA41Q
kh/0h6aUrJL1Az25FSm9bfDBHma0TGl7X1oow30eRDYH8WrKgbsbU7xkS4g8uRI416sP3vB1T1uz
TtxZ4rPlt5UQWpmpzb6H8qXDIFl2t2T5Y1JY7dBjEK60GGm+X4RMNvmf89JVv0NAxdltvq1CrsSG
KDJ0Ksx32IniTBNDULhnDhwEeKRItNQyzp9T+OHJcFH74hJ0GlL+mhnY1odL6O+VDR0EQ6YnyJiw
mwummrt8xwG5um2w/zzz+F7iwEKv3hnLX/RONAoNzJaMFCKBBZ11Pk5pd4DkE/J+rVzIjr7gH1BM
Bf6KUtWA6+BnCZsr2FPgdDQzFsNdl7/FSzPWzRLp5XRHv3WlL/p3W+zyzQZZMoITRad7orKi7h2M
Qna4TdgkzRi3XpsngMP96CC1n3ItP4CHojdFxLr2FHvJ64WAi0BhcfaN8SKvibQVeN3GBdzsY3R0
khr/vZJCG23WLSwiWPG/Z538Ap7AyZQnDYDJIDdR7b/ai1nhG8IhI3KxDQ8kofhnpJzO767qY82D
VoTLjXxoS341nI2Md1srZ1GhcLw3t3yil5kHPCUdSicTGUYLbmP2uCeOQQRUhnJppjA+c989ZDT2
XdvU/ZJxt6NjHI6KfmeMEyIJtStu1wjbVcA5de7hcwzR2FkntcPx4Y1bOZhKogZdJqYTPFjTsUHT
kcLpzeGEd21GG1QPAxsMiEHiCa9Hr8RmeblIYVJuRO0QnOOB08Jip6wovZsWmIpX4Z7hj2AfJ8vS
ih1F/GJwBIlolh8mLPkl3JdG8xqAFf0+xWB9XwcFeYi5w4RFBwtE4SCQvMDluKk5xrtuXUZ5cRSP
encdTahjN87VvJU6tXDi4WUC94ANju5lew7cSKCl0Z1nv0DpQ/nsLclCPRrKwXtb5AcY/ECb5cN/
Oh0s7vI3Fg62nX9SbJIuQqeoYX5/lCCSRYr657KP2vnsb4QnpyD0I0XaEljak8FzfoBRwpgbLI7b
m65yWsb3HP5oKWjDx3f16VkShA6P4vV8JYFr2HNJOLwAZnQVfRRuBdL5e7hrRfsUxUFsRqk09oLY
eTSaUu5FQ+xbU0c6eW8mGP1GFDlwxWOrTpP5lqHvHqMfbOlHX+G8ERNLrNADabhuZKHP7J3SUW1I
PafO+XTE0OBp24dsMdqgs1OLMz1dpoE5/lPEjk+66xtSWxPngz7rAYDEggug1txWp2eR/MZ7biZw
zopx48E9dJ7GxuS+E/RZ/gg8KipS6qIelA0G1v+mOTMGNum0xCnIA24HlMN19JPFSTx8k4Hs1m+u
3Et5Eay+ZPdJ8MewsaPiJa/VsDsnKrEJKDz1FxhxNa+nVmhMyc4SZR+yPiCM9omw8KequjNukHFd
1MIyalQ16w2Sn7lFG0X4izTiBJZVKTLRG7L3W/R1GkXbXJaxoCUITqF3Fap/7DbkLJYUZjRSz5d/
wrYG2VIcI+kNrGbaGcQAf/lUGdea9bZ83plGuocQ/jBk7/C2kXOMSXw4ONtTIfi4pqESLNOSH7V8
wwl8LJ6yhA8D6qi3UMK0h6N6hE+4armWgSsGjwq6vrns20iPk0O6VU9DCyjG2BNL6WnDbA45PtI7
zu43PG8ojYlt0h850ASRsCBwzCMjLu5WgPkV2LIz2vOcMbjseczAQsJX+9JA2P1K62Bs/aKgMEWS
ICPiVGs1C2naNK9+c6V6aySlUKuTjV9qJSnZJpa4KT18AnbrDL8qCtqBxUPZR3gEwZ5WsDUGYzsZ
6lXNS7KNIcy/Z0fReoyPefVXtvjrjDmBjcsfQIcRnHil+8lOpa/rtMIDtCFCoeMLvbL80kIeeh9P
oYeTw2V++8XKxAs62tGT1UBKnvPuuq4QWBlDmBR7/7alEMlnL75szAhdWRuFAUoiMQi/BoNYsMem
uYja5Zwvwb6+74zO4o6+Ao+Zz5V3LC/SPgp5wGpdTi/ogKizUFSjOrPrRfwLpSIsGfCY524A3aYT
CFZbpV2bVhNw7SOa3sVB2DWedG1IId+NMtsx+DkjaIoTYOFkOW1tx/RWucn/OB7GkiHwAz1Ljj4P
TJnWi+BXnhDMW4kiKKCpsJ7QUVTtk4z9/0/x6uhI70wah++eDpLAeANQhXhDx4qbIW1bS4X95o8J
fI6aDNhSG2b4il9l3ZtBN4JgxXCPY6SryFoEPRtlsjuyOUDh+hCFS85T6bvJFjScfNJWtHDDvxXB
IvQynd8UxdfaauUYu1EBcH3xcVNFz+bXiZzliCpijLJGoqyTDtT1+Lrd6Fh9CPgW0P+4nY5qlbS1
Hvy0qy3Dy+X6lJ0NjwkfMl5S970AV43rw/O+uGbamojQiXpIPmgnLz9IE0MG56HOJOemFVxUBERU
bC85zG9tJuMsBLt4TtObhN8v8ZDu6sCRWhL54rsVV0NJM3Wm4Lt72PLM4h6gpgvYjNPWeaShLc1c
w1znH8xLwqPRjoNHQaVfdI8K7B0g/pqayhgwKrAxrmkBqG3e5Flusw1m3BPFhH+cQjiomWNMDjzH
QbcdU5AFz3X+WwItzu4fsVwj2YRrWs5sK/MZsBx0J7dztvP6lhZcqM2y6EsKvbHqLPmiuQldvg+L
b+0EFmJh00hjaTdQVuOgKCoMPzXm09IkobhntfwBVys/9xnBlZQExp4YohOHy0FHqSzoS6pg2DkQ
Wfd4eJ6/YriFYn76vfKmtaquVcO/nn8Y35oXo2AFwz//KZfjQQJNSDZ+CWXYal/7Vi6M0S6Uymh/
pp9wh4w77zRE/df2k4rZjMiLHTxhKH9ArdfTnghTaTga1ts1dmxL2mL7sAima4MBb+DVOvg/HG9P
6oLZgtHtrmm2iabdtcfxhI0RzwTaFXi4vgm01MnvhILhqMpRDO8It+G5Vz6DaFvKAbHpz3vxG4Df
G7sVyosataQcZDGSy1NFeePuAp9j2xG1EOt4X47zQwleozlik9nRXfS0h5X9wPa2dQ/Ae4aaQJHj
XVlrs9Hn+gdZqfPqvy0wzbIAL9GUaBHbyrVi6hcwyz4JxW3ijoPyx2pRvwqvspYsZ8vgcUP6HA2R
JrX/9+FIvZ0zmEHvvrk5Rhc7rI4Q7f6Zo5Wlfr8JroyoBeV4tvXM8ExqNfl8gdjXHdANVB9JylAN
2BL1x7jOy2r/ivNjHo94cC01/5GSPSnAxsdAmi7mh5UmYYCyont50lPFq4pL4Wz6DJ4c9KxJiVNE
qxpZ7QZnwhyzk29Sp+353Cn6TrGl7oUyt5cwU2ONtAIA1WPmIpVQ7NNS6jUgK04hCTEM2XKZbZcm
uVkmJOKeTfGH7ykGU/yKqoq5LRhAoA2siaV7CHEDrZlZdcpc9CSMkhS18SzQg4bHj6Ah+rdypWgd
Mmh+C6AT83LoNI5ZE3PDYFFNGyVt9rDqWBhxJT4H1VZCPlLlP3doVLJTONsu/43CX83FhHiAIbhy
0azHtJwXCnhfUdoFC+LtAJeojenfgqyoadyFPign9zkGzqS8d5oBMXRwhzzko42B0Pj9MsOG+Z9A
j1WCI/6chdtFwESdmVwCZbZjNc6oTX09+/fw2G0gWsyjN7bj1NQRfM/yZI03ZPleNzhIDj04mp15
KlpikXMgq1kqrDPS/BNIwvyWIJBANWNAN5zVjArV+qNJ7IVHn53iRMzUh3cqMyXRMoBeMtRtA4NU
tjGv3oRFvYdsPoe0jVbCUVm2bhMjExp46tQwsQhrty1oR7DnF0JmkFzrZTJZ0XXyHNww1xB7XrIU
+kuDhyoTK1Iq9RbILQ6US5tmVWJKEyQKVXaejtTrC7OuGXZlhMKRGKoVm/g8XOIyOdAnu7B0QbVC
h+kFb8uqEig1zt1vWpLSmDuv85zb9YwMtLVdalQQeWQjJ+tUnH3H3iulZ+vSDniMrtvVrDUEQ1PG
PK8LAtvB4Pk6g9pIHyiCmC69yCXzD3IeyjHcAvKDO7ugtYiMC5zTDHsfJpIC1oBu5LsLhEsGGEKW
FLaMnjX6h/9yF5rr8qE66u5mUNp9lPcDeTbtSTfUYV0mkgy2r88VKqm9Mq2FaRn9O6zLTvejOvwh
4olftjfaT8tONOTHyhfQ2zTN+ZHWxavSOltvY1odoSPwmlX/w3sFr/4N/DBzfExqWet46GW2U/3X
5sH8pVqZjD3vMqu7xtgkGclD5LVvIwLe83e3Qdk/w4TxtAWY0XgjY2t5zY4t3ot+HglC8ZjWhl8m
fxqbTwdNSsA2EBN5DwYS6Fa3/deDtOUP9jLJ3EKFq53szW0KNVbuW28BPbCpXxdRz/uDbk42t2sF
UrgTJKHWu7vwRWgKZl7zeDNr+AlsZlj1ZC24dPMfd1OJOYl5LhxvISjbdD3bAhN7FU77Hf51AyJF
Q3948NHNn3FhCOHDRaBPothiSxLu4mYBWy9Lf9a1WTAhRykCUcHx8neiMbpbHQf2vb/Ewq7HUYBv
hlcoCCBDniBDtu1TrAJV4D65k/WdBN3CxdU9Vbo/4Vc03sQSZMXE77yOtYKqiAdwiHLWjTE0gjSf
pgZkNdkRkWOvILXCueOGpt5XcqsnE7LUbdmOUKTVt6VaIlwLsuflF+h/4DRq3Sc9ikeCHxfKsW96
5MrUcAhp/ljoc+zrqfwwMsZB+ubN7n1q7nJZo+vA/qfcFAyIz4y/D5DxP6fDIN8B6QvQJKr2oJgO
EitEXSw+Ms2iKR4eyB0MzKmj7uj5M22GU/0KI2JaLAirGxXU09cSXE467b5T8WqvVJG5HA936NjN
5ZN0YW48S6jkNUOA7VIX2uM6ZxZt6neRQNR2IN1VolJYFwt9tHeTcF3ar2oQ1tLMszfSTDqA9YRf
4UuCXcWIxvhk+TwhgWdb/6DVU6iGYeEAZfH8R8eKMXoHdmsFFrHC2vfYFlbeeV4iFHi5Ouow74G+
jwoXjWbwdQH4T3Z6hrXIrKd4BdVX58caBMDDkVSZhk53euBF6/Xlj50b14FVOW6g3df+roCVKr7j
eZ3GTIhDVeh6is2IWrJUd2GtsIWrqjl0T8F+eBA/YjQEM/XHExq8v260ljTzHnPAGOpPIQprWzAx
u5/EP0diuzJ54XVdz4Z0NqHB2mozifmSiiM4gE1Meqw9XS3YBe+rR1OHhQtqCw32ITWzFpfMPDfV
oVUw2doUoeRR2Mnu8eZ3iE5kmDseFPC5roa63drhTB4gkRDjlor/VlbfOYAoE+ToQyKd+O2uXJ6F
USCuwf9HUBir8Xxe+A8VOIBpVF6j4YOlDxkxBHLQw3I+KdCliA4TNFFGtMWLe9OmFxlKOp1ShDoZ
xEimztNGkRMnnLMlBSpdFalgjhkC8eqzgoUlJf/Fvd33kTM4mO2saARDSR9mlXxgOJFtyTuToqLR
JL4SKkPiJFMgq2JSKsYU2VUwvR73qHsNbMVoZBHB/lOZ9cpZHM1VzBW/ZzEgAR+1cgSn/hnFGV8Z
4+DMDvOdsnoLvCZbjqDXcCOPwqE6hmJefCJp2ez1BXidFdizqjL2r0oTtZrwkjLwRaO2SnVlXXHf
4JhOBpZoy6Ap0/U4NryyAq/gfaFbxPQpRb9rgeqx+o6TmPyek01Lm17xIEsp00iAm4ZRmra4UWeI
i6b8STF/dh3QdY1QPKYkvy/AaWFJgBJR2HQvR9GkKt+Jzs6g/ON7xsksdGbqTJ6IeWhyHQXdfACi
7/HkMLb833zCdsbQwbGWpMC2rraxBG+bN0aHTw2TyRFCWWlnSrv52DQlKowKutv0KaRtWJANoPfV
wA4HoOPxx/QCdc4nJGYdB/Nr4t58k8panzAUlY5t4bEGvec7CuPSbOsAE2zP3+rvUKFBkAEoiQB+
oGPg1Ig+jke4DIDtrsXsUbMvi5TEDSYpcwLBczyWlvB9VsM+FuSEFdQLg4JvZdIfBg7r81MKvRdK
KWxYXo3kgXF7+f1qsd8NKTvP2ndVv6XhnvefKU73YA6qNu7cMrgyKOs/FqI98wAiwb/1jUXplLiZ
hW4N09CxwqfeOyx9ZjELXCNdrBF3nKLWi+wKHJxtli7EWGBVq+Ex++8aHyiRwDGJ7xQWjJgprm+m
ck/qvbmDWQiBxGq/vCHY9QVAZeHO+5Ez7LwpjgyTgBGWGwAbuVkIHi5eH7fV5WmEk29dM4Jflbr5
9NLsTOQus00izPvd/Z8Y61gbvycy72O55SnCaq2TNGpch6wlm9xF+L7/VR+li9/omAA1fv1xAWc0
M7dbns29V+cw8+uwqdUcXATGXqLqkxDIxgWnoYQC0fXH69X7xYFDjzsti5TyS770ZsQMCyYNhoOI
PbACVFHvrdFCh9Gfpg4xS+NJL+YHXudZrfx/PjWJmrtyQ3H3f4d3Nfzfq880+skncy/bOSylrkVu
63taHUEkQ8HhVI8loERw0Wci8rJzXJ4TnxW03xTfiHm0eEGuITomGEFvqfmv01vGOx1hChKIfIYq
ifFj6bY9yYh3tZGE7qz4oc3VARIDoYRvs9qm4flQZO3ZrIEea+XYiaJoOvyhTMeJ1uxsziyHV/aV
JobVXJD2xMfIh6LnroOVaxgXF7KTHp/EbDdbXJLNX7tEFp6cIPxosCS0PBlG6/k51uznvpH0IWtt
+l/O2CepqE0wO9cJeNn8j1VRZ4IbqepxnqeyF0x4R2nyF61TnXQd5W5ucmYajOsibqHwUZTNJztm
HOMEAaRTZw8Y3YWzNwH9d12IedbmC3Un0jVZWrT1oC+d8uNFjjVGFVEV27zGT+5WL1aqeix5Xj+O
t7urnX850/7PjdplBVtPXmXbbMXtantpwjK2CLBesrzPViaAxn1prTDuMuU44/EsxAcGVeHSmXVe
fRLp6Xh87oczglnt53qovVeTWJkuqJCKJJi5JcrhxUdSUKlag39vS6r9YYqA5iLWvQWoQnuUs6kU
stamrpsunPqz0gfKUgQheBS9IYYCcyoBtafSayY4lIeDVsbAu08yYS79POaXUPgJsin73Gf1/U60
DEpIk67txIzU27t4MYvcuARrfyJX0EN0IWbgIK0gDQ9IkqP/xPUwfq0IYR8tz0yHRIpgENRHvh42
4a0S4Lc3YhS4E3fHdrLixkE7oTimglFevHZCY6xC2hZ1ye7tR8JhnOF3pPehCU5GOt6Mdp+Vq9wh
iBjg5tsBf98Puay0NY21unSBLQhkDbS9o26UUSO2+n79o/UsDpI6DLIUclADrknEo9+9IGEeLz2L
JBtKqCIV0BblEPVMj0C9clxSBkWE/c6/IULYO1whfbKAIaSxi/w4rl6lnVqko+S+7dJacf8dfnkY
S3FgHCM3BIXxVuXk2EtKNQz103dNUZ/fuImGvoU2ufj+B6FLmptzdyCkDEPb6mccRMpxSLhwVxSt
iQ/BgG4e4ddnR2i/1gvzgkEA9IEpb6Gt+gISfOxXyGyHLtYCDjHDBNKX+FH5Gcat9UmBdVRWy+Nq
92WGYzx71IWzkI/cviY0cyUdlKzHNChTXijgiKU2LiPw2WL2/jH1DiLQxl5QfYv/1sQkIeoJcxBW
XpEfz0uuAy06m7yHNRbuVfFXOD+k6MB7WOH3kubyVBy9cFKoCFP9pfqH0x0Ut67Y7DylHZXQs5LV
ksCLimLPEiFy6J/mIviYSonTFnyv3OWp/LCEd1n02/UMWtt2kGzINiQheG49/+qXq+Wli0A+yYPW
5LdeZ8Vs5XY1Lr3OAmsUvvL16dsWUo+1b2Cnk6L6jJddiNc7PqYHxxBpeo9/JvFc9LRmL+3ghQzR
z/N1CmgIH7tjBkVWeEjZw/2HQeMMi5SECDineAubPCdKk9AxAe3z8g50TNB5iPbBxnk8fGDq4Tix
k8j5+gX7JRvzDREo6BgPfbVUmkktFwlpGZ8tDr8q0DMoYzTo4Q9uezqOGChkTjhVJjDL3GHg9+Sh
VYtSZtfJ9fD4qwRKCXFOWyqaadOZZFxgh3ftAKq9lT/xfqmKmdGG152TM9VzqlkgGoawV7xklD8T
n3ybwmkY8Q1MoMQuz2TeLx7uK6P2du39CpeIcqjFfV+8TbZSlcljtjcj1lpMhf3dwHxD9decBaMc
hFyuI9eD1S2qbFNYYlrlC+rWYsraQzmXysTkkzRcf0EEt61AvOOmaH/yvrvLzu94NJFi1NGBp+o2
5h5TmHDgcJgJkWkeFhumhrAsenL/wCCA4zQx0Fc8yPwBAeEjA4Kz/fr0+rff3o15UCIxxAe0gMN6
p3rGqffFgu8voRe2Dc0EngGxCCHnqmfD/WZHzXF76SMVq0CgMJVRgWOyQEtaJ/E+oRUdmtte1Uxy
WEzDol93PKcbPKIkDyISVOFmVjZ8QWOSaq5mFQ21kp6WYHZ9Z0s55Q1D4vE/LRpwJ4grN3XRMVEj
kn5rQ8Bu2YimTJXnnsdBGyUsrCzaDUfEXT+Zmhdu+g/u+OyLAd4GgZblJOD5bLOpaaobA5FNYUKZ
X4xWyb4QMo6NFvNx5zjc2leJT0+gDvsCFoDyomVe8FSUeCDSyShumVi/+d+D4NHjk/eYjUf0qaNG
beT5NiqNmWKdVjlC9XaY3orlwVlxlhGw3y4H2f0TUFQejjmeZj9Iav3c/Iffc5Tk93TBvf3d7PgQ
Gn/W27Gi5AO7IZxn4N1oNdunk/xNyd4M+lE7gWo0XRe7eqssr8l/eDewjFY2XdAbX788qcMVam8U
ciw5FKTCXNw3xiqyx23PWPAjiwRMH6Liyx1TG/xbUc3KgMe0AAHuBCrpUP5xlYMVYTq2i/sqOimm
5FkjAYlaf7N16gNJGjRCsWCPB8b/sfrfNITgxStdGETUUrfvXBH66hZ0MjQWJWEKVUq5ud7iyFxi
dpDDqofFOOVEKwVRqZ56QSynKYNjQZFML8gPi58oogD+2u5GEqIBE32ip5IVSBKPWvGR39E+OBzX
VCej0LFDCKAIsjODvrD13rjxY+tM9oXOmw1xoJPOXrWzSgMyhw0FdMSXIboHFDFpzUD97qI9m1yP
JKYuB7pCQ37krII5u56cJsv2PmmDyX+oZE+nZOtT1Kmo9JfrQSzYaIWM+Xg7I0J2RUk3d0imYdUm
YmH4Qy2Yv9G+/z5VgPYsNRKOUGzo3mYCxIBSmSsKnmKdvPaGHOgN167Hv6ZWXPJyQJN0IULf232C
768TKjXEnlxNpJFHQ3lvY0RPi/JpQaBxR12G9kI8G6DfO845HYDCe21afBWNDTaT0YLkLNsT7MV+
wHjFiResv8pXPbJeTsUvXrs3glJ+OEzZJTBahLJvthPQsmKZwws4WntWYxOrWbr+6i84aFoCnTwD
7lJFK7ciOQsRFpBuUrVrcuH3YepFWhcfWx6+XR67f9zX0QtdLorOx+WbiEgNUothV5C6Yj5McNhe
zEFwtrMxM4kENDMRNGaPeU4Jy9wOHpQvU/F1jH1IgiDwp3NffxKR+29gRZIABOxw8EkYDHFx8PQC
Mtm+xb0rnXGT/CGb4WRFhhF1dkdhw1xBSHVt5kQXY78qPyC6kD1nTP0TyTNgymQVhTD0aEVfYvtP
OA+Xl4gZRKWZD4HoX9WNYYi8O5qri10/Oln71q3r7TV7LLeNISkOmxXXMNUqnwyKS8EWxtNNOeya
2c9F3PoRLaAlyfLqd7cmOI10ZRa/7vJlvKWieUD1ZBW87TpQxfYg8h8k1TCk62XIQ1mN/Hkx2NDs
8nghIy2YXuoJMt+oTdtcAGBaq+mUx79fcywlvzRS3tlEJk0TqY3anzgD7GVUruIQiUPtaOPjA5pj
kx/7EXNicKSumbSEFh3kEPW02mMn6fGg9dx6rpZEmtRbLoYUuowdbX4eJwi1bpjPXq2QI0u9MVbI
EJE9+eAZmXPPCJQN61hRVHfK3yjFHJhv02cgRQLXFWFG7frALvcFmcyqRqcpIAzVoLsYv/Osk2h+
zgAuXGDHarKUZJ90pVzC+F9J4/fUKYsmbsI5ED3rr2l/2VyOY36/ZVOSdvUYIWAtwdZ/Ll8jo2A8
94dZFAh00KKcC6oeioAiYykviu9VIV10V9THXYUTHlETdfkudP8RSmg//ci/2iJCx6vatYjlLPt/
Hf+axJCxStnvi1uJ5hc97sN1xMUzWomVMAWjcIDVJimawzhbQGyVTiBl4U1YzWleLpDmpLYaa8l0
uVxzfzYl2JnZxtRSp76Z+rWUTMV2ITCT81arkthf0n9DCvMvW0S+xPIl3ILN1NZ4Y96LiOgiKvtZ
zgrQxBSspeQi3Y3+XBsmSwIFGzZoCxA+3U4O42n4eICRhauV3HeyCbNntpEVM82uF8s2csQXpiml
GBI4NHZHrxzuo6RBiAl5Q/zZS458+faErOGZjoRgdnpOJukO9PSjyWZttXuvipa7RncdFpSaOx8o
rqlby3YXR5L5yC8St5BLBEPoiMM2Y8RVe96B9cIcuF4lORPP3S/C+b0w3jC/ku5byjzSNMtpuFkw
ClW16s9z9K+XbYA5S6Z0IZGLrMNh/Qd83uRfxNYAkT9blnjwwnDwBPB/6zcuPg7ia3xYysxdZzFM
1/B/Uqg6SVep6A5ew6kVGNZM42VTqjhVi/R6gwLnCHRhTtrx6nLsGbGPTXfmaBsWsdg1CHFD+ENW
LkCG2vkv+wPh8FVL3CU/UF6Ib1WFzupTCDyeHEXUzNluKHeAcOIhfdx6NHKe765mbp/Bu2qZak5T
KNJXZGMho/bp9ZGLPJm/q0ZwAV29Kv3nghidNtpWXoucYhQ/RTnwpYJVQiJMFccp8EgODO+Jr8Xw
J5Bd19EUpVn7SFor03eMz0DSdB/ov5OyE5gRy1pepFAQ3l0mlh91pqbdeI/ZVGnG2SVf551iyJhs
bzGdPIeg6oyFRKOXC8WuULTSTiMVppZeOEnGG6KuDapOPmqsjuAPGow1NkOOHULIkeSAfIvRb7op
2gIEg5eJ+mECbzf0zbB0mWzvkUDkieSuUmZmSnGuTM/4tNPOux6OGhhqndzFkjlzI7cZKwpguSEm
yj6ivMziNWKN2e+RiQ/pPTATcmoshYZiDPVtp/0KtnkaHjeSKe/PQ1AmL9DLeSn6Q+Lqs0ZEViIJ
mqyOC5YNImBE6Ww+v1VV4g/fBQLYoLDogfbR0QdJqkdxWob/xmYmgN8vSfqdY/+wVR1z1WG+qhus
FS6KDFX21Ux/RyXZkAsSXWms8furh+mFJCbJfrmXZzWJxwa/jUw6J2i6DmAFaQ9Qp5XmZ2OqKU/m
ZLUbAChukngtOJ3RKgkMG9Ynth+ELUA1oahW9ePKWiDy8AC7Ma23/L/Nn8b3Enr7dC/PT0RSgvhY
4/zKFrhoZT+ZF4IEYivH//ByGsrjqS1GEGyB/HhbBwsDHr8UTeX2oee0iExe+R6ViKxoTnWZPlbl
bf8QFE2Mp0lg2rp+zagnwqDbDnhwvO11hI0FWYtJMr+6L5hMe6HfpG5YxEAr+V2iAaUJWNLkvzVz
n6jZvX/UV+S18LKtKWUQnfyVsL3Y7Q9GojW4RqYClz5Y43O7unsRSOlpLTYjek/aJM+AGDBmid+v
cU+S2xmD3rd+Wc2ANHPdwS1AcQ1L9TseYj/+QZfBG7sJtEPAQheSg6AJNoNRK3We9b5lFGNn/Wqj
3ro57bd48N/DoDyi6hFUSr/Y/5/YdO3MD7lbFg316yJkzuubwEs8QmRbJpesNnbLZOxKzwyAW0jR
X6b80xc2OAvTy+uc2lYtsVfBlZeGrycF1w8GdVQf/aR8vaCuWKeFh1h1wND1gzeDbo3yB+/MqIlv
c/mjWuq9s5LLBEYpC8GCItggiAitZdoqH67kV3REal7wJndVDjgxnTxRMHAKQUbCj01bE5JuZePl
BolxMshXxgXLOzHhLKDNGo1/cM5Mrzc/WDjEHzBZVBPG6h1R1vqokO3b2aHyEesSFDpF+e0aodTo
R8Stj/CRKqOS54IMrwpiEppu803tDNqhXw7OM/DQ0fbsBZzUQk+RrvpmvHGh7+DNtzLFqf3JYcNf
jQbsWJoNU9BozmfXTK0Yuc1Vb8ccrH1hKhvyBu6dvAHgNj9pddrHFY7C8qXELthcQx4G6LnMeVnK
g+vRZ3NQi/sYJhjkf544rA93H2vtyArrEMc+L5cPYYn7CREIEU2IByTA3HYwTMsvqg28n/5Cjrwm
T75lx/xUSmAtgqvNz7/X/2IJeBZ0ikQUoIfF3fbbGANBs1P/W7kaea4ghFibFwaU7JqLJ2vuh1xk
p7AavtuH8t5iaXMtSlywmF5NQFsBFa39itBQYlU5evB8J/0sI1NQuPOAWJG50oDkVwVYbI8BoLJb
XOPoDtL56JcCgFvHJm81Jv3RdgYlxA1clDeZ+MjTz7jWMSe3AuU4mS2vbqoZowZidv5KEIyk+klK
47XR4hYDC2k0HvT7xnvsjP590O6yGiO/10yC2pWnNI5KTonFvVgBkobLrDVdY/gTd/FORNrHsxbf
U9Js4piUhTlYr4xTBJ3UIS2iX6iYFZj7z8tfZ8PAN3wJTlP6GFQJ54CQRytEXnGq4ZNMmyomS3h/
GtiAMddtzQt3uEN/Ul43HDESKrpr3YEwq2pqPLctv3KxMv3bJYIanCUUh4QO15muGOIo54XvDlnX
RTXXUfAGO7OD7INTrtcjIuHo//R/0I+9aGX8hsQokvbT8M/iOccHBRMavdcS9B4mae2cSFpqNEEc
sXoNZGeLnCa/B66HlAqj1Lj2ycgzzNRWhP4o07ftKX81+UEnmTOd016ftHv+89owcfx13gOCjvWp
PhE4M9v3lUtOueTXCutQ7HRaAq7AEY1/C/usNvhT9XOX08xu6IJIRaL+CdKTZKE2MUgdQymW0Dcq
Z1fLEIfol/VWGOQ+yxU/Ts4lQzy1wVXC1+ZcuBsKDJN19fEQiqm6BSwmo4HdD3ytnrMFIfRoHRiW
vB2vNaC3Ek3dFoufus59AVFMqxRA63lF/HyFSPO/5yZlATO8e6xFZqNaw8xGHGTcIeeTF2ih1lxC
VTQ1ESQCtJv2PRRTcmxqGa6nCl9PnjANSnelUYq580BUGfrbRQiBgO2xF1IMQi3ALsJjZkAO6U/n
5ZkvX0+aPsdbvOsWVkLt+4p+HTk1MlOxt59aWkAf6UPvmEhlpfgxr+E6PCgVjJZ9LrqlAGPX3BXv
yOYWnD9lii/YcXmK5nWmcQ6KRS62nQHkEHOQotKDkcsa4nlaNy3sl95voSr67sSN2O6eND0UjQmg
HF7KvMXMP5mKHgZluOPlreuMmmHxtccnw4l41aSADqXsNDHIO4x8FoPUgZiH18p1f4HfildJZT0v
a7nZcmxaAB8pyPX3VBYR6OE8d4d2Hnww8jSmszsTKvpj6PHlPjHrs+7bMCn9bCiZ/fT9RJvkDPXp
xF3s9LLJiSLRwViexx3kzjuiqm6wkgfg3ZqzBXiJ2FIFoUDrZ42qWt6ZKhITOByGMHtCh9NESE+X
KK/VjVztQZVAqD9T8LwxD8yqID6IFCF/GwYLm7sRcI/NQN3xAnjyrMyT5Y6SU9zH9qyraS1Ob7W1
h8bWa2QdiegsECAdGnYpa8QmsVjAlc8y705EL1Hu3lqf6Uwrr7UWzcW4SAb72GH8MAHlx/rL5Dhj
v6TD1OxwwdR+Q2e1udtC4Nt8Yrd2eKFlHZi//VgKzXQKWkUTrsClX4eq3mqdBBG/R7HbuCgvpvAV
nTsugdh9l/9QAOp3vK2CYgMkuSLhmtSbdkEUVzTSxlutaWtMEQucMdIVP/6tEdWjTPV6iUag9zMY
FWkfF4xs3lb5vEQYgCSAG4MDVw0gDH9+c7vGRNuA7eRt+N5DVGVkuIGuTfsJw9s3BsczyxqOhThp
sM1nX+p4kdDshCGcpSLRmrwRxMIXIHFALME+JTpcYPT4STx7h4AyHzrGInQx5Sx8+l0TL/+WI/Pc
G7Hln+5uUn9nBdQpnjVmODCBKjfwlFQi2c0j1P1BryCN284fLLZr3BhcDR75DCXdfSTWtRBz+bxg
NB6Dw9aww19TwXfrdnO421tzSP/WNW0/zjFR+MIWKUpkgebsQ1X431iSexLpOliohZtBhFUFl/Md
QYoMhwQoK68zR1M0OjUdzlv92dVGKqjCUwQPYb2bz8zAXfeiB3JEZUo0PIo3OAe1au/dq0fDPOWw
H89t8t+aYBM0YGzv1DIJ2Ui4aYn1KBV9671u1isMNmNHj6FPuNNujAcI3eq3XIFVSkWidvPWNq1D
xOLYEeTWKRVL5kmSXAQ6MJ3pUWjz7wYqNTN58P2wp1xD09mOBNQUW2UMeNjjec50o6yMfTi2YSAc
YonOl2UAAg56zAKZRhd9YP9U7L+nR+PPMN5BAAvO1kJ6fB17rU/NkbVO/1ObkEzZqC0fdIDma4Jp
s6pLvKJ5D2cVfYWQffIwsJKvDsaKCIZX/TLXcJ5oZGRScd+gylUSwFyEI4fB37S3mduq40BcKVEe
cygjwUw3DPn+eNlqrbBXaViF3TKla9f1GBOFT0O+zQBnDEWau9aQbAo+wtklwrbVUoHx8X5zfZuM
Dygp2WtheJf9pqN+78XnieeLD+YBvKzKuTM4CDNMbVqkS7oIKihd1kygdRel54cELaVOQMaMCJsV
ZOpZGM8erVWjrbS8HUnRXP+mpNqfz34k7qgo8FyvIPtzREUdVcibRKyCWdmsujJQGXhX30zCTsm2
NFkmqFlAEKpa+t5SPE6quHXfi076LuhOni0N0OAE2OvWttVGWqcFWBhofgaHgHXPskhXZSEP6fPz
MVf6tHx86Mcc0nHHyhAWI4+iFlETCGOABz7EYV3iiuvtT47zlgfkVsDRJsYSdv/Kt5yl7zT2ufwu
X3ibmNydKtnL9q2vxsFHundeSWsV6sDel7Zs/MaTegqVYGjF2MF3GpzjKclrWRATxyL/G56P0SHK
3N05wggJmCufMXnWT7WQn7cq1vecIGc93iuNZl8XIzbXkwl49MZslsmqhXvkC/cqFn01Gno3lZiv
9AFgFY7Y+k2xr6dHCUIaX4LKQr/qSaJCeKm6CLFCs44hntjodV/NBqo2NC/1sgn3WV8ygIpsrm0k
J5l0Ps++eaTW0a723gj2EfXM8ZO5CuxQWpl5zTP5C8QphTgwdFUbz4SSF5tuSwGPMtfsOb4PKCF4
hq3MKJJ5PW4tQe7BNto3bLHbPiNzYIEEGtnKhMvDyX/AZhbfZ1nn862e67194o8NecafHIa/zwB9
s9nddPRgWCWk7xQBq+CbgjRRqfKvatdR05aqsHSft8WRKrN5vYRX7Lzlcrv+S23ayD4vgGPd//gA
Kk4L+aaBrm6+1lJdXAPvNLtwTxGaF+3sSPXPdfa+YQ7Se6BT3fwjsIDs6Ia6MnV75x8EvjreTVoE
oDZwSxQSY3XwVOZC3SS3Oa+/UAOocUyl0JX4dmBDpMwEDm+eX4i1keI+h9rxOMCPvPlQguQRxGaw
tyk5F0BzbXTz/X6uSCYSCPq0PQzA4KQ6U/Syta5PM6Z3ZxSrTwFFkun3MmFK+HBYBUsGCXdkM0Zt
6rO/RNG/fwCz/EXI0A47c19LNEDFnAdBnWOtOce89TzyQuFPD52OHYGtSz6yHhDMEjaeQtQZHn7B
dfZwsJ7INQ2i8CcWvp8X87z6dl/rp3e7gI0BNHdUN3trACKWEghDLafEdnkVZFIoMkzl0msTeRB7
MRvWxoEE9foe1Ndl9JC7niCmUNMbiXSyu0oCzs3/Hitbb9Tai6kQFX03/fUe7IKD7DUWZs8Ryamv
Mh5+jpcoSzFMEwZIGgYc4KkmJduL09p+ziE6pcndpqfGpNWAFTbuZykDoqm6BthnYYnFn2CO8TQ8
9FAFiGVN3e9xyfSL8SMUwg5k7V4XqRZVcC06O9MubrL0gP4apuNHRZZMRVSADfR8Hu9HxFHxaYIx
h5vIg/zTKP9a/62uhgdIImFluzFEQ6t3CQ+28a4X0gVxAM4uOMB+Ak315lkyZahtKfa+JF2cLV3e
cXQeMqWWH2LTbP3Floq4cmrd+iBBddOwJzflYNB13XjCcCLOooWMzM/YkQ0pLofbZHOFu+0R5xbP
FjEILgn8d+F6nYugdcdXsgoVcscnzXZXd4CjOWJ8wdF413MEaWcUfhazFJvFpgx18dEkwRuyoOq+
Ng7jxKfVsVrmS1dfQShxKphARn3BRedwn/sp7qOISNbHo/ZZBfuW/CtBKuY6FXXwWQ6CsKJIHKxW
z+dO9RWyKwJn3iIFKWhLf6s7TAQVylTSJ3Yibd9JVZireym1YQDlLrvYi3R+RgxPmAtDymPvDsMv
4/XItTDZYc10i5Cgpa0v8X6S7qDv8//TVHkprYNXOHX36K8lqCNQ/4ka2q7twErNSUvwreI/yTvz
EXcEiiNU/RidfWmRClJggB54tZN/yBW9utnuA6zLpPH55hNnf1uWGvVWp754qdIzl5lkWvaMnHy6
Bwji4QUQa05Q4GDfzLJrKC6rRepC9ahbE7zb1ELxWLhDE1PNVSIG5Yi0eGT3LWWaxZTyksdBLXto
Xo7+KfyvEQJuW8Umc6aeGwi25b5RR+V4ibNOzy442z9JaLChnWDRbsJdrt8veUFQZ/Jhy114b9rj
S7lo7a3n3mR8YaFu2rXEYPTFEp6cHXh24KOdCOdPB5o0P4RmDH+kKPNFqbsBHsaj9NNgBX4zB/71
XZ3ABE4//hxQ5jMu8BbSUIskPcNA+FjNdzvFAyIdsy8NmiUo0iM0KJOHO2G36GCUe3xPUr2/JHen
lKsLDsSBEsTwaUoQT7rvJLY7QVozGscnbrDbDxrXpy+/csVEcZ4xLwn3pzjzgKvPoN1CEDvQPvrj
EPp3npzQQSZE5ysmfpB7bdCUvkSLy4+uRv0XfLcaBoTHgHldnutC2SgC9g3I065VBVHoDKkAUPUN
yRc9KaNGRygnWOZDhTkgyHZrWGSmiZYngNXQxRhWEjO9cdQgnII0/sgGRHX6TeurEOgA2EphTihr
fRywcWoMmTmV2YD2ifpDj2HBasGesEG9hhztklnbZTGJ0qYI/IRS42N7Q8G0GqPDhwQO5kHa3rjZ
Z9vQDXSPzuBLK2ZHHDF9mW+EXhAGlXm6XbiIsgMc+zYphA3PJ0c8X/pwbWLY633kCMEThc/Zzfjm
WlU7PDcasZ9BZQcxCClAtXWHS632+4URbw3KAZXeFTGB6dzsMbh7Erec/fYVb63JaleKKAEkzYJA
i/Qh6OlB/YD9EITdY/NsGDVijkofGARvEH0HiLf67UmE/5OUUlRYUaB5buA2AsUxqFhy5NCTofuK
ibIoh74sttvuFP/jv/9yL5YvOr5zoltWTtmtD2EjTgJ45eVOsF+clcvdHkboaHqhKm8sGG/XMaBa
ipqfX3DblRaghm+EI90NQxzC4vZCabO5hDi8dExE6LrwN6ELPbvga8zfaoZNaSE+g0K7Xqmrdgzt
ZSztEdbIHAe5PmnCHr2XtDqJQWk7mKu42e0SfBsMzwia3Mi6Go5QIOuSkb/qVBA4z5bt09rv+ysp
nDlFxEGop/DZeaPSpS8LYlkGv9CwTEaPwfMMNNjct1b9PFIdkUrbVcS2iRAZeZRtfmse1lOH+Pty
VV0Xw6w4n/9LxReDCixEKLoGURkywhae7JJeUAUJOKfeJcTpKwx8JJRKlK90YNXHheXz+sxbAz95
Gi0DSRZfBx25Nvom/vpNA9AsdMYB46jfENTlqrEXlQBLm0seWMN6bA/1Af030Q8b/ALtAcpJNOly
sfjGVp9MryrNalTTuiy1AIs0o1NnkV8tePQvz+Qp/CCRDppRqppbnShNCZWWRcu/QS5RyfIXeFL/
c52hQ1sg1Im/MYN0gkoK3rWQo70yhwY84viErpgxiSdYyssMTihu5kxVJsAQGTarbORUvptIKxYy
0ZF2ut/y+bw3HkD9m0nHjR491eOhkyy4cDEqwJH1MvHD6ddBx4hNeM64jQTzP/v5TzamR/z72Hdl
R5Icpy2Td7QYjNgmfew4g/1SY3CU13JDxKW9pWU9Vs8HO8JjPZSt2wlz6Q3rgB1mg1k2avmLrPRt
38WDv42H/ecSwYtT4V+BkKwHMNFbRV3NR9g++vw8kEBOs5KxDiVCcnt0aNEPVKzhYYbwS/fNkl3Q
pa0aSGAvqCSRfB88rCL4H2az6/ByrMzp38AyhtE1dw5q0vjmBjvTaN9tk1f7n3Ifw+yRhQvhfggL
4hZ899aeL+xJDb+wA3AG9P91zwqIT56gkb79ADU5QAuwq61y5XT0bVBbQMsOwEz4YBc9CHc9FiMr
eB/coECnMRu8NIUdPAg+aJcwVMsg+dvzsD+lyoFrGbnHIcMkQWA024mx9RnHCbizdOb1o9vkvZT/
cnOYQkP4NxwT0KkvUCkA7jkb1LJ0Trvv1viV8nklOVCbH/QWRKI7//t99Gta4xQaTq7RHgDqShoW
lEsVnyOKa+nex2qIbrszkVmk4vUkSke3zXCcxU+I4B+N4sYV8N6we/pQ2o0OaIlNubLXwcSuB7Rd
CEjNqDkteAOfXFgpeCIJpu+Fwj81q5rKFkkvDOYAnxsj3tiM1IynblNlArqaSTU5QwkIA9IuO1Kx
Dz57Y4Cq4shNj895XbLSBrjswPAEIpEh80nsL70ugUzinOFvWcgIWIDSBb1wYzlRMHCY/y/BBhmv
Md5cJ9AEccQjSgB9BG36OhnCAxDM3fMX9id3gR3G790EIYsgMH64Qgidh64d6BFv+2aYbq7hiGMD
UiWObh3mRfzGEfNKDUdhWsr7KdwNrIvzmRvy8WNDYrSd2+4yAMqfnNkiIi+9+LhkVnCqdRc8gyAy
XpWUTZIJ0BDSU6vmTxtybpA4oVuFQS9bAhkfLzX3J4+xEWHDu/Couk9yrPFwSCaJP0PTCh6TJXgl
awT/fxuzeeKxivAo6atMT4SFVvEj8uAXa8EPHzK/wTdPsA3fUSFCtuDWCKtEpcytRZuzaZYo5vKL
XYQj9LkVk8rEhFPTrGuTV0hAMkkzfveTFT0rr6h6jvRgBq4dV+REQzBb3OwGIbWl5w5q3phWpGq1
qJFyYm9rvdDNZz6ltAOyfxZJO2qAu/yw2jIt7WFhdekznfpMk7+d8fuSYDiyH7TQqrE+Lq+F1wbX
Qgt9SGn8uYHbnlqDjwXF81aLAAzMn3QQcpF6KASjmW+gFeh6FCZUGA+mf+v2TVP+aPTLh6csExLv
w2pQWydoXWq4DU/c6nCFZ7xkJ/8h+od7MtJOBtRnUCUXSWJ+6bJbOMK25u6bf8WN0bwz2fzaXndR
miEWlfdTy5vIka7tSqJtXKGhIYTh0zQTLEDmU02RIUc459SU9LMhUtmJGTkNFQLZn2XkwQz5cEE3
03aZiBnubIJXol5tqw+t+4cJxyRO/tckADZQspdXb6EaspS9wYMQ2WWlG+osSPwCfIG/hKE5XOGv
XTuHiOIt6GKBbAPnMgtbLBlXnoPd62JpNq4dcMAp/eXf7uD3gsPCAPRQ1owfBULO7qwPWwbtlFau
uqNEjDE6SnKdjDvwawHYA+AxZy6+RQkJd5Q32g5sJotRM2iCeXgE9aVWYolQZvOsK1GTxED7EV5f
QKLJXM713HmpVCthKENH1gcvIzyT3BjBTfIAvDuhEDyPsgBSCmdrvjafrNpyfUP8ubss3Ug8NQFb
mJJvUlWj3BZHTicw5Bjhm89MukwQYUeePZQwCp4wH7IZ8tzx2p892SU4T+3thweWFVkP/5Y8+6ze
QofbeYU+YYScSuUEW/7DtZRpXVworRMX+X2OrZWm4nck/0KOAPQryWtL5G9mRz9PdCp4gaRbLCIt
EH1PAOjc2+8Wmj/if+49Aj027CfjAKIUCDmCkvz2PNaJfBJSk1JlWafZUu0jCK2Dx1WzeWGczLqg
AlGtzglIgkKN2+BWEhq+ZcAxD1b7PlX4wbLR4dfVaA9ZnFxAv9eAgP+82iqQ9gUlMJku7A9Q6KHL
PztyOy3oMVnQ7NEzJXr1fgqrsi5rMy1bEFEl2Fc+OIm44/6zeG5vDf441ei1XiAdJQ1cS7cLp3bt
OhUfHIOkRf8itCEb4TwZvI9pAQ2S1oDog7fVQBpzFu5LfMHEdfScRfUkhWTHQFO8rauThPCFPvwf
bs/GJ9NZjtU5/NzXGgHSD0dkxceEH3CllljU1/vvYKwMyc1jV66lpCUxfhw7WoLFLbr2i4QXUpzk
CxSSgl7+NYxcKLNduOy1Gl0Pv6xOUmPDUoMELMz2+UXAUC2wH9X0lBRJHVCsA9Nw5iWkzzhG2Y2M
INPZowiD+p8gSicQ5aaGyMiEWGMh2LhY4NGu5CyAhE12HQDJLekURtzMRtMW0Rd1AHA8tIiI6yjH
5kHEkxECVduAWp6SoarOYaE4LWfC+4fDNnWFBYk3Zp2XHP7I45uE+uuZbi1bKww7ZrWe5kp+kFlC
iUsNeBmJhxiIa1c5HL3APOThiA8Y8hSZsY/vW5qgnFjS7AtZbcb/QwZLyN0V2q7GMy24a2jX0VNn
o3hJMqrPlZ5LiZr/yDaX8ROpkTRegsWUTPLmKsacP9n4fuQQPnlmTqUMf49axVEQUD13o7UfCVpm
vNh6JC8eY6a+fahQ73CscSIjOzTizIDAkcNi4ojKTlb2h9KDyLSWLHkWkX2d0pGrhkwuTMfbdp0V
R72+k9EI4JxqcoP/YGdcuOhhqwUb/fWtZW0k3krHlknrMUtFwO5dUDc+o4AY3M9NC8LyNJB7I368
EDXE5ntB8tzwUp2r2mQQjDtgyBvtoMPBNbN5bsXMySYDHI+yJR+DK8CSu3EfRHnLxvHZy0k24xLE
t2k7BEdnBf00wS9oNY0MDJkAp9qGqnS/VHNd4W3tXRRJwGZznsQQfrROKxa2zF/ChFWWLa4Puj/L
MMDilafvH8kKPcbcGGuNBkic2PM5ksa//i1yiIaeaN9z3M4BFzFeCQ4ZBZuRws0EJd3OK//FwsZb
Dd4ySNwcRv12yA3nQBnI1wWlqB3Bw/Gg4ZEWNcoXjcDiuOvzT+tQavE7Ymua8vqN+dLl/CNUKrD+
zXmG7UfxnIoSWQUbIcRjrWcuc5oDf/C5A1KjT+LsgTShc0ctb39c0wQ38zTBYnF74yQ+ZrlPgUYf
OSvmvW5UVnuzgqorkXLdGT7I49JKHqXlJlJDs9o8UXv9FHD4QcYFuMU4Aynn837qmz8nxqM1I4Zr
0ZoHY0rmBYofcqrbHNNsqW4n95ij1ansEOHiTcmlKbaQyL2uPCll7B+wjwl5eXk2jcIC+x6fUHxl
Dlf5DVCcXGPK+KHhqmDogeD/bsSb1I/Dx6h7GvW5jQuMK+wf44UnwUHXfStXJ7aiiSKKJnwzqi9C
ng4jTfZWmboRSw501/8j40kFzC3HyqFjptTXRZM2+8zWnwNJdlCxSnl7YUoxwyJN3KRnTc9+UVB9
m4a6E4gZP6fD5bCjevaDHYQZHm+m2NC4jrmZiQJdf6KYF4K4YCBRTqPdVJbrpgKdNEewcm6F6VS0
btOWGmfzOixdtnjcEZ3a14Wz5m3e/59meGRxLRn3d/uZCP0gosMmy9eGDjmYfDDsRWZUt6JWHNEQ
+htfW7s1uk2Vxri+w6BVkNAxJQL4OKXLrz+A+DHVXm2a/8T0FXxiXKnaDinfQcSHbH0TA1vpMuar
QI0HLgeNu43ojvbc3YgDrJsfAr2/gppZU7e5E1okmfPoA/cHi7gkkmlE2UxQdbhkb18DKqFfwBQ3
1206Bp4FvIsXoKA1xEiYQRL7IDxpsNHEd/r0QxhKECgEknKD2Gsuq220fHvbnxGXK+G/3kqi4atP
159pg/KSYlkUOUO/W+sUJKQ23ZEC7FYlSsiSoO2j+KYXuiZLp0NXTuRfxghavtxCZA4/vRRRejk3
ZzkO0q7Z2LPAQyfM929VKpR4VYh0TfGopF4ZXWvpCjbVd4nNy+RxS7WpDBiOxMs1A3zkDmfbo7zA
qpewibaQ4CysEM0FlQnbuhNvC1yqzgSVoPLcK2LbIsrbs1bFJanYtUqz5X37SLy/dnL52z0+h2YA
hQ/0RpDqEj8MDHRwIqez+4/80NosWJNITYmjJm1fej95d6LS1gPeVthWNBd/gH5RTPpQ78N37v/z
byQMEI7J7lBnRzZsljoLLach1ZtfOjXF6rx9E+zySaR8bFYY6zmCDDr/oKtsZX66Fbu57meosEpV
SlhhVuxAuvtRFM/Bz8JbEjugXCQMxhd4X23nM+xCpmIMSGq81VRVudljrPE6XUAsMGkbe8uDcZqb
jHFLnwqLhtsrnrP+7rFCp7h07i+H8aYEyPGFOPUzldhTKGMYIU4UN8NBwBC6wQ+tDzFmGZVv/i3Z
nmeFjTgf4tf+Vwi7/4V4JQ8uV0FxYxGJOpryqqm5OKjt2SC9LNBv0SF822pEAk4LjtrkTconGHZ5
bQ8sFIhCLBkP5/2ZzyDr2SZ5Slt4UUCh5cHrKC7fpyxrX9HsWlzk3BwOR7Q4r0ZLelhkELWeoUBJ
mQ9ACqsoCQcD7k0vX2bNDbPNgHLpozDpWv+rtnmw+SYG4vZDO+cfddR6gXZ9xfBbPLetrH9d8cjw
v6hKtullowi44Fq5jCr7SO7Phwk9AT9o+4DyklQVMkFAV7vxOTt+yJi9LBd5lrBTZ1EuB1Ez7FhL
ZHglmChHTltDbwxaAa05rlM9FnBY+BNPsIeV3BYV+cSmCEQg4i+SGPndByeYKK8XzltVEZYhD/zS
XQKtld4frGBCQiYrkFTpq1lNE3ILUiiISAwkd1dwZ1bDSgTAVZ3Lt4eSVowPevzX8olqI707qPDe
VYnmLIktIM0c6Jx5vr4HMYqWgDCERqco/A++zKTBhNkVI+jFegyrVrjzGOnRCsVsZKKPNKfs0VND
1dFtyXMlpC5XvGFlEjnsd4PL2Rj8yTQ/HmPOzurR+QNRd5UTIRPrh6KUvffb12NoY9cHRKQlbSoB
9lBbn3HBeFyclLdQQO7bSB9zVz7iSQDcFg8DnFjrwEfIJN5lg7yuLPppiRzxDBs5P0GaCVioV9ir
a2L1RiqRVqNlIs0MARktrhKBwcJc+bPcVwaTFMrymKCMSCbLgj2M+OJ+kKDI9iigzyYHmIDUNTAP
GYQQjZgFNqgBbO/6knLGb8P6imU4h6VKRkWPPO3qvtcKSbV3aOdBPUc0zGaMLpM84t075OK3e3ic
5/HKlKgl5iYYEeBW4feJo0nT1rGLxJjcnKrZJ+dcR94mYV6UZMQmRiADv4MD7ChaDsFjouw1e1Jo
B6nBY5GmV7lnUphbcIrj4IaDJEeS0pZbgi0X7Nr9SiX/jyKdd21Ub2fLyzRQYTKUpHDQP3eT1iJu
ZRJddOOclbo62PvtmalY1WUUWgnxegR+l+TmSWPeT2AXg1e6g+H5Qs351PBaY4X4f171QtnaCmFm
RossfFNX7PsKm7F6DuEGbMq9bQBKV0efa83XlzjrAn+JzGv28w07cgFJdFNEjaLT2yWIIab9+tQG
xlovMzm5pdWPZSnOV+8Jputvccmfah8itU8j3FfQ6ZzdCnyiv0qMBbbgP9qOP5sr1PJSNyB1WQW9
cMw/UyHWDrqxY4mTYhBFccUkI43vEx4YYIFCk0dXwu6wJl0aHJkqnUNyFIC+mdaBl3mnUzd1z7L9
5FQCUA1OZvkaSfugQpiOKmbHBob7eB1lMAGtqq5TmX7Nhwj+1Azm1k6kTewQsM/MSaHE4OpExx9M
p0oQkqTld6MAbPJg9ijUknV7zS+wCIP6zRd3BO0R1CVyHiAfRJxrnlFYwf24hcTnQ2iClhAK2jk/
UeFEq+hweQwgn7MHgFCtCh0XuMC8jNzvXKKa69pQiPw+TI9tM4gc/hhUprBjZm4Gb9ZaPwCSq6GX
mm1DJDR5qHF5yIaKbdXXK/6r/i4IT5IkUfh+T+GLoWQOULQ+Th5bQ+q7jKTMlDVGHD+auxawOdkN
YvnakwNnN+S55SIdBQ7mxLeOaQzepLwx2IbCqiGIFF6MrjItfdeKklZJEsewClNolleTUvpGOwwP
aVWvgyR4kT9mD94IU6zMODAFEyx/dYbjk3mrXtR1rt4KF5mPOT6vDFLgQJYmwOmCGkwhSLU5YolJ
vogjntAKelg+0/T5GjIVpSxicGYlXz4v/9jkglBxtZZZpdE0D/4Eo9Jg65Yz64a+JpD1AaB7X9H8
sidjWOGHx6OyV78vluZrv9Y7ktRhR9ugYAY8Z78bbV8JI+anhaqOjJ47as+ycKAHhov+tvpvfnXU
xOwr9pPkcx3hm2KmyesDNH9WbwP41CELneYqaMn8LH/sXyDFvgkUJR3Pso1RQSrEzwMH2F2QjKE8
zBwDxZ8tTrqVkerqqrIuhGDF9+Hq0rSoFtYFNeekYcDZcFIu5YjAM/o8jskBbjddNjcuiU7dYibs
niLSA5O1J+ZeYZtOpH5Cf89Sl3k5FSrOCItB4ehmW4yr3u3v2DirTl/CgeC4jyAEcc8cxctv1IKf
gnPrkqLJLd6vPJwc1AX01V62E/oxxOM+pYcLPBNRYgpVzlk4TW9vRS6uNjIiRS93mAZhrIu0n20c
3DcXrTz0N18gkoRxrNY71n91DYm8q8+KTK0M6F7XTbcoCxcYBSw8K3VVBav7U5gpiBdb9/+4n8ig
7qOTD/Ma3/+ssJguIClgdo3AvwcEplwKcg0PPBhAafY9SkV7vStV4WiChANtjNYQ5tMQxcCvu4zc
JloEEZuA+OVZ+krKyhmDcFGgAvzPw8lXvCrI/bnVRzeZYnr8JJKkC2VoXzO/BP0SIyJVeoxPxVaL
OLWpP9OLRKt7E3p/slEnsYHwifxfpQchPO6ijsl2jeS0kCUA/mwEbV3UrRcrqAn5VqdGvR7g+kXx
JTj4Sc1PTyiqHm/FNRxMN4LRjB4HrX+fTtarvBH4DxOl1691j8CR/te4l6It0LTD+DLRkAcRsbxi
K6dy0nO7akutMZYgh4Hv8eQuS+CBXcrGUlj0iTuzON9K6mlg4w405rmfUcJp+nlE1+XHWTyqJR33
m3HqbvpM50akFeMYtKlpyFOh1g2HAIAqS+315O3KaguVetZm7g7jmCxngfC4DDeLMvhqpnLPhtgZ
Gfub2qJPnKtWP8XsBRAAd8YNgfJ83HFZOqkBJBUuJFqB3agiC2QaYbVVf4zd0L4skSY8UNx65wiH
2Nkp4eceUOsXSpB9YHgEhb1VfqZ/RTEUCjIvIjXOyxlCjD5gmxI/diLl+40jpfSnIURV2LkwOOng
sETcahRHEKjMLpBc7n0Ob8xoXsOcvgVXUym8MElvztOkRfzRy7iJ+BhgMHt+q17tDeBBkaz+FKWu
r8dNfPdWVY6nptbKIGSr+lC1Ss6ILeJcx+VtHUM1w0Mgy7UTACvULHy4yaCYMrzTFKF72B4rIBSG
Be4oQwxyLhQ7pPsvmxeOVGGSKOePI2m9r2asxSwcx/DEJY/KMHXwrdS7zM1Zfy1SKplIg3ApgIqk
fV1sSiMT3p4FwIATsLRoFLa8jlWNIcMLavot2hBu/sU6UYAj9rkBtQtxvEe6MNi1fs2Q4R1zJD0T
GEKWqnLo2TMSunXAGUImHNZlN5KxpaFkY5buyplt+nJol5j1g78MRfLbxMHrq8BfPCDFG6/Zv1hb
5lKM+LbA7xhFecjzyf9vovv5qnJsAgJz1qtfn7NWLc9qeBmenxfhyUEe0XTX6wWQyX9rNBcAhmmE
8oRAlHXvvMYOuFuBZx6LW6XGAaxB6PVPLuzrm/LwX65ceSz6lYyc1DkLBRjk3iKB4CQZ1cTULdkW
5ZcMwShqMTS9W30eiF/6Cpcaz/RMsS7iu2ZlYUMTMt7LPVmwsM7vto0S5Ola9UlPEbNr8nFtcRmO
4LIkhZH06mw+Fq9WTWVlnk6Vl7gRPVhhbDEOIQKqvzSYhmLtFzbJ2/WZKsAmt4QY8UOVHXN8xRhj
RlycY3Xybd14bNYMCyoLjr0kBzGiomlcR41n3b+m4SvKjoV4tBgabVO/ssWz5eDIkXa3vqVFXjZ4
8qTB2jsq458Uoj3rJhoQB/j0zaTrcBYxceSgvhA3sSi5/qcWkhaKpfPQkMja3yBiwByLVEU1KrPa
5FDkydgDP2RIOv3FjuZ+PBv+dbnqurBPpA9GE6/PYmVnl+3tJ52ZEqVppskF75z4gbQ1SdD0cA2w
a/5EzLSbRV1BwlTlEsLMyYSX5XD8KdUTg1/82aUSzDanGvF0jAOf7EELr5P7540WTcMX8xxXj2GM
kWFGBKrHLZP0RGpo1yudjVmmtDak7ehAEEOhs/9F4SsBAjzrAvi6hhVaX3qxycb/3LXnEodgTnz4
sdWLgzBonJJjFsL7Ov8WjKUSIZqiAyOrOB2B4B58VsUKRyswTtTpkFlMcGGkN7pmr4j5Mif4XRT5
pynEeFRovFpuXIlGzg1eoijjVn0xAfMpL5mh37aAYyjXZHt5M/6U22HhglBXe0UmgyrS2MagzifJ
XRtdJ0FS9h/NlnGPHGYf9YwpbjEjaAE5v3Uo9lU9A+MIIARsc5S/trFlbNck9Uu1E91J8uk5T7PV
FXUrqoqD2L7DyMWxwxVTVQ2CuMs2C1WNUsgyLexX1oWiiZfsKKiQbQhChQRJdkq0Dk5rCAjopW2l
1WeIO10boK231vrnhQBFDx2nGW+S/SHAr3RU6W0rV8idjyhfEFRU0n7k4KaqmB1rEMcOF+6RBU75
4Hirq/BtTdyOR1B0VgwRVPESjZz+mD54fLrj4yQLfB1QMK6iQR+g+ZOtyjdZsKSIZB0aa5TKHhh4
J7lybVYjhFns2OQZxduh3ftpTS2qCze7oMNb5j6MOdU67FFAdpCgrt4tV8ZenOqlKx39KYgleRjE
q4UckjnLYozxJNPTYmJYe72MqK6uR3tk3M0t16L9dUHUyP8igrL+prYf2gmO+ZJyRljuqf1hkJMb
l9aUr6w96FI5/C8FF0WqxUgQs/nRxLjQmYeEvViixYRIIg6L0BrwdaO83/pv/JxA1FCYfiuGw635
DjI67oTpwTTZqZ2dfg62XYaEoK8Qn4AQgdV0efs805fRswJQvzvGzHkKzLCCViZqhUPd5NFOmS1R
vsAbeX8KHdJoab/PwYBtw6fuqqBcA740m/vxSEZ8w4ONpToosan8/WxDSTdFpXSCQlABPrbv92Na
yMPIXPQJmU1Wt4IKqGKU0GIXnpbDVWgypcvUf42Vgvzk2rfTmxET5w78YT7jhg7I/3oiMEuIRME1
ZfKAp71cQn4SqunMzMj22JkQplauQ4qrifwN5n38NMWTH4JGMwW0t97UG3QhLzWeIglw7XVIA14z
7Pzo0kUNBA49zVmm5r2ztOukSAxRS1IJzJk47ienMcWDkHOX6fSfcrnTr0yOvNYoupcckAdXqpNs
xcBa46OljmWByUUm+q6Tht7HcCaTaQdnAmaVCF9BAi23GP5tJfQKmwFkt2VwizIfuMRP2OM+2Vvg
s7Ux/Lvzr+zP76oPnqDeRldS34bFfWY7+c1fiGm7oWM/V8ObsuXQxzP8F8z5Mz7X0kv74e2jOAml
OR6qJQLI2PvMnPfvzy8uLf1/kZJbKt32hOke4/yGLogsbmKYyKDm6GD7CjhwQdx2wI6qsdvvB2ww
2dwhGOQ5UlPZ0QRudYloUVPvEwTkzAYPf6fcHl4lKSpxBj6v0NHR04G/Q4VkBg7/jafJFuYbqFDM
Q5VAdSM5nBOpTzHKlmrunbbGh2GrCT2RAfFGjfduem38xu/OmVix4h+RtIOEjpCsdMu8N6mOCrle
1nnKwMV+rpvzJYe5TOswU89x6XTYCshOPJ8TTRmXAtU1PsCFu+4yFADXWrAD3z0i25P5GCMt4eXJ
khpgqEyZlzLtCOV/3ZQ88Nbz5Ab+hhN2XUY/tkf+hj1uQgKEDa+biAgE7Nuu+ifIC7HG89BqaLNK
NsRXV9YV6cO/sTzZ1CjqYromCzzA2kM05/lGUXiSMcKq5MKjASPCVM5edd6j7wCq29N5Oh7AFJLK
mEYKy4ZAu+1BVGFMBXne5ahCACw4L5T2KpaAJYIlefaFE+pg7vlxV9p/vcE68tUqao8bfl5l+lyk
jAkHG8TMp/yB/hCWWb4slxtGRy0x89Qne83mQoGPnnvCWPo5bQ4YxcLt2x/PmRLeghd6mCejVyes
l5kPKo9OPSskiRrjArQTg8DXrbk6DxgEjKTuCk3440UKwz3vM+2qqGKBz4mB0+Ue+SH7ERL9dB4/
8lrRD0MLjNcihUVbrUks7BHk7qRKptOkYTJen/ahZ24Sc7V4yJHjgX7wZNeGXJrBIk0svw+Hp6EO
HdVa/Gspsoqhl0tPRW+KGua1IlZaibtfv+hSYSx07Clet7KPhFVXk8e+SzqGDZjBrN208YJI7ecl
zxsmtqj5HjemhPsB1bJHE4+eM6HIMMWrjg6jKcBfg5fcDIoTUjBM/NmfWguETslxDOhUmYsYcWHN
BOd0ZtWyHmH1pBH8c2JKOKaC/gxyBlCjThAlzO9d81oQrqsRopgUuIkwR6xGr5EyiyRyWFeF459c
vhKBRndlOPMCYjlh1mbrpzcjkWTxhLOpSxWgdqTKmERJNxMpdt+DISkOsaeBHKjG1l6Jkb2yt0S/
tFYBQRJfnpBICWK50+SkI3NdCeiOWqMOARIG7B4m9WrApJpN3qwhHh2PAcY+OJ2fuiu+HTvuT8A0
Cmgg4swrI0qPdKkpQgGOd0H2tyvmitakFQuySE2PRthFOVpxn+7BT1DibFdlY6UWtzAUpUDCBJB3
8aCNXTRv2whEmyiv9Sr7JzprQfnrX857twuEbinjHdpk4O9GIzT3EPCbDNFkTFed8Z5dFmSwRZqF
cWMpsQSHVsV/QG2NgC36MQzfm4hhaNf+3vU2HJGXz4StCxNCduyDAe5H/CRcUmFegMN+9fNwjBUX
Rhag1fyvg2ofFwDtRvy/0bhOMaIUAtgrQZn1c+VI2gcBHlDsXUKQA53m5xxkUGhEltne1BEWjPSf
zdrj2A25oM/unuvihQvqbG9HdsxfoCvKuSS5X5F34cEbU7wr6XYr0Zku6Zu13k1CuIUimYCb5HGB
Dx5LM0pGjPDL70KaENgZLYjjobzJevk4WAEd1777HksslzgwcT273ZCurxQ7ItEmJEeH4pel9Fhq
030dLbdQhSberH/o9HxPAo763dR7zEEfBpXpTn7AWRjOQqraYSe4LSHhlSeHESlNd4d18OQuWYIB
+p/CxE6wBfns56CuTPTTsQJjXPRuiXRviB3HidFTXQQocNqtiKf9phTLhsSUl9Iby1YfC2gxVrDX
XujQj8CltoSKJmTany1m2H5f6kNb9UHQRw6eKX5HCxLnPwhK5AZrd+Do4N+YvPqd8Dth1kXjBvR9
t39bUwjbD/hLmxuKWAZsCGiRrHV2XG75PfbGfBuLwFSFOfo2EsDG1/nFYzEm42YlqGUCdyOzB9Jd
RPNnThDjPJgaXMJtlWgPb5vJtxo5KFouBN3m4wL4bfgZFBBnAHTI5gMXTuhRIMSds4P+nDLaGDAZ
XpPNgyxNr/XOhyyESOFyMkhyUa2fiRyEhsW54xa6eEPC1rXytUu2OjbuQaDXrEQXgEbIBVoliNqd
Ly7t/t5rVq56wT7mbbJa0p8xbEfui9kMAFk+Yb89ol5rGFtyBsBMmu39cRMkriYABb/CGvm3U0fa
dmNX5wBuRUOXAIZyF+KghEvOoYHJnj3xUiMQIVvXysDjLo6FxYoUGHv+orJFtPcYBWb/LJuS72uv
Xtr0xT83ZX6PNSJ0lRHo4iZbDjkdNA1CgcOCJbO1FLEZm72Go9+wUFfPK/wYfFRFPJah+ZuiQv9b
HjRXiofvZl1JkZAYHzhzTLUYHKTKrX/gDk15xEN2RGhd/x3oIFCWnlr36n4wNcN/9HIep2Rs64Gs
KJ91E4HzucwvUdUeuhEzNE4bUglE/oIB6WUYhBDy6Q8lpN9ct5rkSJeyuTUrwkDcbXHDIn3sitlg
KLkJKu+B15JI8IbVdpPoUwuJ8lLhCLZLEJlCkdMP1itXCfqUvcT353esxXH+Wyqos/TcA8Aoe1UV
JkEQ5UTqgPwBLu9Jb7SwrgLCT521+EAi31IhU0B4XPm2bXGQY9S5/tziztlDDBviDo0nvXSNIHIS
Q+7Ywfhz3lmkH8+uGN25Uc4FqyTj0T3484YwbPgFzZd63xjd5kNi8R3QsHHuIKRN8GfavP6Pyui1
7TuBeipuGhGGyRYa+8iHbGKPNqWt6oQb4j/5N5nA4OotNhDx9njhDi9OmHETCDToI6Eu24yoYuk0
Hqa4rz8SYsJYRDsl5tBwk7txHQbfAlEHYn6WXMX4JbqFLoT6xkuor+W5Wv00jOQ7uJnitLgAk1Da
MoIDs+8hQZ4Z5YxEt6Hjmn1BqEqBdCYTiKrXQXvWpDceAfDMbHJ/w/crkNCS1FugCWAID8x1Ei5M
PV4SKl1i2jIQyrwqmgMH54qj3SmLUhcb6pzyQjMqTFjKUGP9P2yIA0hjfOSpHPF4c3sRotz+8Ytj
xgmTMM/7vquDf5Ad0r0Wpc/bVoZAEnKOt0eheT8jBkQbtlpgKOMxfOjCwAMwvdRGRemsdbKdbSoh
k9mIy67xtpuCB+FkHjcoiF5feziYW6ypGj+onK3ib3q0eQg84NuJQqr6ZcdfeNNkAyraCsEAPFx3
GqkW95/j5Sb570DQnFoVTLu9+Sji2M7Tf94HspKsA1l3rX39eQQ/4dbyWU8jxcxED8a8gQn7mOI8
RF7pKXdTneexwvRjigIJ61wVawn+gkSsat5JDQsENOg1HVFqlVh2ZX21rmoEn1sXW5JLKYetL/JG
rH3Iw5/pYwsfdGZ6cN+nG1lKInEZ4u/LlcLtoHiS9gZMLznZe6eZDitYsdo079EZG280UzjQpNbE
Syg5h1aM/7Doyki4AL6UdFZU7cT0yaRboZCjso9SaPX05w8rcSJgfVJrKpuwvpAcfH0BBMoBQzuW
5lkRGVPOjJZ88+OCCl8nPPPnXwTEPnrV0K4f7gzwAyahKfBosbqd5kgyjaE/zYMlQrmTyx8gszLs
8HPwbYn/DGW6pXhuI44svZ+MHi8H4FnxSZZoW8Os30w02gCeggceavr0PZpADLeQAPVnoc+tw/y+
qakDxCX5S7wVR2q82eVEX2a5PRLORicKNiGG5zCFYSdfFbhoKg9nSb3WFTHnl4oo5NpowIC2E/hk
wLwC8y7WIot6TTn6SMrDr1MOG/+Rz/dQMvr3BnKJGWXUxeWnQaAEKrqd4ceUA9FDMzNm3MBYUHnp
6ZBWko6+0cleRJ7HPK31Sald7fMfTLUCU5HQMTykWQVJ5r3WM+1L7DJdHxXczq4eYEaIqEBBLanu
Dsr1N+AZC8XSCtnCfmOdaWQh28KejdLjp8dM2Qn1drY9iy2mGySU4w0FgaQJMTX5u8+ewNCKAncx
hzNm2IHNPspy3QQvWHoa8nCZ4l8uPEty8Js1Wb6Ek805/3EMusyeqKCt/fUY6MEgORFo4ftpRqfo
RToHc6dB9bhrYjmcZSS1Y6Mc8hVO/TXFlwiIf+Zex3kbfIJGLzG74/2J6mGCmLKFyzoDUVHaGfbq
styhmo4rXsfaQeop2lH31UbCXs4rJVHwAgXhqCCvQ5QL+CFobV4qg8RjoSs8sMrrKggojVtNI5xP
kKcdMikC7719Z7S/jUU4a+5v3AitknBQ5WhizdcEnlq5F0cJwa5afnKQMywFll8u9mwxnk6rNjcz
2Q09h2WggzMDzEXfWz4RfhM80xuzkE995Cn2B4ho64Pt+LSgNZvOiuPFcP01nOA73s/K3tSbm+8s
hzUCgD+kchzuk5+dANRHyWhATZZ14RH2DvVzUSsL354ELoukB8c3vg37LgG8GvhHKEr75joRAB7l
oOoH1VB5W2BSHgm1zDsGAHVrEj8hK/RCiN+gPY0K8feJtRXd2bUzBajVKtMGJ0am/RB+KdfBOVTV
BU1VNwzX7EZVAPfZml46mrkxL4OximXHZlA1nN99Zvx5BugBeRo/rTTK7CiUbDiJMX8NGcnU3yrm
PUjzgvvntkMtUBSO75mfuMpkM3i9l/Pb0gNYvCEgP1TJ/evY8Y1W9Uz4YT9VUUAS6jfuNPo6YWRp
nkriawfO1+RigBWGAE4VVznRPkwHtHvpyziHY5dWMgNAvgtDyBpDvil6nuMRWCbJ/cPYZNiuuUW9
It6SiGyy3qVNq+QosKdpqg8YqiD/QYPfuoZuuUJBEbbVn8GfRmIjuUZxRZuDtMPbcqJNH3gvDiEc
iIjakYl99VzPHIxUe1qjbD9LrEIxTulBiFx5vKI71kUwSCEwrAnnCDHiKJOBgXh3OC1C5Y8rhPPv
A2jHK5fDCZEsRit16p4SaDAsNb/7O1m8MhMkpA8J8uH7G6hsS870nfBfRmb1iF4YJC4CaKFa6Bfg
rGtBm3CsC9pwz8KQjX7+zkqMgagAbDvIXNUpshglo0n+AIcW7DABoRMKVJLOGaLRonJs5U3tUGqP
9eVsWqCVwRCXyn6D5czBNTJmPz4nPKqYe8HRMp0UXj4fOgeGgSvtei6b+rYJeCCf34xgbbcjkCJn
fHl0x+531sa7q7snv4kRYAeSj3LY68v1ri6o0SbFkcuFoMJZnGCMYxaSB/K9AUqc0ARDFw2CEQ3N
vvXV+auJoQ0iBj8eWUehKy7eZjg2cXx/XXJNsasldCe5h6GIP1iJh8G+jWkFCk9xN9xPUyhTWDZb
Id8qLYLU/xLLgQ5Pr7mIcDM4tLZ7Uhgt2uOxrgrGuofgnvCuXH+qENZS8kJ5NlUxh+v+9B0JnjCT
SG8fnhEYOr/Y6wouJ32ZxTCXu+yKAWBnOkscQe0IjGwELWCXY7mHfLPGj2nawlxecMKiLEceTPtV
M0Uy/ZS3hhDQlKm50kylf8RpEaJgzBGjwAiS8gxgV9VLlCiSYgVsr/SBjp8/4GH5mn8F0oa9+gn0
qrqZnrYiLqr/gQoRBH1Ke9xBYFrp2y+o2kH1bUf35dhJezXWuoh2SKslKOKXFGzcMuFqxuQBKz+7
XeYc5DyRVNcz/0lt+pIQd81j6kF1kXGXllHbfqV3CZ/dSusWluBnsmaQAqKGoirle4Ys+rqzQbTe
eVvcgDKMUN9LRUFNMx4du+Aqo9CYgUxzPK76/gcleVuunCVsH/gOXLN6fbg9NZ35mndznR6rjQbp
x6jWRuvXErZ36JdoN9GwpvW1UXmNSmA/TVSXQE9TF/2LLjyJ9fq7rVpYhF8IxOirQS7S6jLRgMti
HWUj+flj5Bz6XGAvLB4i7dzYtyuDE9072poDdgXf+TDGXV3/UOgko4Kt4pTvOpqHWLb9CujBpew3
7LBFkmIhvrnlKg3DFtkIrLlGrnb98Kl6+ZoS+HwF16c1HCHTs7vEQLoj1PMxjkSBEoSXdcjEAcQ3
QaamIM0JkKbrI3QHVOkopE7mdEQuPqowpKau0KCLgTLcLpj1B5+OSUMi842apfcHE1cjYegYShNQ
JGPuotRCZRmEvKMQGLRAGAHwI5QVZatHGphGvXHEXSZMWPSPUP55cnrDMDVqCeCGAewJhe+3MbkK
dCWcG3kyP9B9oIvl4VmjtGo2TtSTiytuGA3/S8nPEbpcmyXZsRKkfuLqZDIaeGgOtj138rqecrug
j06NGCddipJu7Nf8T3osAHnSq7BRKjz+2+lKSu6zVeho+6hV+RfXMjhLBaY3woZJj87B3yXLpLit
V8P3N+JTVM3/YGImtK52wo7Nlm3A5T3ImOhLOFwP0+LTdchfVxfvVoEg8dhVQ/IMXrkt/CZC5BaI
2zLX7S7XCsTN8dftvy6zWUS1p2BzF/Co7UDxy3RRr/zEpJoobhLTPpf2/LBl7il7ytkpoQOumJwS
KIqR/gl+r6iVX2L4RRn7pg6V2gueeIXAAhhENQJY0jvjjLmaQSw5fP0f5Qs4cr3P0KNnHnsv5dVy
rCfI8vegJnLjcU0Df0ucUlVQZoQI4Jh8scAHH8NumXVEEPK1MOLz89LjN1k8A9RaJTYi/ktQXWjD
4yVQ4qRmkUddRDLZ84hiLK71z0O+7oXkZ8ucQemv3HxRPJHEOVD4Ezx38tNn/H/uXQSQTdZJKDap
qv/NcB+WIk4eiLYK4W9yB+y5Edcvxvg0fXlf2KsQMVFxzKD/Y4tf5OrZj1vehlqbkPXfxfaf9NQF
bEJufx43ED7KZNhJQGRI0i5D9bVjLMJzrvC3DSah0LP2K+YdEUZf0uv+ZECCvD1n/Yu0j+6QfBPq
JMQRBjWIU9rei7B/xP8GN+8F88mlfP4POXF61MxQKAO/hPnBMItPcEV3UqHgbyoo47plInZEkh7k
4v+q0uy/J++Rne/BjEedUBY/tVP2JekD3q9Ng4JKwPzCj8ohaKHIRMvx63sb45BIYgp9ixLqqrQG
2unWBSgqa1jbUTDKay4Uxbg5J91UDpwlRpvmMEXQBVEFwhsv0xj/Bn0PMMckDsree1hln0C4QCfA
GQUKG6sGxH6YLOvW1up9m0R5lsonPcF8fBiYtl2BovneatjFO9yf1janJilGTXC8bxSmOHEyq1LT
7nDUOVuoNCvf7/PKBdyfRW1yn+oKp89qX6Xg+Aav/0KgJ5HUwnE7iybnUPExsmxHr0PNPieNxEnf
tf0tgX7ErTPBZ07fjGppH2zGoC1Q6lvg2QgW+TkdUSQV2yZr4BasVbjhP+QKAnH/J+Vq7Fc+21Jw
Ei4W5IlxYSyLS+gzMdhl/vmdCMOpu0wKLTewwRf2LD4N29A3sAUQEHQtkx6hDxhEnFCdPZYKDZqq
V4KzYm6MoEF6KQ9kEuzbOqFbaiFa336FnLn4Gth5+KeFHJb+ouWXg5TDwHVADUL5Cin1kV9Nlwjr
jf1VXS4pDb027AXWBFl7aHkqOIKrxBho+/bqkc03QKqZupEIOdG4WBxK4QkwWVGO0Nb/8ElmDWHx
BLlNzUnqfIV7lFwsjROBtwB8LoQTedYuVAiSJyrA9beDXAt/IzsB5ZKudR2QQL6AM/OEqJ7Swvsg
h5bDOwrvyRjpLFXyhz05lbhlNiQMCcXfb0aStUv+7XaPhM1iSdnYsnujXHK8W1HoyLWHm1O9ZJFP
CNdYwJCSmW9tMaiM8C4C09MyvQ+lnPLtoyBx/7J7G3H+u0K5tI6RNMAVv+9ug52O7sRhlAJveC7Z
Cu3ZsGb2hLlV3TRBiFPP4um5fnla40gfLj3oF56JU9/Iz+qo2EUHbzKHKKTy28PkC0kJ+1LpGHWW
g7jb8FySpndTo8C6m8s4kixsAW9XHKe+AmVdVqp3t1ohDlCgCHJY+jyVRRqPjqQVFQzy5rouW07d
y70/pkMKzVDCtOkrXBdY0IfxcNgUMZD4T7TFxly+svkSrldChDLnZpztiPqYQlC6JjOp+rWsfrq/
WuVilio1vxjSw0HFt0sVZIhT6t3bgxWmfeRsjvpDhHAo4lUYrNT+iUclJwVSOosznwKRwP638kng
+OEPq4kCRd8oLlxPR6vYCTwWMi7Np2oY7i6y2Rjt+7B9uro/HuIC2z7XTMkXyupAADAdqj5D7vmw
0xsICM/p4EI7ZI/nm4Wx0GucceWHFRSzGqVoccSutwoSgJWQZcyLFhIdD1Jkw6Jcau08lhlU6HXp
GOfd3jycDkKmqKMyvsXIbfwTF103th+oWPnFkAys0WSIguNC9PQJUqBTgM7+98Ro9pl3ZMcek9BW
RzmKjBk3o8avsuITTeudJMh9FVgbLQH4A7toeaSVKhQkBdkk6RFMTvOvQNFhNRmEqNR3zV2pdqMc
mnizuOAEAiJrh6q2l5UIERtVOUDPDn4GnzGfOxe2/t2UEE258buSUWQ8Wk3oon02MRwFVTVlWA8i
H/ljnm9dHzfyWROeSlYHxQzX1b0C5cPoNaHx5kfH7JDJrYl0FmQ25zpllUrh8ALC/3IdBeSY9bvX
30FCbr581PqBKOJOZehfSo6dcShO+j55zYh03wmhLBmRp+Z8DTqd/C0nxwvbSmyks/VyBSC2k+8Y
MOZhY33INhtd1kc629TDH5OVvS4vdR3S/j67bmql/ipBTE/oiz5bJBDJen1Az7u4fXOMPbH/vVmd
RtC1JfxfjUMP3Nmh6KdFWRFwUWCfEUci1dUAwU6bURC70JRUF8/ihf0umIgbFag+4oP/9GNdhM9W
aiedwIKy/nwL5BeLgcen62CcBqkBrgbGhi2aTLGT+x4OaLSIWMnzmN5devJKA7knnAW2sNzylGOQ
wsBQFLruXmvxLhbUyDpS7qfl1xauQdnFA1YF2Fg0nUqZ3/6ffv0Mnoi4rkmkiTkhty5o72Opa/TO
Gmxvc3tSZvsvvYvA0KmUzawOTX/iwyT4fNZxLJlRGZ36nvuMFUolGVX5NvL6rqxZHYBPaOKK9R+Y
STBTVdZPPPq+M9D20S5P+gNmR/ku3jxazvwJBYm4IGK4ipp12yiVSoAZkQrGQdnUSW8ByQOmaJeJ
bM29BPd1xI1SHR/emkCn/QQfDvGa4fJbWCt+r5hF+PEFocPyLrqOBjdTZz6wssW30s4FRBSa/bx0
299KuQgMmlYyZ++BM+WDgZ23O3pkUBtzOpoDRwiUJrPqhC5420ZFx1vXmFYI8PbQN9EV+hDW4NB/
XvtHqIZv8si7P0fyEGNyRyaAU5be3sQwoGjhw1SD1hQ3GQ0S3mh3j1/rlvWZH0WcqhcVPoVMtd/u
og02F87aiyYcoo6oUOeZ84pnKrQ2Ur/hIOcx8Iln8ttdGmKN0xbr13dywjlEICMxK3xn9YdHbfaB
qoWnLYPzdX75GSrMH+XJUGD2m+7JEpSHoNCz5dYT7UA3YYX/nDuMoS3EqOYLtoXzP349KeTPuusj
7fFeq3c0hD3DQP6j7DP05M5RujiecrItN/yjTI8JwMLI8B+/AI2DSXR/gj0KkW6jaoruAMpG6x+0
/n9V8DUAZ11wgTQPQ99L24oasCenrdadreI0RyWpwYxd83CjqeyUPHJkq/Hf4Wi5z8xdrt8HrEJ0
jzeF7aE+BybVBWu8r/aFyw3ycz3W8btOmeN4+QBGQtgNrR65lQPJqjFbMaizzP0BqSfrRUADm64M
RV8xuPWCOlaC3slLRGUaB9Ow2u2XXARilwhIxLMhm7kvNap7FXXZKabE32DomcoabLgdUjzBvrrv
ooCghLwazkMbVkRFgrszYg+eiUiirwFziYv6L7b4Nk0XLTHkBSAG4Dmk/6vxYclKxz6DzQwZCTJR
XoWq/5sk5c0w8VQH/xofYyOKN3iPzRlcgXKjy5U44KrFTgOI6k5tNhbwSBnHLW7cK4pgMEPYaVUo
62FhMHcMUctwjnaVIIuSwn3pbgFIEBP+3DILxXDdYeLd5NivtBkfvUVr05fjRXpuxclVTKzk2GcG
1dcDfErbIwDExBzKwTVCCEWdZRlYt3vo+nVTtcI4OhsNjeFfVEj0fbInvsOW/eQ+fUsxxX0u44Fi
nraXzeeqPINIMjWbkRcfeQ5kJ/Q6w4dB3TFuPMHt3vnePrDk0o3bu9qn6zb/I+xnSJnfeZ07oR+e
xM0KJAi5nFtcZsG4lXJ2G0dwrstBQD8dK0deuha7FnafznB1gqqT22PpajGIIuyn5/XA48NEYt7X
CfnrZl6lDINriyMdXD2XGneef6P3/c6H2H4naAkMAJy/L/C3bHHyPkzOJ7p0P+5iYh9puZuTOAIv
nF9Hsxc+7RmmgdtdYyzFluNJrbbkFht3+/CmjJ06jO3bEqgwqBAxI3DaFvWklZjDs/95FJkd6T81
3VHhW2TM2HthXmdm0Gf22cXEVzJgxTPns/eOd5+ZqKfPA+CHkbArQ5aKu2gTLu2v1khiZP2THMqj
wHFEFvtjgIC63sZ/MVoWwjhMKkMo8SYoMThUlByLFr10fuA2H+CvOQJbRC1XsRuBalex0ivEydb/
4ha0hIbE3MeK9NC03N1c8h6HfG9hgO5E8veDGXrV3jvsKU3ZMkE9vy0nh5XmrnIg0O6RvXtjt96b
ioxqaLi4PiloooDgc4nJ4uEwcuCSdTJndWd7JNlXcIvZW61UpQL02i45z1YEHyBgD+NpXOQWvVgg
4lsQI31a0Bwe0MiZvSQKN9ISM/0fkulDPZNZnm2sNH1dQ3utufF6HMSsJ9sk6vmYQzVCSEfPylrs
sEsuv0BZeXBSuyG4BMiHddzJarfNxR3hm3BkpgeVusuOxVvPK098KKYHQNQpqKBbj0Ia2AIu1SqZ
M51xnzMEamsRMsiOB3t7PQfrlK7B/5pxY8rVccVNinXzKoKxCaFu/I3CFM79JI4pMmxiViVo/z5i
pU4c2FUS+ipc2bQQxg1543w2j+J1gANMYc70NoDxXDcbEr6ZGTEBFnwcYjr43N242jP5MWO7N6uM
0iHKGdg9rs8VrMaGAj7CjYqLnEh3v4m7ZCLG4LAuzU0zpCOOXR+T8R2nHJXqZ77W2ERJW8xEiri2
BtN5kcjScPmC9dko0mdM7HY8jDx5fUgbphLKcECSeLR1Vg60h/wusFUwBrATz5hsSy7ttAoHisE5
DD1O2RIbFBGlLvt/j/TWVZClEfn55mQvI+yApBvn9uQxuDdymOzSv41FfdVQNDIKojZR/OPICM97
A1DVI3jvFDrNIYSg/rOlqmEufF4FV++AhRkLFnTz92xRYdUjzFanMtxMbGTR2cnUV4ob0fikX/Bq
qKhqBw7a2xA9nPuMiSfl8CB27sLRI9vm4CZOq5mUb7iAnRIZvFb9UiqHtZOU+n3CkvNpO1GYEJvh
yeN6QM1abAk0h4DppMGzOFt3+VnhlHdkhaCzMig/9SIuP4AIIjJK5TsskCUz5VsLTRHi9J2IKTF+
70x6X/QzAeGpPCBR4tMA+nQ3m3h+l2ZAKesZzKCQMnKqYmN716CVAdfdwq5ltfQjN0QNx6bz/hlb
bqN4LKzAgtmFJI76V7/Sr7nn4OdS16o0hs+cBYZ9PQnKVtNMOQB2UA5+GNiv51WluUfo/MzPJvQ6
VtDCAgDs8uZsjCmOudPEfxb4UMqc3yqmLErZbsmn0yClLLVri8G6MavHsc/OHsSLkVUNXGfh0doY
S0T2va6lhsxtDHyMSA5gzbZdspqHXJxws4CrJEH5GKuY3fQsNnnI6nPOvJCwWlp0xKtWbhcan80Z
q+IGnap3ZbtcEyuKnbGwprB5k/lWTr2EmrlcVtRNHjCf0C4IeLIProT5rV/xnCwTN21JAHIpL/Ka
fKacTlmdfA6QD+Fb20z0bSKJsv3beiuywQ+tuqaw3yHWUBQN9WrP+R/HO9CRZcYAJK1HncG8HCk3
cGGypSnDeGUPvUP9QZqNJLG7mSR4Anx/2JsDGMsSZRWZDnkiSmNh+iZws0UUyo2zuIgj4jF8FzaN
gi1bDx1RWsgPNPliv7uyQI5tOdah25tY2NT+8O72QkJwxxteyKeWyT+npLelIgiXYaXRd8K6gAnr
NwcStS8sH18qUHgjFW28rqDVqD/GNDW5AnxL4CfNuy0sZ3sa3CwqsZ2eVKQrWd7fZKP3BSaxnicF
pb943mOgKlhBya/FBTy+rSri0g9/GY0HqS4lrsHA37fj3sqM8xcQupqKIH4u1rWS3MIkGrpu47ri
bPsBc/pMja1Io+NYad2CsNPLP2urTqeHhfv4SdRHp8+icDlabAObK9TzUo2lCepntRGE9UgsLxit
IICR2sD7i5bBdTnhGUbJeLJm8v1yl3X0pIz0HVgW1vdWpOsDdLdrGyMTMO6V0F7P6Ve79utn8var
Gto5+KxyiwtgGy9qXUe9LebmYQytFSySl7z5cVziPgj6GE1YNnq7+tZBAySbzr1ibB8JruvOMLpc
s+PcEPYPdaBHfQwp3B+wCO1BZys5kbqTGX6qyr4ftQnfrsdhAhUPdThA9h4+dnxbNqG/petT5DuD
cqiL6ej/mEWlyLY4fJWxxf3kULhyvNn1w8puyx35fPlGqGyqxF6gILtfwo1Fz9kYtHsqljxffaKl
GE2B8o9LaAvpUMjH3EkAgQUtvOg0Ck+h4E4DSk+kSwSdza9Uj1itukxrXRHsF7uehqzJySnIrr3B
dk8i8ceSBdLI48T3o7RzbojgLDjLwAKBuBgjU/GWxyEQtUJgpnoxg1I9uQjmp6Hz2l0MydNJ/VJv
BtvBL8rWTaup6lZVwzogILYr9+4RVp/dlW6M3BNuQ+Z+dLjpNbAy4o80O3SDOB3xKZCcM/vM1SJ+
W1HJKBuX2TLUfX1AQ42U67UUdmtaewjC9yuapEKl7AEeFE55RAO85MTjK7j6o+FGyJASG4dmYDY4
2XQJhAjsUj/IAcKyE/IWLeuzzrJyxKGan4if0E/j0icLXyY4LG0Y5DfpkTjzVW6d0MTG79RFXGwW
EWcrPDf3vqwPmHMwy+DMiLrQpuwQULHzhDvvXyYAzKYM77bti87rC8EuF0M+Y96/gow4ZVjEddp3
bwlk3UtVpAPRp1MIgDQuYrOd6wXj/jlEXZU6An8m9pdojgrW2kOd0s0wXvFsYLDDpzsEFfh7lmmw
ZKKq3Rbdl2tDg6Qk7lfMbQsJN5mo9e151ugDoGr7l4ZFis63fVkIaM8zGz5gk6ujvCA0IOa62Gkx
1UTyOIza+RmPPQdXroKfjknm9N8dlOsjmSp7FSjG49r7REgaJVAEyAbBzCI4Hi88whlWsUC2MV5j
v7EJdP4gxmCEnzlCLOrOLzz7q/cyls/SR64PGb+2696JuxyCqdYRNLqcoUmKsOEXQAoSm3anVOXD
xG09Ak5/lcBtQE+796l3/Qc/zi7eIPI5rXtQOdC40QtaoJrThLR/2ANYRXIbBfkydQAfuZdY/Wc7
iA+G1UWVrD2ZeZtuFzNH6ECLkSAas5lim978Nee0aYq6gXec7WOU2pfoCUbzVTXlkc65585Bp3OX
vLAnWVAoyCIyEcF/tE2FkvElR6ScccNXvwgFQTYtiy/9ZYYlXuD+XeRckrGkeeWZuzUZSb1Mh844
5EKSnsIogJ3llmyjbmYkCJeptzmv8MB7+8d2Sfn8N5v6IddWTJAjpB8Wk4AjzS+ZlvUFuWgcTaCx
UcXmfuXNd5E6NxSjFTBdwYIVj+kKWSbQy2QQ6kxq9iZJNlflAZsq2SMFeRDD3irxuTdi9wKOc31m
Pt4c85nsHJeTGWRr2FDQPFrnLHSx/x4AYL8GJH1Is4vaFZKXWqxhAUmZjr5hi0Zv7kH+ckQSbRX+
SwXupHOE1jXaBzJ+CTvrxaFuz8a1gOPq0lI6aPPuFrhT366e16Ki9t2LqNRx6oVzIjNpojBOsNFe
wcH7JzctkmCOrjISifkAuCFX8yFo+2HfyaritCDk8+fCovt14i6s8i+zdDbR2r/iakgEP7em1S4e
QPjia5Gdb8p+9CSNqly7rCUPOcGRRnk7qmsK2kkPEI8R0ZablxUOR4Qme7LMA/lBHVI7Wr9Rgg/c
6Ncgj82XXYeuKJSP/zfL22o7YCOQpMxAA0WrXnomFPPXcRGtm4jtL6xNYmU+0Z8Zy6pWNjVumaD0
4PkRqV3RAGflQAzMmfqBUx2lIXZwd3I2wM0TWwTDYPOo1poHXcyCCgBmf0yBkApwsUspw4+Q1R8J
hJCscfMENdEZy2nmbafW0DEKQ8Q6Fmef8a6MI1teoH8ynJiRKMT2ozXfqKTdOfDdXtNUK87yYGwN
ORdV17fe2Gv9YKC2DoHzkDCBpzMhhda3p/9KFsCCot/ydQFhwHhCUEb1Lqb7DufyIbwEtUkJtbsq
BzuF1RNGcylnoUTI8lJJPzj/t9wt7xcQ4y4eC4olV//JkRoXmz9a1M5LEA9zhnQM4xmjlutJmvxZ
wyJdFPII+0qxf2oY7MBUouvK0LQki99csKuZftD65isa8kN7rdWz7skQ+PWf1lq6wf+Nl1ntVsR4
UY572rlzASrIQ5cDXXwa3F7kwISd4IAmZHx5dxhLQZ2lBNmVeUnva6+lHdLfH9dzK909QIcCZA6p
ebcPYvFh8LR4wiwoRYzSdtbmRxWPybvF5pWSQt0N+Rg+txu1y2VgGXYblhGUaTbJX79CncuapCrJ
cYkSBNKZpZbMvo0Nr0RTP6ukgMOcIIiY9me47FKPwO0q/fPd0FxMPmr0q2mjqiUNeSA8y+yuqw7L
AesaIZ5Kpt7PWuAbuuzI8wyCd/gb757bIZl8TfEHI0iM8sug5+IrmUY6LDPBNtXWwbQdBMYJGYV0
ME5PjE9G/QwG1ajJjhy1stoeJSqj9q90newTzNsxWghdRnzbTuiZIqImqqvY7NB2sDWodOsCP2lI
ccQf7jsnbczUK3afA8H3yT+Oz8zhFKAu9uMRW5R3+IQ/g4onRH3v/puJOGccRKJmMagUNJ9fFwl4
97xgDv/Y5yDFuwZ6sL+xDySY8n3Zk3Gh8ESm+PVWwTUHoXV4BgpDT/sw3BpOK7/u8hIfBVCcVDM6
Irqp3vKSph+c8uUWrG8fT82z+NNM87rgYPH0d5BYCJPUSeSSYsrI59MLs2xAylkxUPXEqwadvS47
RlLdebXPvQX3MQksgMB52sm/Sm6Fm1ZBGc8Qyj6hNPkCoRa6DQHjkFbLs3rDFMiC0sKhd4hUzjj5
Lz16ADVDgbKVOXv9Bnfs65Jkw3ARq5Bi6mEEb1czFdjx5QbfgOe6YLkQ21FmtMPPsJO+/2bkguVO
4G5Xuli/VZbrMEdH8eiITpWgFxKQr2XioG0rnaKaT2nImNVltHy0EH/ITFfv5s8RZXE+SFEp5Oy9
5IbzYJtJ3NzcRKMGc8MtOCsQjbyMKnHWumqflsFPpyQOB0fELRtKqxt0bcf5dtS+mMwW/mJV1geq
jzKeMytR5jefKAK9CdpZrEdyM1WNJzuFm0Dd0wDaynPXYPOaezEH5IfLJQbvFNnk7yvhA1WVZnSH
T6z0yXUy+sal79FRk4nHfGuP0YBIbYR/VOWyNXAXZeTsSTXWujyjxQYevlKV2b0dK0OA5jI8xdLV
B+gmbuxgYAwIWgtRL5be91BdZ5caE7/jZQWFltNV2fxukQuRaf0iJ7Ag87Z2z279EjRpk/dVCrXR
cplUarp7EYAyP1BYios6ASGYplXMONnSKt5Cu+Zi9e4L229rybj/ymcdv5KF4QxynCc9/0rL7Wsy
x+FHQKOUExnXELsnx7eAx/ieZslaL70HL0wbi6u7FnGaPpJTfhVtyFASMMoe7x9wPodbR1JOtpwP
7jACoFcZu+izUlxwY+VsK8TeiFE3z9Ay2ntHsuythNP4T/o5hs89YYX5GOouNWq9dmaVy8C+rpFV
RRZyl8nvjtnjTMG0oez+/lzPRk5+mYqieOSusVF9GizE5LkQM0eBniTTieFaCTzlz+vhRP9Fshzl
wPAsjWqQymU/Xgc0F3YYAtG2wB4M7JA8mCvnuG4UU8BWkCMTWNAC6j1v4ScR7KfvbJgYyXqlM0Bj
wPIp60EdaEj6Gn+MrW1rY1wrAH2dNKKFKXtMJZ8RfCI7aUWqqkaULFwTVDWyuuFgWguu6nw1xkQb
UX8W7AVewlVYfJpk7WWm5GvKgOQ9xuzaKar0SSMH7qzG/VkAjwXx9DUhdsuO8W3mZ6rOWLapgJZc
A0V6rB46n3pGkQMiQfxfwvGyQfu4haZo4pQCUjPfFxeeTOqFc2aFjDFLeNJOogPcK3crDeqJdESb
KhVd7+nMYtw7OOsERtNaHWoTL8XQlaScnrcYiWAu+OFbCGJG07IIO7k3awBJJIFnlodflP1rWNni
f6mn7j63d1nr3UpB1GT/oBr4b5ZiYvOxsp6hKLDLqd4DRmKxyQyiy7V46LLlXnfulQb+k7F8aZg8
yqAlamrwjH4v7RHOG3ugfKNV8Zvl51AiukScya8kxZre9jWJlufq3psWdQBr8+U6zNK8biCq1ifD
kkXepx5LbVQTqFkVGa6shAiXRfa7dwwKoU+8bdTaIgq2vRQ8AI2dLj/pECuZaqgiklX0hYGBX+Zy
/Pxh0pvXbZ0LIO8R4G06OVIfMbw1PO8q+HUmVzUBMJ+1+fcJFWsl8g2RJvy9qbz+PZd5kEVTIIor
0VsURmKiE8QTyLIuTQJL5iiHmqDIKXshAH1HvqTctdJoZKIAc/k0O32+sNnWGcvrJiL77J7sNus8
IGWhwgVnktGekErbpYhU4YIrdMPdCqkGENEsWD1gGELY7OpEbpRq9ypGOkGP2ke8SqbdLR8MMqbd
cI0kV1zxIVfRcNPTdZZA8ucHueUSGLSIzEQlE0rr/SRPduknFRpJ8WisVERIR/Lv2dT1b3lrRQPD
jpRx0tRezrmhiUV0jKEnkOlgDqU7TF9e59aty4mVRwm4tr0zC1qqy2Jzn0qSFZIz0SgUMmBfeIR0
hGifqNi8PMp0a9XbNtbAQNq9hqM6Go+PfFH1NySZ1lZ5Kzvjj+Rs6SRPbBhAQZyI6k/wF6DqBgBC
Rr2WjH8xjbhyFFWHQplzOwUSUlYDJVdPlnrWI7lGbaLdh/GVDVX0dUkM80uzTOHUYgffcG601YTR
IxBcd3REd7GpQOZChNY+ZzjuQU5a+6qZF68YvWP2XjKl0DZiRVkt1zkf9+JzIjJjs64MNUb2rtOg
zRRM1Xl4tf8can6yrsUp+IS6JrBRAIKMxpJu+IEs22SRK6iZ5wLUCDPw6SQnTqT7YqxIKizpPkmR
9ehWBS2Hb4hdiQSVl1/X7ADsy2dRgUjWnxLWaqAesO63zFFnJ4uZvAg02k2RbeTwqJ6wnZqziHz7
2BWvLztigGabrYvMamq+kJDbmovArftqFgVuA95Wv1wq95c1B7idaOc1/E8Nvhkb22dlJ/d+p9Xm
y5aTUfVZxWjbcIRo+7NIAPOmq/4yOUV+tLpy/ZUvRMxCZwAapy0s2lKZ+VDqpt5iNBxWi+Rr2oko
8a5XQ9rsLSCy+qeMAzUTUc03hlp0dvFqXBIMMP0Zl8EG8KbUxipIuouWUlt27dsdaRF+pLBuHDc+
KaLt+XczGRQX4UJ/YRFMGZmDqfobAJTdk/ryyfIRkHRmPQvqznTslF1984PU8kdqUdJY/O2OeBQ9
EQ2nMu9ovKvgrhTdEHf6sU1VGMEtFCy3FgNUu4/9Wvh/zmAU+nACHD7kOrGwTpsftPSnZu4OArlN
+7rhCdMkOGlBc7WQpFjMrK8sgpVeyqX2hKSq3IZP7F76/PWGgnPr0dQnZMf/E+pKHudyeNJExcGq
NF71oSZFpD7xYThoDxXgf/U739l8jkGATo5otnTkOfC5Qk2bWtxssU82+UbYVSoZBOdm5fnC9+3I
TZPZSVpNiXHGxjVjOEfwDNLRoPXxl0O7aGJeX0r1TbW3GhzhvrEPtGpar3Rr/E7rb0ZhIxiPcAsj
b/ihhhfedyHk0+UNx2mWIuTEa/fXDLpG8d0n9xJMKP3b5BLc0dNcfbyn2+Pv/TuO4k0NK8EyFP1S
MnyTB9/CdOVcMHIYS+1ej5FO2Lbybza1E0A6uWHWWLum/W1psMqmVFxp2DYuon5HGJPb3/Haa9Oo
tj9mgy2ftPBw+RggFa5sM4URbzYE0Y0JongZItMFhzV8ncduGC0xxEqkI7jZXcT5L4fSEIncj0oV
jTtNTicaY19rfji5VSIlkJuV0IdbpI0KRYKej1UKfnG1nYtTjBYJkU1AGuEupJMwNciYMy2r83bp
131lI6czgBUCK86jo8TdxRtatWNKthPmwByu9/nbhBE0GmzfSMaUpMbx6+u9Apyvi1oASKxRsQc/
twZVXbvPqE1uORah82/bGtxTphwkPr/u7PzgDJkKSjSqaRM3p7KXzCayVx5Bb+pGB/g3FhPjH1b4
rvRH9eBYqexVrBgnCKW4vuGROy/kU1bTlzJZ7vWkzxP4Eoc+xAsllk0XATRIfAKdB/aGyArwR9qb
LHZ4Nlsj2xYknas2pSo8zLcdzH1pIxiDoxyP/XmmRKP6GfHrjgN+OPaWh9WtMi9FxXCU1CdG7NGU
rSgs6kVE2q7Bt2o5k2FLKdjjYXvrZ/J6b9h5jzakiMQwRoI6lHuBNS+XGH3ZgHA/cJFQ7VKHqo+X
OpTF0+Ld87jIShzVr7L7SljS94cKsALcA64HYP5YZwv3s0gcOAVT0KgOJ0+qL20Wtcpcn9NoUXAU
srIjTljyq+EIbro1eZWrwkjVG4p1AZHbjkq22QKPDxL8UKCpjW84yooqKe6c7RU7ytAeDMb5xakX
+Rk+LWrgjp7OdFwrU91lIJTlRQTPFraTyp/7g72mUKms4r8eoWWhp9uIrxcxI/bHTNihoCXzl0uy
VBlUNGa5NnLvbiMiVBmfj7bCNwLBIN2O4tNv+GIk8Ih+JNh5kYbB9q+llsLivLw8nsxZxfcko9sG
E8uIU2cLHKuCmipJnq3/4pJkssTlNEnMoeyf5J37vfJWe6BW8phbCKPs1qOdZpghtEWqR4GuC0Od
O0WfLxegb0Lyg8TRniyIWu5vmk+e4JSXjNuhglh2RWTifA9VoLKU7q4bHXY05Gj9eEXVIN9YDf6y
1R8Qgo5aiDqZ+wD6TLNo7lmpwtVXFA4ZSWDQTKTlEgnsi0sjOXJg2epso8WiDpU7TSpwuugvpOH4
FTZdbDQNe/I66nKBNHXKDxjssYJw7sbSCs2B5dN2cif1G/ltjQXszgmPo3h3ZcfBBwEDWGGkdGba
7LmssGjIZOEkDP9s3/H/N9U3mDmIRd8liVcn1AGJy7Vf6sYcV0MYHr5N3v+ZVLdGz/PWBfcowWs7
yV3/wd7ZSiV8E8iLoDBAGiPNGHr6nIJBXMv4mD8Y4+im5dIc94bC8360J/s+SpkaQgTxXR/+yTer
/Pz/vkKIYaYXKwun3uKSuYi1hdGF5x8qSGmOacf+wSs6VR9s+YYWrpl+2P7nXS+XroS/rSudEog1
nGprQR2iQmr6CyvQEQQtAIQy+NcmFYQfHdt8rOQwNjbucFt2T/ITdWcP7pboSWtDPBN0dQ96P0Cv
OCWii/mNgo+J3PvBcf/J9o7IczoIaQ7rq+85e6Y92sXwIHPvtx2SzTlVzzJCljMQ1QOIuPahCjcQ
4cYG03u14GcBNlgChBcohkZy3Y+zvGweDryT94eaH3WfmCL5gbhF1JRb9OeqnpSzisIkCHfztMgk
gVqSo7ADSGW6Qn6oU4lU40/DAUzwpKRT4Izx2aPOlgesAcJ03GzHkXEsdpoltrm0H+dXF8WYuXGb
ek5htYowqFLC+iNlVYGQkYocXa4R/Nnk7WAVBLGOCRtdi59SILXvW7ba45l9l/CNdmMU4q60/JXU
g5BnyySSWYlXW+wuKBMSnmYT7V6+Bte7VQGwcwCXsjVLcGlKNWBxt2/mp7dXz9lM/gUma+RjxIAD
4y3vKu8BgGxFZz2TwEuYo9/J+qpWkTIjaoPZIxeoqGFi//PPl6TqDjrcoU2L97zwngC3aK6rcLm+
7qILRTO6nsfQ66bOpDc5CISWtsSqyzvmgAobP+sLTeuBRRgy6iUay6v9QoQIhRtib8IUjpbSfYJV
vO3ajhiNQ/9KPrN7mjUvscCF4r5eLsajd/ADpUB9VVChdBPK62UKDYdsnzU5ZT9NiBkn5oQjpfGe
PfssrtiI9FF4elzc9te6GGyQS60wU1rmn1qSy4XVbN2t8A5NOjIuX6WPbjEHAW7zn5ulr3e/egWd
ks1F2CsV/R1UKqCLDTJkmJIaPJM44BK7NkJSL+1qDbOhmMwhNioz5EDRcpMUaLI1nrkjJlg288DX
MFZwprXrDzv9fNeigYvREPpdxu8PIJUh4KcsrxWgbDKWdAyYqoz8fK89U2+cqmseAoUfiUkmaHav
Ip3jv1shx8cyjTbBYw0wXH2KZL3r32Z7bztiNtO9QqXQKuTVnowyEvEqEAdqnYg1XXgbXNTLWRUm
rYwbhFh4/IDyxfYZkyyCVmU77y64JzwbveI0fYcipdH11CJtFYT57WxI4f5mFsQvMeWc3LGVM6FU
PfTnREBLCNdYCfonLoCGtd99OYCfHkzLiE/UJWB90SZa7FvmDDDzVhxCCugSx+MohlRf0OZ7gOaj
AH76i6Z/2ibGHhcoGW73Yz7l2BFD/edMisxlIY0e4w4djRkccKRgXGcO3DELLXzaRfu6OQM4d/7o
HEIfp8e7wWVgk4GHKIz8IocS/UI3AVKBHFzRWqugSC2568yBlmJHBhGoUCiHLTHj5aPnptr/q0jD
kBRX3pMzdN5unpwwRblJ/02YBTCkYg8wq415OXTt1UdvWAVlq51BXgV4r1fKIjhG6Lj0mA8Ov5Qd
VK7YJVpAvVuEto9ZFrP84YdoGeBVBfZ2fRmI89ftXcwasEdSyp5lbEc2tT8E02Tr9uOLKwnjnfE2
D2PKFyB6jIvY36R5NbiKxKGQeB3YXc6RdwbDu4sTayP6bnyXj8mrz8Gfcfff2TYoJIurhdch8lDo
03ZENDODu6dOESwaD/pRNxwcr8eaPGU4aAK5raLA2CM9DlYjZoyBSeGIUqaCaZYSrbGIolUde5fH
OIMqMnL986/sTIknTYHW6PZSia1VSYNPKgXZndsXz7CSAsLu7FfNBPrT4y3F3z+uEvS6unBW7oCZ
7R44d//w52aUHRB2zhcwMruFfDSplEK8vQv/Cguqn9T/dyrMLvMrWI38Rf8K/o519Rf5SGir2IkO
FoHL3dSOhJOlw228kV4Qz2lYb4m4rAio87vjgVm+j07nApKorhwMZRau62rJDzuPCT8yKvZJMCH4
6O5/3dj158GZVDpOGEzX0+LtdCyQtpZdlcch4jKezuuaqfZ5HW4H3yPY8RiAI2nKPsvtTtK5OfPD
jq6OX44SHK1mFBKcYJSK0RpJ5IHUoIO4pBB1gg1DI63LEf8KKuXxRGJj5jHNM5GGsGZJmJIeH4Hu
kxeOWaExUkZbOokMYACchpKLS+b9++utXeZcTTbtWNLWRTiht2N8qCnBta/YMLrrEOVMmjoK6a56
6f7axqNTk+IBUHw5yGPZuYKbpX22TLIkvB/VfmTFqDQFMzh6IDP5EtNwqUZlp9HbZHmgl9wY28e/
qPRsBZr/tTXfI0mV3cR4pVOqE9ae0ig3AatdOJZCNOwDOnhkrNfSChhYQtEhIhcWiO97ASZeH0q4
bwgqwDicqbi29PNjrQEW8+BFTXAElUbz4r5BTawSanElFL3Y4nRcpcI6hzFezKUHNEj9Rw2QVJwI
Lfs34u38FrJZAyO0JuEhioP372eGEwLdqaFdc5lBxNYT8EolbhbIlQJEphmq9O8So1p6+5jyAfqB
dY7G8+gRUfMByPKTfFXsTaoodRvgCceDVrYQOZn+gdV/xnyO0IAgocWH0RxKS4GPKbpf8nQPGjql
lIH77jBFbuzGC1/wHFd6ZPtIcmdolQ6815tpT6FTJwGlWPB4UK2JqFRsZ/mLZiZ4h5ivOxJZwPaZ
PrCxmmdYNOKdkB1gC8oYW6p0DnL0Hod97hllLDoCklZwXp7SHDxzh7cmTSU786wZqfnuPlbvUOlv
UQ7Gw1EToANr8ax/KCRBc02V3ralvp1WbAoJePbP/TVco6rNh5F5npYIpE/tPLGuCwKa3MPpjLwN
LOBw/n8SR28XerYf4MQj/irKZfCCkXx08xmuHrvveeP8+q0bonH4GqgB1NQwBEue/gw0YQbJ/B83
wLs+9+dj4hT5nmdYFfk5jxyT3exsihARjlCjFgg2A4s1zvUWGokhNdvKyaoyfsMKgJCIFjYuqMn/
VEFqG7YwxfMGL4SEgV0Zskep37yOHk1KMyxhmOBQEa2E5zUO7SROHQac4DPRt3nq6nTygBmPosg6
hKMhmsUQOGQ0WtjSnmZUnm8aASHhLFikAV7FRolwvKY4dSn1N4KfHE6iVIzrgHFwvScFzf8+eaal
dRGLWfGQcYvKCnIAYNGGvfcGEj0qKWAe3DBmFG9TWdmMmGBQzxPyzWPNlVkb7NoHlfD4QYj5WCMx
Biu+9S2Eytxx58xxMc+zFui2VQ4m+QsnztxKDLnOMAp/7z2Rjq67SARPJmeORVT1duEyfRpueOd9
y0obfWnSgtfAv/Qrq1nKeGhmWooKRi2/3JsGqMUMXNRr8vzUPO/wDSyn9N9t0Pxfro+VVCb/xRmg
G2PVv3EeP4R8SoT90JAN+4MrM239VhSK0OAsjmKlIFEtoUGLLD3+g2BA2TP+xtVB/4l7wu/8WESC
2q+Ba0WMcZhWjwPM4eMDdkkYvweku9mk3wBMguStye5uvL+otTd5EJop41urQWgrXqUubgKnXtsF
KozA4aOtxahGZjSn3sCJbGZR4rDMTTOqss8mbdnrOV/mUi340qua2ZC5+fhEm85REAKV2uPblxo2
8JG2a9FOxT/bitKT2GjS95RIoLZsAWLbrei96Az9H/sZAu8cGI5N3qdIR5/h2VavQpp9lbqPp1Rk
2my2cF8FvT0XFgAol6lZcwXO36u3xL8OJIxkHBBg5URQljGXh0pvLv9ZHiZWGRiYNBibgMwU7OCn
fXt2VeqVhVHfBFuSgdugYt1PrtiR/tGBnsxR0vO/CRB/RYaEhS+afoIdn69pQdr3V0goNNhtHkc2
OARYBm2xNl/gh5fjbwMxlRI6fou5XAWkcZd/YwWBHxFZUWdG86lRkLw0jSDbluExe23olFiuj29x
bh0wm0yU3uvUAV/Sxsyxqo7jUZP688IwvaluzFYY5gSQeJU3O1bIEDUb203ShAgbyFM9sz5LulMz
wOsTyG05zioGS+hPnUKUeMwQLVmUhi47RaQvuqM8SqWEkyfcdtyeVhkGZzJzmOSJRTfpLaqiLxZF
ImyY2+VdRLSai4Vr0YnyQf/DDJthdjsfpvT/iMeo+fdw+zlJY3QvRW64ye0M4hBBOtKDvvQuvPgM
1yF7FfrIX0adte//U+EGWa8cmfxF7VGb+mxIBkTex4bWDr555zoN7d2HQd5wNp+ul5ciWou8DfHg
gjwQL3kNcyYA2D7AJuiX9O7UXjBtoXCM75D+Gy/l1JrbYv2vsINmw8Sj2+6VNPw47KQRIO+PiixT
jKUe2CObl4/NH38S4qHckzPoy+H5ylA5LX16BJGhEosOYJ6rWPYBd/N/k08DOcZNMF+qR1aO9UDe
gekepo2ilJfMjK0yULoeWKFwoPVrBYV8hySlboz4HowmZF47bHD2X+CFdaND1/1Ru6GdIew8HDWq
wo75ni9d/zAKI04DK0x/iCM9MrziYe/xo6htdRvNYSAW2LQilzl7TwI/OXvKdBfZodwgkuF2KR6j
gdpp0CxADw7mLVcH2pDT2KMbJU/VSLnfmEXvsb8ANTHin77YuwsJOMG5UhJbiYl/CN7cxwk3A5uj
A6YrGLhXj3lJDO8wqW9K12PlTIXUEeSV6Gtkw85GMejep0G+wgaObZUvRhR/NJzeECdbV1JUUZb0
wvlN8uLuUKmSqu0vL/xiYZuXy2TIUmKSLm+RlU0Mbzu07XhUjIw6y1ru+katrjUN/gi/kJNIr4lj
kViRfZWIz3IfzE7SObBXYpSjsoMRM4TD/kGfoF78XB7g+OsoPqtT3hVgZFzAcSncGzoeUs67q3cs
xc34bFM+NPJENh0AMLoKMP+vZm1JBu+6rrEge349lN69OSt/v+muoP/icFE6nDFKU0fxT3rdBJA7
oCIdn9ZCQPBLqDqkycQ6wlFY9md2dQVtU/U5szmP+pPWLiGUA8FHV0T7zTrHBWipQ7/kDZA5fi8B
r3cas9oXXCCyjhPNeNDOi2cR1Z/QGLdACLwasow90brR5vvPjCWkTnkpBYIbIJT1lq6ShgTgXybw
mquDvTpBmAPzhXcgR5EZP+IU+QYV40d19n2tnGukHg56Qfl0jafVy2FAfVhgPXwZ5ivGzDH2ZERE
+a81N+P1nuyTXOBslSxFhiGoWhoU2RVjQ06fct+YOb4brQENZ4C4qQQ0p4XhXzRPuz2gObFxqkGg
PzL+N16sfO1gAnL4Gtd2Qi+ef5Mg78EX7ueZZL+ImulGmj3Wwke5dg7YiXnhZgHWezspLJHG1rlP
jYd2mSUJmFA20dQGRVYDwiCe42CpNKbPgvrcO1fikPW0dmQpXxEpIVv6b2VgOcqvrMYlK45ExYkt
PcYdmQ2JytokenL1lw52nknnO2KWVtR7+aepb3SYxH5IIidUfAU+zif/U7kYYfyCgTRMRUkOsvLt
l1exXoxUJK8Pg8AdXarG26CgBMk7rl91I/oV49gurlR2osmAZ6rElW/QT3ipGyfaYMzV/MCfcZtp
JDbqok3rls1vpPkgvvL9aYBeCcKHIQm1POLkbE5btIrDj7j4wyAfBtdFfA606kJ70oIizNmScNRx
wBMQDv7t8bPjvZSxOaNsDk3P2K00ig+vEYH3CNtKIDSoFd4L6Ag4jita9Qgiqlo6d7JfwtbZpD6/
XXRcfwM1KFPkiOn117qHEfhw8N1DDtTTxvuWPkBHlHXFJ3YM3JYvxnJ5bbiMU/HmaQQOPTsfUAib
KKPJIAz4WWPAX7rXaB/TvQvOgKxRnaqp3FleiS65R6TDDjlv8aycwcLt6w7JIga+cxEbqetdqPPg
9qVwy4buWnSZ2AFMZaQtC1wiXdOmcii39oFMspyQvMPrt77nDHJeXZfwPWEkfEHWwAnDsQuZlUEg
WwJW2xQpcMHa14fv/+QMaazCInxP5kdBvJEfpFCCtt8q6sWlsHMIZj2NkCjG4AMVVJKbylO7zuCu
kyVu9fitcSiz/r06TPPauqTtkgDNkwc67avhTXv76abp6wubPoxTWbUsIUlfA6cUQhYCt1QsFjZB
QJdm5RRWtzxmXfJsKx9g73RBig8GoZwSzLDZDEfgNUNJ5vFO7QbtRZINqAYTjHzlVDOkXg1A33Lq
hYtRUnjYfFHEyTR+6GCcQ/KPpiKi5C5XMrvXE5Ix37lcjt4OMViRKHEl55J+DCDxLXHA3CUgZMQ3
BbKYSnW5xkgp0DpVtgjL/bXYyWTUL4JvHXeRWw4fJFTltt85V7tbTElnVM5PnMaDlq3vA8Ux13NY
uQ4aN32GYq/5WZzTEpJt/qQJQzAbjyMaR3uSxNlvfun1NW6L1z5khbXON+IkhY99MJjr1hwGLPvf
JIdfx43qb0t/6Gf+bR2YcqL9QOg/NCZeUoz/gMbNyMs8P5B5/lZWDaRbtzFUYalXi2hr7VDAwtbX
q+s9tSEzR/Mw2I1s5CCF1VM2ZYb7y33dLgqZzV6D/AaFd6SByX5shUOtTD3sE0ggHCbp5VVNTmLR
XLL/LHkDyXKF+oZMQhS0BeEMw0UOiLd8LbxAcoyq154x2FKyZYd/3aZPaUJv7/Ik/8ahKU3skybM
MEcThXaaEzB58iBBE13VctRwmqw3zGCkylLt+KhWXriTNM4V7yIjm8iEE7S8tCzeR/Tc/Cec2fJH
baKZo//tz2vDFaf53xIu7HQAhNSMg2D227PGkRB40yVebIVaYnDtjNZPdxPGpce3XZUgiX+gQrjx
9dLaDEeCt0ugRkDrJwK0MLmVxx8Dqe29o1rvdnbguUcKs26jpDxw6oRxWKHBdzd9rK/fhevUdXOj
qkOLWgXUskXB7CLo3kwCLBNkvWNOnSeKkqrkVS0/oSlIkoz/D7+Az9IqdtuCIY3KTRk5zmJMORO1
tnha7YyX+82ALrUx15wxVXW1olFrieABesmnMDn+w17fbY0q1SHgOUphVdHVl4XUJpnrLjuIaAap
Nx3lAvzA1RhhyGJ+yuUSifeO+AdWeLIbkeIQuATMzxNy8x39p+5nekT+h+RefVbBMeOr7JuQEERv
sAN/UrKQWcNy1pdG8Rr5w7pEXcdy58AEsLMF4YPe7Rt3Gc30vkeQGhVzZn4lGmcmdn/dTadFWtG9
0IKqyKzPn9etjkTPyY25CFASSl8hOEd9zmxuyay+G5EubIoDd7QG9kEDv1VaIqtltPVLcEZzOELy
5CmgVcAMybGKbwbGAAA6UXHXxJtoGPulTRsFobL4yHM1uunwyirFaZVWGNK0h3Xcdn1+pS7Ev2KO
saL0bWTwLOnRmWkuKvmw/8PQae6+FvAWtnPJ0YaSypWyeyb37eQrQDxfN59kZZEMxYomsDy/Vo/R
uB7XkIzdp9U4CfdSWgOwSUOJER0BfEJ+Z7Uyj1+wvB2vSPzSHjvXhcuXLK/nbZ1V2kInsfzogUHK
9OjirYSnURQW1nMNAm++eZbBpT9TpgfdfcL3NaEi3fcBP+W53i3if4pTc62T8HRPR76Gc47Ck/B9
oZeMKR8qxpvE0ymui6PPImoDvBLH5pBpHxC1tJJfvyeNEsxpElkBPSuE4AHWscovXgqI5G2McqUg
A/+Z8napb2CeO+tMlz2eZchikT/6dYIoqbVBJDuS/D+2VU1bP11WAgKWVDKKrjeDwO9ENe25/uN1
2u5RgHQctfi8kyfZ0OHczR0h4defJg2ehOuyLmksAKUVeqvlrCZfhTkxly109VZ9jUoMLcacpM13
tl6PCmaz+neRo8FAV9FOH07wX3hOJvkfjkDwbQsjqTyQRaEQFASe98XJUinOD4pdgy+UNjhpyp/w
Qr/gIKRNHrgRn8OpWcoS/QKo43sSu/f7uAvMiyk0qybasHIskTA6tRgqYEOJsE1YOCjE/StiCJHU
Mo3UBGBEtfimS7Tye0qs9zOfpQbvVtfsVU8sOqH8rRvXsUbgstrqON1jXV0V2cQYf3vUZUW9HOLY
GqDhvNqLUil4QBMut01R+VjRlZ6QlpO6QVTrWCZ4DR1fBPWJnR/8XWuwWinvUXHgl5Ni0Ku6TtxO
8exc3wNHlD7Uuohc3Wgx0eI7ehnIFAn/GcW4yArgL39Eceq8m33h/BmzFGQ7QQU0rx0Y+vi9XQ9L
vjcM7UAp+rgaD4AmVy8G75bE7NYNHKv7iVR+OhS2pBKrXSBtvNpewJFXlqdksXVksEHVDmzoGZni
GQj0xcBbdejxT3ILWizsEruaJFPtywcHxQKV2VE2bJVD+Vve2g0n7gz+h49B4A7xdUEtYcYD78yA
XMNbHTtA2RO1/sJsAKHeba8buqU6tPh1rkDJjd6nWFIlxEMsNq6J1DTg8GqYzV25fB/JkqqlLUyJ
4m5ixqK2XaI3lGYjU+qo2BD542YMmJAdTyZxBoUK9CPOeJoySP9QQSnaq+3ODYxjrM+U1MHnJUIn
tZfjHafj5fgQJYtXtrp5VzLDQvMgjA/Pxdsyt7tfZ7FPjI45QdIsSEUKFw2EV4dF+wRh2tC6LuPp
80nV2GXQ46c2+UIaMsyVuCaA2vnwKKmF2WIDLw7OiJB/ox/P7yLbx8/R3io9sMUTN4rvPQ1K5AkB
MlWxT/UmVTvy2FJ8jYJZv151yDnTcIP3tiHVXaE563iTlZYdKfAbRsAbYP2VDmPxCD5fMeDqzAv/
1jcsGjXtwU87bWs/QRBZk8ayHI0Z/de4jzzfjGwxVEjTZoIGgag5NdtUWebFKMrVWT6LEqCjN8wy
AGanE0HAivKX4canBqfUQJQnmre5xltFM6KEaqEzME1nzYoFs6O8PdcRTjj0Xco1a0bc8OvPCxAB
NGrRx3kaJwGCaylL8n3GBllxEpDk4EsS21m5BK/eBTsEqjABybd7Xtc1mJ5BEVyuJj4TYZWRZ+mR
g0yihesk0gIUO0VmTlcEY4UkMxkjjs+eXq5ROpiPR8J9MdOY/vxKr19Jq0u5xMQnMWCpWUrJFYnP
yOJRyavUXx1Zhcko20me2vQAAr/Y6aONgjTPrR4zBbrOVJJImi8ZkRKoDO0H26nilIFOpwTFGMRm
MGzfzxCuiHmCE/7sReL6h1palOrS+bPE0brsh2Vzx2W2oo6wMKVBcMIMJqsX3ZivquWRr4D2HLR7
zWtSlk2g7fXaJGBqPBTu1Vz7j7JukM5HnKSMeDN9OpYsmBpH67vo/4jcQrS9yiFpGFC7uZ9LNuN8
wnJ6Sb66J61ZpoCOSRmzIWdPwL9FSyejgr/QVZ7pAwZc7Qehbv6X76rvizmrk2UZ9Y5I0Mz27Beb
X20ONzKNA6W5ATmi5ub9hDmdv0rSk8O1LiDwpataKCjWKIpRAui/U1HR0mJee00+vYnDODUdIrkv
menkb3A+Qyds/+Ma5MF2r1Miiw12m49pkZL5PcBaCGoDA3/Y80qd6t0BFD0Pn3Pfd4dNYq/stHHV
xzTiU+Nc2Q2voRKjoZJ0onuEdpYqdtOR/c9R0hrCYL+YM4Yv96u2JnNBFneP8OvuUW//rLkocl9Q
u/IT0zmWW4BN4Dh0sDb8Z2aZyz588O/gsd+tSQqCu5lLhze12ta0k40Mi4OXr07GO3SH5GJg2CXo
cwLjD6fmsSK5wK18/7lyltIPY3j81iytv1U4n7HgIvcLqABSwxYYxgwj3dInLGcxV1qdx3G1e38i
Iaa/7yPi8SaXq4w1rM1m0iGuxQHTl4Zmd9ZR+FyjbrfQbouT3s6yZMbhWPOsp+Du04YfAQ+He06j
ffS+FZm2p1JghYYUHZV6Qrc34fJePnzE3UHUFIjF7hLcFHnrJ3BYFbg5JVnuWCl2bK/H2//16k6g
HrBc0lXa6xXK7wprNkK22Q8s+ONg//PIE9PXURJgLRKHwy9za1mzYZfigU4e6XBYYksBuRsyR+95
I5wR3UTWc9n2DtDtzUwzbR/OZ7EYHceYcjMCEHgemIDgAVkKlGgGaH0JDs6ludRVlxBR/sN9c9Xj
5zjtEEuYgvuO2oETbbiskIFsPromPtYiZZ+jTGGwKsyMlr+01qzomoy7NJHTmVPmHZdg2OlEPAm3
QfYKUT0zck5S9gySXwphgseHjiqMlnbSRZCyCaOdjxrTFa5KAeifQLZ0FYPjxeDVBmKWThhgwM8k
9F9EPsy1C0qedzpec3/YrMT7GLXo1XsOVf2/3OyUoCOh9trTVpZ3vih4o7gRI4X5k5rtL86GFO9F
KbOYpLjyIVxmUBegc3NF8rZolT2JJgexjvrD25CsMSScux5pIaao8PeDk8HiHdEVgWXdRxWd7EyC
cNY2e1pwVS4Y474pGzmLs3/oyUqfZn8dh/l8Cq4erNZ0hcWuHvrj3JXpS/A/YN+oohll3v9Cc4uX
Fp7i1TSSdQxbdmHsyRwksLxPbRhjx5/auQbQsQ9YEcTJTplPKpIR/9+vRANpvF0TB/PFC5ssB2jz
S3n2a6pKv+puOY5l+iSeAeg9IOLBS7oKWk2LcfoFfBKf/9NJanCpULIUGFertWIeU9jvi27HSDeb
wA7vIYPbJjqGv3vsAp1sP4YtFvvwoVey8BJ71wXTDhU86wmnG3rK9p/zF7XfKjOcjkuEPI2SvpSY
VKnTiWcaawNpDUuqLelAVyxobvJkAS3rlOOlhSPk5Ji34d7NBqFNyjcAWwldMqPEx7JnTYOJSXd+
pr61Nhv/4l/ujj0h+tfLE/9ufsnNew2rlSqHacOsDGp0DgUvLk6Y+qGK2DT3nDXjTcCZJ0IrMj1f
f8DkJe9WcdNKtA8Y0j2RW/Q4s9kdq15balqT2PfCd5GzL9Lxg94VRBTuaPfrXFryODoOrkdK6yEw
cq/ft2Lfr6sdAVeGfmUBVsZtGUyMXLJ37Ycn98vrM2BTuIh9hBik7hQFd3XmnMtwaqpR1rqVn4Ry
3l4YCVsi6TGWr/FvpF3Mi1yCAIa21MZj0mvj5XNG9uDuy6uEg3cTCxcffkShxN2IryredOUpAdCO
wWziNM5RlkCOfnmbHyWT+8J7prl/rAsi6OPWFOncAFKnQ55XZcRJ7lN5Q7pi16s7zBxogOolaAuU
DajQMeb+2OoH2keF2HPmNeEK2s8uq4vjjs8bP9lVO8Pod8ZccxP2kFuzDLWOSwULFTsea3AnkivD
6iOiyPRh6eft44CrNUuTptleavA4rRH58B8m1/XtNAeKZsGIi624SbUVWpBqMCKm05DCE2Fr+qSv
2yR0m/RCoab7pgJ4ecRWUESW5EbPWAmrRVIvqcEHMNli5IlICvfaSz1W5qaaS2u0U61NjSfT1FyT
5PCVgx2heMEFP3tjVuCnh6J0f+DhWziwjrSA23hJ7MUcfpYOaPjXdrH1P4ylH3uZ5p9Ax1/PxAPZ
bjvYF5nYBHdZ0rQ+MzCYB3FwAMxzlQ2YqUSbcf/2ARSKwfMmfX7sOK3mxr/BQZHSK+BsZ2VR9/EJ
f4nFtx7AvlvEPPHEfIP3SlMzrrRzDhVLfX8Ys0s/Y+karA9/Zi6s5x0G8QyFJtNjqDg8CBOphOnL
z4MpbtlP9dMEFrryg93eEVpfB+ZiZ5TbiCpp1NbxwfNgVjz1qAGRtpRS0T4iKCYPK6pI48OPpP0z
DVauIcoElmBuz6/hEMv/HmL27K1lNfqApNEMtjfMR7aEn8fgXWiHbVES73mEZPUFldD8qx4JZWXZ
4GQQEZNeFQnZyNSoYASdt0PbyZdbQ6ylD4fjmxVMjLJzA7/eh2tkdeAHVXjL9vRLjV2MpVpxBpGe
B5vStyrWimkb2FWQakBbzOxqKBG0CHCDU0SQKotEFVpnu0aRlEjYD8VZ/lJs8We+igAAejAyOx6g
Jh8zezo5bO0eY/nLys6aVpkno7Se4tzyaSLd1xaj4q9Sfel/WBLzhTxc88Zz448pKHwHpX7xzVR5
Z8sIWq5JZ4kqI2cyelhqbwHRzl6UuGDpXLtCsaTfohE5Vvyvs0PYhiVVYreTKEbUqkZ4epMFRr3d
sOOrTbrCdT3BQwnTqRDYEbheStejM5iwQgVZRRxEH+OzSL//GL6MRLYpMn0qPIEthtF+rrlhQjS+
qmS9OeNi9HPpNkk8P0XMtqI4KdQUsEqGzS11gQZwx3F/sInPdvtetMeaxzp1XGJ3VOjjpNHAwjvc
aaZ6xoYt5/s36U3vUtSpn1nOhPyQl/pTaBRQmDDtmwqGfqp3I9FBBGnvIHVHpuk/xV/h0C+yoQf6
SeZszliA75MGvxJWaZS899Tq7pIYoY0Sa/CtefjCS2EEBZcGLeqOyCQqhtDrSPyS0xkDDf+khGqF
c3TjoOLuK2uuA/vKQRxte9vBinmC1V66jBpsr8zkDzxl5OhTIwUzkRaq2ytW32yqfLQxOmyO//wR
KT8KOGxvic2Lw+EI5ZniUe1sVaL8IkqxMDjI27Es+5kqWl3u5fOgVHDBlMqedg8jRYlmZ5GRkHmz
UqlZFm8Yk1d1ebsdmIizXj8AVcvIbYnJhij6ObncMT+G+m0s1BOUeY/lSxr4ZT3p7I8J1LjFllw+
zlKKiCy9N68gXJI+rFaODdZFwiv3fwcX25xOrzKqfgDBMbcwm61sydiBdqZ9uuMc+GkvckfIsyMM
x1pVUzfmDLWRmNvdq7qKEOkPX57zkwM8g7ctlMu/2RHeoRShOrlS251antgq0gpW9RYFh2Mx8pTN
Kj8lvH8rIByHSsf6ZAsAKU8xUjW/YVAODK58TirxeKq1+9FM/xFNtgRRiQDSjXtUbwNrb0JxL5LI
KDq55qvN8ul2h9QVdZnIRNfcJLJ8JuGQTa0i2EgKACxFYinQ1hHbCGDLHSNiQc2laiD3enFayts9
3KtZx9rivu1UbkjFTaBq+d4wyNRRD9PLLhd6klxUwUuHnVorp0dBitoJEMmjJvJhuYJy9P1/mJx3
EuboPcDemSgK+e2p/lI5U/YXHskkMvhkz007io/FO845yZPyyS53yIxGHVNd6yVFRi7OpZQt7Yz7
KLL9iEgGWj87Vtn8TNOT7jGPtBvJ3lU97Lbx9HoUiGcuAC44Lj5JRrr9gmQdmc2bR/PeF0ArzTbO
Dh0NIN/8czrPm68UguekEtXzMdZGb4ckv/d6l6Q/klgHhJaa2Z0XRBfRNGjvakt0oO+Ydm7r4EBz
FAc/JoMYGKbYeMw5LC9VwYcVk/TsQUbC07IpzY14L0iC0yXJseQzHdC8xSyEF4QXXWGQ3loS7/ob
g8HVMHUD76tbyddoWMpwxy29EuLIuY0Gg/CzyaeBEWayJbaHtbvnWqrDRa9uZAUk4ksSeuTjlX0M
a7J+VgmKQOuIx+w/1DoEHtnIARC8W2ucoT4TmPP0aEXunoVAkLDrtqNY2lqETFlSGGed7cPOZzTV
YREY0vpZqADELDzWg1KiF9+KuRKZiUgHATdV+yspNREsjXrzNC2yX000PgKNUaADnnefegkMr40D
azLmb38dVvG/QU5OANI5YE3qXjrH/sRH9X7ttSSsfXTWI9m1knlULEEnv3EDZmcIzlT4Q7zJlL0I
+Gbzcs4dDR4FXMlPVW0A/wODkQ4Y1kwK7eOjc9l3tXY1s/GfUAJ+MpW93D2C8Kub34mUDTnDxkc9
uiv3mmTzcK0gYbKKTB6zW5IvRBNuviV56+pUxZYwj/awGt+rAHix/EUABBiVkOvCx5Da1rCgr+6/
tZYOHshthJ4T72RfjT/PZI3W/+HRot5UHqZchzIbdeSKA3s3gpW9Amdy4LtykLX7shAGp9wRSeJJ
/2ZzxYT72Lww+dHtgWbJBsTIHf5vuoYjUwAeVy6wzVkCGfLfGKDdXnUIL34d1LsqfCooIABL8rwk
NpXUrKwZJY2bi2J7P34P9SCu0QaMeg7SX8/Uhl8tqLz5cenx14bP9vYEziyWRIBI38i5ZkbA95o9
BswzQGa60eQD6CcNkCk8zhbgcZysl+5Z0WdEPNXJlXGjjT0i08la3J+sQrVnFCsWPeoPo8p0OhPl
ajU37PkQlZQ7LKfj0dqdkSOl+bS+IlI3QuvPny24TLwe5FGI8RHYkGy8PnvCDKRGerZa9lnQBetz
ApjkzXiSjmSVJOQolr4xLFPvcCh0QgSxOKU5et8s92hcG8qhBPyJIASZ85VAEZScGS/fexeCv9SV
Da2d43kFHOqPrXToSNWgGR1s37Kok46Wu38enVjPIANvugL3Gsn4eGuTW38HBCxk5MRihuMPp0A+
TZHGvwiQQ4iOThS0Q8JicCMhV5HtiACWuRJP1SQknwsSXHYHSSP4gpV3S3rZXOqjV7RGyvkFFUNa
SNG16UWLZCUIVHZMtZNlyGuAWParmgz+qQxDphkZWJ1+ZPpMuNno3csd0xDNJ6+vM2ppzGLvlpGx
yz+ao++/eZeW1bYjwBAwryxdBAG+TwGlWMssf4Y0oMf0n+upuvnQ583Uy/4pBIsf/J67r3m8EBBL
M+MRxsib6PR4s74zeGr5QB2NEM5lGK0ijGstInB9ONtDGEHhl0GteSl5NVuSmbh4txZikXlaYXF3
TsRpVfhcAfKmRHpyM03E37hpFK2YH+yVOW8vm+lP/VNP4Rhjdc70BQI053SdmMQJUt0a94630ocz
mJAoyEvoeAjPQN2EPwWQgBAqkWC6n1ceJcCiSPnpTmYAYCLZmYzL3+jwrCxHX12ostl3IagKibwF
OKXmj/R3tS1yBgjmgQq4vT4N/YS3cb5DSy4AYUXfEAMvk2z0EuvbyEWhReXvrIFzcuhhj9TSKf6m
GIfrUMqyjiX0sZIFoC+K9wkelq8NEkinEzNjjYTSJoC0gHh6nedf0cGF1bfBSRi4zOQ9MhG2F5mS
+JQ7NYFbe63f3m9CBRAuk5DtFrQdKdgiAse78Ckbkgmrvm5WVr3RLIqQynuSpGmLP8cyAR/7wv86
K2n9827G67mJeQo2xM+F4kGmUSV3jT92Q7RftridXrGeiAIx8Zjx02q2VTmhqFv5K+aic/wtsm+M
1pFTM8vnzqxnRKUJ3cY8MRLWX57jphgFaIiNOwqFLtLmORqG2Dejd/AwuOXq6y3Xf5zhBKLQf2cX
7qYlAb2sfbFAwLBbvr282CEpXEljjdEP1274vEnBfJqh+aO2m7pAGkc2rtx7SZctJAfeIvnruMHp
s0HD9gKAxAZefapD7fAKL67BqzFr3CUuMax8Qp42FCg5ORriaKwtSOTxXehZn6u9J4zO0ap08LUv
E9G28w5SdnYqCKANgk7/Uh+wlX2FJ7eDotrq9yxd5sdNNlw93VRdrIkMdoXu8xtjkNna7N/xPZTF
+ubEZ8psHhQCcz8YPqCeEsS9PE26syoUWyhARj6JGUVkYeBnl5NzsWjCtV8vFdrZndVuOJCnPy0y
X5dcqbxJm7QuW55X/gHf7YrIpB96HCyPUQzD3XZysipou6I2kNm3W8L9aYLXYKpc6kdqyxhAjzo7
VtkYovPZNW1otJwsYoNKC8/Wxj/ZaYBcQEW3v1MvtiPLyomR30GS5v3scspMrOpyjYqONhqOAdl8
hdvmoLAu9ZWsH6X0ExcpGy6gKvkRvpC+AbFHUPZSVWQiFqHQ3w3fLvyv++HSmHIJ9HzYdbhrQJqV
AIFSSQyS8Re5sx9T5jV4Z1f77zlwHRTGNPNDzakfL8a01sUSnWptXkAaIg7Rab1Bo2mlESWzqLKV
sVLyIvXfmxxv7uskAoOvH50rDgO+jvhKQ8OjQj3QyIgtwJPpDXI98pPUTB9MQ6QB/86np8r1P2TE
MJkvJ/8pegogaXddmEhOxwFRREgpfLFmKGsqyww9yonjNwv60j2Sl66SMVOGePAP2EWyFbG7ezxb
DCgf9ZlXnF7Ypcm9CJT6Kq4l/OVmR74FTk0YX7+pMxIpU3KGFqjpZZNil0ZKjQSXol2t4Zg/vI3f
I+sG6iUprfAICfI2gLrMh1fLZ4er+2E/JuSyBQ0hz+mh56CKj4E8Pn+fmzLccmINRaH9HDMtLxIJ
+5EYOdKtlfBE/8iMMbzfczVjA5OUjisLlymllDF1Jc+x0bg//5pcqGex9xbJe1zungU6m5aeGUMA
D/3Cnn/OHm675r2RCBy8PWsMjTtLRVU9ln7JGxb9u6cbBkLSXx2TpIzxnbO6dSFwTvcFTW9gV0gP
tPmq0ju5It7pHOl+HKazOLmDkUSKdhIl0UAiYvtxNPMEWeXmGC1NmkH1dKKGnGPHjQOwI1kzm+Qo
RnLLwLzVO1/qECsXsMdX4xyDLAArD8jeiQ5cz8P/V8z6dHLTyutaGDXyLhiD8GDP0Bhj6huHZA1W
p8GfN0gj1U82/BY1ikYVzCtFsqSsbyKd/eUvzJa6b9QwuFl7LTAmQ4t5jvaQcKVweKTZdsKI0SJX
IP90h63FIrjzCiE5vIQbOCcaFiCDGhSOYU5WDuQK6+b5q/t3Jwe0bAQP6hW/+VQIesXFaxnxmH+R
v25+x3+XtImRLyOsyRSLys4DraUhBpePGKl/NDVSF0+AesFzWV8ZSvl1nXoeo6RNHMwJXcet7aPb
0gF+DX32h7Pu4iZPf2dOv9xR/uGcZVEM33gMSq9MsoqRNveqmRP/Du+58rJ619dgX2FbXQKFZ6iK
TAseoq6Sve02BA6QGHt4vK+7FMT7rmWCxjI6EU6MCkxgOjcHypbNXRFVOfad0GsG47fGzRvZiysh
MOmFgnR1NIvGbeTN9GTe8opsLOhrcd3igotbPUQMu3Ffd59cwxQUkXmH7IgktFT5GOnMzau7CFzk
rq1hupSGawVExdliHAsgztwXMW+V33JyJmmjnXTGMjfJR4OLdA0VF1szM9CLG10uD+x5yHEPwCQ0
c/f/4kzr8Ph/OVBSWwRZQevog5m3B44UilEX5d1A/h0GJlPIRG4hRcq96YhjiYMLXDkc721O3Hhx
EogFdlMyntR1uQMxjABxeMbLVzuRL/IKHBNhVnZHVQKjba43C9nNQTvf4xaU8EozSpv2mfWBqZ8/
tiJ2XqxTRYm3pAtd/rrzCpDccproUMk3zTQ9OAcR7991GqjG4/L+v1YvUClyVZ5TyfX7TQ7LAIE3
La4kYJkhxXB7jjqlZmrigyaC7Mc7XI6IENt/u50zxtv8R+hqZbWuOrGzeltqizkTdm1fp4RdeON1
R7XtebrHGf7cw5aAYRKmaXtECnKpHx6UojuPycaR3FLfCvJjIO3y10VKIMqDF3TMbNPnmq5Zfq7K
rgrFr3dtiBsPZnykeA7zOtoTKhAtApvvZwYFIu7/OtVRvxXbUNaIFQINcbtfclGlwLNZR4niaXZ6
l9/aW133tw2QhVAsUtiUCsTNzxedOvr1yrfGm2LroAALVDqRf8r918qpJFeH4mf+lnaUIy2vtcCj
Q0jdC/b+SvsRJDp6lqhJZ2ECkvXnkz/dy7Ii34BV3pOuBv0dp4ITggA2LQYiPOhha8Qd0j97S7RF
snYIYkiTUSPaJdLmagrwaEVajXw3zzUtMm91NAtb1qhFgOe+vF+mzcTwu41RERS44igHpPEWkRcG
VczAOgcY4NSal4HgO4dhNIT4wehk/5jXw9D7GsfeZSIQ4u58tHk+dXZybTdyVeYaywDkAmSQekh1
YA+0dfcO7Q4MNVI5k/r5kBv/92y3Hfiyfa281LyQL4D2sZzvOAToCXyNZiDnsK3PaZJ5TgeNKNJS
87PIrD0aplvGu9Fpy0IvozH+JtxJSuSn2q97BMQqSzO3Cx4yQxgVx/ggA+LnwhUMkj7pWNlVzuFW
qapuczHHb0mK0EwCCwOlnXoOX7cDxM5622HZ5ZaWdCPXoqx4MAriofDUuDo+sOu4de9eEYJtOWQg
Eh9tIaIIv7vsEdUH3ZpeqET4Vj65/9qJ0Jy8qJjTsObJIpf4UfrqyrATeIcgCPCudxyd0OjZ+Jzr
pV0ZSEzaj2ngpC+GSSoKZKird6EFya7lA25QS6jrVLjK3BID8useu3GQjqI6Z2StRt0j/VBCPNmw
hvJG95pRk7d8XjROQ8oKwZwiixH9A6Dz8R7NEui+jw9xFcN3+xXL5N56yTgooeQUMUvFU52T9Qy2
U+DTVr+6rh+VZAvzZzCS0yleaI3aXxJRE+Oqj2wE4Wo1PMh8aY7XHDIF3rd4maAJBb66Ci5XxMMJ
Sl4y37F8uICH7Wh8lrCCasE8uN9tqkrcMZJghqVjtfoFp/SMmtxOSoZ4HtJPE+lfTdtiBkWVzFks
dC1Xua512Ck2pJ6HY1xaJhb+PH0aK1wiOgQEJPUTFdjWdu+3/tQvR21EMhTWQj/ocQBJD0AgyPdD
3HXK50B9lNRVM4mq0BfEpgtd72esKvLtyUacuO+Dpo5VHMatWRCy3L3nG2ssUqTJu0ZQHLXjrDi1
rQGShIGQKAn7U+FtdBcfo7xhLyBDosfsOSpcr/CVgIbWKPncbv2RGmBVCdZ2gFsX4RtqkykHs/Hd
Gw+d7368L9ub8sB8ofE+w+Aod34kJBRzsyAND4C3r1PNLcmu1E+rDxYoYBmdJAoP3ininbvF4nzS
N+mSTa/pavUvgIEwXhZ89giRxJVIDRD49O5Kyr+OdjAvA5hgL91V8srgkbIv1FJthn0i43Rwu2b8
jngzER5Us9fL4MOv0Q5zUOWuCKMPfXbWpzqHqEVeljxsMWOn3Oorf/MyncSrgMBYSRqpklL0T5Jt
lU0fu6yyKAzaySIneCwWq2waN7x7Dg51R8Kke33k+xpNSD79pFc98qD8qYW9UTFwSo4jY8e47oLv
q2mjI78kNpNSUZh3oBLbeNekddSYbtA9G5w9j4b1sxn6HrnIqQVDZhYjINQSYf+BLhRhrPzbssNn
joMKo1Qc6NXHn5f10nLfSKW/gze1Xaatdt0DwPWZu+ysv30ATu4GtPkNcnC9xJbF1UOgV2h1b8Y0
U0Ir5yFM4dTrly5Pe8GnlRWMOIJ89coHfnhfItDLHsjeE2FI/Woe8u+aZ0wRbT1Qm/LAXeALwOLH
MunFdfNw2GY4hlQb4iMBe4DApsrMLI163RCBcLFhO/Y6U0qsztSAIRbAfD80VguKbV3iavrHXqY7
oG6WMXVKLFd4wJ8yQrhvTFqDPx8fkdBe1aYW6DCJ/QGrj7PlB/l250Gr1fZN+CRsJoUSl+FxKxJ3
mRwn7ELAIrRyxi8I6WSfdls9fOCouNVtjjJDJiyAsDad/5z8hTze1Y/MrxbQE8rsbZOtNNKq6/3c
o1mUMQtbo2pDPJnKcAYpTbqlzsGxffziq6MF7q1RuUTGMDRk5f+KN6hHBAg7NjzFR68gZHIm2Z8c
YzuBQrrJhZM0yRn8IBUNpkIgcJ5wJ5WIelElRYZ4kMxN7mxxFk3a96RcBTjWCN4RUtdMzz2HcvkP
dtLdEERcJjR4wnXXFaCK0LFSqG8E3ddeB14J5xVPJyQniSfYs1070B2LCQB8P0IjZo6ULiCgt82B
eydPI45rWO1ZJRbVJ/HbLCa4R4g5Q2/N2v3H6fFTpSYMs0k6r0xAix2LG1OeOoeGAbeJSA42aE89
nje6ZquL6NtxEBqNSUDYRjTZqjLUtw+OowGl0+akNaZjI6OW8Qvg+fo5RWCa+jzBQvnp7/IyNMZD
mX+8HKfURtr5noaRzOiwSeuwfRTeMsEgmKzjbjFMearMsM5MHZQ9Mi2PWIvDHXM+EMi6aXEvT5Bc
/G6LJi8R0P5Gh0akqD8ACKMxXUyrCf7yqM12AbW5Cz9UN2X3yeUuzwdhxvwMnDjYUwJVcwXy4/lJ
C3+Ay5UMO55fN+85SPwKjoJ6joAi73hoEdhiSoD/7Sc7Q1GgD5hSIvxQjEGQhUKvkZh56IbuNLxz
q0iY4JtmdacLtIZrsfR6myjr7HdoOrCaVtvPrWxU+R/Zo8CduzvaJkiiL2+tLFk2kb/mydj1NUGU
dJep11YIlWWMQTUOM4z+olkh6sqRl2Cm3V76piHY8lB6l3tJ0gu4puCBXJzVVRUOc06DvJr1BGD1
kLNNJPBudwOCR3KcT6u5ovq9LH13/ggmp3Q2FfFGTTpePa0aZ/Rl62PGUHuq1bsQNDJPEsUcMiGd
4hFNkogoLRKgPKjsxHsZVOuX7vetZe8d4xF+HjCp7+SeiXYl+l54YFdEPEkseFEHyyQ+D6jvokee
fvzQSEGaghI6xSVojkPu6/d4siMMbkLudk6GVRTDMBJvraeehLfY9k460kM03bWIGyPeGHw3C9U4
0rN4D0E7fBoXwRI+cgWI8FBBzsY5gF5ukAj//+UKVYpv+S2KFYDQFjZIN+3HW39BH79cCeTGzxoe
CN0lUD3bu6x7BT+btlWanrLGR+NrtczuMrTo5HdJ71lKA7SSxCzMUftIK050oJvGXqmA7F4PzXnI
QNS5DbxKxFM5WKnFYBJsc3le0UKBHNGmUUsyZgd2NbXfXg0kbFJXyVhFckYSkz8EZdcmY7CvyF8t
0avqC4aTBFN3DLMqVfQYAR4OTYvk7QDiOWtwHSQk7huNAT3xRwGVIWz1qVA3vEen3MimOJqFPfDW
Tai9ID6LthWNtyiOiJCYJA7Q8swo/ly0ZQkAmdLfgflCGog6J5bs46X4vdkU9qj3yEnjyY203IsJ
M4PeiFb0/4KBi9bKn1loZp+QNrvOK4N5z8AzUitJElaGEZiVE7NwYZhC0zrSI1WfSfKvPRk85FW9
fSCTs/xPV/QdG34kBEUoR6jytdsRDhIunoqJubH9dEfn5tENm6q7VCxTdv7qfa/EoNBkwlvyczp4
cHYm9h0b0w+kbD0Fw5RfWjNup234OWmvUwHnRWzViugz8Wsb12RoGDKY00C/czt68fe5/rLQ1dhx
ek2NmPxRnsRFyroT2BwZ7lqgzKU1VAan3yoscD096MrTFz2R48GdTEbrm/c+07aTnzn4h6DL6vcG
g6eZCO+IE6zN6X9BcEUDThL1tgBvAtJPuDPco4Aq5taYBTepTLm9UXlDiFyiiyJ5pRdtoVHWJm/Q
Db1J7VPfez34b+72yKSfnkbhC62Tw2SjTpDJczKwYNEdYefKbLdEMqawK8Sejzy3EzYjGIJgfIcP
KCkc8OFm4MIQL7U3OX/wRWNjvHbAxoyMwRkQPF8s9Pimvc2VUUsNcKe7qWoIvxzoWaOwN2ojWGzq
QaSEM91XGHFg4bAS6SfcCIz9VRB1O1CvBJzbrJTjxeVA6CU+N5te8y7IcHRVPCnGWURRH9uCkJir
E3L3OZ8p4lzu/L2X4RdvYeEB8Ns3XXXksY+ktgw0HOO03Bhrz/Ez4Bx1UgD0FVcW4AtIqOuYSqwZ
Lz9iyQ3nWLc628+jBUjRo1wvayYgeIKKRHwHZ3Jfv4E3DRjvEQJsKPjKCFL5dm3Cz7JqbfnehOA3
XWeHv7PY400UG53OIMcgp7vtbL6Gak9QO8nSNw+ttae6frJ2WsxkJxBX2z70zkOe/rMrD8PzBJ1x
jr0IB+nRKquWoHT47JI/z+lgyGZqOjdBFcnLRiPH6UNyOo6WRugId6q5yse0ozRTcVF7jvDkoSL2
qKZ1SgOznNU41i5x7PK3FzXni2cNbY96Hq6vf7khwvL+k7Lxro5F9w7y8whKn3Zy94JmHU6MXiSp
cOQ80VvQs7JpMtP/L8TfUMBXmjjGgXM8Qkjvsths1my8lsv6/8p66EtI8F0hM4eiCQ1tHaNIZ6Ud
fQiKjs/KSw5+ZD8guGx/ZSmudaPdJcPouEUeqXNLu/SI8Ch7gNRrb9Ndi3NvZMgixPSCD9kKBUu5
q4ZKS1+g0J6bHvDerfD+6HPwJlYXQpzn1vsG++cYtYDtdYmoK+zmq+xcpUExU0PCL8ClGjx5ZEI3
bKwjLWiYBNphCSebLKOfStM9dV14C/vTI1i60EhX5q+dnW/5pwG7NuH32nglv4+D6Zsp/RG4CD9r
vpCyNNxmpfo6/Hh1HFvFu3inaDVRqxko5xTXi9KW2zHShTzL0k9q0xSVplsFkzFIwjL+0Iz4WqaI
3NodexscBGg949wxdIYJ1kXatC2Cavnu92XcsBFAvjk09CHu5OcKYZWaFkVObmxeXVGY8l2tYi/A
mWAWvJ44pAO4UVHk8Ey6/8AzbP8CNhcWVMUEbREIHNY95m4uxRm5cBRYRsK7cRenbNPQeTQUORI2
y4mWzx1RMXc2HfH5ocxZ2XqW0ys5h6vsc25OdaEJ/F5Fgh0XZ2WTVuqsw7O3j1MNg+4ALhHvxIFa
8niIDaE1+PlG//G/rTN46Vu/0/OWG0PULymN4OPseeHxnvVGgIVjE+TDBfasNkP6YmA22qXw6SB6
UX87/RXpaPvZP5C/koKZiIdkVhyZVqcQ+xJCdkYgvqbcwMiVM9IcAdcqyG8BGi8L+nkpIPAIROt4
2W8DPKQM+11CU4sHNXdllcJKeK6LvzPoRH9jrA0WFEay38z1czVi+ry4mdf3YzipUkEWLcV0OdxW
leaBLWELtXCw40HZWSMGMmWXVQ/fnwlwvCijVbpWU/HTvbHu5J4CZg11cuvTkxD/DIVwmOkIHJHC
1wBwV8G1Pi03GYGRLlghhC6cLIAkJrx/NzFhWHgifXqWDQW4JNV4ofqXVZlEnnaO5PEZE/s+VgS3
pfK3JPaJ0Rie+BadTZa+VU7ECOlFD7l27QL+sbeUpnDbc2KEGlH1fjuHJKoBMLd9OMiK/gBfRwDe
vLocHt72wZkO0IWIW5l656oH71v+VWSvhBe6s3Ej1LUMarXAdnGq04zjyoqDxbzSMwwoKnbgpSQr
NVbMbphLC/X5UcfyLH72qD7+m6y2w0wAcBqwRBG9TZe/IhqVgmOrRHxs3d4XgtfCdrA0ysAiZbV5
VJq2Ar71qmNgsnMjLWjdBGVCGQyNR6bMZjXZXOfYN+/GPcOUzGIWm2UR8mSOyt6oDQx1A7ZNX17M
6s6BZ+1+VP82KfisFdaTGYsHaBj+Rq8QbjVtf51L87pig2Xn7QGrX563CN6vhQag087QzdltfR5i
fSg+s8Vy4nmi1mvq51zO7aO4ohh0o7FB9CWu82pmbbuvBtp0AkFf0Nd63oDgom9lE+YOiO8zcyDf
TAccsP7Stk84ujamCLPVZ2EFyHvWbGvvEWP6ZafNf/+IkcmwpQbLn0zucYRR607mOR/zEYeJEBxO
7CkJfFtGdugsXULarDlOUEI+z9ZTKaqvanPzqlqmn9IaS7OumGiZTPpmseQVXxcxs8AQf2PTBIxc
Szfr1F+lTFXHGLD8ek96ME99DMwLThlHGqeeo0Y/HYpO/AiW1QiGHwXJjj9AEgGr35F+C2diR711
VsO1Han1Uw+QJYUdwMxAhryIFvJWAe/tZdw4dQC/785cQN/dPGGrXoBz3EOvPtAnbQqL2usN/RU+
2iRlFOf2j+35JPo6rogIo7mPPCmo1cS/rlAwz+Cut5w9mrRhdxUwEdI8e8jzaaRTC9vOpar1ClU3
a2vn+qx1wcOiac+eiHjEIXWz4DlQGKW6+y22Sn6cAJOq7zrRZrMhucuN16MwCwSqJfFRHBHtuifn
1XoVsurmpLayO+1JQSp8jQn6o8Rmf34saOlHO/TiXhsm9YLFdQH0eTcPZ8SmC4T6Mufk3zNvdJGV
hdzBao8MlXzlhvvDpEdXQw2gv4XWRgASyxrULJWXkSfnm+E100jCzQKCNdT09ECfZp6bYUMp9Aze
A36CfPGbMJfOig/xnPQgmN6eaRms9LDRcOBTuEFvuw9efiwV4ZoXHejHUgZZvYwrvUknZAHnuSim
hP1qFRPQGw57CZUBNWT1odY84pyHDf5wOTm4PuBz/ZNdJNOV/daswqq/4YtvdXgtRpo8dNZRK0rf
+0RODRtrR3WCwcPeGkstieCgAEV7HL7Lfq6tuaEbRLS4hcu/OLEgxMAk2fHgAmSDlW2amKPNVYIY
CW6KuABfNayrnhuWTU/8qLqDhZJxxzqz6oKgxZQs3ayeSJDqBFidhohXcNZyzTUXbCo6uQH3dAQh
53ED+KnR6p2yzpc7419atgYCl+hADKdvSqdJzNS6rCUNJ2rGbjoQAag/SxOJhFVKo2u5AP44dyi1
Roc49hGfg9JjjmsaF0HphM6TKwaauCDhsa94aTpjWXw2PHf4zKPbASWA3PIs6inf/AFCWHZe6CXF
6tMNEyUexBbcfu1hLnCQy6dBHLFWb3qf4rQvFYBCjMK9sfGs2Gip3snW429EV5yvKIgBwaLVO5xt
AW4B/9GieK1BD97K746sw+2zIHcHUe7IsubcehtJrcpk3d4WFH9iCyEwq9L8of2r1ArwvvD1vd3J
WFT/Quyt9pmKhAmCwwdA8gPbTRjxrxvieMgVKHEMNyjDLsGQKhZS4ewOr+4/LAykDfDN4YfnhaS4
i9oes7Bcsp9bKlGd36XzKSpoKtufMRyJZf7eHwCKkn6AtWlRHpFrnrwnKbJ3iD6JrSNROe2Hl/wZ
DaAzWZ+2sGdV+EuAiYhtCyisRd3Ue98FAb6w+2UOk0rBjpPIpHEEznv9pDHQG0kz6nxZmYQTf0wd
zfS696WI7d6oxbELWt2PxPH9ol3eQN5j1ymPeTC7a/Jr9ek6bcgLWQ20+DdR6eF7Jkeu1CQyBSzX
IW52IWhsgYorGCjswNvnZhwW8bWWLXkKA4wOmJ5gAQhAiyeMtiraLFtOU28xWRd2Wx2NHltrd6K1
nS++0pSly8aXLYDXDfsPP4JsmmuEilhu5w1YWbccVCBtgb9uv0Y+0q8qBtQhbLl4MPB+8VcZr9/p
mnm2ozcUJwEIWol/s1sc3UrBpp/tFwVOwmdWVL13Y6RD0liHxPBsVvZwAQf5s/Y5NrxQnQSQLnAF
s9g2Gsnopusf26gT7QCqrvr3EPNXwwmdkZnUAdZyDsti8h250ipmhE+ejUz+0GHA3dhPgjDWn0XJ
+M8JPoDlAo56zJ2VnpMvK/NMJXvgApzxc78coxhiAC1H9LmjubswwDp5COWPAu7lDpbUU/GyeAhp
ZcGUe3wTrOl/xUrwFYRAe1W1YW0ILO25C/d6A8y7hTeAO/LUbY3C3LataJIw1quYSPuAFDKvPv9a
fSBumlNMYNIY+ksq++mSMJltVWwIOYEEmeSi88wgeAI+WQOAljTX88LSqcIee+ZMrE8gDHnEvBgi
O5FjHP5x6EOL9Kz8ZT6Uvl2Lchat+9G8L2O+emCDplHL8TDkL+qJU96T8LHY5q3cHeM7gAreO9nN
mLS9TKRJrcWO+78S0rr3JNv00REAu6pLyGkFAUzKCupRgrH5WMx97UYmZ/zGjeBLF0Ee5lSx7Zvx
FwQ31DrQfwq1QRKfyqqGiv1k53wTPnPcu840piR9sdr1zkipTDuWWeAJmlR55OJLI2a73/xxEW8V
L762GJFRs9arTJkM204MCrRsMdise7wh+efn4q6FBMVQZcE1nWOzQu7XXp0sp1+03XcMYJBM1w56
DHQSN6xf3AwLCmn8IEAK08a6klF2k/fIsc6kvtPtslc+X8rSblvoXTrLbQdCo5LWzug4U3Cp+bYk
JgGgi7WGBWMdT/KTF3voa5ReSRzwf1qcjVZAmcpwycji0vDAUQsYK4S/CVTQXNqSSYsAgsq6RCB1
IPqmopIDZ9Bsy9LJu/V+Kf66aOof38SYF+m8vuVXjyuR5LiBvHgxWfmWeEJVgu+Q8OUk0dmSAR6t
A0YgXSrOhTpI9N01f6BLC7NHWohXhagc5h8SYJsuJhuPDo/T+R7i+abKjK84JskH07/Dem4hfl8k
uDv8exH+kbXLYJfnvoWykN0a9eOnwutnaU/g8iKJF1Ho1PlH+t+tVN6KtfIQXRmdMFSD6mHwviNJ
HXCawzMG25BS1vsPEbTIBeeNgLtWX59s8xfLq/dZkQwwST1YPJ780EUhDcz8+kL6MNZ2JcdaYDxf
x2rGAXxFD95K3xE3ZeBXvTSq1TGY1+/kz6W8Fs+ZYWgf4xYffvueB4EthOCLhxpxnxAAWNJZSfiD
UcQJV6llBGzfOtuxCw7rAe0eB3k9iAWy/8QNLVhcJcysv9WxQW9RCKJvZOvPDMBDUXI1URgcFROo
jVMHyS2dx4Id+HtkyqriHG2M1Fp2HrpXKENhJc6+1cSG4tzhC2mJn66ilWchrCLU2hE2Rr/Zuldu
EziADHmijeuIjnfEWdmaZ+2M6hsFBsgeNfdRzKZYw54uAJ+e7BrBvNHpwx0IQ4TDD5rPvodB8OP+
cGUzBEYhqVBxcW+/v+4wx//wjNHp21DLo4oXFUbE2FkNM5F+KdYpYeUvJXSZjOiisbKC6CSE/1AP
0GQSlmYVy7dLrW+2DbekxZHxUCuhT9QGlKbRn6ljor+JO6RuXldvrWIqpJbZA4UR6jCmozqFh7ji
918tUdGlZp8a7xdh+x9nLFtVMBZd+guy438jf2xzagvdlk21h5UJmwMos3pFzmY0UzWD3cO2zE3B
o4UsFYEl/KPIm63zJ2IIg/npsJ1O4UiAJMid2KoUWGq13Fvg/qC12Xxm4VG0R2e3n2Mu4lRrr/DD
MgfXY5Y+6Njm/UpIc9jlriBv5a1MPyXozd7iKkhbXv+4NcAdZ619g2nj/gVdVqo6zdy/wsDooSI6
9jbblsouHggdvR4cfo2PlbwNjGIt5BmESLl9ChBGaLYj73MLt5BZ5xsAyx/xUTAUPa+WlziLnQtD
G30DV875P7JCK2ql2obEoop9MLt0kYxard/WiOMDrJiQxMMZ8UVxp0QOw1ZV8glIPs4VvoWOodzX
Ehbw6QFdZ0orlanMcUgZzfJ3XgFtYOUy+l0VZ3EOCA71qMdAJ3IzJcVOk+xb1bwHGqjJN5jjlfb2
7sYvAwhaDWf4jKIW7gq+A5JjojgwhxPWxcBUj4D26/78zjt9OgfIOS63cFgUjr7bumQ4mKSkMR4F
Pw2r/iu+Ae2D+VKLUa+I51e/CL+o93x9Hyxxv+s5Zov2rnTFKys9m702Gedqfs4IyZ+DKQTwD+g6
U2LtQ33CoxraKM7kRSAZBomAVCBgCpU/TVvM7gm8RerITmElfeNwT6PDDaq3ttdjcdyLX/EyWY2L
tCt8kpdK+c50KfiCyY994KBnRkfhmiKJL+CAVPPwgmmnpQgCnhlTD5ayG+fzMbP5eZpBJKk4NonF
3rup8nXWivl4Xwzi71QaTcKUrNBUnKG8KIjhyyZM8/Yd09cztZNob4PQXfHWpUQDhXThFYlQLMZT
uSWPgFSDWiSFkKKyrA9q4W68WN/v/oxGHvNNrxmycYBi+yjqXm0lot6UYEdpFORSgAulLcCMMNts
jSs1Uh7bsA+VsIONTqZbgBAFCyK3d6jGC07pjODjUJ8oS2u0CI9W+nXml48kfJFm2APC7KtWR1Qv
VafCHFaAxeMaG8ubzckgmA9RK396lPtOoYfKOFTtqoaK2WuyZfunpe1IiX2F2fS/QSalneeYYybe
AK5SG126hwlXh0K5USWR0YemMYi99jQlD42UQ83unC3vDZ5Ah34x3p79hoxCjWbq+ZJJOlWoZbEe
ssGB3HP71en1rf6b5liXThBVvQjrKVh8WvKDCwzKADMH81+mJQuQUOx2hy3l4vj4Ps4/L5OxMJzR
5H3X9G4O3Z/kr2jj5etcg0KGD0WqOTptIiltZewWrt30VwKpZYvGbp5cgRixVGI0hE4AI6JIsO4a
bJF/ZsNo7AQhUC7GMzgvYqAFn3QDNx29t9DizPaHf1DnI+p/MPqjVXE6zBraiH6QxljBtPRZ6WU+
y+zoBq/DLJeZQ8QDlPlr0YsaS2YN3/0TNWy04trX9qDXBtp635PY+oo4YmtY13VYqUr1QkbkodLX
MHN5zMd9utMmY2zXznGuEhXiXKWlCAygdlvq77MtEVUpQrF014pZgtWNG/TWFEhoNdMg1WoA1P9j
43PwDirGWQe1oDzH3KnWHqV+TEA40Zla71YNdybjL64BZIG0NkUGqAPDkRl0voibZYco7Mre6Ek9
QVdzcN/FGDAIv1Es5sIfuJtQ15TgdA9BpfC/ouKvRYcMAb482iE3ZGXVElg5NdUujhT0udCUoMte
0rVQQgatuwjRQNR7R3YcSa+V9BN1Ea6RD/MSLgdwCfjSLI4RkW4iGkFjGj8SP70KEJChR43TfYys
m0ojWQRMzs4enx1SdVLknxjm3A3OT08ajHVDlxGaJK2KWFe6fZ6F8dhtoOGm/NlMvlle9Bspa/1e
so2vnniQIOfD+wKqvdiJuV8VXf9q2wDRrBuwIEQnFk2/RHKrC1PHjBTRgsx0mZhceH/QHYazKsa3
FYvsOQQY74bPgQAoqzlNQU6c2GpDDL8vvXGLbsY63kYpu+3VorOA43KfcIan5zg5cJDAZN1oSaUk
fDGIiHBhkJiVSlH7ygxOfiSuH5OYVBlKg7aoEvwP6cX30ZE97CG4eHmSaNU2KtsuttWkJTxkZqKy
6BCczj2RPOY3uBAiX73wnxd1fy/w0qdE/gbacaAU3Qzs6CPSZeH0S/7nI4qDlj9NP0VJXcuTGtpF
m+KqJoHbZJPvaaO3DgOvJrjmOex/ZtQN4eYLifoteEhRhdRslY5btnBGMeKBJWTdrmDMVSTCWLx+
3tKqSbFyM5ryiJAnyf2UHTVIk8fjgBddbfNhPHEpSK9O2kam2468KKW8dU7WOaW4IaoMFdADvj/j
C7xQoavIkqf3yFxfExdm7QwzJOLvUJdEN9zHMveKsL3V9l+wgdzyB1zQ45YR9yxhi8JLC0QXGv73
le3CdV1fDg0crE7xPnqMfVTXlgwrhLmsOq8YcibEkOvqE2u+78uX/viGHcMAbjQ2oaATptr5mapN
ReCRPpl1jUayyfqBHg8g4dBC2JNVuryzcTXDaNKGWnbCv/0X/lrVE3wXRVSR0kRGbzp739nVtOQy
x9FUBgwwXzF6rsTmBSqGtGCq0K88T/srj1NQKb97Y+JmTCL4mgOLOMAi86n8SSPIGMT+qTdfdnek
kPtLQe4OAlaN6d3ojdA0F/SBrVU8AhysDoF3JIuX8GDSES/Ap72l7nv11Mg2Ent7tCPxRgep0/be
FEGyfruvjUyx7rLUe0UyZOQgx1FV3G8C/GJEV7lpv89xHrT8/Kl26Y3CXx2Nh+Q3gHcNZ0Do12nY
DaNXNUblMQpPkh7FDrvoBZ3byyo9YrNq49LyFwpPBy0Xu8IC77kgpDATK0hzkKa56seYU+DdNwvx
RBBXLUeAp8Lt1WJNnwi58DdtdRFKsGP/8TWca7xNEeTYx/IYFjm7X2qinfBxuVBKEsWuRc90VTRp
tPaAwsJ4cKxqNLhZCuecjts1MxRvLmDTX/k+HTT3BF9c+zv6g9ftr2RyeoDRTtk/cwNFkHCVPzYg
ejPSpXebF2Rz3/xwgL2Ij3+HAmrCre1UlpbGiC1YbZum5hCmt6JHLzasmejK5flqdJyFkmHoFkpQ
XyZEQsFSq6PUwsqoTvwlPOAvHQG85alMyWTVewHzTzQ6g/rL51W/IGG39gvvBnKv7OWgITJBnrnt
0RmvCkKS9oluB0Nlal6rhilEcvCdDkfk3xIpQh8NJozc8d1LR8EYJsfL6Ii4h+u1pMkFsUZNyzcL
NEqQ3c36hslJBOdRZcWh7F5iQioilzZCkGiJpPCg6v9sF1+2dIrreJQxjROZDkl2DjMk9xFKpjdh
JfPH1dBuaY8A3wB6YmIyOKbYxBmwa85K6m7/QaBn5NA/pG1SFZlz17mv1Ueka1zhXAcu+fPv5Cb+
jyKuU3C/LGI5LF1nD5HiW7QtDPcEtkXyZHR96pV095E3grNZ/x9EjtDLB3mVU1QwgdnDCAQOZrrL
mRNBBs14RKTWmBOtgKk1OkCZLEON6dcyIW3+3G59xOHKmHRSVufzLG/Kw+avei5oDHuNtjQyOLok
g/LFhmjV47S17Mt1mRucz3U4DgOAdDTthPHtBy0ZjWl38wu8Z/TcOFNws0ZvH9lGTYTKI3aLCymm
Ah0AIgNBWIxM48vZiAF5wJSNsgr8sOPqXS97vXsQ6Cl3CQTlRkvld4qKSKOpHj3J8O0Att2tFp9v
Yvhl215c8LZPW7rnNXp+jmgt2O6Kyw14DuRImQkG69oDLmymv+G84nanHkW/yiM79K4jRG2Ql8Iy
eAJtNjK+rAWVoBX4BvmNaDTzIQUsnNWmtc4/Vl6wQp6haor68OSVnRGGyd0rL3y1nSr5DjPRGnkN
ZqrO5YkGDtYFLoE7A0TnLGIQt2Q/ltObCpGrCys5my5w1JJE0LNiajV09WBz/JxGNbIYcUChUk3Z
1QrP8IrCBHtNLKSoJd5Vy2Bv92sBX2f/tFCPQCH/BMpb7jTDWydjDe0mGPkIka/gC2YgYWEJn7AA
G6517OKsXRTS+m8RyYa5hK8Dq99UdTCThG3PeLOxKHxCFsjD6A9E9PRaGtmkwc1Vn8Cb6e63NXRt
fW/OsWxrf41Z+PV7rkeBlMicu05x+5DTEvlmg29ZRQz3mVmoXmQzT/HX9blUxf74luPMOKjt5lCV
I2vN9TFt5Hm+bOn1z/eqjlZbUYOiQuDe3SjTmaywWujjWPysr9uJoJxEFnkwIACCKD6TGY1bngTe
v1nymDQd2ZEy6glJusmWGCvef5AjxVafPweaYMfnTa+JIF719/+DhkHKuDXTppAUdzejlY8LvfjR
vzAunk6NlUHnTgaihHRLRaxIMCzlsHHBNhA4x9YkGQ1iaY0P7VBIsFB9cBE/2ippWv6P0AtxX7az
aVfy3tykJ7aHjfq7w5qLwPVo2mdku652fh41oIR/MbWd7De4dkjW8SUF5ui6q5hMa5XsRTsDtgQN
PcXG/TB1r4QXUD7gCQVW/tugz0VnG69ok/l/70wNPFUwRocvBMODUSlYu83RVNgVYJk4s3VCwSjU
oVI9W38YzM/icpLg4498rfrNXV8eyNVdLM/ZvdmsOPXwX9rF2oe+ySz6fr4LgIqBxaejIJvtatwo
2HZXrMxs0xj6d+DZDFpYowp2TRRF6FIh5R8ui/+fDhY1YfWQydkoR3Pw0MXcKtrPCrGnSvGiWwkK
+vVXBR36BV2oSbdwAk3/ssT7i8NrTLGqsP4kmtQzR5jUlNQTVXpU47ASCFt1ZrmQ0TjhQKwWZOBZ
TMezi2CpHEjZ8R9riXzcorJjWdPBNI2hHKkKdcFszvcz9PD+s/dMGSzuqZqUeuiWPriZtSL7+hjo
naeDRZvtSFPNFsk11IVSh4Z/Hc6pl1cKuYacnzYQPRfio2FSoa7jI4ANAd2UUaaAIxW8Ro2+gJcB
Zrc5ZGUpPNvlTz8Lz5o2Pr8BBvhZF9DbdWZUyXbuytW/t8PZnKrlzf8RjE2G2+Y9kkwyHhc0+bgq
HScwgjZjKytmgA/AvGpCWlhAW4Npm5A+uWcJTECo9mcpHefY1nU2zrjDzX3sz/hnmKAev9bUDo82
zI3soYwEE+2knePv1P/KzdV5R9mdLKVbj/oGzyPo6hlk4Xd7KJKq2L6weHL5boCqFqoZiE1txVtS
Ws4QoIY1BedHeX45wPEZsJT0AMU/Khh7ut+xWEF9Yr/5skxf2PSifiH4nGDE2W8ySVKb2Ikh59uo
ywT9IDrxDCUvewckAvm8uQg7BCAJ9z0UVFrZCtUGb/whrMfH/35mULN+Trv4r7HBBUNMw1qKB5m7
mw/gm7EtozNsUngCR9etCQ8QTX/zyJD0ygZtncH2SLJTCsFDAtI8v0kN2MPERc0PdBmd4a+yZ5D7
+5P1izpKgjO1aHwaeEIX/2iw3pQW17qz7rtgIplB1fIE/fV2D58M4lqAiFF+ors2LnWpTokUzUAy
k3p1W3fisIr6dck0QujLYHkQAyvwbNxfABlLd9xOp215pBuosGEIathelMvK63D4KncjaoU5ALK7
WSS/qLLlY398kGpVJh1rNGkIAGHtmLjnoLDLuvtS9he4WNNvX41O83Qtqkql3CBi6jhtwLFBQ3QR
qRIXlQ53kmBBwagHh3/aClVt455hRXf1T2nV5DLJLsl4ug0aLXoCJ9zJdrmjb1Lo7tzOr1r3IBUj
2W5sRX1YhFHhoiIqcV1S1TfEZAHMMD22jkRXGFT1ZbsJNRoJJU6m2YIsnQyejN3zkRN+mQIIbQ34
e+TVT9xpyTKmZdKunENOe4QrNVRYxVpVJaOgQiBOg+Rb/O7xKz8jejKDxTjLmS0qJtoEaSIThi3A
kyFd5hUiGQU91Wr9cyrWKYs1hQCPgF8Z+dCEWUbEsTPu51s27OSPqtTY3T+0QIIjGsj49K8up+wh
GSaAJzL/Oc7q/F9zoSlM4GBbJ7G4roMJsNYS48osllyx2eXG3QRzqnY9ZxXgK7OUZkPOpmuCot/H
6/sqjx2e9oSYMRiBFKEG4njs8rDvgkTVmoD9N6tAoaZEVTy0w4GbTDd3Q0klGHvHP9edLlyuhXOs
FKNbEePxlxykKzw9aMvJ0VyrOeVk1+1DAa6CvZ/mpA976xkLNDdcSg6VRKc8i8tGceJrmz6qkVd0
9zorbJ6h5jCcJey3iNlKprfcwG1R00vYbkZv+OqQIYwqdodk8Mkp3d9yhZ79NLWNYSG+z8QypzEK
kdaQf2x9YrvAocTAdJDp+erI78R0YbYp8oXeznk/xA0KasyIa4oSwIDSoA0ZpSOIXXN8W7T6Gp6f
odMp3jAQ5qw9OTNBFIe6LhOfF+Ss9j2vL0PDkbQsBTEX9vm2FIOTAzS9oM90tBYPo+0kg84fbCRD
9KQhQSfzyPByX4HdUv5L955zIPJLha71mJWx7Aeow/WVgiA8cvWUT9ZDYAE+fIF8Jjh+vP9X/AZT
yBZB6KAmw2/H1Xqb0vBbvPIEStr7KEPHtwlBnl9HXV7UDSAWKi2f8zc3bPY8NLd31wzx3QcTW8BJ
S0iyAgAUNXM9JnE/BZ2dwryOop0ntH7D1+crcgvJ7UsW01ewBn4QOqe3L3WP8Y3/uYxbCmV3NTzC
fTnW7iq+i2Svv5Yl/jQdopzGwb5XP1xW3T5nVnLPxTTfsfrMhbqF7iYUwaOHt9FDTFkcUqN5Zczg
3XtgjmsBpdzL4YnsAU6k7jXrS0HYYi9RLa6qjMlakaGrScUcInb/mLJVxNnhiXNAmiOzDHH9Z5Wx
mgDSG+v4CK0otequO6vxGLZbuUonM+uqOLrz/p7HZCBqEzhaHl6+UewzeriB+dvtmhyf9qBtNTC7
LF++6V1pOloR8tgb4wjnOS4IxoQp76m0cgxOMj/Iw7DcUQvv1wzg8I3+Gmi7SQRCB3FdHmvty8Vh
ME9dt9emD/aymu5TL1bMAFkoVMjktbcMrOrVtjWUWbIy5WgnDifcwi0/z35UGJ/hJfIlkxB58Qsy
jzm4NhoDL0Kc/G5PIgH8Z745tHaWnQb8Du6QuEzgpZgDAfM2AUSDQr6bVaBP3gWakby5Hv0+pf0m
O+SSu2ZcZnwkLk6hSbJhk60cYG9e/OodWdS2FVKeIDVZc0B8RNPK0fo2IqP6+MEoiItPP+HmlMXI
OxFVPaOzgT9ZvPnjkGnvdcDnHy52T+mc9kh9KC4oA3t1xi+NncKotlFUu9nz1RR0Ln0uccNVz2uU
FoLMFWMcSpyVlpNdfgMDc1SJBPkWdq2okgLV4LcPyDc33CtQ0fF0itfOHfzHYWRRlZkjG3jbUdu7
km6ER2x9bCFKk7ztXBsSp+PyrsakJrAo++hk0aacHF/c3tkSBmNNbyClGhA235dBuKatC/IxXh6y
KbcPpnChzzYgwQhTYIhSsCEKPxSiQDXYxuLSVd7QNDrOuuCLmwIRZCnI2ldGjZtR/SOEprMtmCCO
suyul98HcS7796VrJ3XYuoVeFP+F6naX0IomalkHFNHnccxapTZsgFApG9ooe4e+dbxlTefaUhsH
gi41PuLt0jnde4J6pbesfvF7Kak5oWOwV2Upuxz5rR79/iIQd7eNPASEDOgayHoezzDYjk35yKFG
cVuR5dBvaej8u2VRtN+Rtm5Dh2iu9UPaRAxe51HJ1N+rUpoXL/4nu5JjW87QWjtSmexmN0SFyunO
du0PVC3fRCFW6QCGTXMdx5zmQgN5sg08HeU1C0bY5f2FdeSCU8jT+aabPivO2gAfbPYIGWFxNa80
TQEQyWNvKpHHehLacOqrYaDywOAEb7+WQcIASmDS2U+IyQPn95Zcg5J6Xt7xCI4RG9P71ErMcUVJ
dxa5FVnBRIA9rJyXXKJYiRXKjqC1biyAV+tUpeBlV8TPNQ5eMDXSMSZWY0FPN9W5jmQYxWqtT4XY
6JbltRZzYPcUHpJYnoBY16LEvFF2EsM/v3TNqwyDsRj8AcRti6x1p5EXCG11Wm1JOiA3hMpmEIst
yFvHs2TykVCu0VH+g/mmD15JYiLAJ0D5/Mpfx0RNzAZ6fa/dJYxTB6U4QIbBOHTHGa0FI//YXQAK
D4Jq9DTYgexa9GIkbWZkK10UoigGkEskoSDxFrshtz5x4RmqepJn//I3VkLxODNmzJ2zT9JslEHp
eAFu1QwVWd2+JqdQis0KCQXHK9eCXJqVbFwFOZZk8+d+zT6rYwrcPdpIrdKQCgDyqhsC3rUMpZU2
9n+PNe5ZyH71p+5T3LSzZqzewxfOxAKXCeH9IRuY7pBJlCmqXqxuHgLMYXazJ56ol/ayxUsqvObw
jpVC9VBDsgDl28pbCPFZjzFZ9kUGHb+yfPaIF43mkHSzLoSFY6nwyj6GBka/59rztKrx1IPzWSip
kSOr5JYFUGQVoMuJpPwbSY8gOaqIqJkLIPJM3y6oYW6KpBlfNNaa/ZTqYCDwgDX43IFgxbsIyxc8
sKjV6LGS2kKd2CeyEsMYkBcpWLP/U4P7PQEG0OyHZ1K0PW4mwOT6OOb/bIaRxwRaj96zhWyphosC
aV2pFyqnm+d7ztTPrkpVh+eziUPfcURA5VSJb/BsesoBuzkgnm5MdlNpfxHddi5ggGy1vEhp+qcM
BcwOY88FOd0RQ0BCgj8cbY/KM8GXvs+cjUVlOHV1Ct0qiKdPPb3hhJ2bLqIhiniqBtbHzK/dGJgt
fNpwNjtimpQrq+zYbG253KEdTMoU/wYSXU59Jay0aLaqxQQjfsD8rkEwE2k0dE678pqe81nayM1V
Sf+fBGbhwM6RCUz5MYn6tOcMzs+0keCEu+JFOpa8MPq6/sA0C13rNgcYM/0YYHhBYD7M5FLqcVi/
00V9LlKlql6Szoa1pmj76RuOgmFli7JWhhMgXPlJ7FHU7TXzTmtnm+cKEnMNLciKl1WD/pG0BQz5
C7UHP/AsMpxrwjYQZYa+d3bK84xGcAFKRkxjLOHinjcd4vXPEmgpg+xrhNYpwAF4Ruu9FX2Ci/bP
zahtSjofSkTGkTUO8qeFuB4SMKwfrOLiCwSb/rsyFgUN2dOJei8cZQffWFSKRAhxVXkeKIQ5TCXp
dakvd1fiF1JHL7rFy27GS3lvLfLF/Uga4/hgqdovrdQiOegcKjBwyZlsHvqTPk2VWaF23N1Ixf+b
xzmhU7q4TY7kNKRjq1o/mNcjwxmJTlXHB0SdhGcl9gZAPR1iCwSOKaOU6qEQaklwXFJLBf3pFntD
xuoCaHPebQLZ0poenOE7jvzWyPb25ZHslP/5CG7b6BZ2Smr2m/kymx8uT0APohuPRivq8D9bNHGY
6VHzD23lSFbuPoEfISfSbWBbcVfP+RhoGtI4tKcdCKmyj2C9y5s7Czk4LkLJdd8CnbWxOg/aCm8U
qf7J6I2uebj4kIrd/qGrIDdADM6VgiIdhvDET5cTAIIkvab8W0Au5bKEdYyJOhQ8zYdJvQDRlR5I
g7EmDyadQH0n6ySMPZViXwg+5NA7EdjPd2TP9yiSJI86UPQpKbCHd6TJkNgifWX22w9uy85yxttY
x2H3ifDEUmJ1/zHIg8WjmtM+xSNouR8BaouDxRmWJ5hwP/ldJtgvKr99tBlIMPhufC0gZANNPLnw
GUMJCs5VFAcoRo21EsQARIzn4pz3MTpQPfZ3FlOkViVTn02VflilFCGtbqEVtXagzblh2ilX9kpU
cmqlUGj2qnn1N9J1xfgvOHA3kQ87D7fPCFGfX+Ec/UMfZl5owKgETIhv5LtXhxlHLZrGrZpbcG04
xw3mOveiM33FCQdVbn3TIyToxmyxkTnzi9wSukaDTRaelSvmNc8haYkb34DG/P3e5kHMMMuZFYBn
KoS2c+5bjqZpfRqz3Euk3ACGwUhfaXfHiluRwRbljU/PL42Z/RaustOtRVXAIXYh/0+dPkjkaAAT
iSiMXW3QzbWCBKYLVgKDhdaZGxZASS0lHjLEr7NujDrgZuszvU191rJhHekSikNOZKn347cT9MXn
8ahENsoahSyx90X+lyrckpR+dpEj+DkpZo5QCbZilVwDbD2Q9dqjmwnumyi1UPICGuQF/l/W5sDO
KE23HhJTEdfplO5zHW4HsGLOXHRxigJceKQDQNBcYVhp9bXWnZMh/EOCApP04Se2Ml60xc6c2vbf
c286EcBf2Gq/+b/JoYWQmeHymhZWNQ4sJwpk7rVbWCrUv6xIUAzrtGlQwPkF+yXWya7v4c0/QI+V
YAQhmnkIwEhN6nRDEBM4fOuRe+GEdTKDxeNw4oskGtBlPpHeF3QGyM53gnTm2FgaKNEKC3E1WinE
+Jtzjz82GloMFwHqD4Io91i+KpvNy1zmbq+Nfv8YxQGtZPfkdKr+aH0AyUgs87Uq0T16hFypzw2e
EUWeSHQov/YIzc7eO5z4WpzcBm3opEWPJEqZCH8LiK5pNNL1JNmiVcQHOD28zmmnonXu5faWiTrB
NdxK0WOWUJGzuhZgQ+RUZlp2zCcmkb8uysoVeapCjqo++M6iFCdW9O8/cTnmp3ZbB6JiLMAROGGo
/BHoIr2rvaqVoZQVaGRWmk8GdxHFFUh5sOPMKY2H3BT9uRX6OoNlefNf+9UNGPaEJQDeINkn8TbN
+q/1/v2B6/Azt9bkRJ8g25lT1IkoZgVFa8sNRfi/HOriqt4Hvh4wjRbTxZOrzdoFWsz/t6zI7i51
WHUNVhJ91Rws+aydYqRxh5IRVjszvNUGnMpsRYzmfS24BxRabs7zEqG7jhyf/tcKoHGK1YxuBQ12
DiOuPQDmqGCvK9woNWH3SYgGDfgBmmUCUxmrw91uEWzce/NiuKUarScJsRLQQAJTealVd9jiN0Ge
uBielWxKwZZawC2Uy+QLD32yTUp00BCqtIkXwRvA6CwpCcf3I+qIjGIcEuWTWhVvjKsBPFZLa2dy
vwWYmMWM9lvTOjCJ0hLUlMeaGpS9OGzts+30zIbyqJCMlJGlECzLHXdAqjQ1QErVWwgkkrOQr4f1
wWUC+6bGdhcbWC07HkJo3Qz7eEKOgDZYeaFM2L63O+VxZ/10tb6eFkNTRj/zuZdDmdJWGcYmHweC
DZ2L8YMkU9QzjGHDvMcsxJKp5XD1rIRL7r7w3XYQxlxn0DQEmwKHchr0stsLK9FJwcvKxxlplagv
or4A2hWD1xAw9DpaSDag2eyOzMIkMInUa2eU/Oo9o1Ma8aqqIhH8BEzdm5GwnzOndBWJFjECLn4Y
6puVMw2xy9FfUts/DGJxQzs9YVznuzXT2S2Dl4zcGWm80n1dfBCd1Kfqd0ypsjjhW/IGmw0Eeick
6/sl3UoA/ZzgnpgEuJwEhLY/8nOl7lXS0uby5trWQ5vAfXne753j03hZRzCwB0Co4xFYTj0wfE4J
g8JEM978eqkZe0MMKaeuiCLGAauiuJ9s7bF+Hgh7Y+H4RiprZqlcsdqEl1MOYefkoyqG5Y6ms300
NuGn79wNkKwmBJ3lrrTqcdPh6AOrrhj/HIzhNYyNkhT5viV6Z4nafSZz02jkIHvB1VUdecuStUQg
g0YWsd801bWMP05Ms7vuo8DQGgbNEHyIEYjVTZ0gVQNAZmRdTUsYeY6g1dPQob2hnx/i16HBZoO7
Mu00jSw1m483q4OA1R/htBCka2g370+LLMe0GjzK9rRZeND6XsYTQQRNJpwhGe2CX1fV31B/4ruJ
KFR/l9ftHjWmq8fBJOcDwnxCsUw9/pDwKkDaygHExFDplitmYhykK2+s/o7qwY/Jmn7A4aJATVHp
xlRQJ6yITlrt2LzMwKEP66mR1ZDVO9SmHVeAA5MylCYwr3uR1gVkiAnydEUaodNH5PnwW184yqJz
XQg/70ryOAmKiFSsVdChjP5bo0j7wBX4Exv0e7gE9aLcTVHPCen+8O3aT7S9IvA4HBwy7oeemOGu
77mqaL2rZ0t1bvZ5Qu83oFpt4+HkKW+s8DIzlBzR1RFh2ossi7czP2fjnOPzBD2nz8wJeOzjjEr4
Wdh2ZAzDuha+AzRNfkUpqcrJFvuWqFopa3aGAyWL08Hn/s51SbcQntJrkSjyIDlaiehP32Z6KvdX
QX/doXuDfzIo/5F/Yl2fxPhYl91BunV6tcSW61us63nNywB9+ogGKAnDj+C5izly7wqsfu6v103S
QMx34ANq+jdVjA+nc5jJB/KhuVfmHi6W1Z1+7KFG0NxhJPCXWHNLlguz7Y408qAB2CxFOMCNhl+m
sOWkv5C8lceyVrCDv/4c7zvTBphpKb5QY8GfUwfd6C2TTlpi8sjobN2vDkTD+UxONm0ctpT2fb2A
re+rGXXMMPvchxGpGaRl6x5mpy9Yolut0ZZFYLCn9ZcDdGPG61Ea4Y+4WfP7hw2TRoiVu+jjqH1L
uRLkcnBRwG7WV7rfWCqkrRMT85yaRCoVq5ID/alfy+/yk0bEIORhnLBIQa8B+RCZkcLeeZeHBuh9
DsqLctI9RV7wRHQ9M6XIZFz1qkYp+LvgHRGR6ChHHTERsQ/rMrH1fDqHXVahY7yIvVLw7j1q9Dr5
FVYr4IU4ZtQWVg/Lqb3GtezHCP7LYy6ozTGocPFqFgpJ67gGGnlvexXp9u4xhFSdegGDYiNQa2M9
YKDSoKasGQJb4PnDnSzQIDJox2lq4351J8BcNeZWjQaPVGZzv5VZxYCXUI1yOpgM39dopk382FLa
dj18brhIQMZt8v7a4HDB8pGg2Y5FeDlQPlzH8SID1GhsFPBO1yMXs3j5hr/LgfL/p4JMk3jWWTCn
Y/4jASGPidA7iIoPu4bJbzF3tsF4y/Qv2wKHcp3uWUrOtnsLZgXLcDmP3Q25voDlNQVks3tr2jeT
oe2oG3dYSU++uTdpmg+yMBTc8icExF981far8kSQOcAZHZuphHBZ+AkQY2ThVMCQ5CRqp3B5hvSF
UEH8gI4QfgHx1jiVzvmB2POxdm93+NodtcOcE21az519jSauorrrg9S1RFc1fCIwn5n3kg9v58kN
ogTUGQtj2Y85kkmfDN523D94SbwVuFEcDdWB3uiSq2XyHZzKxrrHDJ451gG1hkgmOeQ5mxrIcwAe
76XJ+Rbl5dfXoYPXiuWtTRfTRSk9/dr9+XGkX8yNc4r9CJlO5nC5SH7xoH9YCE+5foxJqR+ltP2w
I/H3squbUmvhGZNCefn92/JRO7B5gZa8DrIJEX28TjJQIcK3r7rMXA0UzFnBbhotQMXsIZGZotCO
BHUx6YfvgQiDRi3O2RVuwMuRrVL/ST/Ah5OeXlWwRy1cc19tMwvM9DpXTFul73IFLz810nj9/KLx
BvxIjVmE+Sa81y3mM6BkBQ3jpEoQiFETWY+ySogecP1x5uaYfT464rRWcROgUQ0WvRsK2tSQY3xZ
gL8RDXNA1oNz3LyRowx5H4K0MQ4+U4X7njG9wwSdZcaNbYvIjvYEjyFWvqPYUR/DUKzXXw6Fn4We
bhQ09uQhVPYAQgHIlhlVzw2aEZdVjPvWE3NV4MQA+yR9qnaRn+UBXsNBtroPfTCfI5PIq4RC9lgQ
Ufd7XvBmUlqMsZBAS2uUZtmwX6vrtWVmQW7ncy+MUw4ggWLzDOqRq71nK8UzY3+YfhghJL5OCu1i
IhPT/Mj+cvNhEQjDrOld9zJGq7ofcY3iaoIZiYLceMb1uF1mwWj2WQ8vnjpoU7s08vMHicMQUmOC
3GS9GC4Rt6wQGmriUVNYnGxUNBo11U17rPSd1Qklzs7c/QH+6fqhOaQN2eGrBQWmnrhKCN8V+Dqi
Pma8ZRtyrnPzo5XVMzV0EJBu1rJ+AEPPnabPe3PuDyoX8/ge6LiYsgZR8kH2phcmxrfWslEQ4ZIe
pdqVFuftiMdFglbEz8ZQMgqwSxalFzmCoZOnSrG2s1EyV5QbVvg/Z+gcJyluETm5crqJdkPM5WZ4
Sa486pHSnELgK1yXBDx9yKhSDScpw3dJF9Z4JS3Vrg7IO9Du4w0ZTteQ3H3L2H7/5hyZFm5dYt/S
XFaQ9A7Tcbt6JeDWiR9fWHGlvVXmkZEyPMXeRiAEH0WkIyN3UQ8QdT6rMIs3/yKtpj8x+W80YjWd
gk4PLfUPoNFy0Ph+1ZqdzGqdwWUfJZN8c19eTg8j030jbxLT3Y/a23bohQpYF5fvDdKMPbzTu0ch
pQeSD/+uoM7os9PLaNKKRBEzJf9nW21rIqXVzcRFwOiboVFYfWBHe4UEtouW1/4VvKfKEZSkums4
mVAZtYkBX9ZQgv1L8jJdtHfXNEGZEkrQQ8y0rieDCAMW5YDAAgv1o434719irCOpBdeLdKR08EU9
31USmjMtJCM1CDXvaq4trizmdU/feGnkGPcJg5kvJ6bQx2GvY/lcWoDJppWeUDlUICG/tk7+vxdi
FqTVBnnKWqRebnnmX3rsMDVIMl8Joi/uLW09VntKwh5Wr3Yb5hU9aag9UGnql5QdUviIMFdJlV8I
+CCvMCgmPXoqY7T3ZWVTe8sv5xVwMQiy9zR/MUF0bXA29GzrloHqUYUcE1KDLX1CZNkAmm5Rhe9Y
KVXprPKsvq6eBoFhpMejnZdU4CB34MtAUfwpu2RWFuPmKoXRVYaF6ssG/xhfMMXE5zE6tyH1EfaM
q6HNKTQ6fXbjtFSpWN7dcpZg69zWygucfyUhaa+uE22Ef5xpPTGLOOdYJ5ANgxV9AW+0f1KHJHP0
aHYcj+9RtjhQdOiiSImCL3pFa6dIvlP14iMG+RjLKMvO/j4tOuYlOCLZVfHOn9kY/7IW0Pyfueuk
ONV/x++WVcVxJglZnrdxXqMxuDwMAk6ZBPPN/KDP1jK2nLJb2YwqmaICpVFMuTok3J9vB9jFopNA
jY5U/FUMVfhbY58pLBunJx4TGjTGwfY9rS1bA5uJfGCdImjuWOUE1XiKITTexJCHnmLHsssPcWi2
wVNa8BuPtWSG0D//xpN7Ymr4K1mvw0Z8s+khgAJd+BYahzg9mxeeJqI+aIh6bl4JYksoFYrCvIBW
RCIPI7csIdDLhNf/wXFBdQARCTTWejcRIGdNJAtMH3XEqqYPJ8yIALzRTEZPjyN4koEvDTmHpdQP
FYw8Mppei/jP6LMdDlduQncuLwYiVfGKo+1HyWrJTbiudb9FI8GtPJ8SCfF8I5CEA+Dg0PAX7avz
wm+zwLAMVAru9xyL4kUrrHSdrLOhpAx3NZ++iFI7M3Ab54ice1raESUNscx+4XBs6g+DSD9y9uIQ
sx/kNtkXPcmms+446AojWITXpLkEmXseIZot2Fzx3gJygLjf64fPC02GZqvQTVDVaVuZUbISRSkY
0Pbj6obPYkwRTQKjRh8raCanZ+ZZ/K3goiFeXeYaBt55Be8ePGfqrbCR7v8B+cXSCbHqu0/8z1oI
IVRNKdZy1TsbX9A6PIJSvXUSp9QEVb/GRZeVsFLGfe3bfonE/PYPogyWVr8SB8p544yq7r3z4jG8
FePx+2LfUw3MEKGgHk25FcyxRkb7KNWDXDP6YQ3df+WK/UBhJ4Ob6Rukj0WQzmNqlI82jsJQWgLn
y0uFQFlDF5StErFeHAKdEbZwTVxOEL9DIO0QCm279xnC/qEZnaVQm6LGqGbeiUMOLr9uLtma9id5
C0zldF6/isCY7dOKYXJzi/D3eMbX5CbF5Fwia+WV972SkTP2fQXBKImgFDAOwGQ0IOP8CQJ/LXih
TA7m75aF2N22keHsLq41Op1wwOCqAKdCLaRwQGJHwoEEh6ExIDc5NPyrjfY1s0HWpe6lg6R7IbxK
G3cE0K6jjZiHhgL8zQ2mVAFJeQzqugukPq/d6SjOpcqkvxQ5EEhw9tMeKi4SXS0WCs/S+01eCM3F
xs7d9qfgbIl64kxxemgNyCOKTpU3WMTUlNNzB6L8C5JRL373e5GQPUBU/Qzi2ZDZ1+qaW/jl9uXs
Jf6dqDqdF/vUrmM2vQCl7n+ct51oLy8U1LUSEi2KVG5IroKXkvV+y0ENmkHJkalFzdyLLOxEnaF+
z/z31gaM7SPByHJOwof2S41KVVhpZFZN2glyVL1qvk9IxNSbQOdgYrryn+sKibsversIPc8PyMP/
CTIcIGbcVO/CP9G5LuHBz/9Z9wwVBdJexediq8zXeW0WTqrdVd4fBim1t5797XAc1iOgqs44bnUL
D2D0yk1iIuGt3pyisWcxIII+jiKQ0Y0xj4FJX+ZLxVU4xX+7id0XOf50yx9NSN1/EHFas1HQvKx+
r6zPBJAGlgEO1+rH6LPMmAlBY+hMdYXtKsvePDpuzlLUJ0c6LYHqqB9UQ2PaeAQUiXtOZ9YvsUND
QGXDeby939/+IfDxvXrYoL29sHO00uXLVfb3qOfH5sG2vX96GhpW6GfY7jVPk/oj4PqLvASQTOFt
t+3FdGrrTEIddk5DyFvw8WCcuP6AKS5BpvWx0TmO27t2vGICv/TgiCf7IapD/Gov6wmxna7uSlCs
c/S4phPj/VInOcxJKsw8S+YRbfdMApbRqSbvgXPyMlMY4dqy3favfA4BwuGUUuVvGEfO0SYl53Ew
AhH4q8ntaQ+PkK6hPt8QYOJZoE0E+wrX/Vn0OS4olCLc5Ci2HR+gNOj7beAQ0pMYH5+8BqIyO6PF
C2pRX3YfevBJxwZrgkNxs5Nw0xFdac3uYrdE0spnDgtDUC+n7TVfX2EmJO092k4b2EgUjImoIOC0
oQdBSPuPPfmHdKMr0eJpM4GL8UWyPCIvxBfqJS91kH2vGMqku5+WVjtepiODTXUDrtSNQlgcW6bw
Cy7TlZT38fiG8CnvKENWu8dMBBWBcW3F8dw89J5vODtqBbVOPFtEuR3qYYhQop13Y6MAaBU3MUc9
Gfuous8PGpHbSmYbQhrgIXREZDqnTBjUmb/ceEBoCa4dwcremlXJkXWicfn/b2LsjwK6g6wJaXKR
Q0pJpOl7FZvkMJTAZLdj7Y5qe7WL8lwsdqaixKvtJaL6GarW5iOESYoC1MmUqCyJ54fIJFOxEBz4
NWnxfyHav3mYDQg728NOZOdueeBYZodBtZ/xWWox/uMy05FiFpW0rw2JUDcB6u9ot5V268qbZMSE
WzZQpslSfU/Bagwo7HdBn0HAfSbT6ZAz15i2w7izL7EiIDU1Ed0Q+fZMrycYL862/UyjJ6YcZWTh
18/TveGzsJME5PGgSmP4paho4EfLOLF7aNEa5jY8DtC0LV8f3rVClJUlrGLSpVABXeIpoSrqo32G
o1187fNm1ut7fOmXXa4tg9qqAeU5bdpG4tbgXQYnHyvuGYHCzQegDFzzKFYdjg+DM15VON8l73Rp
znX1gn6SblterTnEyAXgR8k7KaIltlUMc/JAsMdmFLLqjkU+lT1AcPYYuBtZCnVMbpZnM/EH50T/
ixrn2aL6UeamCw3RBUv5tBarbJb9YTHjn4W4yDBET0SAJGFEizrCIttqufAMBH6x2h53/feQt0lt
4GowMEVwIwuMH3zL0AnY4P9r+x4EC6L6Wlyo1zH3b7y3nAD2W/x/HY1V6+eat/Ydbc7rfUIDjfua
t5ttZtCWaJVEtr0RhcSIAcfZZjnmPdGkIOXUBIE23+pUhRS/KZ14c/RBlRJdJ/Bkzi3czYXZw1u6
v+TXi0FW0b0KD9FoKGqzwq8uwsI8ZpNWcrygJd1wSyB9gaAODsF3XNHP3E34TacIUGBL7+2J7SUP
aSSV4WBL6QQW7xq5IqlqGOgEznlBpmUVDcGVMNQKdc0/YzK69afjXFVEoinbXHhy8SW1dn+3nvTc
z/qjhx/iXEGJGpkz81yJudb3cCOWvndyx76pozD+NVe4iB7WORa3jpySLXITfa1eL1zc89aAhTxV
ASRGwAarqZWpV8wqOQ83m3Gp3ujgM+/VLPm0JY/c5aTvyvquXi32L2YSC/oDWyteIpBMufeLDetL
/FjVf+oM+i/TRZ6yoJu3voeQXJymBVdfNrN1yQNnC6VaygmVSAPiPBZ4piSDIJ86FNHizM1sctXp
u6H/1ibPikvbRzElFn/GH6nO1dMpwHA8FLDAWyOIwnG9ELeIDohqPNueYFfrV+BvtC98WLuaKBzi
qXCE02bS6OmHn2u2Lc0V20bjemNxqyAlqpcTOXyiRJlNEL/Ud98q5dhcsI8LRtBUg9ZzITBfv4RY
7a06XuqzKRnIJ+4K9ys10takrgwV//+FKu/Ibzn/OQW0w8OA1KcOGrpdpd9RdSNIFFNVxkNa5amt
1G5QD2nXpuJleoY0PJ7gxkZDQIi2kV3Y9zzSiSCQU0nwfHLFx3MKZK0shDS4GuPRBjgzw6MDkDqk
TEa8bDXAx+dH5Qz6gSevp5Niaz7y4kimaPTDLp2d4aQVlXn/0l4TLGdm2UqsUa7G03J2e26ui/j9
mnSACzPiHhvBaj4kEb0TIVOc2Mj5kIt5O+PR5m+no3ciKhH/Zwpn10S5Wl/VTRwW/uOP+JxcExyS
Gf/HOvU6OgYl+iVrqWTN2Jt3Tc9cWaPqu/8c2EnC+alNKz2u0NH3N4OO++9YRjZLvzbBv808/+rV
4UY7XMLIH04wMdHTERN8AGvfZPWNoMCIaqLSC9jb8D9Y1Mc6BtyfU6B/ht1eX6DecH7kFVchbmeu
iZfg1WZsRC9+aZcHH+TNJxChmmtjaEJegdAxB/YsKyROmskQDJdhM/UKKBa78g/XPgROFmvrJtGB
9fzczVIKN2ucmHHCL7yT6jMpq6/QHswyGoYHTPo6MsI0dn4g0eKgSQIEAdfQ6ziN3DWcwQ1mYtKl
ZZczAPNZE+YN6n+LS4bSgJ3hoRnqhR891iKSSUItfbFxTX5dHazMoQG6H2r8HovMoH2nIegS4GES
8OkjX5OiiN+Kn5ADjsAyJ8HXLc7sD0xvnZK2hwskwj3jYKuOCNnuCNqjG3bWYUA1tMvKxXcPjr3L
lfNaTojZH9TEk8jZ7kr/Q7mIma289zgbKHf4oRKbK6a+HDYo1YvcWm5QKa2Mf1cnwwrY4s8Wbsz3
TA6Tmiszqu+uwQ7TtGGTNryW63sxNkFbAFymOaZ8HMKeBkBDBfXhtD7YvZ1NZsNi5yaaf3BNKxWp
ctQ2EQy03xm5lHY4quyDI1NKoUF7zyLXHry8/i7Lljrq/ZlpadL4gmASxKGeWsa8VG6/Y+20CKcZ
jELfreTIwDjbz5ii42tjcQgKVcuzU1PuWU+mFYCWcuUi9bG4+2sae/rtgCQH+nhTtX+0BX/u6UXn
28CEaFdnqbUaavmPmsX/6sbll9NTOeR1KSs4eyE4hArZ9tkoLKEOTDmtyQ7yC5bRUqz3DnSg/esd
ytTQ9+K8geS/uClKOaTgblCsAhgrYHxGn9BvgS8KvWI6oR+Mvzeyu8FyxrjeILLMGXuc88EHrApi
1Y5wAuldAj5r6B2JcJBVGlbvDOYPHQEeJ3dUtV7hVeclKiya5CwWi9R5lsLk0rIwTXswPjvdAXin
iZ5KLintyCp6Lm5Yhmf9P8WqY6sW3TyRKm2N1c9KnJGRm1C1C+AE2GRFCVzIdXoAukpaR3L1yW0J
Vf5hEZitufcwnRHCehPESga+jreT0viCETzgKwhV+7xzAV5kqNopmoCPGUXiyBiculMyh355jZtu
Tri8hfMrOBN4Zr64UM90rMlfiIT4WMMmSF/Y6DIqDwaT46gUlMVy3CMdBdBXrkW1gut8zo1SGifH
dMiqFCJY7b7AGCJgQsbNlRD54axv7UZCP+QXpz4Nzk+u1ylewB5/m0KlGVBzTpOaEww4IvlmWA7E
fbH9zIXMg4Uo69xgmhcPEgJTbu3NGayYv93/rFQDfg3IHPdxHthI//AJSjuJw5Dcnx3jzYpdtV8j
rLN06BvkxGgLN5D90vk5sbvGmPiJ5Czx4iaYwKQOOE0VSyDCFxvMxn4c3DeJ6SX0qQWFBW5K5aPn
3RSG9gDoBBAyebxKpMQjyG6qhBWiYAQe+aPTvQnwBDHZd9yHo07vib9mA7iwbwM3D0R7IPGTz6az
mfoj6pC0B0wMzIKsmv2LPz1wuYHK+bKTqgQZJ7QHiMimEyQzO9D+f/1qGpBsi0ydwj0WDDoeeGlS
CLSe7mrXuNKu0kU66FV/cOVykQXK0gqQkTvTpP3X5ds03PPk+l2+UIM7wkUvabHgWqK6Ms7y8jm6
Ix+DucTOCQI0u/R1ZvbfbskhF5KXesQmrK/BudqWAcYU3lA8PdQmQ1I5lk1JJDM9/mC0D2HrTQyD
mRHIMzeCU7YsNq8YbZVP/QAb+I9ZW+iedUC85yFDVcbr50KQHiTvIYNsizOo75ZkSomMDxuy1yG5
oX1L1ovOm8zLmZQSqZM3MyrwbGzbQg4OWx/CL7ITCaasRv5iNoRXxkNnjGtirR7PFvgFNQH6bLFB
13EoQKAg1HRbhaLg5DkdTwHmHDHeERM+bGil9lKR4HFem6HsZjMNdvrIMbi3xL3JA96J5fOT6Ohn
Tvo/FGXaV8VZlgqr6Yz7hnCpNvH5wxsmkFCEL1pDn+F21WbmdW9y5lJV96MTFYEaWJyuAf2snc4N
vhJOJgEqVkq6yOeieVHVcjqfmZQUtQWkqMyAZrDMJ9i2MaLdYSUtSrQdIFTdsoIhWqsAmTkKFFAc
/vlK9DskdicpfNuruy46+DXu++9lzy1Zap/d6cg+sf8JGHK8ohdfmaFPfnGAN8lvP9P4ZmC/tiNg
qO30YFBxe4mCfXyIjwQwkdO44p4SJe/jGDkGE3JOOz9E/PPmmlNlZyfrcOleu6yYEcIj/Br/BscG
8lk3LxF8RGvyNZ1vHRPLHnCkKovhVM5/+ta+ECFkQ04mLFIWog1nq6/4FTj7EfYP9Pf33wt66h8Y
SUb5cz6QaxzCjXBBZUB9cE1oNXTXQhgUU5Qv29OQWEtv/4489NbRV3zOEXzwkoQNVulPEbkEiI06
kiSNg47uHJUes1UKwGsNXwKeXD97USvFUZKQdOThbjuQnJfWdjmg7PBbpHcCQ/50FFkfvq1p3vpI
vsmD84l8PrqKdVrQ3dQitCWgy0hQJzmKjebt5P39mx50zRST84OD3mBPUmlfrR3Nr/wZSdPIZF4X
tVEVzqfME/IpPoboMnMWWLNheNMcd1K2ho/BigM6Xp4c7zGmCMHYAx0UDU71AOpwEXG6zfYCPgXP
fitTE6GNgkcOPtLMWTSTTAD4ladBCwjvLk0xHO02LUZV1tRAlihtYKJwnEl9ePkByC/6wIrD/OFC
1IUvZDRvWB8d44cw90E1cZWWmqEuXYu1vSNkElbYjkTr+wc9F36Ao10jfuawExrfUc6RSPDtAJfQ
zNYlZowCOu2LZLOyo3pjKfFmSdI5Edt06ydYxOjFpBDcLRjYZAT0dlR5ciFJFcidbMUfNdB/teYR
VrMxiGvrhRBlVCaEJyeveGMkgl4pQvrVsGTdmS23PJ4CVIf0jmNcsKOHRG5I7lRJIUPg3qVeRuey
G0yad77N2Kbuc6al84poO6ls46F8gA4YTnae+5H6ikhY/UlScuV8Zx3Z5gChz64rdN8O17E4qxAs
JYolNMp+kq0Hzu7WOfnHfpPIyxO+VIHZh4gbnPgHtTPSD2oVRgpxKZeVpTH9HYz6ZOBDBhym9Yy1
SWp2ydJHhqqK0UF+OnZ3Pb/vtF6u0A2nkAG7eFwCqQbMEYMNtE6Rvv+fzGOHzbu1KE3uYcDVcV50
GHZJndGwJRVfnL4QXRamNnYv8GyPXUtPcxZAB8hdTdDsFEFb5AO86/DnzuEjJP6eYxh+oLxP73aY
gfvbCN8FQpHMbBoTHUyhINak2ZBqapFViNwj6lZU2Gg+A3Crz/NuXzui48B/HBbTc3UgWP4UqK6i
O0yZHiCTdvVB1R1usAXERiXAhXU+BGWMd6gCh/3cbL+y/jwQ0JMetcsBClsTZgCXmjrpTvso/YnD
O6HgZ31NHlEdxj/m6Z1XUtyGEjVHAjCmvJhjWnGUQksMxxZkTJSWClkJurHmwDw2YsW3YHq0Ch1S
w20BZIKjx9iUMyiK2TSbCy/izns8sfKKOmkBp9T4GykiYCq87SO9nygIT8py+GJ88s/00dgBJWSP
cimtvQx6kg4KEtH6sa4M2YhL4vPn6Q/7d/5lRX4sjT5FHNRCnM3MbwMUb6FkPdJPVD0XEu466rIU
igNJhw62CHav2Ab/VaLgC8aEtcroHanodtee9BplTxu6VLcB33VQBtgny8lzCI809AwvSqQ8BKRK
zysQXd2NP0zdB4U1USxzb/QRrc9PNDN5BJJDkl/VVs0i2NhqNw4W7fpHpY8O4o3WQw5a1UqlMCS+
mB4Rhg9TasQqjzzZIgBGF/7uk+ej2ZedEGM55jS1hdUpbaoFGcIyA9WEi2gvDpcZ29+2lTrEHPEt
yI2oywCpWCLLgAh536cBtj7dP+s+KEzltYZpstXT+jwppNckvrAJNA8qo6tIzT7IgcTbf6kXev2g
bKDN82ElRTLmJeDkftLcG/eN+rlKLczoD0AryZ3EXavGdJ1AX9pmugYvn0YWW4KZYHrO63KmRNJO
vns0kwidwwxNj2daeLpcclSPAzqlbd2eZuvlipTEAPikSkkCvKRsY0QODVyrzECosNBiDbAD5bVO
sHf0X/UbuZbeGFw0uNgaW72NAEKz+IhJ8n5lGeCV1Yvhh55E+XgrLosKcS29hcTpEYCUOsaZBwW7
RhTlyRzRUmqaBQ4wb+yC3IovDP/B1+AtIzSZcIEVzS8MYmvnT1IA2vEcJdGRTlBluNjx5nr/FkY6
y9YgQTUf/WhPdmQp09c3vvl7chtWIoKatJXL9862LTgJxBnY6pwgLXKbdj22ftWiOG4uqE3yz1hz
gqFndq5cHqIvwJ0RUNX94TDeMrgxNazd7dt+ymHMj3UbmIk7a9Eqr7Qh52kHCTWB0538i0P93na7
8SIX4V9xTWeOWoPRyejcofq1yUxivDhC68LVFCtq4BZvrsMgiiW0UlF0EbVikZUG2xsfprXhHVRI
vnJYjWJZU7wz1p0aUiNvYq0T6nTqAgzj8Wj/eqyLqIPigtL0u5HnBx8vbs8hSnFxso4AxZ7m68aV
fvwMSVodrMay+ADpBGtYRC1SVbyucgaadMgKnGnVZqZiy8hz3YWAo3ItZN6+B7arhsWVL/3ZGphW
jMrVkPmqTfVTS9aj6Zh7SdGcY4cTZyUduBfBVpxiLaXhYjmAWvrqYeqNprVwqWn5Jnp3+p9S7aUn
Uufvdow2lrIwvdLYPRr2EgejD/fqrxJ/EbsmCK5OrVzCH7kUeX1jBAFwxQ7Qnm9s+c/PWCSvrhSg
VnwjNWoHgEysIxixVjWqqWngc18+/tTdgXUm2o7Idr//ICilog/cFiZBKH8JcDixSBzsTj7XlHjk
jtMwcrG9pV5TeA2C9FcRMPAwPy/ysBioNRaVBeHJm1B7UkE/f3IflnFXEmxJGTowaavexHex/Sf1
T+7fhWfgebUr9ctqBt8HruU8A6Ws8xaOpmDsE8tpJ98eW3ppknAkoZYlNgJY46yI7ElFHr2WtmAb
cfRXOwE40xWkA8cSyey91R5I7XzfBTr+OxfpWZ+jOb7VFDKl+sYg0oR+NuNkZfszAuIkkUjQ+pOX
bsESJPaDrxez976tw32ovaHxnOBEQJjZUT6U4zXRkSELP6BTwtepjqYY3FuVdO0i11qE8sXXvehI
iDxNnuhj3v3dvrRXpUJSvj5ltnIAOYlC+vYkwhA9+AAlg4sHDVRZXx37F2kJSQM+ok83veoZvBAk
HCkRZV7J98KMo5162fExtjXQ3Nw0XDXMxbKqmQiP6OZ6/DalQY34n4HEO/RrmXyKuX4BvaJq9FDU
Bh5sby0t7sd7UyGaPn/d8PaZUUI3JDfBx5Lq9KU/Q65m5/Wk1eufPLRrFokO/hHqBuXqJGCp7BNy
4z65fjUHJqZ3IMkAzkDjXHdA/FQitnp+E5wbFBlFAmQJ7iEkeYoQ0o/WTjNTJYhcsATYR/v2QRmL
TZcV2lk1T662PX2fVM7vpmo/pHzOuF8ugCTXZm2H7qCI2ET/wgOTQwe9+OqLVOnRvZjQmZHaJMZp
87MzA73BAWxwLPy63iMBRjpJhOH9s4OIgVgCGyzrvTPRzqvDJCxWxygpi/wNWidse7sZb/2BbbIe
Zxv4fViFRsFemfMvKMVcd9B4YtO8wdc5cjVOgZ+dGVAr5odoczpxcLwqKGeITbVZsSV4o+Q3Fjz0
0N0671PNQ5OSaBQTnCqxFbSAovOCLuvAVZPITZVCUk74OBn5dZTgTZcVHqCWHOf+wgLv/7PJrEc8
VcdvOYfVJiQsS04WGVUwABjiXWREWD9b+GMB4aD7yNBwDqMNEILMgU8RvSQzDEgI61oO3j9EdaXf
mz8Bc/40/XiclZznrFUk5BTBTJEe4nrGBpPCK4YglxxpHfGFQ4Egi+9khWCc7q/Z8hS/aqz1izGA
622jF7Wxf040GD3gyrVgQS932DqVsc6NbUOa6/44FI9YoereuepiYfjORzK4nxgK4eAj0bsFNWxt
Ks5gLqHBLyXgTV2KkL6Cmi+EDy2jDBJ5tj8jsdYrKbI7A5d9b93/8Vvk8J6zH3NB/sGenptu0P8D
+rs4pawnPqKA50RCx35HJXprpp8DYVpV1tgnXgI9BkyjJY3+WYJWoxkDwhjjXEM0YsZP5OzH7hgr
FfvNDmEdaDgmMp8+cUUJ3Dm4qMT6xqNQOh25gTXplcfmaGcP0pRv0dgIpkaXDEpnwQEBRZZy/yNR
EVXq5PGyujRzGfsWdWfcG2DOsigrI5Wp81nTWSiEppYSFLxiEXqldVdVBzjqKyYhgGGA4k2SSYv4
IFOEBVis2SUlX7S9lwtOTWqxhdML9qZDTZaWsCxorCYmkRvLbSO2joobHbbY6sdoAF+wyK1cT3pz
OooI5U4XpFl8vS8eoaWdSvsSaHszJ5OCD+ljmb/pm9+S5lOX8BYC53WCIRXqjqJEsU2tD88M9cjt
NgQdazJggiY1gFU8ymFW2q+nweUq+mpYKG6vNlt10dP/fSyFYOalNKn63PYmZ24xNBOGaWX+bnto
4TRE99nOWMQhLqb++HiEyWv4v7rtU9FtBP2TJPx8zULnRkuGbKSym5zABslX/yOEkZRJaRO5SYgP
+UWBGr+Woo8fUBSRBmcJkG1W+xxZO8hjTiaUtlZv0oK0QO67BO7+HmSMYG7WaGi6zRN4ZhAmHL5S
fGpFy4+UQs7CRX7VxT7maN86yAP3IhVjqQuMZZVMODiyJ+CuoO64sj2Zq3N9yOAVZDvl6eAp7zZE
jGVF603q5vYjkcosCPO1Ec/o7LG2Wn7pTt86hZESdYnfUOqEH+mu427F8VzC+SAMFGGYV7VQWl+k
daEFI7iiYkZvUcazMHjpH0dnKBnjb3qw4clUR6RhEzLfPTFXbB4Q08GVgi96TbCkC5dnejDLowB3
aP936OTHYhveV0oyfD7QrrG4UIGR7y3r99611cFomxiDzUnEky48R97T7jo+mImjl5uwk7gCToUg
WCAcr7jiZX9whCdKkTNbN+7rtsAJbvno7n34+c5/bH2zTvo+NMBsxPInMZqlGPuvMHMhjffDDIgf
2+2nQAIxqBAM0GHm1B4qJITqPIXGjU0lFNMs/sg0RTZN/ob8ku/ojr6w5BgkamIRaiLLgcOAblWc
6i/vse//K4/IqXmeQ0ZTyCZecvh3RpV3rJe3khdoDMJFy9S/tvnLXZeAhDN3J45EL2P72i/9nFVH
5b3mI7yPhL4sIY3a7UFPq0B/9cnwl2zA+sJg4hXi8krSs1bS1c8MKeYR1rdcl8J03PEwPhCfV02c
Ww4vpNjxP2w25aMSy6rCnK9WJrksHmEq/Qly7Almylj/o5qZjPzWt5O44D4P7wV2oEgBql2hdivA
N/saPuJaOkKcLCYJ4+wH+IbIAw6USbNdGy/YzEUpNRCmXm4X3oEns4RQ1g4DHILnejaPQrmQDaZf
Q0q6mfFG+ppn3qF2XVeGtg+f//FU4j8xqyuQ2nH0uZ2POy3tOo9kGmrcgRMbIpX6FDqcn76JzLhK
oN/JyQP10gUB+48vVkQxhiZVttKK3IJSyT8oyogaOiVoi6r7urKcRshpEHsTAzDaVI0T3V28E5g4
jz7kSOypGi5XPk7CdGI9U5e0Aw8FgWJttoyNJNoRZk0ziV+xOcfmJpsYoPiipNDQjrdwM5y1GKcc
0aiL2ujh9FcCva1z6YQTN5mTnmhmXveMxaB0TRqw6B93h2+KhFm/AFqjrwOpJ2VYIYABbJy1GAdM
m6gg1MAnuquzuSrtPe/qBavfo0cK0OkbDwSglf5deDTMQ6J3w+xGc7wKRPd3xlLUAeBtdnDyFURx
nPIZdJIex749H00LqTYwl2nBO46otTrUUgA92MDImX1KGr+zBCt2daJ3L1P27tb4A7OVnn30hw+R
To18EF5e3m2z+Kux3Rm19SmPDSMnIcYWTJUTtrNZ3Kv5DAsjD2nwhD1146Fs/UIoE/LzJTDKhLkO
7Gqslh79crXreCIMYA4JGGnmuLTY8PeW0ES+iszrB0ejXCALyunIVvFW/5QgCNvI35p8bjUsrfLO
KnLaoykFLM2uElZyKqwtUJOMKZfie/8C05Lg4rf7hfVDOmP6sCZU3Hxrd8Qn8qjUUu5BeaHaaEfp
iyiHY0jtskh91+RSl5VHtRfpo+7q3h6TrO3IkHdUKU/cN0JqrzySS+oJ+mmvnpLjQEVOEOYOqLMe
Wi99xgEzfkHs1ooL0uq+pcag2tWduvxC6mgmC4xLeCWKH3SPJXZ3r7CKeIDe56ipEC+r6lgrIVGW
7/mA6JNCd9yw4sF4k0avaGjp/zEWQ96yEYGAwPbLU40FDyclx6ucHtsKVkdIJkQwrhlS8kdOrjTj
Zfh2bKKx7zazeDrPYge2R6e1G+WSVQX/l+CafoAnKrQ1YVpVhuzvR07cWSHhENwUS4RtTxvVVTrQ
WU9AlYWPdrcqo/GjzwZYd4kcoGqd8biZWw8DK5SVWaW34Vh0rfhuv7MCHt4m9i0QAXp29Q9jnadi
w4Pgm+CRhOOClC9PritlJ9x5xdoaLqUQrC6vGbLNX+y/a9yhU73pUoF2urQdsajhzBfI4HDSEAc8
B0s2a2h2G2Ihy+CmD588fLEwVUxr0kpplJitt2HXTZt4+e/2APhNbGkBFerVMOotI/eK15BKffGz
UdtEZwapHfwqhGnXqFWIgLsc+yvcIVObNN/HTIt33GmR9YftBrmnGn8eS8yZyiRGmSZG8qhgkJCU
pxqBrX38VbK3CVH0ht1gSxX5jSqg05+Vz9wxmQmYHsJTJONcFHqcZfu8BwrRjd50Pf6IlvJ8olFU
dgIcQ2tA35L+0096N681NOVm5VyjCWmT+oSL+QJ3RkAmndzC3O8AAhop2BXPv+77w0zUppC7H9tB
5xqp/mUKRbKLNHRKnNh0Uj2rR+SofIbGJ9IQN2ubLl2IVBedDBJ79+NikQ34cwTseZYGaZLsn+wV
QcKTj8VwFocTCbdlaR7v7YAKxIBwWoktBRwZPrrcXo1vhLA8Mp4ynQMv1U8Rzmyj8A3G5TqURAHr
ExhRLT/Hysne4MRp75KcZjOwle0XQ+ULNFmL0KI5uSoSRUfg9JFiSp2wl39HZaDhUtqVRuwel2WA
ylxyvBws/CV/Autu2HEjmsX3G1A7c3s4B11p6N7RMl+a3RgeSmJmpwRq+cdTs8AZgFodXNm6CFXp
1n9eRFyE/hbUXNhhWdZhZPB4HimcKOwb8hLym1vJTm6qDef5AjoRKQW6UoYt6k/5DYGLENGceDtq
O4iconBnwf7jwAhXdp+A+VX5w/3O2u8N3tI5zE9HtHnOrtpLx601MKNT/5riFIqiuOyW0JB28D5q
K52KVJiUOELrMPX2rnKit/uGSyLKgPoPho2p7n242b+SLwLRUHWa/kaVyEfdW3Yqu4Xh7nIlFbfJ
+YnfC3UvV0hbjo327T6VUPWGDNVcA5eIQ/KqxjgXnLvR4m1J2WB8tvRbQIITJLgcPvgzHGSpleM8
nuxc6S2Gg6xYAPTJif9shmbw/EBxZA4qYsZoqDyAJ0RH5ETQHLDnepiItjkuMR4sCBBGLr8VtBH7
iR3NWFqfVmsY7T2I97dABotkXhutMOdUCkUGGnQfnFmQdtV3RvQhiCyn05cWj1r3tbRXLzjBqFN1
97vEINL6KdXV4D0MdlqrwFUNGi1cJnByj9i0kwvB/LXkCVLlvCe45/2gi1ua/jZ7WlxlYVzw4V7Q
/z7abQO3lw6+Ix0boOvx3ecDYFD8+1wm2hmRz4HX7kAlSWwRI0n73tSKzfpNqZzDNAK88lTBeNke
JyDdZk1DmBWv0xbNzdnishFnSUX9k2lPdq3/4lq5cAjydyJ0caqEb5WckLlgDq3MjCsliI24Jey5
6Q7iaZ0ucP8+vuDJYLYVCUxzzy7EbmpoYQVv0/7hTwuhY5LZa8cVqyvNCqnzf/tfXtk6jCZZ7xBY
09h9UP9XQ1p2H8yGlCO1+foGkJudq6IQ6qDwsOoUkgQziUJUVLxNmeN7YaJqW3VciRWNl/BITDKZ
MHD6DZqX5M55acO4v4Oe1tkR4ep189tv6w2fWln/6nWS5uYEGvDVmIlbiwInu6IGKq05Iyhvicr+
eBPK+j5GNyd1E6vjWNS+o33NvCpe6SoBZRD+2pxfgh/NkAXu41ODGExNABqO6TOaAL5XU5e6SkxR
2QHyCvhKu4uPCTYgY7oESg5bpcp7zAvenQ4tJCE03yvStDUb38OMtEzxWql16slRyiExzBYwW9kr
+9CzyoZKLhVkCkZ07OmL2nNxxZe6zXOw31i70vnWqSz8KcEhYUFpU5TDON7qaFTQhQXJdvfPMj4W
84uWLYHsY3IUxGtc2gqKGJ6Wvttr5Il+Gr4YNL0MkFzz92qfrec2JxjNDlZ0Sv+Hok/VPTnomZuG
QZRzAb+L3vJmut+Y92owBJycCFYm6a3owhpz2OS5c822cjpbfUWRgVWhrpUdmWRykQZHIuSQ9GMn
Ao5VWTT+KtyJzUbgjS8rl38kCcCDrZfUoXygkOgtFFfHLSAKVmnuGeoaoG3yMi2O+N6LPBcrsdN7
jPLtE/u2spIq0EGzBPQoqZMWsp5I0vkaBahXd7uH3pQbRIB7l+fPA1TWbXjB65M6M0LehX1BTNQd
dX9ciD6uHjfN9ublNmdRlNHUgDuf7MES0PCNk7tF21N5WoEOk60xIap/8oMf+1+ad4O6SzVkq9hN
bw9hYZPlFNQQR57NQsYLuUClhU3BHNrDkADXn8bCiNSdF4ryvjxUOqdGCt0sEUrsHX9zqsX9+EsR
zX4gVvPdOiGrzz/MSdTGM58cqxvT1gGskkxdQoZ6sgZBbXkmUQXBABF7Ofym2jmV7osR8Ck1KYnS
XKvTiHNCZiSbF8aRZVZFGk2c3+z0Tb+zZ6NyfpKiLc/EihJJtCNvL1LUZhCsKmLUZG05ylNq+BGR
NEW0cTy8MVstaFKYvOfJNmnvCiNqpBG9Mo+NPWzGDvxuBQNHuYyAxev5896SgYsKrq4a8h9Bh4z2
p/vE+FWKOrXY9xjVzrsZOX+wj011KunV46SookCJExKVCFpwbF+CVu5bfMcf4dLFeEArw4/vp7qx
erP4wIHwYpeYZuhm7ferAeKp0kaVWAj/UWDGNLkCSF2v5SuJpjLGaMct85CuewihGgGmKsvzX7Le
rr8vpKZY4i8CdEG7jHQVzT4FbD1vvZEgZaOKtvKbRbU8cLrzVaxzvl0v0ahuVLHH/bzUy9m3UOlL
HgnRdy6XF6JmurtlT/vP4ocQVo1ViqB2ICW6TeMi4TLhTs+/cckr7S+xXGV9b4hwSh3KhoVxA8Gq
pNSIMyOl7dbmAmpzt8dO4U/6hM+2Wag3BqMARoCxbWBg+usBiUfYeDDWkzFw472lDmzlF3Ype6jv
iop+26z6ypCYJtNP/m+z+rBRY1b8Owf1l99JHJBKqwfBkMUfQFVfCFgkVSQlIMa7jkPWuCav0PjL
HIZ6ZG4TgHPFKQ1Gr1fcel98Jpu9wEbMS3ma/X83qY9n7dnmDz9uV84uXVhmB4Fe3Ucu+1csKuoZ
zHQeZwxmHc9HPf/aOyi1eMhtu5+pDrwl0ku6bmR0TCSXmvbKDLfrkHCTpMAq+jBpW6BvndGoGMjz
e5YfgJVCPALK4LIkOQ+9MSIiXUlKNfa8+AyxAYn5EvDND5h5cm2rR7N7z+1Mf/PaIM6QIt+bDbKg
iaXfgbywjNOQxvfqwZpllwlsLvv01ih0rVfQw7CRvDjizxkR6bl9T/qb0U7uUE6TZlzk6MRI1vvI
xjAcDfeKY62FhK2DINm4Xbj0b0pyQgDQWaa6prvNQlkXaKXBqd5TNyeHnwe9u1tk3cDWMCV3b9rm
s1/jfBG3qnv6I+lgONlhaE2xYV63VVwsB0CGtoLfc3xbQce62gcfXZQShLtKVJzjI3jf7YvlF7OS
KkdW+A/6HEfxRJaLNbCbiUINrAq1vKSWUTZjKTLxd2V89IyKdUB8Pz10ERP98dV27ExTuHP9dFkJ
V8/d+qDTiqVEzvbXHMn6+XvuGf2UUan3SyOuKBD53lhP4h7ikyfy351cQaLeWnhgiXmo7lqUomdV
hvTY7dk9OFz6vNVqKMhhyFELKWIVena2HecKzlujTO3w7OKj3/z6H2jtGwGaDEba8iDoA1AvpvRf
AhJjDO9lPFn87UMlDCH8Ogg0pigIPfqICQwF/JoJPQBr/gZHUKrskblMZioXY62fbTG/ajNWvaJ8
wsq5ZFk/N43t9TgRgpObCUi1BnOPlEXwxJ/3gYfyyE0BZ0S5Cp3qh3SCUka48gSJCMglGXgX6waV
IIBmHz/IivkfXQacxP5UW7hpKiTt40UhrDZRKD2Vofb09GnMcCzYzEgMUnmaysqmC9rg/nzryCCa
6DVW3WlxF38emvTVvKjMqkDD5AJDF7WotoUMjgO8fnt+Hpl0omN+keqpjpKVPqUyqKZzQ0XkkdEt
0T+GeubAS6/o5Oe8KJyTbIXNgOysMmDDsZaRNc+YPRWlMZqTLAl+JYqn/zZPZag2vQvSqM/5K+I8
8ESl+QpEbWcJUd8KhtI/hA43J8/T5n6PW/KFu9rEk+FmZTevetn8mcmt4ZR9X57AWqUIdaoujxDI
Bnxr+gW04hqxG8C3oj+WrlPulocPdcImizqs9AwIHZl+Rc/cgXHnqBMntiAnKkhw8gNM/KZVqY2w
2i3gKGMiYH+oR0h99G3UnIfNTGp5uLlKRhnw3vET/ne5f4vBS8zVdHthCgX9NZMahjienpsxfyqO
7VcZKVWgCX+WoLiU9mvoCL4+pJ+A0Sq1nKm5IXuE5jnc4w8dLi3ff7oROfCJWW4tessdsr7eRSAy
VUUh1K3K6U/SAbDYildbbrDRrbhaLMPFmHFJzKxJxrmvl50WIRtWYc/XOp74TqMxy3QTVEbfcjLI
ksOtJd+yamFP48vqZwEtrz2FkhABksR+wc+fzo69m8VAkGYRCe5SMzQmgfHueP4fxq935yY2HhR2
M99Tfd1VwNHHbDDFKXQeDt/al8Zmd9qED2kQXOw57yUdvuOIdJ8enRRmTTMhzABNjmnR6bBJZrGA
pQdVV/kN8CPx/DEaBquEHqJpED1stk341ZIoqtwurNLNgnIHRgGqUddqTd0F+XTE56sRDNEy2KeJ
OqtIkZZZcyFP0w1fFckIe5n/34/ilbjyVVMMyeCiH6DLRId2SDXF9tNi/pCUFGolPCUxGXGXAJBI
N0ZhMr3uap/DotXubOcmTk6FbTHd+LiaJDgYwyI5AfVvYIrLsvp38LmhxPBy+NVpWcp8hMFWGITx
xJfEP/lTocpMMvu5OXiHQAQXbigLDnVi2BXiWhqTIUdjozi1/OvCpzLgzRgsjB5CeewsZnpwpfXF
1u3nZrCrRZsFs0qEu6wLyybHPFODLQodnnX90HufURDsVY5N+Kmj4c12nSLfKAGSbm81tLnD9Y+l
8i3gzoP4wHbOJ4JzFkfEQOe7zIw3Ez79jy0tIqKFJF9BFHZmpQJ5wgApxthvfGoFsd3zgPzT/ELN
uX4pgEDn0gYdihookvv+EOgJbPXlKNORNScsHS/bW0r/wZSZaa3Ci4No5KZOgvROf51YBj5uyKdt
4suWkGiQabeupgRGkyIJvK4gAISRjwGbx8fnLNDSG89bvmt4CBq+fIsP21X562PjbkjxY/QD2h2m
bwmLzRvF5vzr1opXFDbQSOvnllNuNAs6Qo/MozV998oRs/CEhRgGWQ0xcgEwcbMxJSCzVPrOb5Lu
voqFLwG66VEP7IyEI0aQOJZbg09IY5eyczb4J+NL5KOVQ6Q/rvuGrUKPgEUX/fMnHW0ozJ6GkgVB
ShqfYW/Cy8pGiD87T/krCLqxyoif5/jdV13p4FMGtQ5E+CJj/sKqYOvnk1CkIDIXhD859ItxKx+Q
f98sKpeSFQkqYTD1rc6en0rmG+EWPZy7uZuEMe+XbvE5skasZ3KUz/80mI+tnQo6s+9MFEH4e/eO
KKuoWNigsmS7w1tI55VyLT0uOCvuFWrbWXcV2IfZtld6yZbJQIe5UC64k6WxX6M+PFUrYFHbd7d7
XLqgtkFIIhnATiMEskzW3y+QGqmeZk58RG8O24pM05O2lKwjXRTaBSwGTx8BTib4VzC0Xl5GmAJx
0+QpHZDej8hRiyVUjT4lALlDmjmwa+uWApv9lpV1WBjfFkHTzn4SY0b7ac+LRuTBwrJvMiKxiJRr
Z+fPi9OnS9sQ64NVKxmKr5uibetoeYY03mye+WXNcDXQ3cspyO/c7NlcG7ag98Q1Xs7yc1SDPpx0
UQRMlwnU34kom7+/AAH4DJU4bjjGHBecYZktJnMxPjnuCLg4sDQUR5E+CsnquKRhgoqNjgYvlc20
15j+TOnd/BzO2uqLWzhd+ZDazMv6xoeYXcjS3whLaOudlPke0zSa6gsIaALTwkAO0csTOna6e8MI
42zM7O9nSwd5CnNXvTjE2i80TR+8guaUSP6vTvOoOjsT8cQayl0TvapYHUSttLNICAzxj14Wimwx
7fxwAD1RQT50pYI8AN1OAohNZ3rUGZbfRgIG6mxYjPrUaJdhk0Nm8t+RjN/mAe+41jeg1TbzIALo
kBUgHGrosqz0FDPuY6h0oPWJmI+ZODc7xiN59/JdLlagOVLDdj/F+/+7ICjIAoQWrBji3pwlixkC
4NA5gwOEgw9DxKSVPDchNFVhLRc0AN7P5w9QJ2hKkCjKsbbrjlufj1oESMKZJPRh8hHb84vjBFgJ
l4R9NIur4N7XJfr9HtMhMvPwXzcLkpQHQMriztSNMWZPjgm7k4fBvkXi0dpzY0s2OsiUBZRHx0ep
3ACtiJ9Q2JCGtR2e5D9wxWxZxj0RFYTZqgoNPvdHMw3Vyml5RxvYPxoyELIqtK7ENj8Rrg6T37zy
kVV/iZXgUoSpJxrutNFowqKl45mA9xDBahoeEt/VgcOidFaLiBCouKSO+8Eo6Ap6Dn6NPZtGAjRj
aXsk4gbG7T2GPFiLud8p5YaYOM/WddO4wRLh4MR64WAHjvH56j+eSswCPuybAjh37C9eiZ4aiusN
19+qxUbOiNm8Az1+3uk4Cedjqjz7d6r4qRqwSe26HUm3OEy4MyqlhaKG7C7cELE9CGpiq5EiMgYL
XnuCK/Sk4NQHyezOJd9hmssLl9M0KVCrOTqEiDdN7GI0B/LGQ3vlqam1gIxPAAGti8w3EEiV/vIa
bVcZdTueySSzzbPCnWVWjvKCq49QLMjMT2fljJNPotoctRtVFqsToJCs+p3r4ejgIN+cRK6NqQts
81QWYHEYB6FFjwNAfCpuwStYfKScCxU255UL6JE1yOJZf0SpCQ9542/xXnQQRpRVpmad8BPTbLNY
TinWof8+4kqGUlKY2tLesxwJwBKzLt4EraLFm7bu8I8IP0EWR3o1wIQBM3JOvOulYLCbRvkkP6EW
/NPvMGLlr/joE1f9QGsfAkj/1cESih0wVyV/vrXei7Ew2eE0zdYJMhtvdsoFr2eMMzQ3jpkBQVWz
WVbvBJseks2kYVEe0Fg6yI6yj6YIFVcsnhAQIjJ5xbzzAVNc9tAOlR/9ixus0tq2WI1EML7ec0xT
lxte0Tx4HlCDKbvSnYpfsyaS86AReRicAedb8LqXmh8647ehdBSonr9Fox1BYY5VgdZ+tvfT3pz1
sejhetvWZvLiKs20yO5vXsp0N1yyiHxz+7MU4KSppmwsDsZjqaMdMsshbTgGnwuV+Y8xz4QocHd2
FyF2+dv3pHe2m8KaCvsD4aI8/WFgAaohfVa96bLj7J5538Cczg8lkF3rNUkW3J/fNYbDWYOJ0Hjt
YY6jAnKCXC7xZZs1Tb43qZWfVdfHC5WIx8irFHsY7SSvChpQaviE83pDZZ56q+uqnnrF1LzSDIH6
IJWtJDm5om/3Q83BBIAS9klInfYbuSAB8pPiFl0iT1R8+RCcrv97hKV2J2+cXXP3kUG1Fgvh4XYo
FSlqqaAWqHCRtpQW//HNxz8GOiJcS4fpviE5XQVPeOVe8Tf69k1loEXhE6bfrPFXL5O5DhyghD1s
1lrVcwZZyTf+9RRsNIlN7LXhF/s40cDOR8Tnf6eLFY5/Sd7QZ4nBIPk2susmMaLjnyPzxrDQ+7Sn
OouTWg6pDryJ6jDsr4ariXeR+CRa14ws0MX8D/toMGL32ICd+ox50kNJCorJ7j1KGwrbAkegtjlP
mKS4O6VfTajnVKKJNTkk+4rEWjfeO+i+Vezj5W765xm8aYaF+4Vmt2iZvUT4BS2qZ9vPhbNVk9Ra
adJC0Oq1ak7neMjSAOTE566UAMDM0E1wIHtXBf64/TlYbOl/9PXIkss4IuTzDrHgpMJ1B2kWwVbF
uvVDyH8d34Lb4CGIe2oxKmnWrCiOxSU0yB2YZIQVWjTLu1JNqhUKPIQ3Kv60hnnA4JPRAaLF88Xk
0YH7wKlmSe9GCujJrY9KDZ9E5747PBRj7/YTZX6lvUIMm6dRx78L+Gy4p9I5RtnLKsSCTZ2GzWgQ
+Irr+9w1T5DaotNFLz/LdIltz25Za4v+eLdvmk2l8bPCe8UCTOYEWI1u6PLtZzWW3FT0RtTLXR/F
tZxgkUmd3j4MsUx+hMEk8GS5lV6+/crBShWMW35ddtrlZDXRYxfWfkKcRl0N/+CdrXOaKCEyEsl5
ayU3EFY+ycVERnGQ26GUlRKP5Jw5cYciYRqsSBuY1Pnbx4m3xbPPiLOtEt1GfHYNk9gAfpzJ6L6b
gEeFd4kNsaDLF5aYUu+awA0+KFmSLjUVd22F72ErXZ0MWkO98c+PTuw31qbzReWZM+5eslVirKqn
Q1wFyhEWOO4EByP21lsGb9B6JDChNOms9xYM5245mGvQlVnhaLx3zM83a+c/V1B0NZrWntnF30E3
wIktC79HSbUOBg+kuIN9+OtIxuLrcqYEBjz61tAaQqDARN94EPbGRdNoA4jkfm08aTPwroEGJpGS
A5yqyPvIEDQbOsNr3kjA0LHZOkL1bVR3Yhic0zpU5B6pxMZjzSGYvfjFJBe4afQl+kf6uAcB/+nj
y7dOKCnTYwySV0zk96ZbGhkZsSDLsXdcl+7nmeMGbLaZvxdVq+4t7Iu+flzWG9S1lRECPQ3THiCI
wnSr0gLfetSy89D8ptiH+G9KOJjr0YGVlUNDmLmqi4NlfQgBmlSWWwTGxOyvVzoOCFYNDLCO1qhj
UuKdfn4WuVyNC/w69wNgVc/bWBHsuyV0BzYiSvcEvESXdD0/jQdZlzcfsGC+B0REKrM3EGTcUqT3
etEGLBCrjUdny5PoaCPVnrGYcTO1mT7vYlejkR9UMPmRPPmSH8hgvPQuxp6ekuSK6RCUX7AF44LA
IIvBxq5lXzcJ6xCe+syOljnX23z45OKJaCT5Inhrdh+qq6HH9b7oBFzbzZo5g9Bp4tsIMlaA1IHK
zsGXwe58jsSP8i9JFABjDKSE6HIjt5Tp8/UMoAPOF5ebs1ydEi9+/juQLtlH0LGGyz/hOQltGuaq
tSpkzyPNZ2ZJE05DoghLV3LcR5voXXyCY/PN53ylgoGPTMAAuABbTsXD4CSESe1Izyfjo4ZvUJNe
7OMV8daIJ8aYzBPpSGjNPke+o/iiWNmPQyIJU630PL51ElYGNWY659AT0H8BnAHYqBGu9R8FbC6w
MD5srCa5YchPfUckvsy6D4z4xxeZCg3IPkjS9spQz55eh3vUMklsl+ahlf2JttQ1+iLBM2fo6tAE
4DarSmOeg85uhbbCULMuyQARmt4MPQy3dHrGlQLSpTDBsYdDjfLC6BqEqkUEdbsrkemd8QVg6UKF
WG1odC+6GrXXFYxfLo8TEL03zl5TZa1wBPc8hNuDS/mTFVj6bz5HCDmjVucdMzKUjEAuiZyNOnoz
2caxTQj40O5TggCGcxb4YYhuy/7BQ5NPj1FsWWySlUK/PeTRpAYhaZc6FoVJ7IMIPt5Ee7XOrxu7
1WYK3hkGDga4T9f5+tKKSRcKEIF6V+7fY3oPqTAj4RCI2DN6zRRMynIp/WIFJ0/xATiJ3iN4OkO2
BYaajT+wHTRk+tTmbfeQBV/14X5henYvlyuZ3OQSG3TQGB1EQhm1VTP633MoLDVMOUFe7mFImSEy
wvCSFP0iX69pig9hLPtXwTywD59WEVzOCeuqEa9W2Hd5Q+r0ppHFfmXB+IQOOMzRMq+qBUxi7wrM
Fa2V3m4GNNXuFVXsjzUeYLJk/X4dJFnaRzVNVXFNgAqD56TDijCqafNrJavqaFdHx4Smq0OKgDHI
6FWVgl5Dhi9PajH1kj3Bgc0E9gu2fj3ZO7djqkf5kIUyQAHgdVEATpdOcCkcEl4JeNc5AsnZQY1e
tNFDunK0+3/hybtl7e6vOi4k/tga3wx77wIQCAEtyVZpIfDbIJTJVsmM6SKs6RH3NvO653iNiXMu
9ke/BzTRbvVnYH3QeHxi7kFNx0uoIEIAFUM7TwqhL4rIHEGcu/a0fiZn143y+vAsPYYN0bz1Hw7+
HjCbuehmd2mpFwr1i9OgufR2F1hcO+5meMXVgCFyLLDv+tYhyjS1Ia0NaFX0MxeDZKY6DGyWMm5z
zRhJr9pmoss3xI+3yWwD2Am1gb3jH+ZoJbR4H8m0KzMfJH2AYZoscPrFHChFibl2LV78Rcd2e/oP
E195+x4ZC9p42V3fyOSpR78IF4A02DdT0k1qK2EycZfADxCUOJwerHv4a+GWaJQv/bUNijptTTJl
hCH0Ji+yp5HF+OpxLoCK0f70+2hT5pksIvps7QZEbi+ek5L27BIbx1kqHEAEhhYfnZWh8DZYeYPP
jFBdVgVMPt9Dk7aLvAUTY7FIlu3GtoBA4w9Us02h9ohdyOwGrMPdzUY6Ki6L3rhE4269t6k/XbLu
GB1IcsA+4MjIsTqJO8Hgo6y33SrD2Sz8Rxqn6AU2o8jXMAZzSXcu+eZNdnCQKQCX7xis2GbcXm3x
k4IwQTd0ZaNOiWxvibYaO2dz393ag2j7E6ralBLC1MnyjeITcXN1Ir6OAI4bbN2sK2hyZmBPtBfe
DsDx8ddjpp6l1XByKH6VNlbTlIv0zeCPoeUfkAWiGJUxHF/Jh+VqIjwUxzb7rr0reJVQvsPpbWRO
NCwbJAPB+VjlxYib4y8gwpML/W1r5gQBUpXr7Ao8MKT3xRb8Flg0ml10xoUwfLI24UhfgJYi1G7w
6IwBo40wH4/f8KWRAa5PEsHWKhbsKiW1vh16bBwprxiEy4dz1KBGsAKEwKgo/7x2I8sD387jIAtU
72EsFUuKr62ZcY97nhhy4gBGiTIuPUETEXLSTDboa5uN1FSzufW1iizVrt/27T6NgNTE4jtraJNT
lKO5xAFZ0x1u0DOVvVSdymAsNOc4Pyn2v8p1nD5p9tj/V5uVp4WOAnnC/jYxX64BVbSMlGEWGzvm
6pjscNtMfz+SI5INLlRm/O3oTACwzP4iujPoWt/APp669QiJZHTfYlXxxfwgZDMBVrWcNZrC4RAW
WXc7DCKjekfHZXJpWysxWtxVr/+MndO8FCYYesu7FjFJo69MU/AFlZEf0BO639ESFXrtsS+PBAKa
Rnjq/AKuxhpi0w5I3QF1mS41YH9UIcT3rAcvWw4EneaT6wsbfvAM4KxBSTMibV7MM4XJjCGR0KTL
zVkjEkW/vKuv1rNLIqmnVyRbhaw2iqM5KqSg/NYnFk7rJCKgdAKcwEQ+HS88eABV0q4XF6B8thfK
h/JbVW1E0VwDJs785PwxSCdn2OBI4uWD+24j/ti6oYKVE1IT8PMcHLIGjjn03L/QfjLqfkI6BQVe
21tQLcN2Trho6P0djlpmWFs7UZ6CP3oAIv6kcaryD3RkNjuG5JKe2As/b3J0HJ/Bgo9UvpG3UtRY
6gJqwCyh4kmoaEsx1ovWf5Bv4BwXWiP9OlVEg6fJc0n6qg0j3C9jJJtcNQKITRCpxjAPJ3ksajI6
NR0QtQFB+Wo3R5xrwUr5AsB3kf7YCs/6r29aaLIhd0pS30CMAY2Wle1SW8dU24ndm5QTCItTrYiQ
9Cb9pjYXSQJAHzXIZTvl6QPdLH6Li8FOw8/ai7cB8IwoT9E0B6b1NdIvUad87wKMSk47pKMc7dQ2
SA0Hk/KFS9VCo/eLM6ipai9MuJjAH484IM9TBP7+Mh6xqctjzN8+iBATyWTI4HJFXAZYyqeTZzMt
KDyl0wqE6MLRg9X73I0CZH3yXzLTDh8OfpLA1OyDRheUvk3pzA7xdIUco3Hn+n/qiXxM5lA4cLQ1
5GVECQkNHUvABpLDRZJNQVxIv4ijaMeytW+CoxaH5II5i5uiH2za2cfFboZY+z5qfWGD7EZNXYbr
TMJelUFKFtdvmOmLjlORdjLknM656fWQmdjImIj7A1Xt8Kria5/PLtbrdQz5zlZBVFUJEkAqPwmo
5oB6efEWXRiBadiZcM/dx3EcFruRkQcXuLH913XVOsOAwmlEyCk1YnAr9gS6+GQP3u8aFG5HBer7
5aWW6PrLVcWAwcfhz2GatBMtDZKPX5WTN1jOlW/tuDfNx7bscm5NSk+SIBWvcxA0zHuD0TLI9xpf
w/sCj0M7Pbzo+7hzIrDfBeIWTfYr2/bCqAj6P8mImiu4wjLbw8n5BDl4QP9i+Sgf3IxnLdmQqF5B
tAEAJ4+z638/Xc9cugF/qpq1ebYLl2S6KHhrZpnGaplhN+PgrzbSLARqk/aBnPJ7TERmjHN3ZkC9
LwhgMkBqKq28BIQEXkHuYWFWTu4dDxYAvo4XaH6knEzfC4/4JT+Nmyi1p1MftR9xefk62GCLiAqE
due33a9De8CzQhGiuYnGhjBlzvbJdB7Ij8s3jSz7LOFP3XTuUnTbyqpzW7e8NX/qbGmMy6fHQZgu
3dxZc9eKh/Z/cBoiz6+514nSivw2DyJJJsGEgdn78K442ehu/0jkxQCmk/kedC0iGFPyYRqvhYAy
ODKMY76l5ro3pQJvdn/tqXKfMsGLLXGS3wtoLV9P49mY5rX0moiEsxdWrMcTPqJPP4PWFyaiRDD5
5/7fVXx2JIiTfac7iYxKQnIRo7Ce1oDdbTVBDZqmG4UYBkNz19KFOm4u8Glh47kfDEH6PtR7lT5/
ozAMuMo53LZ5hBByxQ+/61BisRjTlCVSpI4yIDUT7ogept/xWw6bl5msVmAi7Dk61lDtcQ6jGNn/
9U9HyJs5XgRTYtRHpT0sVzIqPVuMvBzoRokMprrOrsjlQkMvTn70PAaggTG3nTSxDtYKwJZQeAnA
exZD+10AQkhrPhFTU+RtJYsHkjChF89jNorGAVWwCvICfx9jAmE4eVb9N8L1IHBpPu/abaZxNN3v
gCQ2gCd8mOdDPI05L5Pq7peepueOC64Tu6MfH/6+KL70vJ7uZnAOA15bbfnYR4DEAjWXRPa/2aRL
dtHKBOdiK0F1bm6PG9WAWNV3YOHlp/V3iPbgpNi/wvXyRdpd55HkhdoLMbJNaKjdDif1Fjght1dz
6S9xJZnEqjNZZ/f1tXWBkw++S+YMTLkhYIXsiEmOBI5+cGfxz0NY3rL3GaLPFBsvvL+t4ECB/Ozh
NlM/rqXQkqcMmPjphBxz/XLgPdEouOyw3qP/Mc6olDvtjW52pIm8yedQZwksQ01TCDgK7pNyHRd+
fGC0J4fonaf9VrV/W+h0W5j7xv6Y7zaY57Y9FJ9Wr8llGSAcyiuYDO/yXekzRH1y9YqUeU9K84IF
bUqlhoOJihPH39KJpUajDmgI5n9LTLVSRRIIcWA92MF/L9lAJ6KBv2OgIckDLV35Cqg1TKadfElH
pLQ06GllIsNmEYC7fMHu9uyQL0kLZY0NYVObB7A2ZJiin/0lTMZRsN6EivVQHTyihNDJjNnHkDps
Bjx3yEPBps2cLpR9MMCsHRPArEj4I5jzAV6FAWrmdXom7yR39Fo/Ri6WwqPS2KoqIB9zh83j2Ask
/i68Ik171ascdluzaImQm2wFxijP50yEl9fcgCaT8brNEXvHgAkvnPBBRapufxKAJluOpEYgVms3
WsWdK9vw8Y3PQzOc64neidGxirtwYJEqCFCtQcpbHwbJkEdEiN2tR4pbrBDvLqLqP3iLHoqag4C2
wPoQleeIin8yHjAR9uiW4O7Mh5AMNrL98RjWhY0/Wp7Bn5fDthiDPztQzswWsh+wNrbzLKHslRTt
9JaQ2YuRptmdJk9UBYS7IaKZOCw7EesbeG8LFpGZAb5G+e156yVylNLUl5hIOZMIFLGvJgi7t/Ys
NGaXh0D2frnxDKPoErNfQ58RnOsJuEroW83d/lckdGcpOqXs+ebMnJppabKSHvwiH8eN71BDAgPK
nBmp7KLkQ4Fsmh0mP+pYeErIzRretQPYVana9Bme0In4PCrxXD57PYajQGB5tvEG9M9ROHHOYgF0
0AikRJdJUuuqsJUkAtj3hDIKJbXbz3sZ0HP0twdIXTq9vkkf8wCMvx1vOZUK+LaR100Y1P1yymqv
VyPSsGlL+P3VnvVM8K3531Z0Ij1LoI5L86eGPhObrDoWoc9x5jCG3IxECsM18s8kWYDc8KEmghPU
VOOhBAkhwriV6jDjP4Js/Sj7aWzf5SguufloNYmupMvhNH8Ct4LEB6k3ULJ3alBtiyqnfKZZZOQ3
nbX+Try5NrWkc2+1pUY9LNPjqKfpqwm1SFDiNzy8cBC7uJZ9OSAlpECWJ9PS/8Xl1d1QzxHpuvIn
kRnqqxX3fSH5jUVverpMJQ6g/OpBQEyccEtH2dyT8Rusu8PmodioHSvpzb38IcAvfBscFcQFT+ph
NnY2XQblxqZXYl9netGszpWQTw7dI0UZ5ns2TOVPjBF+wXmDSm98vnBciMGm6tL6BKeC+qUvXTsC
PBabN74fUnUc2A/o5nBBWIXF7HHemY6/zIvkZHdmfq01xCUQQH9K2YQ6i6EMEev8Dm2evoykjBDx
TRaKWLrcBaAae+MN2c5S4cYcWUGqv9nOi5WVX1IAmntILq2bw8oG1Lp0CH7SFo+ZYpbpPxoO912a
WKQz+2vPT1Qy6I4HqFWAYdlb0uV86dpDhw/xk0DvOrYhtnMlIRdI/I0pe+OhDXYBG7t2aORZi2F5
PbZXQxEwxvS8+3NUGwwv6xy4wtsQRx3QEVFcyvEFKIL/I8JWaQwcOvQ475jen6iBy/GtQlUKX5Nx
CcI8g4HjwHSihrJXtw9VBKby7+TKQ4O7r1cxYjenPhN64l4neHtQZd5+srqGStpUTnp2MzAK0oXp
/VNynPgyefjyz6ZFG1ZFIVm+ct4JJoOu0I5LOeJrgtnJIWm3QyJxG7aH3QX+DO79pCDHOXaVxEuC
CKqrQinf3KxS8Hv5pAfJDfd48PGnLppV2H4sPRyeqa+c3OLNuiA0a1k9MQBR4/7GgiUpru7vFTae
A3e22mlHWoQv/cQEQ0QTQ5B65prcHmD+AoMzocgkoeO8M2u8UC7mL9qr/gwruPfqSmF2j2OK/zTl
kUTZkXLeQArOz7dO2Vdd5LPLrSDLsuesCcXcOs7m0wswkggNYdUMb4ZIbz3/wUHvdmt2A9TLhcGy
tcrGfDRv/Zg/X1joPepO2yG7xWFi7rnFo/BOS4FoVt6KZ8afboU2MYW1NGB2y9aA9c1jNhnXEE3u
1x+n8tWyGRgL5hbzqW+pKPYVTP019sVK3M5lasmgnCWs0I3oz4cHLLPwruwv1zWb1JYTZYzf0fEQ
3rELSail1Zq9OTLOAp54tGNgDTuPiATj9B3FYXDwLv8lmfF7DClppRGcZs3cJWwjqYyJwv9eYRV0
38YyRk9FVfvIyN3V5VNoC+PHFiM0sOVUzwlPNLTRhE/0cWw29iEf+DbrpRkeV79KWeC9I5rCxy/F
x2N/ojCC2HCxRtKgqUmk2dxWh6YkpnPQTPjPCydUzxLj9Q3RxqAS1CvOnppNspzA9eQ1eONDI08L
fFcm4+mDBJfPjwA6AuZwYYEUF/yNI4TOe4EgI1yfe3jJ9iRJ1Os6nMz4VlX6u/dvIrz7KlUawwSC
zle2vvsFWF2Ts9/ur3tNqRpyUab0GsLg46/cFWowFCQroWmiMJjTPHNdyh69gQTOW3QqYlWMUFYP
KQaGqiV8i8e3x+HQuzT47uK/Q7mtfNMbgeGw9PTdhPGgAmJ7spwTpZjtIbAGlE1TGKG5rVAnbvFr
Q/F3+ViX5hCVwSyZOgW7bPEudQN8jBnPXsEB2B/gLIJbrDnYigvHcVupeUG80Mbj/injOWMWioDL
3ZZOBYFITn3Su77jMhbW85cnUjQ39H3iuya8+knooxFt2kedvHxzjDVW78OTmNdkbaFgRMwWBsXR
P0Ayt3pyxZIAsuTMt2xRlhu0dLH14xydUDTmY1y74sCeucPu2MO6eflxS+Cv6z4D5qPGJDoPv40Q
OUJ70fuRp49ZWBZ7e6NewC34mGsi0nEwkMLEsHwdT030C4kkzskYwoUFsEVWtRABXzX/fYdjgXZK
pcZOwxSKOzzP6Wlk8KEL1qrpGYl4wvZ6TsJcVXZrf7letNgGpeDaAavmv4GxScc79bdqCALki2j9
2rwxj2KmUTeG+/wWirZpy6d+nRtsuLQUytWXTd0oswS2px8fgV8CLP6P/NzcP4Q4kCg2pBp5Yj4w
rORoclrlpZvs7XF113HT4BI5dsCw+L/YbYdigJvm4GxhhUu8hRk9g9p5rreHXcevWRAF68Uc7IQy
uuIM8Q1Gok6kytGF+cikrGfJ0MLTGp2xl5uY2HN3mUAY6USqjq3+ToJZAAWBov20jNCY8Ht8oIDZ
kTAERoED9rOwzEtFQF67JhJ20ZSXMyTfyfY5IXbh1Nz0ljuAX6OanFnBYQyHGxmNmeizZSym7xF1
/Vza7Ji1Up1b0aUg13O9N0aDpbb1CvFm7DpoDHTbU4a0++ZHbw9N+TVBLKma46Ev2PfS5IBBfq6I
sXmrIO6t0UQoyxgyaF6jgJdyaoAfHV2DjKDtsHaXrxgw6a9fjKlVv8ljYmV92jadXr/Ir2bbxVn3
hPaTfwXnjjKiGF+Qo49OR6rwzbeIjvIYrlMBut+EuV3PxQDK6UGgTC5hx5uBaViA2MZoGDzSHcnT
hDargVuycBWsxwCl3Vk4XqlQwUKhTdZHJupjjZGMKRv2v655WGzXuuYckSlVZLQUf9RpV06HkDjU
eFuAoN5QEBZr7Bhx4HW+dhqmUG/Iiz28XnRFk85DQl9YfVdQpd48oXFnZ82uNqhNKDatk+ZfVLyX
RZLccqfvHNH4qIf96L4fo28+6ak4MZnG6PJ178Uy1uARyWjqnpBgjStN8Ly7OemSHM+hOUfnr/o3
Cie8vyjxDiLn9EDfJkhpI5zhgVDbp9IBLVHFTbF4jwoVQE/nPOMzUvP/gIZmj8oLCm9lJPMbn8DJ
42Xd1WMg0M8rnlndoQv059V/v7BymjuZ1hKjNs3/LntvZmdwR6WJk6KO87NzWicUPn7cm/fW49Pj
XThM7f/0gZti97KrsXpxDCMg/P3irYuacylKjMcudCgTPklkAug5rE5gioWkTg923xfsLW7BrMUg
38VCxUpJnoa1KtlTMH353XYIKyk+XKstBXuzeJ1UW6EG7WdV5qnZFvHczn/3WIN1Tgic54Ba5bsT
XOYwy533o5YcuACnrR/9JfSP9oLF99ufnEKr+ALRRWbappioe2vvetotGwOrjrLstV9vOWYxXJlp
nk00+jgKuaEbd5ue1aEB+HRzvTvbMTI1Pk8uiTkrWgCKpJk63eP7MJjO1f4fapiAIU4sIFHJl7Wi
5AV8VMtWDd2Vi6xn+AUGj8brLKzmB2COurskBpbUdqtRU8y4kyhQM1p9b2PnH0omsalwgwwF1dXK
KYwfDXwAHQADtlnrc0572DtCZsalUACtDMda04LQXZt7ltv0UOa5vN9+xF5tNMfI+cL+mVYUP84M
f4kJp3I933iP4qytvabW9JLLGgjvzVa/rdVSpvtSLiGVHwAhBiiFfVMqYJjaTsoxq8tGf2aWyYyh
dsW7wgK4pgvAVMiQ7VcDA1XKR7QoXf2mmLGU1K9U9Et2fiyqJdeIzvDno0dL8pqZzVt+YIn2/V5s
9ORmBEY+PvJT+IGfZ8MsQ1+UNISd28BBNYAEP1wctdJRJWmvEAjnWWfwMK9K79RQEBJoFvzatELI
0l+mDwE14OVYYTPDmD0fpyp3CkU1VmLfeZyekFk/Ni5FdOqY3b2oEUtAczEiVnG5iNX+SN/vHCv0
/hiXcxF40i8pvJoAVcdsJ+yhm8od7LBMoi+3jEtjx9/RMSQOdq/hJLBEsI5LVuYtr1FXbW14JqEk
Bz4DuBbb8UGECxe/oiBTeAU0x23WzqeVkBH+SViMw9IMCtrV5ky8IrA4eVzDUMFB+VA8r0uYV/bZ
lmNRdUnimz5AT0z0IVh9jLFn/CC7KXxm8scA6a0RyK5RrubyyK9OFeR0MqoFYmDn7IFc5BPiltM0
0hco0ILC4k4aKsOBrj2WWrjK8GzxCxDm03ZTV7dV0Emtxyhxa2rp3R0IFKrgHCaTeWN/Ay28ua/i
OhFhRVbJ+YEOWK8alugFYve9Q2Ze3/RBUWkiQUnFwU+vSB0Xae7g7PJyPEZRO8/hgpBBtdKgYf8J
fpk4bRFJ5MkmZ0Km0x/VgHX4yZwphyr0uAsRK+l5P1Ni41D3n2YReIL9wq0sGqO48enfCj17kqe/
ygqz2/IpU701ev2SIxP+6wV9eLkidaBkrjiIL7PteBni0G6ryZ8pQc2AbEJJ9n2rg/iODvdkCeWb
tXssy4DEW8jMULqBb7xUQ/7MsI4Ymt0OXpj/BfqCbaIJARk689tA6oaEuAMGSO7aU3P/RT4QY9PF
Lus4/Jj5fa90paXQLI4274KilCUKNxBYr5Es3nzIlbLP9W6qgHWJiP20z9ak6sD0Jlof2dtzYmUF
QAIf7HA8H4AB1xTiVOh+psFxl4pLKNPHk+FxgOd1Si9Fxh7epEBOhUrmCKmSfdSLtZD4arU2x7KW
4bCv5RbeGDabcempnPG3u+Zx+tm0ZCO3Rppm0LoSt53Pr8gFF2xF5E6ecvM4xM2ud4T3K0ZCsxgk
3WzM4cCuSxdV4+SktCflU9PnIhJObzOm1+h08LbaNsKNyGd9cJPRDOOewjdox/OefxsZ62A9sf4c
kvtBkc3UXpv6InUPXsHallm9fqRFp/ifoXiO5EjznyNFEUZhb+7J6N2yA/CZoRU24+c6hYYnvdye
SMLW7dXw90RVxQJ9EIixosWrkCDkf6/EK8VlwSpLFwIUb+Pyh54YsibugLz3df5KIkY83RMpCmEw
gC4CmlaPYHWUrOqn/iiJTP7kntcaFIqxysI9Yjfi3hDZ2rZmeaAUow37SfmsRgJQPcUzd/Z7DzEg
Q2S1guNwIuO2CN/AbhAert9u7O2fXx3rjbWirs45FuPAUmdHDFI0Ill4PXoF449fPfmbymmbyKTn
fXCQ1JNHFuRsi6WyiI1b/kSySCMA9aO8pyccvqkrpSySU2n7F+E54/h4ZXX6Ha+uX9MzpsynkOaG
E1Gbzjdeu1ud07uGZd52LrTah+OBZ58Ier7KuLEAPJb/PnUe+1p5Z4pZ9x3gOANZzGMQW66TwXhN
TSRxBy1li2UombURqjkzga0WYAfzYsGMxTEszTkig271VPjGkkc1MDNi9rgNoewUaCAXbvePpTno
p3qSTVbjbtFyE3mj9JYWQPYvxOTp9TVBw8CgwgZrCAQcGv0NTKiU+sU6LPUvwUTUcy1HygW1aLt1
gtWl8FP3ezkydXa71WdJDeKB94TIQO7h8jzdTkD2sHoapgh8fKMGik/cDBr2s9wJbApi0K6Msyf7
Hxw0Qu/20BQedzGPeJIeXOyW6j1LpUa/19F8YlswGggV/ssb7CnZHYpgdX+AYoSzWOvoKidPtDmQ
Qid8dcmjLF1VjH4Bq5Hm9G0jl7WCCaPKs8d6cK3GVyXrm2sHSv0poawfWVj8lrCekLsnUpwIg01J
ffBdNFtZxTfqAlvqoLnBV4HRlahnAeWLwpr1r/yGXMAD0tNIGA+rtDSAT0J0PjObjiwPqpC4WRxZ
5pMoSkRViJkMxikYXIOYHGFjc7aIh179ZN0pWvtzuNhnWxYyz7XYjBr5qi2jNAM1fRPWU0OWE4nW
DM28oS6cKWat/3zAiWTfojSrV32NY0rcimjBGTmOkTmy4muScGuNSfURp/bBKyglZ/lXnPnTthxv
qN6vZaLto/PoILYMETMDhmDsxk10qCCfbuKg2FXnXq/RyZESqgpG/3H4kDyGsVYNTBOsEjKcyyAZ
QBOk7nR2U7ij6UgxjKojjTlNPbMvD0mMSWahyw7qMh1Tg5Hk6qE1FQdDkYM4XVbzgNL5N/cNUoCD
Vxv5wfBTFaShqfSzrKr9B74eyRkiR3O3R1wIJDAVjKC1hhohAmkivHIsotFVDjG1cWZoDi26IDs8
8nN9qm93NYERELw72+qIj5r9R1Qo4cfUA82d/X8xWZDjTCb+awVcLPCSD9z7Y1KoiHlx0cHx8Djn
qeuSM6BcGV+0GWFBKnlUeqtqryGDDhMbFswkULm2iHnpxIIfg1taCbvq03QTxnT3Q4NAJOcfRhgQ
QuIHygUp1C9j7Pf50IscCTKQLAfAjM4neDDAoqQb/vqq8+4mWog4c2P2nglr+ue0XKg1t2QRjiGp
4WA24HZP5eMhRO8oFZHyhdr440zirvVM24J+e19ETSQt/QD3lWXQGJgqe0i1UAlPNe/vjnvnr1ZG
9AOXly5h8TI89ESP2cM3X/mieDa4h1P1ugKESqVB/iiP66LE4fvAysUrH2M0ghH45lbLQfk9/dHl
M4/LFMsOB5a5KCaxOld+K/zFMoHlnpJUnX1QJ46mkYisKcIymgl1CJYpbsRW4BbkB0xsPSBeLTiw
MGFPdJLlPFdOhomRG0FSmQna+/Kc5GJ/5DM0bAHNnpYpb0k4gP9ukUwOBwYQBiYtsRfyF2LSzuGN
59GJvfWbEiMuyWnr8MM9Y5Yh1JsoHCSDXISRgbRqp5nXm6qmtfuC98qP89EgSJwUGU9yD4gZR7q9
+//A2BJJYMGarSBfF5dLj7A0y/k23PSDsYUFZ3H9YelHAOz/cu5y6pokwNOfkha0yA1B1osKwjx5
smI6fKOGTDRmN0gheUwt5yVKgMxZGTGJDafnF1BeSiSnk0woouqSZTDOGbtOGI9Bv+FpgAPECeqh
K6Z67EndoqgsF58rwoUP4HlFSpigHxhYVn6i1Ya14xpLCa8AWuHmABN3uYHJnTtuSErWvQ6hX1E5
m6HYwtHaVBQM09d1W5H+ktSg8wVGFtN4XjI1pT+xgH0H9lllcTrtYa7jp0buSt5pjG4yUaHiwPTh
ub2lWOKdsS3RA8WShnSKBD0YR/iIoXCCXOvmKr63W5oDGPjISR9Lshmz8r6WF0azXiUmztYRLLr1
M8bApCzBE41Qc2dCXeXCYrnb6IuRGB5xyVlMm4l6KZh7na7vwAISsLXcHXhFZ44haET1ECYriCjQ
q+7FlgJgQ5Jil9NzLhYTQOdSmPEzFzbsN628SzC+S6R6OsG/Ts2QbOWKfN3TbdKVg55PGOBHpv9A
ONsygYSnLA718Ld0gvPIy23/RTCR9pWXYuoGnW1pRhXJl6YuEkSjRq043k3nFQQjr66WO8x48FKV
f7Fyt8iY54M96qF97ucL3IavNoIR468wOOg0B3XqDEygOxFhk4U0UTZ4s3LSKcqkjnL7OeskI0kG
KvrVemLXVG3rrjo7H9JbL6Nm+DKE1cvRPE/KDi+wAX+OUK7xoyylEKQx3WiTRECr/85uDb1jHIJK
ie9QMCzkHkY1KCv52lwVSSbFY9uBPMnRgJTVVJQO6P8hnpe9hiWGRslC2eZ07qxbFPH743YIuCGN
U8E4mFe0WfKiMFtSCvecjsajFfwuyKjJl+Dg3pH+077/h0xEDHX/y1Ik56ppDUudDOJ30qhibbAS
w/GBSa4q3Jf7JB7XrDcgOqz3zpny+zp/Sn0rRk6h5eMTa6nVIKjDvJH9R4l3+on8Zm4l4C0y9GBQ
2tp49MXAUETDLOnqIX0qjB7wj5zlvpqC0gMOYrt0yxTAEaMVNt//Kbb/F6qSJ4Br4MhZy66OLmsC
necZumV0v4Y4dzOtz6WLVJioIwumEQj+4pu9ZfQIgLU5mflzwP2AR77Sh6AK95ZwSQIwsEP7vwoN
joCFTQgUicHDcwxw6FKmqOiz1ssTtuR7IgHIA1AB9nsU0Fq6kIadHMOWDBE8qLKhB7RpchHMOQQX
Az2eyLr3m+ZbvpX2ttBW0JaTFcVTJlkcmEc5ORDnMfhUMuUe0LGslqAEfYDofzDHCPTRi8w/Lx3Q
YYXB1sPhjE2bfWIQCNZYxNmVxVC0XURRJLwTC5Sspqgv5Mxv+HTVM+aQP5dBAFFsv7xwDdQEuJo/
V2xIuX0wjE81pv/LVUT9XJbLhmKPjDLJSLwfs11oTukANN376njYAisbcuSW0oEz2JUI0vDJmPdJ
/dORuJpfrnkTAQVnWOMaljVdt1RNry0c6A7Zg/LrN+euYTzfjQQTyYBi5jjRTeDO9Sb7MjIGikDi
Fi79oY3xuobL1FZ5OPYfyP2STl576/FwdaJPARGQo7WcVL2LgGDRfutsrNsB+lyMHLGOJsinhrRZ
/fH282IW5tHTVHWjRIL7spzPqrlJQ63ITRmxLOnk8adKuIjBCoqTu5YL/8H1zctf5auRNdAA8SAw
0c9Oqp0m2V1Zok23lt/gfnhUBBg14FrcGiFMfCk1gWmLSze3b0jC7Ptrhb5UVtqSyRQr95/GDGWI
aj1AQZzi1Dfgx/ydFRGUv8bIGc1e4m4x01PjzvKcDqArx1goLP9KYtdDeChR92u07wXK3dW1AGOo
WzG+TPXjtUKk/l2AT83tEKoumVB27x0k3rBHsuY+4j8un8Amar8KyoV3xnAjyKUzi4YXA9n6+/uI
5XCAGAfrY2Y+cvZHZg34VzB9P+ExFU/sSPM+1V/HrsXI3F9bSLKvWaSORUarLM7kCrw62MjKG25q
klvaiK7V0Jmh1PQe9q4jyq8G+Jp4c9QYtm377vJNbCSG3EJsVOfF8sZFzI3XDRir5VkLMY69pqZN
0GKbRGghYtT0zlUQMkrbHoXZCnKMXdey6k0ECBQi97pU+MdY5xIgo/T3SlHHpLK00DZvnevqPCr+
xIzh7vLHXAm0XSxfG04mqMWir9UKk5VVTLO8McE9nCRDQufGMPIFdlmIBpnL7G2FXppz5ws60Y7G
3Wgzgv4fAod5B8aTrlHb+IqhUku8C00/5B9o74pmHxeUUJUOIXb4GYiagLh8aYH3bjxzFqOuJg4t
Hqz/r9JKwROHXVJr2F9CanfeTHPch3Ydp3DDHY5Bn6FJ6p8+OBYC2fxmkvQeruWtRCLEtMMZsQHE
wZ61nkROZHFO5qwdgHf7LgXDsRsQ3GnwI7reJDiJ3auG0hH18OqYfAwTuxjIIMT2LqSIUpTYxlMw
jb51xu9I/cE6ZSerNxYRqBJbYc0stNE1J3yE8S/0hADztLIYTzw8atsDmCtDKibpTvkR2gbmRS1J
kmmtOuj8v8hift4YXuW5Wa5XV+EuaN76KbkTUcGgxv+UcJIgY2gJ0vD9iqdJmDuFN5W6abWKDXKM
xa403yPt9bHHU5RC4yJwSCAdTWt1zrdXoVO+hxj24x5Qxh3nVj7hA/YSNEmk04kGNSgIu5rJwOgD
uicHhDlUPtuYotSIRdeVsHk9J213SFXe25O/yFCUMC2ej0cDwCfv5Rd7WeNw4PGLWgBtgbai5gvd
MYy3/4ESQtDnOy+yuAQGWzNYYdsri65ZmQ8QjBy+Ua4H60t4jGEzO2mO3GVJMhjBOivQJlOG8kYV
whP0+MnBAPZhbq/vGQoLgNh2dybvraytJ1fk4Rlmh0ZNxFW7NV/4QfsoYgoEd4Guftc06hUw/94j
4RZW7oZ0nPD8mhfVMwKiLkbJ2JR3SgHxlbE7/p5QQrir/LpY1qG8t+6woyFlPPFPyIBOnDRqBpsM
sJXwNBlC/guBgTUHMaN87VZBDHmE3d2egrqfku5aBfumJMirp8RkLog0BQJkiW+5cOoCRXSCwWpa
eQVoRvKMWeOrb2kWw1YHdS5S+eoVG2NFQXEblNZPCMm6FIdWUCJNaJPKJWhzsKw9qhv0ecDqKDKq
ur3TRKTjvWqKVahsu0dqGk306pUMOgyqQxWzMMKeqVdaeZdFTg4Ku368L1LiWFICGp/Ah9KOdm1Z
LWcFFcnokK5n+spoLxP62UFaGvSa2PWxndtMG6ZHyDmerQVwPJdDxTJflzHb0NpftVB6r+djmQ55
NYC6mDyzVQIMUoPRv0LTCLDgifkOz8Ylert0ZfW/9cYSvGllz+Iacyc8phdJRSJkGHr9fjpXM4lx
9nrAkXTQ6TitGB3AoWOyDh0/d8hAjiKBw6S05E78RNfb3UVEE+JGOOeWdxQQ9AZJ0V3naca3dxt+
aSYaAziX5NhpAtyyrVvcsFYjhbjeaNBD726jPfyFuguwmHlJh/YGLNT1isspAWgzmGJJGCgrrJn5
JfiABRZ4zbmDg223BGCMwv7HxtaeeGmLHM1Vte+usIF/wUS1AGQd0cc8taO6UGkqgMOZmDCdxJCS
XWWvg8DR02GEhyJgQGJtpUiFiNBLOsrQF3C5KufsY/HZStsqsC6v+08ntAWmH1WxKInCwVXWz7/3
lQNluL38HHmT82ng8AbFSws9ZQW6bBAeowX0jWq5/rVWSlzb7KfSE2uUBACmgCUqnI2JygI8lN02
SV0S4Tbfl1Yy2g34JVyvp6HlTuAiITckLSCEjiw8FKTtmIiPxOASV+iHNhDIWXZZnTNPck7bDh1V
RohG8FcLxNdmn3SIKAy6BYyyRqFCIz4gt+HK+nfb/SRodF72EHrXEDtYzocSNDchgvEkpBCEg0LG
nfbM1UpCYdx31ebjsGPVTluO28CjXdKMe218vv8ZwQlSCI5TvUX7ZHRJBy8vpxFz52keZjNfk31p
7kVQiauE9RSOadgnUrX/Zrf41Pr/i1BpjjsnDtqAyIxIEhTBtX3bJdybdx740vJcvdy/W+z6gVhw
jjZ9FehvCDcDVPcdv+Pgc0JcdfF9sOR9+OHsVCeL9eeZbcNVfOE+qHQzcB7XiYyGvjOQR/cFWXga
QxgTYfB2fp+lBTtDOdYogG4hMcs2tjtVCwHDMvA+pnx0khNm4OgkeFp8AgAG/DovtWnXq674f0we
BgBJbo4A+oWMPj4L71MJLeaobBqk2D/5F/BLPLHSthiJo0gU2QG0sk1eB3+gecdMQ0VfVuO78rIO
q4WwlAh/QmsfWul2IsAX1x1cwOAecztN18elBS4xkL44xAXLvpiXC+Phhey/Nn24BJ3pYWJ+BQ0o
IcxM/oJaWKAyONuzTJWZj5Uit7DmDyNgDY+Sq5P+3s81qYEbGxwmF29HWJKo3Wi1JmXxvyuqCQqs
nYf4Lc/ZOs0N4oGMNX5zsi2n+wUw3hiMyp9iF6YwcVSip4ebHnm4/kzheyL7km6e66hKOGz6btIz
fJRMYaq55bSHHZJnyjmY7hXRO2IGAaR9/zagUjt8bCktq9+v5CUA8E2RvkJITe5IsN8ZMxhHmFZE
R4L9gJ08tKqXVnEetw/x1MreqBQ9AHrnenICqkYMxUtE7FsTfNqq98rpN+D9KMx0P5A7FHU4FZrC
LfIfa+xvbsxx1mjsu4lYRhJR8OJtYFlOQ7sKzzO6W2F5pYfa1SJ1qcEIzjlMtZYdNtEIo+i8kE+C
NytkPlCv/U22cGNbLtxtGiSErue0iW20YKsRc6qEz4d+DRukO4xdPanojlzAFHCuJhbTWpz8Sx+W
OG30FI/Jw+5vAE4IYWheTUM2DoEQFr02jLK8Ss1kIj++9YTkBniwhoCbs2Ol96O2IFRP6BbgdqmV
bbMmiCGEMDjm5aom2uamRwFlhg+/Yp8Esh43lv375PMnT5B2M7szVVkNEle4mTcvDHPypEYpourY
6EYxL0iV5Wjphfv7d+ZB4Snu+kwc9atd9EsCyu52qAOI9bJJ5g59rSGJffZ1PWQWH2ED2DnyDP+k
mJcY/+GRWbGQLERvk+RKXtCH6ntkEkMVTq9jMCAxeHo7zgJUm3UA45++Nb1jjHKvS+ras5XXg2A8
TQz4aH5rI17eDxOZqVVFmQEXd7V2eRrN9J9pz68dGBwL/0I0slmiXWVQT8on6HYcsvZXOAWFG00m
KvpE4o+/l+EtaIQK5zs1OvSt9TEkYVyp2O/vmzkv5irc/Nfuznzc0Ru+DWmSXZA2ek7842MB4UCM
5ymMGzH0lD2W7yBM8knUF+29CUziGCAikjyB+lw13QTiP7coNtlVoVa651jLJnIMvEWEpgIiVXf5
1DOcHVSpZoU//5MniB36xUiPnABGF8/RLoBM5s8ofKfUTtq5cUCmLSs2QxEkOc89lW7ahZIFra/t
ArmkC7HVEIEopcHr2qDxs+hwmtKq6p5azdm3rBi/iZfvYcIoXut4TmRgaMjrUe+2esJANf3RXqep
cSxu7uyXaYHKRk36eNfnEdMUCmWT8wSGaseFUp4F5Zmp8NmVpdQTa4vk/d6mOtm0EPkLJJyYWnjv
WdoewQPW7kKNEmSiP9fAQWRZwJLRaqFuBdM9mccLVVVMOdStFoZ4PxWn/29KJRFi7stEtIlRLBML
H60yfbumhfrBERcK9y4iV6plXyD7htEu/wlnWzzZYBa5qZ2ywXBnC9nbxs6I/h4ygv7sK2Xe+2U9
F5bCy88o02RKPJK72roch/sQ5oVhSVoZiXa9OUx4z6Upv8aniFQ/S6KCg2sIA/fRu9FwgmOesmZM
bgcAch8PauM9VgVsK8AXJ5Y/sF5BDQsYtLj9Yu1rDF2dxzzhevo+O3QdpUff7UGQFanK1S1PcwjT
Ikny8J9KZ5i1N25PpSEgzIntEKQ9MCeMzEeFG9fH/2nBtVFTyIb8YKU8FY4homkPMz+sKrQ9gz7C
Mq9MwqvRVbEHSVRfGy6KeUQZyUOMXU+RZ7RzQBmvXLpLgrk/ej+PmSih47dLQCPc2SQ3MqIf+nSN
IDuu8P26iRly2qjeYVzdU/rwzuB1jbTyvERt/tmDlfWkcKJh58+YMM8JUXQ80WhYvKdxzMLvh+ft
K79bwofmgxQE8vZJKECAoU2OnuAV7Xsts4QYqLpEoEgxqqRYZAVgDC9INmlVLeuRyPjfosloA9Yo
4bHt74zheR8VZVGTDEMb0Rmi3Zpm+huuGnPLyAwf5KlGCzdOrbko4c7Ahl6g1D7FrHk/I027RJD/
C2wUH7PBFAWUbzqdZ8kFleq+WOe57wE9hK5XqqyefegxslEJzKvi/zxswzggPpzfxbRovdJ+aQ+x
fH0WNV2N/KXQLl06WCflWGP/5KgXPsTuJUHF4KM62kauxybjlkGOX4xwZ2nM5522jHdrvLGgyj8l
4SyhiO/WvLdU7NVp0U9KPzvjFwTzMRW+fR1TQ/1fJpkjulhawHpS41BpDwz3zBAKRHKzCPYXWkaz
6vuJt9FzIlpgvJcv0e/qRO0p5VfWNh5HXHUW0ckoDlGTnBh1B0XXRYrijn+hbNbYgKEv2VWFqWEA
kVDdwPA7nxdsBrVFMt3EZs3SzvWKGW5mRdPNTzQmRT+yrR0G/0UlDEW1z/zXB6j/VeBbvQKMD2hI
kfBRZT+9qqAOZX3xrN8NXGrhSyaDUR0zVJcYptTg7S87tI/V+riaP5FhXX1advwXvPkj3PH4Q9Pp
6IYFWDz8X4T200FGJAW6EryT/CtvxjLhK9ZMnxjX75M4gfTsNVbxin8VPhywksCYXAIjFBkyi+ri
aehtgZjhWBS10Og1INQnFmP3gM+/VThSbT3s6n09LT00i0u1eZT5JMi3VDR4zOhQ1YImqiXoitNn
qRARWTUvs2HRcPqfaHjRQH9pdH3NxUBpjyw2h50Q50Al6XaFTvlGXynW61ucl/75ySHajNg7jS7M
LOGJEKOGmTlgXZz5K2QNka23sitllkPf6oXoQWQhJdAg6QxMPgxH/NcrwooKUsFHBCQ1pdj79dvn
jeZv5v7Jl1yxQCPn8Vu86RW1oprxC5pGS96s+5FgogGDOJFmk9I6JXKB1OPhfTfJbuqxHRZR7+nt
UFW7K75uTPkEHSmrtwdWde2PA9n0pNcQxJ7XRH/Z+6SPeIYV4yRXaXUW86hphqwHDB7Kl7hXqmOo
NyjbxIVVO1d/vTpqFT3DZZ9CqZDPDIiQ2r7g6jgeGXqRYs/SwvVPb5gSdeUxGArnqb1J95MYG2zM
7UNOP+yEcrrHnQ54MUhi8XBpzoOgiuIA+gPKA/sy31vJcwcZWJEABilj/MiXYdN7N+Y2DWa92s5u
n3lwk1x909dNKJa2n9Wm1b1QiOmnJsZNeVsiIt6bDrWEfhKIVZY2lz5AiOg0W5jXvagUGFJ+jc/f
mOajJfriKGQ/STNo2voxFzK5Ji1crBm1g0BkufaFKI8nPO0M7dmok9u0WzkyhZRCvP1m0RKfMCNy
352yOtIn8FtApt6N4LMSpVCrgOGugTtOO8rsGlqXyfl+B0VyN/t0yPEJd75NYc2UVI/p9NlpXk6o
/s9zMeA4yt2foGhTkbKLuvVHlpQ5lJUsL+KWcGrWYajOPA3GNEWPIO7VT9rot3ZDQVBDjP7vtNEu
93jnZJRIJCCP26EA6QkHk7KJmuZ/uE3SYtA61bWCzDwVAdZcHgGjF/fCL44Jrhj9UAnuY+AntyW8
D00H1+SYOj6l0H0zFLcgNA+sDDQ8Fnn2CJBQUdBPwWoPPID/B0jg3+JcRnnofdar5n4bnkXA0xYs
FHQaUpX+E/NlTcXdrShbbvltminK4DReVblq2ELGe4w7Z2MHyH+RrH3bIWidjuAaujS18OR8A+XE
rydfTAq2WKYe6NyzEkn3LFiRPhIwwc+UXreF1A38/UQSmhJjTj4VgLmQesazX4bdit1VEqkbYPxl
adeWrgeKSWZdmQiQqlqHUfFRkJk57bBgfA5eblcAPcCc9oyyilrlylkW9kf2EhV/Z6aUgB0BmDFe
JC+1x7C4rklrqEcRw/CQfrdwVLIwd7dCFL0pCtcvwr2XkXY2AgOFaAEhfrIBfxUQ6sob6sHOj5IG
QYGdsCFyqGR+6vGegalirGlEm+8asrDtJiiVwEkVmRguKe8qHDhA61GyNTAkAITi5Bt6a3cmC+Lr
dwvF1An2rKWA3RPSVIE5YBY18ZtOLcK8l2HlKVGJXth4DuUb1Z9Ue7vXImRpzN00urSM7gHUJQWj
FFPNjGq2ZEXCPa8rXbnKOKuKez/cwgqqBrfQvty2s+zgP+vsPZNb/cuPZ+6uXqGPRw5QriBHk0Gu
w3o5RCaF/aycWUBWK3SgXyaQzIiu4VAwwMKE/QDancQyl1Hib85l/2FPH1+A4ls+FKI/ugzG7uop
vaqWtTyorWqQxAkZNUEnbUpu4z9bPRR7gJxPCm+xdSa0TKhpp5ZFTC4crTvd8hLnmSu22G18vqxo
5WhDcXNDn3yc3f0knGCw/WQ0+nkNOdQU1MCCqzzkEhe4uryKprUfKOL2AF1GzxFeI8tuIa1CZWcY
nyIDfb8x2b37DWezkRGJKuvLLc6n4L5mLxCoQVr3e20Bf9QDAJJ0qB4Lcrt9GMODS+61Q2MjOSQQ
nz97jO7oKQTNeYsrKUjVyl6PKkpUKA3OpEHdJMsehIPIPkMi0KuhpIINWAiAcTsY1IgHbmQv91Nu
rF5HMjRzOxGwrVvKylIJGTuIoVzZcqXXUIZqtbz5Qj6nEE80aigJvNDOUhB+MWVLyIBsjfunvQ45
pGXs9iHn2moscg9JroeuxGOF0CxTEkVFmuvOHgXVW1cQbG05D/BB+mPrNEmmdvDv9r3n301xbDS3
aydOon9jXGJaPKavvEtfCr6ueDhk/qwCx7ZTZv2m7mZ2fEi18rjKDS8yhaZoKiHze72EQcmfcUe3
DIfNrGlEzF2Y94N2kolmrkIlNzBj8N1H9R+WQZDvtqvHQxZiORNyYaCHeh/j8lR4ErVhl4yrf2iy
/AIxOMmC1CdFNO7VEZl/sSUfmjRvMmNP7CRYPOWOhY5bTYly+yRpjKGGQ3Zl21E6u5nENsOQ+zFY
oC4hZ3nKS3RMYb7Lt9VDJ0f6bXg6ch6JMQndkNJDS2iyNrqIcMzutcCKI+RJdP9ULyfs1gKt8SSw
Iss+YGoVcOfEX/EtihCBiLWiWy4pjDPZxZ5llvRO2f8W6+vQdF5ak/Qg4Zdbar9HlNI8tvlmyfiL
7PS0149VyYj0jO74dXhxUe4bmQuMd3aXui//VKsnBBaoSoVX6Bk3QncFWmYYjM9zXecu/8dHin+E
jQMay4f9xvsjc1GHNGOBLBvFsxQXo6rK5Ki+EdjlVy4j8PV3witOzk45h1iE9f4d1yqAxDpTc2Rt
DDB7KuzvCzzvosa64V26djTabx2WamSMPzjdr1iT4GOkn228Yu5pxy9JlDN/TnRJT88iB7T1Q2K9
1Id9XBMgj/SBtnfsQQLhyw2KeReEmsDqICeHw3QII3O7KgaqJ9vL6nZ0sa4ueSAjYSnVTIqnTdud
lcPHaC9NpOVdoZjwrfJ2a02+gWvpA/gNToJ/f7HiWH8CeDkiL+jEtfAjtl7VXzfTiv67sv+x0Wd1
9qUZm3ASy0nz9+sFOTx6kaKV2s0TZkFF+rkldQhkQaoSFhxoeMDW5WVeVV6FJ1WxwCDQwQsaDwFA
QcG75YYc/QFRcAv7xGhk0Q9hKkQui3F0HRsSTt7Lu9hjwxpjhvFvbC2/f3Pre1jnkWA9xNTN/ore
ZJhxW7vP3ToEFRxHrHrXKg5bosmfDYaX903xUZjdVxleNsX93jrQn4fkotw55Ijc36wqZurz/RjW
O7V5QpuXs02dXUKBFe5VAKQctJQuMqYj0zBfr8z7Rxp6n/2UHPK+t3AQ2ixmLde3p6nzChfiEsjv
k2o9mbKGX//iAMIuGWr1Re3tRi2kavv4nlJ9px4Ep4uDbvxLqPdUgLBnB80W6DKopn1epEWd78kY
sFf2L9CfeSRkGm7dKAQOkYyvjuQx2s5IyCGph4A9aSNFUJB2WfI/uT2SjqxTr5JjiSNaoYIU7eY7
Fe7xmxfvEUjrksgC9sK8GRrbGJY0T+tUCvlpb954N9rKTO2x+hgt7N0tT7MDQ0pGTLjkv9q4CF/U
VlUfMcv9EVNSRk4E0gIs2P4XQ5v9m9vG0DqJdg0zz1oL1pG4VGxpwEOqw8uq5Kf1Yl+n/aQo0Hxn
vgxe4FfOkk9EzR2TwETthyQW6CguQwnAJsfCc8GN4C6b820vDq1ie2A0jWw6agEbt2ECFDijEKTv
ruvIwHyhuH43MSNmpa0O5axMA4cSkiqhk14EluqVNQtSEQu85ULPP9cbyPkQfNqMTTPrmdvAfcSv
eku8hYeQ5AmVl4pjV+8jRFJWPnA3BaFopxMYqh3VWjwfco2g3CauMHVxCWBxhcz364qBczFz/6zm
w2LDFO7TVeBBhrMOT2rBHU4/O+mMpzEiDB1FmwpoDVQlXrA5CZGmdHKTaiaosWUBBFH8ptZEYqdp
+VDFsq8rIDF4p0LEYr/+bXl5KkDwMlaQG8n0XOE8IaM6NRBeDMEVitXyeqeCP6S9vfO7rFSAUnGn
9oAendrc1G0sZ+do5ZikbQsmZGamQfU+WXvOCOUJsWwkiRzKwbonMi3MUBFPA+/djJ4Sb0OCxJvk
Ft3f9WpFwMrhwjuKI17EXBww6YKxHZ6yqwb42Nn7ueZ2ovjbRa5ctrAOQQsrRNieioguz5E8wRMP
R2FyrRqYGtBwvoVd4Kdo8BM+/Gm7za/7IDXRQjGJccPA+YbY4ZQVcPJssqdePQ46bp/5GdVRStu+
u1xnqVPrG2P8WhSU9S17pIszxuXHwn1jXoV3nd+yROFQyYzQpf6lpbeSVe0R3sFva6FcZjzLQge3
r5zU2GCvIrL7W16hgEi1oCqYccH3ZbVwXi8rAhEGXFesJN2SaMSkifKPPSpzaafDc5GkwXCUY8fQ
rVkCtlzC8uK3b8eTmhdV3ThQzhli2Wl7KDtzLXU+RU3zxfEFP3qm/n7W33jf+RNoKEzReYxwapMY
YOieXbiA3CVbYeeCX8NriS148eZHz/DCBXQCiDwF1P2UalTvp3kNw668O+JZzkGO+rwxieO/Oy+p
jBoCNsy9rxAtuHBRJ3V9rs+tiYnnInRajwCN+0EL07dxvDpNLsGOP2uMW7YrBPfMFxKq3C5h1UzJ
NMelBJPpTmFUo8sWmBBrbGLeu7m1zaArruFNPhk/t7QjMG/KLQrna2KvUrKkTQobP8/CesvxpUAZ
wYpNWlKz7sOkIgrzKigM7vsC4iXsnJA+ESZ1wq6JLr6UHu7HGwkYZAOENuopm82v6W/rD5CW2KhW
zrPqQR22/3eRZ5YmUPruAf0+KDCmv+f49Z8mlFxBLo1CkRO0iFw/oktBNKmsMNK47JK4nEt/8xoO
a1TOEiSCdwdlkSkwWhPDOAYQLH5XcFIMRu4u1Q4XMU9cOqrwjGpSNE3KIEy3AJXW+MfkyRLuEJYU
L4WOGfY7PoG+ZzCEtU/NwJrmN8SCcgpAqSxWtc5Wn70cMYk4m1Dg7JdFsrB4wYGk3gIvmga3YilM
LU4A5lJptAP+X6+BrUU+NCayyp201xi4HzI61P+9c1/cUsWLdRtls3aPR4nhFqABP/ZshMdIAxVm
KW2QAav2LKwWHtGsaCrEXTd3DJcLg6sJkQLI67QdQW1w0LYU74v3vP4o9JbQbGvgMaGt+DC1o1D6
yrjf6VMrKhxxX6/o+/Sif6Ln04cHXZ7Z5mRpBrq2XrWswdJJcmkvbdHE34XUoUyeIQSN4EqFaxin
klT2mBDm4rxyc8qPCNF+7ei0lqqoyKNHn/9f+opCvBf3a+qogES1eKuEr+q1IkslkTb5JjnjxUJo
U/+EZvfgezey6irAUuXlmakcL6aEf5lQl3W2seb+sUCfyJqR7WLLdhVW3hLV1yLSt7VY3dEka217
37VElx79gplhEba1fy90kzW8yB93g7tdYKP2auZsZnwbouKSHG33nDlomP1EjsYADDR25LtLdSu0
NtYww/O+ft27KMWzX2FPX0+qTchy1/FVeveY17dhOgDoWwWoI79ivJ9QXa9rGLLVUi35lmgEUdvn
O1kU8BYHMOrS7MCYOGPMNqpo/fIMjcuypZHshTZ2btBz4Cw/g0PgbVIGidLZud7GFrYnTprdvTcO
/zBbEsri5NdS4g5QWlmms49oooHk8L6ILDZM3IiUl6y+XFQl1OGS2SRR1YvpYpcHwCSD8AJY9jVB
lRusxqo5XjiztizQeNY5VNp7aEm4vnNp+DmlrKz+CbiqkF7KoPZDhiS+rsGTXq5QpqIW9YrEqlsP
cMwAtzpRFaPGa8jyxRk7tvm20DUX1t+0NYBhB8gV/YrJ4qTn3yME2cD+TroYUfzevdqIkN1jOkRV
yzinrXrXnfOkIOoOuSwKfOTCsrg/GwAT0KO4dBCkNLeYQqxfL8Y9Petz32uInNeQ+SpcyvxXm17L
AWWOWBMG462yXw9vfABNxwstqIf1YyN3ZFEEULJMmsEYSh/DC30rSrvx+xFollWa3NsMCBa9eLUc
RbM91eJ4B3Epf4nwoWB8oT9cVKWm+dGams8pEj965em3wEEAoLgpQJ3hIlookLh1V3+c5gOCrFDl
4bkUAN2/XEvTAQKiaOexGKo2R/AZbV/gCLSQMte2EzxM6hMZYYo4y1jbyP6qu3sMRNX16QXkHe7I
NriL08IIWAqTDl6JW/+BO/BqEuBd7Ur6RDPdi3zKizfiFmLnphpzjKRO5EFBgp5Ybr0HZjlQamNv
amQWqtSc13MkZBbYhyrOE4hGhSibvX1ZiLARzt9yFh3L7IdqwzzjcKpplShlszax/tm+Qwmk0O3U
rdriXa65rOuNxJza1GZ2mduGgGDzQ7P0nCQ+Z5KZ8fREogkgXwSZFSI5pgn5Q8RkhW1UbxAwJcle
nO3nD/65r6tg++xhO4n7UNFyl1PkQn7xet3VaUIxVsWoYjIljxnX02WFCSKrUsWG5IzmiWs5T9ui
YXfI4fRbYVTc9MP4GnI/q8sfI/kGAfdCr3mVLITXUc7i/UoEi8um9ASaSgVGx8jI5wCBReXwq0a8
mUuuxGwDQJ7Ib+pZtmMU7wjfA8XiiIaGZZgL4uHQD5oEEROu/5Ar04IgKFaPRudlXwQj6a2asu8L
gWa5pdAIsRu+X3ZW4Gv+GMgcOpJkFHnVElp6gm4ANIbQf6l9FUxrhwdWAFWZoXxzW0i7S+6AkOXP
5wZ/PhXPO02DXrNNAcmnWRKZ1zSkdQVMejsuXuVOMTYCl6M25IunGJGyBhtcofLHnoRQkDXR+afI
iMcwTjzmNpDZ+Qj4wf/aS+eGTIh8Xp8HyACyezZlGPR/U1FmLOiFEJ/zyuBWJKkvRPAum+6bL/bE
BBnxDvNpbHcpl7Lhas5tFoZACD0VZWggj6b6lZOUPZS7b6xWW2nMTbl0aafBkt/q+P1myze9j3BQ
yj0oqUFEwOn6CXgNB5TTicXtda4s8sY8/SaQvNXxgPkgorcDHBiyv5RplPFeeWUIIk90bnY54mMS
Q3wDAPXiVikCExkz/SoeWqRVERD/GcrzbvfVyKJjARJB68QE259CzEq9pvMOtmLlAQ8kMS2Fyi15
tdy96YbKVIgD4zO5VJQBiYiU+uik8KTrGa+Ua0TmRjbC67lSQ12v6DF3I/zCwM30ba8yIqYJw1Zc
WylHsuACAQvJgnyhU8AFYo3teuQv2rioeA2BNgA7SmHDZ6X28RwptyVmx9CjgQU1yXqUBzkmpbOP
BZ5tBq+9wpWJc2YqIgkr6dLAf7mcJpB4oKEuAmGJf24vC08C5j8QVceNOJw/zBU+RTMCCZVF7pOr
/sHy+W8vIL6rniefE4fS/e0p2tadKhZ5Bj26iN9LXGSqGfiGoRyka0NQUtSlrZM4m/mYi6SzEvo9
6S5oYL+onZuXxWd5JiyP/brKzyyehrErzfDVwvecvPPATmuZllWIlO/+zMDY7gcW9OKejvPXP6e6
ii1EojojkJAMwE3RMjaARTas0e8oz7dFJwvjTwvWLHm8bptYDzhu4Ag51yNikdnFTQgUbLohrQ29
3JDy9jpbBSiNJz4xvnA2UhOOdRqcrGhJe7zzcy5UFmSgMcJLBMC6f/wcoJ4xHelHGTbKu5E8bJS2
JF7qlMH2RUVWbz1/VpuqsjuG9Efy5doo0pgG1CtBRKsq1Vp33pDfT7TL5hz9KgKnD9QLvIn78H8W
PHJ7uILdaTuYM7m78cspBC4j0zeIptvZyIexvYGo/s956ng4HpPqJsVmIBNCx2rpfCR0vIqex1Gy
SSQ59DptpgSbIoJwcCrC2MmhJ0BHYFIoil4bNRZw/S9z4i0sCMA6AGgDMjKP9SyyVegxJiaDDjKE
YGhCaYklrowAVWY7W5GMKv7iMEQ33qehJ6q0Nc+lW3h/5Dj0m4gk/lYyHUhJ4ZgCSkxeoGta4O5s
IfCwbv+hI1pA0vjGri0BR/1CDSchSqAW3Wdq2ixwaayJV8BOanmKH5zUCzYTSVOQrD3eigtZxyWz
E6ZzZ7LYDTKtdNJalVQrtghDZ8P4/fWGgHMOaFXsllbycs6kDRQwfb8lK4Uo/OgYYaSFy/H3f2Ry
bbCd67B64kU97zgIHWUXlhpluzwa629yt4dQRA+Cr/rN+R3v7nDFD/nxfPS+rBw/gAkUM8dQHppX
nO2rbgdVCfq5Ujo3fAmX85kgLcJOvKoT4ayzGkeQo3oFKWVfQFBQvh+fJjReXZ1B1sVpQt86eNfQ
ILcz4tZNAeK2Ghi1q9WDVs82+/vLVpfh0Y6q9OAdpBijN9JiKMlAlpyrUKDt7hqaXImJUTVpJdZi
+RkjITNq9T4tR3Zro6cI1uJDkQrqciFa8rmNsNmdj20LVMp6OsVDmiep+ECIrl21fYtyN9838gMB
R6PwVGa4SRCpjULssUU/1INBfRznNrvWLVNRL76JdHt7Aw2MVCqZj5Bv69pIfOxTBGv+Yy2cTYMh
CdkU1GVByQlMypSGYQls+SnibD8a/EY94V6dcsGizXNpDqiXvQzZHfw7m+7oKPsmhqRCDCBvuOs/
6zKn6HK+uR7avUjAjQS5viNCWjJFZN0doxOTvfmgD2aEt7cSTTrjDy8TjrRrEAgOLcinU9RoUFxx
9JkqATQTnOvSz7lN8hsDgN0kT55+2vYm+jV6wcPuzEFC8V7GY35FLponBeHyKndR7Uz6DC+25LZP
DzAFGlmaSQBaN+vEDX4oNIQ67Ej3dSoACalf5z38+P3wGBVUKBLmNvymI1azvkLgXXbYYcLgkrFG
JUpUtnQuqTel4NfWdZx0YuyqSgDUhAvB5BG+xu6ZOto3DSo0dOFJ6XBBDSpE/Vw88J9t7A9aMZzr
2B+3NLMr64WLrvAuijbsItyOQyQyiZ//wAXu5zq6aYemCDiZqiux34doEpBAgiI9uvLWG3jS/+YE
eblpA4rH5+qSr9UUP+ZCp7GXOxVgVqtAmqD2bHEgx5jZdvpis648YeWoRlHsUq9qKIqjtlf0NhoT
wvQ7EjTkYpGCalrP82qIHWlW2l+2CjswX6W8IVNk+djX8hW3Q5+f3gb64UpAXg//Yh2ct7aTgp02
wqs0TExg34mxpPJWF+vmlN+nE8QjddT1nZpIkUfJTwC7pXi8QMznknnQth8PzBSP60ahOJzAcOmP
04NQ8tc2Anger0YJxxGlrjDNfRaIw/IQESMCOH0+JhfHsVyaAflinn3CMZVpOsxbH9fFkmot2T1q
v3ghK1vWRnN1stk102ZdOrlRoO23beUGWggYlGPi4mIzLiWwranVxv4ZZU/LxVjdANQ8CCE50YhT
uEMJKAQPGTrZUODpvBPtZ05phV+OlAMWwY3fSnB4hEp0M/grpsTsTbt8uI+M0Ait5bDTegdG8jGR
OFdqBdHRfBSIqvpHYWL7AJuZ+JYqBct59uiZZZMRePh7pdTaPM9inZGx3yRdtuJUYkucyo2OmJQB
WyQA51zT+iYmVDnKudWSOpfqNON/1vXSECF0ji3XUU60msNe9e4onKWRxC9Q6ZO6hXc2n9sX5Rmm
WDIDy0ud8+j9xc15aDlm8iPcpyDHBYJ+mGNcH+MrsWIsyD96A5f1VBpw8a/Q296IXlp8/n7Vlxe7
wP70U5XT/TQGPM40S8VXlS+eGg7XA8pBe0NWkDmBlYIZP7RRhYj3AqbToeIE7a81BA5oH/gEPKv9
Ro+WZRzpKK34REm4OEhXkAuv279EvVds2GkMiewoBkOfVy/Y/98ROzlc/Fcy+d2lqAvCtnEjRApb
gRnfO/6uzELwRltGaSEB7hsvTk9r28y7ecN583XGYx51g6renep4fgwQqdKX+mgXx0jIgHf7CLIv
4k9aOEuYYokRMdTMXx7TIIa224COR/zwv8Q0M90ReDqjj20kdTGXv3Y04BZUVCLKRUoIBC2SF6Pp
GuQA8qj6OQDIbqfkmf2RVOzxQjKLVeKSeqctncDHralkg9m2ZwZLFQ5Tl87bRsE5Znh22O0Dmdu/
bTP+MXcXF3KsBSB8W0xvHoehfvbc2ZEpb6wdxjNmzad2THkYSxermcpupMOUqf6DlrbqO/LFBKbf
l/MVhRA7O2VNq18eYsIKRRITjkdqst/ckFLr53zhw4+A1hqLkTTlfXyKaxy9S/3dNiuESMps/z0O
5pYK6lBuQuvDWrJD7S/QzrCWAtnUJ0WmmxkWwz+8cbEfvr3XzAILGctb/3WikOCJ6Ufx63JvcTSh
QO1P7yBa6sKBdK4ayACCDpEwYD0TiD3eQiqLJVCeD9W9PJFOJiSf9/Rse+KJFE6ayNYQeAAklHU9
Z4Y8Bswgz28h69nSUg75joaR7p10orsAY0UZIyto03gg3twihwIYotL0SjPhG8m1WHr6uKlGvbL5
sL74E3FPieObytZsBWeoeuLtRTzvX/0Gk24Tni111HLlOFyTkSjzrBL40VT0RwWwUXJcklthTljD
BAA3aKAiRaWUm22VGw4bH7t5mnwZoi1N4ociT14FWQJLSBFyPXphb/FjPrsyvhXORZYIIWdb2BgE
+ots+bnIg7PqEQW7zbtP5HWArxEWGl372+WohvVJRceyJRGPKhCJ7O5E/qfV3QUn4gVEWqZsIBs+
tGGmB7l7CSgF8Rm3MtQ8sbpoT5ZrH2/WUcZvjQ8EqXsd8DpEgSNEbQtfSEji14kuQ1aMVeAhN+X/
IK9JX+nbWALBZ+qmVt3vfYpU7br8pXp523Q5TK0V7ahLCdGGL2kw7YOPjRS+WQKij2CfqTc1tQsZ
wDEP7pYfMwFIpPx29gIyg6q5/US6h39k7YgVyTcz1i1exeGdF7/lMkYN1/WJYmY/aZVkv0gSXFAK
R2Rc4rhBHSG6/vEMryIXDCSZKVTa97i9TcQFmBZawt4rtllOQ8NwFghtyoh3zwLO5ZfIzO+NF6f/
dSg41pibfUXTI5chc9Wg25EW7/tjF/yr8Eh6+Ftx++LMFmwty/xQGpubL+/Q9/5v+JaxqaDy5VXg
7yAw79Kltw1ZZuinkjSb//Ug2ZOhGoLnIfPIpoB62bWB50uFx8BRb6v2lp3Ya0Yplw5grWbfyDoO
Om7KJUjVNpR0xH/p9WtYY7munHPs1jwxU/V/sk7qIXgkDoJKu2jobqlfqdWl6P3JMZ7R95MCGbyQ
BigxfBgVteY/rHWbiD4AMkbjntlI+rCEErLl3cjfxGetY1Z7/hTiRn8ZobIoO2GycU28UUqSQsr5
akhbM01ejDcBT8WNpU41aO7K4pU3E7M2j0ECcQpVAn/j2IDIOGSJpd1pyB+IDKcqx6+0in4NZjEG
U4cZ+hzc28ln69bZUB3tlVIWtXc8sz4PXRYGmQQ1e8fLsRZPeWMYCb0s9wVMLJ4AxSqXeH8glwB0
waKrwp/zR4LNyRFbH+6GoowJmRuMKfCq1xF2GDB+U+9icM1LRdEHKTDBPFuSj0Bg8qka1wASjQeb
daEcIWIM1WBAA2vxEf+xugSQsLJ0VvO+o08faxUwiZ3gsH92qjv0p8t3AX0PLBDR7zpkkjHcG1eL
s2dJrNy5R46NVQZoNoyrOc9+xmQs8eLPaviNaTzitNrdRuolhsh6Mjm4A/LA/CmVakl9/Fk0vvdn
4jyfZqmdxMmmqO+IRZFcPUNnvF/P2Hyuf26e3FZkystLczirxevywIji+gOHHQ/DcssL2jv5JsuD
y8TM6Ze+7v6Ceye6UMP9lK7KZcMp3m2Uzpc1UWzmCDZph53xtk3olMyhnJnDqyE2ebC17KjDC73E
xiNd/7D01HCoasWcNPeVSzYV4OL7335tfYIKwABgaoqzyN/gp9/jjsXWhU7us5ffiZB5gHQB1sFd
59+X7E6pN5zhM3TvXkNpayD+XwQZVkKnA9B5QezFBFZSrOkwvhxBBaq9qh1zgsK1HRuXzZWFNrl7
7S3bZs5tWsWNif90dx8bpieJJhwvxIRMss2+Em99uF6Dn1D3MZH0AYc0JBupCUASJicaaIVZbL4f
HYvrguUBP4aYCjthg0NNg7Tx/nG0XO0xsOAIIAHqQyyIa0pta84yAGYX/ToOsPfVAvPAFU814yPC
lyqamsZn5N5mFILQ2xezANV79pTtXzhshpr6ICBRHGv4jDWYFlrYx6UH4rcBVJiuwGEP0eIJ903E
mD3S8GUcAPiuhIwC20KdUa2AHGEExlSkUN0jiGGTFG6QK+UP1FRPZfV+VPQG4aF6lE33kX0D/56f
Yr02G9hNuWCY91dkgc7rjdgW2spJMJp58IUspzZ30YkcYwx4FjT9Urd8+0ofbc8H3kWCAXibjM3F
/AP9jGINrY6VUFrXv7+rFiucfwl0u0WP2KaYnaQmkrWZ+JeuE6w8e0jljXgMWYDrPdiDnSfx/QPl
Xz1BkpIFv2oaO4cj0MYk62Tx1ltDYIGUIBpWe+PV9qBXqW0gRBU/DYryNANae0M06e6kO17UED3b
XztZWJbzAWturwY+VkHiChQwT6t2eaojlYy2wJBz5d9d2nX+cGIWE5PLtm4AtD6QnX+KhCosKahe
FqZTvw9+VgSrO1NY880PINFrQNyIP0IYiTrpB7odIZFWocDRb+Sg0JSx1ddGdKlVOvVA75kWyFui
xCi+35MA9bgx5Gjj3ko+PlKxDToTIBuDmZAqs73XsSojU0rxMxRql+7lLOSbCOJVt/67KpKG2+YW
qiDBPfVNfMzBYYPRXNEbqT7xqn0orFgk9kvbRMk+jDybBQj5ya92px2rA7cZkY3DGEwmWCWVCk4r
cxA4uizUWjBLemkWXIDAeKZCNGKkNEEjvEE+IT5nrrxcZZmfvwUXCz/8Jv0kfKJfQUJ5owhYns+y
c9NCBp0MF5xVomFhoXPGvu3thS9DMwfD2UVd8uxGskiAqjZluOFSiyR6hjW4n+1PLAITlekwQQI7
xebZDj2Gj+GxlW4deJq4iCo2XPWZdu3pkDN+v5ntVPMpnnZYrJ4lMT46IzEnJhNasjf3i6bz0rxP
KgDnhAbVkoEOVtqs3iZ0UPDdteCBZTsTtFKUCWO8FBIMoTZyjOq/2XUSOqogB/CEaVR2cGOZCazB
i3pBuOIxOAvdcBgF3VZTdkKQzdkPUZeg3ajBU5CNWfSes4OGJ+Owgunbc1OCWPgfZOVwIdiNb1V3
OMK2jV0O0ZoToYgxDnqcjL3luO3kiE9oOjtR+v1b4rCHXJNsZK+oy1J3+9iQBLhkgb48YvPTS0sb
q2VsKv8rIq3wdOAX3hxfnLxbg8gJ4LrH+GEC5nQP/d66BtwJSwqVCjAHvJ1rhFXRvHJ+C0FjCsNY
OkfWEcEveNYvSECN/7wwBmQx/eOrKacoFZ6/TnepHqnP8WYcmJKsWogMK0rjxfkSY+PWYpzMddQ5
HZQYDkJrzpWDjS8uN/nbqxgJht+Wi+1SQNvVSXw5EKKM4u7O6pe9psGFiYBuK0329Un0e4V6/gF3
HwIxVpreclJvwnwUr9/2Hv0imJPwghPETwioBLc4o7uxgCHx6Hx3tX4UVTUktEUPHV8zEPWZ90Tw
ad69fgWXTJY/IC96XZ4LXbNMq9vwdP4rqMVuYfdi9QspOT1IRDw66Gqk5/KZggI13SjrlErqt1hU
MFUGu5PqFgYnfTALpoB/JWmxBn1i9sHDBg/6/NsstWQWnHoEEfOAkZODFqnXnREI4+DFymGIf7Ud
I/FZD8E/BPy3yE7aQ/oFIMcKdmfUbH0eRgIWafiV5nlXR+J1vxNBFuz0tDrfgeurLDtBDINDVlXf
O6rE/6rxIYR0DTFTAKcJBi7Z4bmBfmclfESbg0vWrFCcREH23wMo2OzUtCJM57yaC4R//sd3C4hE
SA1pD4y0J2+KY8UrCtQr00ooAQfx7YPIGrmqbTq23UZ1r2nLFp7FeiGnPPfWicWt+SbyjT9Ob7k3
pDl2lSfYoKO2yER6y8MPe9fwD+CIZTOE77JDn7LDAuIZig8iogodYb70N8HIUo7vysDR1mQ1DHDU
Qrp559oygVSdfPg1Ch2MsA7am3eLrLWMSA3mZyUVZlcIlpY27Uegn+zfes6jB+I6ZWDa+JOqDU8X
kSt/Kq/mFb/W2WwNpNqSilk5yj3wLqXKZ4LT+/985T0773dYxFk1PT0NVb1WIUUXPU4LnY3WU205
HHEZlKs45QapCWetaJwW8FOJYf8GbMwibkbtjrUny7CCidX2CR+IOgDLPk7U7R4RHDJZ+m3MMIdJ
96NiM6xLocLEQCepBokLWToOxQHe2hnS4jLilZ7uZ9i4IHtGHGJ1MyOW26MYn9YWWa637cFIit1t
dCeFx5rsiaoxvr3zQ8fyYzmgU7GVq4q/Ikb6+ZG0tzfsfNjeSVxxpD8Zss13F/pJ2InYfSt2+qTz
uBA29a2zsJEDfjBARqgxsFPXciGe4VmTciv2GQaXOBKiSNrjZ0+z6lz4fIna9TeQLPObZp5B4Ed+
qT8IWXOXgSAwzW8nueKmRaMv8B3VvJAzC9zsLwjnc0WAU+Ps6W27qQi1aut2lwPOYl6HPxVqtwZK
/+JtSQXAJLzti8KvdwYLAaLwLgyuDhB44Pcb5QQ4FFW690FjqBttQRyM9cqw0dd6sAHb81tqkxG0
Ti6aFa1/AR+HTDj0Sk/tDTqW4QI4qaicR5Z8FFTh2CAR0U8KwOKNQxx/97dvtRSUelBHowKtzcrJ
eB6zYYwv8ahsyi53ZCSbyUyaXP8S7nQn8+mKdY9n9vwa8IxfIkV4wOx231sWB6XMtjFtVn2Eauy0
OHp2P2HPbXFQACClWX9zc+xlfk01SO+0+ywtxhm8/p0q6O2wmMkr126b93REMP1rW8yfRYitkRCW
FITPglkEgxEPdL+r/o0vJYpBMUTRj1kqeSyGYWRrJR3t1Xi1GgS8nxrZw5ahhHYqeP9XlW9lj9Q3
f/xoARwE0VKCCbGw8jAllyOH2HD4gS0LATUPuaAVahXHnB5SH7NrF/D6eOZKDYR5moekVBGzURWr
BuungST0m/jPw3c4RJoVw0yNGcTZnFKNwCIOLcAS/olTuPDCLaqnzeQRpH5cWdAOmERfLFQsVVZA
odqISYA7tZ4vesKFO3a0jzsNRIdJYJluk/V5MOW/kZLFZ5ufPfQVqgbhK9sP5dPe109ZxWv3QTZg
1JYTQ1emPvG+w3LPt2NTHwHr3KfMAnxAdiuvRh59+TpZGgy4EbT1ne+749zeg9TFGZZxFit12vX9
9NAkwvoPYdsOaJ+r2fIV8ffA5B7kU/XpczAOTYvJQ2SKWzcEUDxDiOpj1kggfCHoha678dyAKj5S
7pAkE0nqQqWpIYryMFc/wCRURLD2PC5QiM11MrkA7f1XXLazmSSKkHpLTX2XaK/l/DEbx+Hgzqru
1eeIB1POO3hlE3OXKnw2DcuBZeQzRBy1KvdR3fBdtiNlpWB/w/B6kh5/yURdj+mJz3rWjgzQErTX
XaKcIzGccQzMOOshqPfYpu20Tm4fg1OpndyPTxv86D8nX6fc0sJx9hh4Wo1G8DdAADK2r9tHjOn8
LsV+egfUJx/YAuGfydAG8sh9QQ1v0MFVaYz6fAzXzctAdNclCAGpPa7ZEqfF4s2kGlFhNq7Na3FB
ynWHg2LC/THFMlzFiyKXuCEdcRZKItg5lmLRHNUAI6y6Sd1yXiFICPhn1vfbivsj7BPdqeD5tk+L
UhgOQ8hj9xfnF3P+dKr3TyJSX1tNPI0lULl5rlEYYDlCmt4YtGJUb/tp0lGJTQBPOqCeEztRjyg/
6zSvaMZR3Edc206NCQyIam7Ni3DP5xWlaWhWArqqqi731bW+BVVJ9u2ShWRyqgoaJm3kE+zwj+YN
TJREKfQ6xD0Q9sxrsoU0hTToDIN6669qdcuQ+sOq324Ch8EL2/C5JKX/tQ3b4TnuJg67nQTU9cFy
R+XE+gNZf4EWEUQOsO+Ale42u1C0SI/Q3TArI2dL8z5boThHD20KOWoBrEFBTPPMgVWurWUn/DnW
CyP3l+lE7W0PnLcbyqFn9yjZu13Et7kjW8uu+9co0cgOeOcQtx4pkrKgA0fgdotP6YIHG9Rm5p5f
byiMitR8p5jC3jLVLhtU+QvT2LvEAXPjsWiO7iUazFixIGTeJbSTLZjYrx0q9jH13wSScx3MlkEc
PqJyqvJzp/aayfn1OR6ylck9PMfR120nQ6G6i7zhbKmFBLtG3dy9cRcknLvBD6VFkzyy45rlPJcw
HRS7am50ZE2X8S34MRVXu1EtndHGE1T9WX0u3MOZrEMA3oZz7sQNeWfvxcvT9ZJbB9yNtfKiSE0R
cJkHN/Vr2+oC9jDp7XD022TUgOKygXkIf/lLOm4Bh6PRg5YyMeitMHNAauVlpJWsSWJhqmKpcX4V
OccqXuYTvVITctRi1+j0LCJUVKIFNtumEaBylL+pqMb9NMoFCOwq8HnyTt5594RGYhC2nDZ2Dt6U
G1WQcCcqJ1wmntHCfPQP/IYsUuS81y9xi9gCddzTyi9qiLikulM9URK1b6buxYXE9xxqbL3sn8cy
NQ1sw0TYFdff75oMcq8WsWxY7bpQJb1eZt1Jqgbn0HN8eoHFJytubXA8M8k/aZe4U380Sz8zHEvT
VhONaHehb0ZWhr1ASnKPInCvwqPZUvHee3dyCb6VYueocEy+VZbxohlbApO2iTvvwjsj6ckfbkOX
XjIXVaCftf7s+X9WY3uhvnPVKzSQ9OdLrqTofyIQ7ryi8TwQ9/j3imfHZVY/Wn4WjqkvUU4gFzU6
Udvrstkcsv1eOxtS2p2za0i2zNCCKMaG2JC+xo9YpzzkVtfJ3C5RmNENioUfp6dS/ROn1ZSKfuoD
rKijetjlLCp6EwkxVXPZWNGVxH2YCNwjS8/z1g1iF6IfkpeANT25S6zPU8+sTof+UeOJ1wXVoeFg
zJlCbQ4GOsWz8wU5XS91mmfW4DFYsE/XHE3oa05lXpMFrmL7XbMeMZOlJWkcCSBDJiCiN5nL6d0h
n4cwEiXnDs8h2U8PfuzWmeexpUwJPBbZVY9QxACjJK4TA8NVUbUZjFiTnjW/QwNcW8zaAW4ZKFWP
68KkovkFrRDQ0MrR01OISw+jMY4e2rX5OflTjqyH2XyjnZ4AynzQJT94UxsufDaHvMHLBylVT+dg
qBjGraYpEoJeP2l9ZZ5RUxYljNUmw81X97Pz6Al4BsYGfXjyyWyuRCWSfY1eqdMYpO0vgQ0e4tPO
rACFKb9SPZvKCDtfxtXVKQxYOmAUBD+vD6R8jjC2UbxgNo4phuxhuaLf6nfyBI+CVS5kQ7RBGWIV
3zMxORl2yp8Dc274F/7Wg5OnWJ2D5spsyUX+Rj++rvE+qoc6PhbjAwM0Lm5uPPjErgVe464DMOG9
zG3Jt2v4bmQTHcbz2WecDOvZTA3HZFD4OGBtpsTI1GYq8EREXO30yJjgA2Zu1aELPYS7AHBSwHiu
R+VJKrTEXqUT4+tq/tsRfGq1Cw2fqCg0vlzoZY3qyeG72eYMF3r7UGyGKwHry6K7oSG04YWL3YXd
RllBCbjF/Bketho81aXBpJDQH/vDRIIjriQ3kvBSs3lKXMGjlpDhG8ENTnTjtNi1FpSFm7RJHln/
pF4Uo1b6FLDvH9q3tVL8lPPiULQwy8Fmu7pfhl3CqBP5U4hj+Qm0MvXwjqoDdsfQCfjUUBino3Yq
jo897wTZYAEytx4fa6RRzNYwe7O2AmdI9F5vD8ZYpLDDEkP2hY8X+v6EKyEq6qNhgeX15HlL4dZY
06gZ6g7VHimMUbW66bPnNl7AuFLfWHTrzKpADejJ5gdmI8g7HwKNnaHEr3d2Z57bb5OLEYmapN2S
M6RsGiytHhZTiMNPrnDhU66wUKFGm2Vtl2GSlMjGEFdxhW+VduQBJfsuHvvRUKEmiZvwagyR9Nd3
s1WfViy0zctGlGQDoXSTtmr5FapXgSiFL/rkORQmZPHlYQFjrE3mhm2yIGUMOMCbr7j9jfa6N/wk
Jsz3INIwBaPQ66Zmjbso99ybGFfvIBDwnDU01tTLVwe/xxvp0com9YychXUoq5F2gX9goEB5k/+M
B3YCJ2SB2mrwPnX2Wsmz2eKOTSakBbrcP2qfW/wEb79Ukkd6zN73HT4tSyZZhFIgmritpD+6zp6E
3fWNb5sO2FeYQotqcm3cYcgRjREpihVrTEtTKT6XUcc8gYhf0wlysFgZH0ObNw/dOXZml33exdS+
jjm/hkbC19o9hQnX55Q6NE2mIGqYzrn4tj0ytqGJftzQi4ti7LqJY3yktFS4PApIBRiXoGrA/Q3l
prqXZGxk5Vkgw+dWzXEwyxkJJjlk45SHFIJ0l6xO31DR2vFDwLDm1JL190K8dlTwAF9k1Q1hEkA9
/S0WlmXdt2oehhL5pVaAiLY7+BGpadroD+Z/vMXn/8yKVqIcrTyfvFAuZxz1ZwCba7+4fD6G2oFC
Difytk5IO7A9OfhcqXiFS9EZ/KfV++ce2scaBxb3lL+9/BprnNs1qliNP6/2RxgDZlMr14qHNEpe
7JWTLEVVieN1mjHRPDru1YEjEDNIdTGu2IGygJrSwQBv3DKRjnnEuwNXB9r76iuKT2+bhNr1XdRI
XqBo8Yf/MXGarceDXg2SRw355/Y9vO7RLJuE9Xznaphhk6OoYjk4h2SuMm6eqFNjx0shBDcPZKgj
0n3koTq8He3+6H4w52r3m7crFSWj5XZq2u9P1hNeaNYxU2yQlze1YwZmYXK4usITE+liuR+9yZKD
r+OWZHJMYfeVh41rNuSbG39sdSqwv0i7FzFTpYDSrvVhLkOtQJ5Hrx1VKiIZbgrPExUOo2OdYrtN
MCyF1dFPiVFlnUvmLIw7xzgm/06DJo99hzZ5UusvIzffvQKuCytuYOlN0Ey0AnKZ+GuPNji3FnEh
Nphfe4zVJHCdQu4jF3dHKFYvvxsQ1zcLOUrWa7rQBYmgbJ1Ki95NskGWSPRfc3K9pR4c5P+yvRus
rClmeiDEuVDQmhSfo+c6kWtXrSJqcaYrLAxWmCgRm8oxTS67dJOpodTGC1V0np/pfkHI6QF39bDm
l56NeYY/Z1QEpi7+nvtBiUxNvHtC14C+jSbmG/Y1A/WqDqgSBrbpEiqqNTjgJAhnugpv/7rIM/io
kE02qM98003PfA12a7XH4xri00q9ac1oVs4gzrpSzgzyk+WS6/eUeXTCEQhMDUdvoeu2+wD1Z9Hk
+qlpwbuwxlJyAsuAy5ki97T1GfRG0Qc2HmNisOawBt4sHk/hSYeMiE6v7Ra7kHbTCq8bItz7twmY
t9lQ2fDASYXUAZ0dF1MZJ0jj+je3ihSVoe/GyCyof2HY2UqfjaswyUmyOAmyyMNH2HuTwOA6gp6B
Pfh0jyJmFTQ0U8YWJR4w9EhnMVyX26TvHP5j6+D6r4KF7Nv/xr+kw1yo296pCEeR+GoINHoDEUmN
UPedX6sICaFq/eEfdCIldB+063JPXzUVZD/UClWB8XuxypjdxxuIBBZ5ceoy3K0ArImVf1ObVo6j
yxZs9deOxmUp9OVIfEZOaKEG/JmWuUe+Biq6VggYtCvG1uEowlfQfnU13+ZjOAIN9scYVE6OuoiI
uTRnKmzaB/7pi/t5MowfGrvvugfp3XaE7OC8dK+Z/5tUcLGxnv2F78hD6IbXH7jDAO3/I6uh9lpY
3ZapHea27bpEv6+V3yJdbznggbHpo7tAORnjgWCAcxIEKZcUZ7YT9UfqbhVQnGZL/tL/qmdd5jE0
vC3sQvDUO+1PNcJgkHoaOjdrt0NFKj+K2H8iaVufDRXRJp8SALtUlnAFNpogYI0VErCFC3hjJ7sa
AsBGKFwV07Ci3TcawKf2oOK21teLS5HBW9GrwxGn1/Bl4oulBbmi8Ns3MW8BjPJCeVvsHNc+wfWp
K09i0yU7kDpYMLBf9+5DMGY2YE5XMF5cKEyAOwSIrUzaI0hDJkqmQ/F75nlvwApxj1byoAODQTXI
3wXIjFYFlU2tizevvPglmVE1zCWgWS+DirXDAqluUZ6m5n60Ktjj2dn6hJnmoWNnQqx0yu8bfQW3
hDEP1U5o+ryMuim1JSj+2lS0/i+Y57iJgBQj1XeqRlVGERBnJsxtAMh3sC3yCkMNan7NTOhatTUA
RjZ3oYHpVt86GVvY5HhhhNp319v5tSW+fpdPU/OsUfawht+4miP+Y+5IKvvG4MxrbUtBmK/jNfkm
TLofli/qTHPpFaAvILiV2DoCZLO9x5+4sVKTQfVCq1LWcVlnsb2ROnklUUKq4WBeS9XajBCxeShy
yZ2DNGTMFCdGQxTzJYM7Cgrt1vgRxjd5KH2qmX3wYSIFkODLopbMM0AlxJqM6TArph8DMrkOMEcx
VE1vM/gA9wWuHRjxdKs8eFHUCCBqfmtsDzDmjloK3n6e9whYwKwQfiuvmgiyH3pZdcMg4opvaEF4
8Alo6W/snrN/IbwIl1nH71FxW/CUOaKIo8peiJ+pPaOhNWFQUX1t6PzOm1YGj2OhnVmEF9Yia5MJ
8cf7K8rZAj4p40kD/oznNwHPP1/xNQAHHUz7XGrKyj/AfDy41IE0UTiGOlxEp4aHMIv/KG+USw57
7XmT6xzD0SxTu6qsotNiAVDSvdM0RJsE5j/ngBwFdzf68GnUkiThfY490YnRnHeS4xRx/zwYdAxI
21mGXTWt3/Fi/9PaRk/+HaOKrBoSbFmnP2RtwYnCLhB6J4TYBOTXSSyOxkykDENzGWYUNOAO/S9a
wwUDI4DjYvarhq84ZlgFnsEpOyeogXqb0JCHPHxGRqf2mU2wH+lizitrBo6ryirXKeFvs12NHH+B
xtkfSC0g1EcYyCIuvq6F/pxiyoabzqaMeFUlsm/vWUYaBLVXK0TjH7uCW73sNQNHSl7txb1o6qnS
TfNavYJ/UE2490XMlIxxtyFzh3lNcquKI5X0Fo5JQvEKiWlt+rhhLhwlcgTMr74HI7IHlOsNullr
IA2S+dQHpWHIn8GYau7lzURaeN8NaJYmL6zj5UA5DWRbaSMpE4+zrnZCNK2EPwA+FSAQDuI4zfbN
3/RfhlWL3b8ZjUD9VAUP3hQDhk2sw4em7FwrMWV1tMMEOPhdg7cwgf1QBJYDlz/FQ0CFr7GIDKGF
2Gf9M4Mh32YjxJFnJpaChOC5FFMyk1C/k+VAgvX4KsfZwGDxZsSZOxx+OGlVJGvDOMlNebN53Sb6
HAsuxs4lU4u0XQxdy7ApNTwefoRjn7E8lqNhS+wVAyECmOUE243BOEfK1B7SYbmeXW14TTiU0nj6
mouahAkZLMxe7q0AfZ5mQ4n/TW4jXDcnQzMNPTqN4Urh2F03YR+n1sl7sKoOQSqzlu+uhmqUXNcN
ww7B9nfOFANR8lq4MiIyAyRqmwvBsvrExrz41whWXXppM6+Y1tI9xHUIz2J/Qc6ipuD8WN8C3K26
4ZTIf8GIbs+DE4Txx5ADWji1bOGOwcCsGpZKMz1JphnNkTNZb7Std9oe9J4+C4yHymhISpu+7coP
K4N+UYXNMI2bS5vB4VOfThlRZDZx0Wa77RCEl1by4rfpgRa5WEvGkshElkk/fChfJOMieP/L+rcd
ppTJS12KrsmQEGziyi1DLnpJW8HVFzdC6rKl/wjYvXqhXfLQRazW4I/v2yDxjzULAhfp5AK7pMIF
Rs0ugV5S6aNLKzk/QdGasKqkCc7/sHiWTgKRygFK/OnL4QV7hg1gQqlVTjcYrNkcoYk4b7d2KQJn
7NCg4BvhWYFLH7Bns5mdB0LN7NKwwqFtLervI3Ro1JeIvusjMYY4m5M8FqBMFLM7m4LXXPTxRYi8
fZY0yM9PWwxHrF20tqQy2HbD9zD/meZRBDQni/2I77eN5e6Nx77waBzsfmDAWQasjalO/mbxtINh
n+f1v0HpzuRlIB2nKoy99il6X8A/plF4obTRZyMRTJODbSY9zotuDSovleqbPx6oeZPm7p9L/l3i
hsc6K72mFa7D137NoKjaw8fcuzFxFuDXeGfKe7bWPDRXb7875eQHQq+aNH+A6jpIxtlR/HKNonBa
YVzfB6aVl+UuASSqwKMy7DqpkfDLh2nuuyw6SvKYMSDwSycatYPRbn8UX1gWy9g3OBwIn5lCYC7v
/TjKQekkuJI5lRkVwgMAHYiasY9cYEkH7z9hfPSYKSwoCgdK7VWeUeh4LKguH3Ig6eZ5z/raVKzm
v2RTIVKUkmnIg/c4peFgfymOgh10iTGkyc+ivHjUlpYjdsQwM6/Y1ym1YWxV/iYVIU5rZFLA2PyI
YQ8E23dzFcTVqx/1Tw4FwgPFOkACGsHQB/8uNq/qhqjRzsxN7zZHzgV+6OFQ0CoNR5XCvwvk1pMK
HK2BeU4PwIMRAGXKtiAxaso85CWK8m7FVQ4P1CnmbProLopWLlitA7FYIeBudUKz4flwHmnDdhmX
NUGCpxpnLP8wcX90w2mrOsWP/iDwg/Mzwdo3gIw9h4g6XOHN/27AsMD7zmFaaTYeP5RmkOUhll/k
WtJWZ9FhjJ+TLppNiDUiOcnMVEhj8iQiZhC0uuzDbvolNjTLLuIKASvp62oBt1EpV8dDgGZeqLLH
o5JQuzm0wyAiJ3x+Jrll7qmC3Xxqv6SB2qcihJhuPhkFwLqkowH+kBSvFiixyGQWSSE85CW2+4yk
3On8BBP2j+L6xdY3Lzz04h5WmqQlRrCA3VI6IhkTtAExoMRcvrdKv9dQozdfnvcRzoJOv/8kfB7B
EYv/7JRqgM4a6+J3hULsFqSAxqj708+cZA/ntOmmD9E/BHzyFcEH+ydu9dixB32kg/9k0TOw/bGC
uBHr8LDdshjR/96y4519MK7kWti8Iw/CI2x1sEnR+27TEuydr2RYLJbaTCewPwfOJNZ9J2JmR4r0
U8Eo2C0s+u6vY8vHMrhErNqxxRKJHHzcLUSCXUKgJp05c7uv1hwdgJciOPlCmZS2yPXIj6zje4CC
9aOqCWf3tJbbNW7sQX4NXpI4SvGecClRKWKSNgqiAgbso7VBzbcoORwXxaHqBmxYGeSIUAIJmNzE
Gc7QUf8me57t5RD2ZDBwcy99ODujWZe38DlNPuUAsD/M+AYbVKahnxrjAbcSgw/gZZtPa0vvo9B/
VD4YjGrfJ8ZVyklyRARnQMBjEnsnkz1lcbCW5SffBn/m6rxkh+yUH5a8VJKiXWMiQlJ4saMeUZiP
brmDK6a0iieEpHD2QjVhaFImwyCrN6V4Ly9PLI9zw25QYf0PFOFe4rgwBpOvdwjw4JffTzkvps4/
Fqd7I3Ig1ppUO8SpJOqrJduPUpyCDCKQfVosl+9wpoDeXY0a44W6bYUCL8ZBqFUnMVnACZKxvceI
r9uahcbS8ki2sVxRWANgiqxRFmVQ13EOotl0RqJbE2HrZsciOTlwPlU9Cuy9jzRkH0Hkctv3WVGK
KaJw4kf8rC4HdEnZ86Ggz7nEuww7agZ1XYVnBoMVx1jSK3l/N5lYYr3Od1q+j4uyYKtgmXqEbIjK
MqZLx6fKVNf73Yt50KqjYwq5Yeq45mZ+h5kV0xQ3lXDj88gib6FQz25vQ2bUB3Qd4M0g1958gCZG
H/DSYMmfx6bzYaFwNw/Qon20mKlAaxMZoE/Sl9fKduJhCJ109/FfHZhdsmSqyAWxhZnRrXYxQQMv
jdsCWyJp3I9iT7AgcViAeTqYbD3LLQjtVIUNbvpBFmMOVHdq++L/SCYz1+LyQJXaqTEHOu1nnme9
6qN3jU/7xlUhtJiUbD3vDR5wI0mB97bAZYj9xQdfRhiPT0jrNEL6t/A4o51vYjKt55AfCjq8oklG
s/UlYbU8sSLYVBHjpimNFFAb8S/Fs7qZINl1Q53B4ve6C7Tr7dRXaqhFbFu86HFD/awUWdBmsbNH
MA2FtgpmnL94KtSmU9LbfKFD/7fr/Y5pEG3lV7k185bGmT+QIfn+IE76J04J0PnQtnEB579ZlOUb
aX5lKKf6ZMJMc1iE7rs51HF7/W1FVizDWzDUsqfkoEYGkfODoX5cSfnYuyiZUMYacIBim4Uogrsh
GHn1ss46olftDdL24WMBi/JFoGEbPcdO9VS2y/JK+/gtdKwYwFGhOf5yG/3PX5mcvMZ/e5n35POa
JvH72gZ3etCgbLozFaFfIPWNYpmuLWsNbyX+a6iRS2hF7r/FjW/b0LyyuXRdkSwBj9GZUvml/iiK
cSW26NR7QeOhDLfWNYazFf/uxUGYrY2ltQ0+SPkW5VS3M2Ubi+SsszZ0Vb8O1hmOauQxEJq4kUc4
IYEq33MQFNAL1l4etqSPLhLOLFZQBNkQBKJ4TP+QWaDAel2Ob+oL/GXk1+5ARJC0l2OvcS/0DXuy
URy+MlsEz50l+n3l/n/x8XjRmIQVXLiEiUGfI3SJVzT+p6aIIlwbgeTekedqJM19nJTLwRzjPXbD
5J62ftuYMFNhI/sII23TNxCCQ+1U+i/8KPgQZEetX4XtA5MQcXMjS3y14b4RtyX+lYXde3KPB+w5
bpAOaDEbYnhOqOoKYN54K7b4SIE4s2qQeJAD/EmmpdgDTKEOSGiCIUg+PzHt5FZnhrkkU+rwEt7C
m3KiOZKrLa1qH2g31d/E5/bTMnsp+5odjtJCvpHR2mZKX4majqgYf0rPSeI9alGVkcTppVXe2gxS
6H8MBc9QrwwAtRi3XHW9FhobRkut8S0GThcCYnjKJSPLkh1dHmTDIyXuoQCiL41YhyiDIuyjY/gd
o7Pe97DaD5vKXwCv/VVsK2OA8EIl26UDWW4jen5Zk5V4upB7InoQ8dGeq3kZT8Fa0tl1/by7HObe
W0vgXJEpK4ev93XzGE91wl/GoFddmk88v440m5dk5+Y6PE+QIhkdaKhwTy8gF4WjaVEufwHmet/j
lQtk1eZyRr2DLudAx8MJQfCiYvbddNsr0JvAbeCB2BF5LK2iizFqBLQZJ1gRe2PNdyV+N9o+IdTI
sifPzWIWt76fcCJi5l6y0bdr9/aGJbm0ynHwd/tTHYRCuJ+aIWEVEQMegYxORSMNoI3Vjuk5fyow
fV+TXRzKnnzJHGz37eaZLu6BYnioMdAwdWaG0LBoY9iY8lHol/yp9gqPHgKYf6EZLzbU1QMKBpvC
paJihnGy7DHKANq22xFVtQdLbRLU7QlQH1xjEMH3AmCY0pePZ8qJqBCzN2bRccoRW7qWqtMMMz0j
/M9HK73L3s7fMfc24LUJSTnaS6GOzju7W26SuvdQ389nHCSqS+hMLiDLWztPyBfUEEknxZily0CQ
ViWg37muXCzhN7BJz/bh8fO0ohGnv5JDNwgHQrvb4p4xftBCwtWYTXDvSame9pkkyBCyX605KDWg
l7tSlJNdrrYDXJe6wHIOj/IaUEQaCfRSHkalQsATTn/3AokBBf2ArtMPhyhwG8zevRvD8pWHdjDy
+SFNOnZH59ZFMsM+6P61gwC/tPqPb6x1lDKxdwf8mCZYRiJyyIj+sy20/K8Z6ke15TPe2qgQWE3A
v6DUbpzR1HRhHcp2j375XPSxVt/qgNvUNQP75wbPTSmt/mMBQiZIfr7ot5Lq4fzDi9q4ZOg6LxHu
yb+Fyco/Qdw0Y70tXO3sQZ/AjomYXa0EYNZVmd/eU+aB2eDgAz2CTgRIMNMCJ0+0uAt5YB62/NRh
XBA/yR9fr17cXxDMSUMxAtl9sggv7cFRibuwPgfbySV5J3zH3cYbU5IeV45kj4fagzN0ePz6U3ci
kSl5hwrHKucyIAkCfXzvk8aM6XSiYx9mWGNzp5ViGw6fC/fqEE08ICIrASJOPs/9weOvWY2S+Qv9
7jJwxr0XSyafhNRScrq4QCZ2ZWh3/IFZmfhhO+cYLuOnVrAc9V7e9JpMOYOM3XaIDqJt5sI7xXQD
PqWfUOc20XYRg8ZO5zvZ7U4bNJ7Q/xAqy4dpOe3X42/TshAg2saYSzWr6yBGMuTEJgQ6u248Gfvr
FKb2MOgcbfQ/Ly0RAZ9a6EuFPxzylEUB8xzBt9ydy2a9WFUA2x/XLqyPcSpv0WXniXZvnCWPFQ9s
Et7ss9l8pnxWaiFtJJdS8iAphaGTQ9lSlZrbP7W8wgjCkoHEn8CPk5txIFCSoE1XLP5CdXFI71uO
1Uei4GqKnWeZJhKJpMvm/0rfTi5CwL7aeVK1CBNXhdPdE2pmIwdNm5UOTS8/4ooihVwPMZn4S/UO
lF0oNLATPLaAHQuKOORoCPQAI99MiKKVt+fQcV4ZTlOsEnP6e4ZX6OUP8Ra64S+qMS+kZ/N5t+55
jJyvzIxe8vBqJ1kEl6hE+K/vtCdmI8nnv0zY25zhMM4N1EYI+yHcQH1LCi9l6HmBXpxOANuavp5H
LQsmW9wTFbEB3youHUpIpzwc2PDH4fVZ9THmmme2um0yhSvjtMkR0MoFJMwbeQKYGosDs8T8/G85
47cSSXPDIGxnH+EvTXdfm+Vwp2U2vghQK9trFgCmWjqSAo24SSlaBlDh8R5nLZVkCFv3cU4F/CE4
yJGTCzboFefgJ8SPKcqMlcx701GGdhyXaJlPjG43q/uACiMy5lxHS/R4EfiikvY5FsnNLNAEdYWH
SQ61YgY8tHOCWXaCo06hq1gxD4V3ejT5v29Xa/NzKDknde2bCt7sUcBevBc7/Y/8785z6vYgxgO8
1BwPbyie1cGji2JDsmqw4pAMEyMsJ16fM/IbJxdfaxqwhNTLyKBit3Er9737X0DJLNyFbWvJi1YN
6/ThO2pwjEagwmbLSswd2SsCPIr86lGbB1TWXIochI5qm3pSb5iVmw2L+Q735vrCzo7IberUfqBU
yNGZC2iHSPUcdBAGpR5XKXr4REyui+PBfmoS96jw0gXCDfqif5EgzQGKADWYx5dUoXPgMBfqjpPS
Q2jgRg8Pg+kSTrGQvHkmZl9lLZXuP9bpGCEZQUZ6kKNs/q6brvTAcBc3LRCjj3u/Q5j/W7lmtJHA
x97WidVkg4WlhVWKKdYjG3p1682185vd8C+ZFo5bQdnrrDgoAGuUxLsmPNJVATBjp7AC1rjT4yL4
ojOZ042HAqt1OM89okWY6meGdWTEZ5/2eoliwCFgVhzkHxKrPqHUGcrbHDp5HfUm15YP9Cn2ZxTO
oYlWJQPxWz8N7rd4/kj0RnkKr4JeUZmVi2FD19d+IyJOk5e6z5eg3fMpMEYLxMDc5GvU2Tziy/5a
D+813Qle2IqhG+SwPcwjR2/iG1X3M0k9SenNzhD3olbUy9kdFmjAntmWGGw3BTDE03/Fq5gvCcYv
ZZZStRLsyfXOigcrVj3HamJtpWVPHBGWZzznromZbslhjxlQWEFTQemw+i9Nvww022XSXYJGo0LT
Ubu4TJ3W0Z2r7JjgED1J1UkSqyT7CSAPf+GtG9Fa+Oaw+52JUayYj9zow2BmGVILBKhIF0z9rYsj
G1r0GjDZtypXb34rzTwMa4SEvkiToRhlKwIFeZHMh81kGKAlW9wpt+9zEejUrPVVTcpkZ28/a0yz
ISkekEZ7wXjt2+256hM9wAYRhX6J4mtKyEbauMNkt9nuIhiFGpdk2MK1HNV4JRVKm4ALtfwpAiu9
Fo4G4kHiwtbvGOeLUc4rLaSmg5piQnekAZ0rZu4Do4kbfR0oUo/edJwx9V5F7tACOwAJ+gpG61Om
FbD/QblQjA2zsZVkgxkWNg7hjacD9+I3okD4lQ+VA9v8KRcLwSHqBGxaWcKg1dsXbmgNrvN/J/aH
NKfxVCDbdYnQjlHCVZalDS2W+vfSrwulq88NeXatOB4hz6AbLVyc0gpCm5TAOq+7xoPcPAMYCBm6
S3e8lpUwPgPsknOuf5NNdtgBvOx3wMwgVcLLwkz1PxytTuU1TIFyzhcaCwtNSCfJuhtZvr/NCO87
jWFViyvPJ4a9++sLm23FbssM5Q/VBM3pQSGzkc3cIPyD78BSz4BVNNwUFACOxtvNMS8KUQO6Ostq
8+IZ58JYgid6LMh7Ber1XsicXhaDpu3jiUCFGoCdUp3o56uDrlkGdT9i3jnjEqdqns3FA/GI8/HE
jI/QYrwvZjhYDC5M6FaN2KIB6uT1AJgnRzJBm0T7mnmTwlSYNV5KcvtTj+kPXqsxshSaymwXRRtr
JZ75CdCSpxJN/+lpjNmArZC7ysut54LXivkrLEVcjT4I/LJtwCYYVue/JaMJhOyuXfb0SlCMOBlS
t/iPfJsyQczyFgTUBzX6IVYOJoSSD+raMAMbdEFtH9wrc17iQBv6UdGvK+5xxREQFz7iWNKEgJxD
ipvwzr6kz94slh2U1LMLb1h81dWbw+VYrUk+BTNzk4lKiwB7LdGvx53r13a5jXF+dJqRytlY0Hwg
JINJTdMfoveXpaWsGDs3Ocf6tI79FE3ffLirccM4ExDmG9zCUYHunxB/2/JE3JTAoJFxCc19FFzR
uojaelTAaznlu7fwY1ldjJTN4L5wvClmzxqQxpAZWJF3QGY4xDe0R2oVCq2ja085+v97RamzYBtO
jrUbn8X3yM4yS9MW+ebyTnuRxVHsfHrVzQTiyFLzV1y4vWdE4CK5VGbXTlsF9nJmXO8ic08uJNwl
NDwCX2J7846u1S6g91nn1G7SWADGkRvmmXIs8y5db7jTVa6Db4VDxIpgGCNmdJeLZMndGsy3nCOm
SodXht4AqUKExqizn6xCePZQdcpny7KqYqiu4c1OtAxV9vqsFlCQ3Rw8fWFFqfYGGXB0U5cC7y9C
Io2gVft4N2oC+kpHVpTIvpyunD7/vlW8ptR+T/tJpM4CLozbE7PBIY4qgftYSTWyJiE6nkwnv20q
czTGZr9EKxkbScv3g7/alXFUHXoUGTU+YCfI5posSNJsIelvdAoTuhVZ7/tfTUXWLMnwlBjwXkkG
SzhTGLmgk3OLFF9WCtV8/GmlceCwD1e6YeKHg0Nu/yO2u73uFzL29RYssJxiuicDj0nkV+gIFG1S
laQnO/76N9yYeOS3h9I/Y4AiTvr4aEZ8UZyRmib4u2NEguxy4xAnUOptyHjoY7qgHZ++8iAEO2HZ
0bX/nnc1OrwoL5iwezSCaPpnr0v8hLU0yNiNPVlHd4uBPoMbTj1QUld5GNhUHxP8ArAG+d+BL8TU
K60/xGmbEzlsIMh4YofmFINfpm44CAb1lIpqQe+xiv75wHnx0g1Jt8dwQtjeJ5R2t9m3D3sOV64s
OPUbMhJLzNGe5YjpiVqtxWdxibTHIJqTx6QoL+D/QJvvhXe5ChYf6CabKq0pzxtoBlzuI3lMTJ+Z
kb4ytIzx01dle+tDfvUH+g/fhefdOU67tUcN4FRiVEMV2HEAzMTBW/6LkHZuATAx3HrGV/epJteY
895SOcu8QqzV2e+nsl75VYCVI2tNyJMPYIX59RqKMjgPoMTx4DHSWNQju6h4RQcqNQoZhRnNR1OQ
uIWGkWzKhbZC6poAEUSoELJXH5X51m5TLarqJo9/pgu4+CBVF19EtN3gNCeoEFKK9KO9gIgRA05+
673lPdP9q2BC65rERAKGqtUfrUhdzvpQhdc4u7TcDT703WCjymXt4uYHiVYfsf2h06f5ygwwkWz6
wjtG31aQwsIJKVit1BkDe7vqu16uJieLtlc3NilHXarQhvipAKJ+tFfvzpal+sVUuNr8NFF32JG7
2KOmefmdR90JkbIIjmfJKSoAO8ThjJy6bMyjRaGd8+TjcSzQ+RugNv7SebsL4K9W/rizbNICbcf0
yqEw+yZ3jFOeZUah1LhfIXrLbFL0RrZA4NUWJvup09Rqstt36kbPkp34dYjoZ0SAX0ASqVw+D82g
lAavxMUQvZ2Dr1VqpJJAO7OmycR0Nc9nwMrMYyJFWWwJYJ5NtryKPgQr9/NvS0D6KH9sQio6eoiX
V9gWtyLRWiHycvTqMNuLJlL5d0Qpv8yfqVVcE6rpdbwA31sS3bNDgi0ZF0IEj4oJIA2yMXGHGX+S
raYG5UWlyz3PIFRACgRJ4FbTVaM5FsZC/LzNvnX+QT3oYiGT4MxamyLsUhppNiLA0ayMa2iuSoTc
PXvCGANRZO1OMOYNKWtdfOcS3jlJUmvH5Doxxj4Wf8+XL4JaTDoJMEqu1F1rWxAAZj9cIenP/EBA
hRnulbvDVD1LVOXrVoYHNBRipXbB2CD+/hOQs/s9mdjZCiMapEt/NOo/MCxT11jknMQK/+Uq9Zr+
bmc1SpVgTcoe1Yp7mc7ojchjOHHmUkaC4d0tZPwvLlmtNujwwCTnXJveWL7H/rikczaqBAdnTQiT
tEPGnYPr36sbhi+TN7g5ByZZg4UxIS5CXMm8KBkGfFPbnmiXmGnhNqkEJQWa6wt+fv9gLcZ5an7Q
q9RvDKmvawjaXgd4iuVS7Bw7OnFTpBFS6hI++jVEkbprPakDtpVtCn7WoTHxuWjJi1X1Q8tZoFoS
/NvlnVSzqHSqjSt62uSbxJuRvEnsKOvxXQ+c++4iwG3GI7Yp/1FFWbJCWUEF0o5k6XUlguLfLeTx
+9Vj4NjVZ4hyrXHYJ8hIOJkw1MVTeoEavw60VEVDzqZKX6rb7H+wxkLJlpIjDogivzof+qqR+J22
KSIbpu7382smY3rWOmtIXSIKTBzm3xWx09nZulKnekdqATJ0Wz1HnRKDqrEBnYu2epuGyh9/yR9D
F/25mb8YmvBuYojWJCXksTty5ftUDnQUyopgluYrtNFsUS6Wc3viTBu31LZ3iR97v7Zq/Bj7/35Y
0QcTM4bMc3WHyFJRtKV9HjIbNe2XspVpRj9iRW70NIZRWhiwRZXP46Zi8w+HSpH9XYH/cgFJ5aZY
TZCD9blSV/wh5FcyKPMbDU9k2524cwoezmiJWTDwJt8A9jNhbGHw0QgGG5H146KHPwZFvP2s9u6n
+OAFy8h5ELzGYtVdyNGeU14aGZnfYqMN9DXBW3BrAsYDmTFAoK+d00PHilfvmi/+bb4VzDBgnWTK
H7Ob7CYjGNhoa68r1c7ptBvYgrnPebXZAHIoiK0P4looUeAaRYeeZfdSKFZO0mJq20tMKe+VN6kY
JpgsOQ4CzSgPiBMw7YCUE8utNnI4ucopWdAHriJwo7UOX5VTcTVyWe7I06/vvR6l9M2kTxB7hTSJ
g8718UhRmv1HgIIq7wkT+oReEgP6KxfC4yl0O80URanbNLr37K6YGTEW1HR9OlGk36PdB653yfH2
dqjLWd0muN5if/slfCQSP2/VSD0C9clU6lg6fYQXdpKMIIyHpD9ki9+MkQxeWlVH3f6RWPeRLD4T
G3ctbd7XmV0K8qP2E1cJc8xfhAou1g6IYBKqPi4DPw3lPF2NhXNvQNchrt55+oXwXWLl8+cnDAzI
n4CI45twpe/cEXkPi4Qslq1d7svAV5ov2SaUn1FeqVTrCKaDpULYzb5UDu+zat1GWKKIVHSn4T/y
obT/4FC0Tj69kb9pWFOzcl9PFOxlcLGMMrxZWb1KL0YWUYfavZ1aXLAz9ylZQ0c01pagr2G7BaXv
WDXjd4vY/GS/PhanSV7Ohp7kF24r/Ebffv1ir4wtGyuaLOdc3jE6EvwSonncGZesvB/DLvtn/rcC
bsaCnBtqxCUjl6FA34WiqvztifLhhTK01G/LF0f6KNzLkcPAPDgk/2uyMMNFbHehwIA/JgxR8AYK
3GpySNOwK0FXx84zDvNfSBxG8btibVLodVM7/EJRqjFAsSexbH+snAxG0lH/QJoEsD938SFiLGxp
IEY5QY+RWTu3+jv3caEMi7RKo1Vk+Hy9C+FcSzaWC4+ZbB9aPnmhbdAD7mZ72NFYfTvQhccKrA68
LhuM4J6Se8Vvjf2qbAWAJ74UYz62kkfQDAKIk6QH+6CK1C2SMbFcAiPe02Yol0eOhPWfsRgdWGN9
/JLCSG0rkGjwsu7bDBjrHyUdMyHrcN6ijVeZBR4PUO/AFmgfp/D3NapxwE23xf5Ny5r4pjXbMmZA
ifiMiq51ptIyb/v4v1ixRwrCrwDDp8qYSZPgiSMqGjkvEmveaWRaBeh43r4EJnXcFboWK73V2RJs
G7Z8/E0kO//mrFbHam0zfI0hHokKuY7ZYXw5pLIdo4DNxwpyISNkGZictRK+Hihvj4pGNu6xsGqS
SQpBYsYzeLw07AL8Dvx3SE15L5W9xFYJvOZMbXLq6A1pjTfnRHve54J7BzUaa/eAGhqBTX4DPx75
Abp6HEVxvX2yjEkMghEqNONzMjbOajlInygvympRglQBlYcKy+LBd2ooX79+ENhu0H+TmJMltrkJ
9uXDScdfRNtDTeq2kDv9rDP9EZMj2NWu+2QqSRBISy8aBc9yuy/jtiZYGOho7Mi7wEMqUl9deccG
RTrh1/oZgB2yOUjQxB3NAuR0lzQPBD2wauVwzO/11lFxIE1aFz3dz1Bh4g3T+S9pKHuppHxO/Eou
xtpQbMlFYvagy0sMYtdnrO//wdpEEXCED4N82ACpeT81KP9aTZiM2FCKAcYxuupfWkcwNHtgw1w+
KqcuuLQX4NhB+8CzN7znAT51Grlfght+eMU5qZqzt/+6MXkw4FdmJzSlWl/+XA6nx9Uzi8q7fdRo
A8GxgCweVqylKuda9Q77ooe3Cle7sFWDI08skALZpLFnLiCHw9F8Mf19xK8k432mx0NyxhYm0lsw
dLLokBp5lq/AZR16mv8wC3HjbwDxcBb/aa6i+zVT7z0fs3vHAyPw5440KJ9sJ2f6BPeJ8xpVvVNI
8J6hVcGzVcO+BwfhRzlk2HebMrKp5pt3pCc1fMitdNPPQWB0unzKmwehFrmIfD2kvKjYbJuHqNGl
X2u/jnnjUtrjemzkAl7uSctnQ/oauL/HWB4+TiOXLnwk3fSqTiwV4yze2sfSXfMwRBLOYebCkShF
6n9mfcnSgzEJe5uFU0pnt/Hq8Fu1A1TkOuv6dzfa3aloVeKk3pNQk1WSVkWbF2LlcFnToexQwQIt
2+JfJnm05caU+L8D21AyQQGg40UsbLAH6OyYksmmKPjZGSfp+XObgnskd7Uh182NiTXRnYBO6sX9
m1IDHb8nNyv1+JrkFhWgZlm22MZ9vMJijX+3nHb/viZrqkpsXFQApCWIK12VfEw1gHaGr970085x
jESZS0IVcOqWtEAfBfC7GmME0+JHmBOSzeNNO4MPEDT4QC3iVkw/S0YK0OgKmHW67IrKCjGPAFVW
5jMKuSZXjwPrtMLaOIYbA0hCFM0jSEpslE6Z9gk06N7jnV670jGugCmO/0NFRFfVNkRUuxZXzNTn
BB9fSgVyvVmT7jtmUKdNDTdHnfoN9v6rcFrMA2NJtDIEeD8rUGW0OoPhwLYNj3tvX3lhxE6BUirq
6nwDsPyeipXGeFqpDpMDiIgHdPz53TBr+F6W9NHH+0vqdnp5FidBEXQpO4sadLNUsWV+yHQ3qWLR
fcdOL9TRK8dI4ffM+W2IVelNJ5r5akZJrQtg+czMbv8vzzO2piIYlgqPgYhXTOBbQ4Ux40NoLFRs
5BvR4ejo7QVpLyBmzJZFtAgzA/PHDyZaLm8e8tYSlL8D2pMPCjzAva5aO0pmCWJirJQKVWW2Yzyk
7OvBHDHN0K34uOfBz+WvoqnQcmA6Xni5uJ0TmRhZqClvoyXY3EOhbdaY6DqHKevMEkos0oMcprbK
pDMCIMbdbgzJ18AlbgGKYmar8e+Leb1jngKISlKM0gieB3oc2ndsiuAUcPdX6rQUtTzdyeM7uDM+
p2QWXP3kHCdmF7U79SUlRDC09BHeUEWkNPapQeN1n59P0xVz+FxYSTB+Knb14c9uCl1lrIL1HXP3
2ZpOKh3RBtgUO43I+nbKWkUWHyH0a7/3whusW0+nLvYTotAwMoR8i1ldEfJkTKTmy/VAAffdYBGq
e2j+MXz+OAtzQwh2eKbN0Ed+m8MA6Y/AmlslNRVs7CW7pW5IhamR2fdGeGZRA8cnMfY0mfyitIt1
KE1AKMkcsDT2TwdnAfKKOt/OKJvAZHgg8NIZBgAagbTgY/L1NPOn5OIPPgICYivfhNrjhVHEC03q
mYePcyehYH/JoEPfVojc/vBrLMfVdinhmSFiOpQp5az+KI5RFMDDcQVTRJrHHc0uQKwg4HZOMifH
N8e90asbnTOhCRM2nHsffmYVUO778n00NdYmdlnvdEPQz2L+ap2Von9ENU26GkOiTmtJnFr/jIVH
Pc+9AaRUDt/RXCV3GwZv3zl9jr7PhEBt6TQT16ZmFNYE+JDiWvFztIyEwqX1SsiSD56kDDCjcNaC
ulXqIXKmCWH9bbqoMkM5XZ+W2R87JQuSz/69mDP10FSvyc8MlohNlsE2SdwQS1j2wLcb24twPt+t
e5cNsVRpiipQZ5MYdeJ5253no8bt8zn9azRQ6jhT4SXkXxZaus90IUuEiwrtj26c5SNPocoFyvK1
vqBS2AfkkL17+Vhm2K0ONHzpvZnzOcRekFKBe8TN4dKXCHfix9g+5DvH4wxaW/S4ojsgoXOgAlG8
bRoPwLcBFqyFoFnaXCJCUf7Y6hCi+wZLlawiB36ry0px7PjaMf+dGqxgsA40LkF9KQtXwQn2MQRD
LUf9txy1u+GJrqfQsl8uUrCwrB1S9wps3HuYZn5aNSug2fipNHAqHzKITHnvwDpVOggGwzQZNn2o
x+b5u7uALLFrjGjbK1nrhfUSHLie4nJwg91EWY1d3ufw9RVQwBrqi61ZOAAxEat38l6il8ipE+tC
QHTNLVj2/qdqpYaGIFkvYzqoqf78GnjkqfBd7E7S8DXUhWjriYouuSZXSeVcbw5TpdIN+TRPaP5r
2PBULH3BaBYIOl7aZi93aEb+oKY49y8LZus8Gl+XNGvqw5ZIQTcHGIiJ+lEsN8EPs8vNeK89qpN+
eFMpflYGbpL993TzNIffP2gIcdJC5B6uXczY9wtl1RqVX4mvPfC6ddhOY98IzCmmX0ot0mGrohOP
sxmL8k4zaKEspw9Srw3UvzD6fgHvl6HQEcjeCdYd6oFlVdrvckryWhgLPomJVmi2/LdlmQbiWb3j
EYVgjFVSkotP7fgQ56neqhrXD6Q4h3gRYXymkiewcGWxi/yI76BOUlIEZ0SlYdvF5zDIkFbEeomt
lj6yjA5UqR6fjWM/oazsdx9G8dHIC7inM94mFV3sjXWie9Oa2fccTdVyZmELAfSCZryaVyWd4uOh
LuweQaeI8nxjElM6i7Q/3AdDu1wIPY3v032Z/NcbkbRYxyDxVmvtGTy8He0SbkCzTRRG1iZ+EPwa
Y35wnSOVS7/TKARdJrbou/b+zoM7fHITPpAqbyWTdLcS+Eu9Sl77TKL5tc4+35HCOnhG7RsDi+qB
narxZa4Up8rez/Ym3aMCr4fNgOKeAvuHY8lkBj+JKlIp10+c8VAScApHK61xFTHZ1EvplC5o2rZr
aYXhtimZRxECVMCwonF0/ghFBrLSPXxuhwexavie9v75kqNDeZNl46hSnRGW+Uoiu9TfaMWNP0tf
IDBliX0DyxibRp+PG4gt4NLDkT6fip8RaX7Qy/B0GsJhlb0ulaEJ9mUunZs4c69AGpzaLatDUSuv
+/DV2AyFgALmO1NL3s/41FvFnTlt9SmsPkbu0XnU/1PK3BHIbjdoP5qxhRv9MhRoFHrWPW10J7qD
yMOigk6/3IwnJDTAxTzmeN+Hiexpt1pVQuZej+gsgNZsHJZziHG6lLkpTewS39aF8NzYzwy1mwmD
Al2EXTvURqWl4sS/6DFv8eJVAgoNBoDsYPsZnnvgpGxCd8LPPqkxm6C0SB42dQiaPCMz8hR0L/bq
UKj20G1vNZ/k18pbBTgFp5HcMFzERiNfd05Nm31C8BlZHal2DAIbh4jHBvEQKB/Ugm374dP3WtfW
8o3xuNnLfE2+XNYwklVZXemKi5Q3YFSqAvF2kda34NxQJV2QXNBJYcebwoFzw5kEYfoq2ijbzVyi
y3J8hbtKVv0ksO1un3hDQKohda4v1JaYvKm/UeuOD/ZXd6Bc22fuPxzsIs8Pu+1dOIZbTPELE1Gv
Em2d7ugrDuDLWSEIVe3LlB7n/jIfmqFhaT9TfEawO0edYRtj+f0wR5vrlTDXnOoBfW+/hIF8Oe2d
2q8YWCbfWvXXIBbTfo8fMsChJX0nzH14OxyjnW/ni+SQF6az3MztLmzD+bZM1/dGYQXda8q5a6qk
DiQB/4I3JFJBVZpmr7R0MaC3+/gmJiBryHJJsTcGZ6v8Wxm43GR+T0qrdgjDocnIY+eD5GoFjDQ0
FJUMiop8RAOzRdEIiXYLRUvjXMAcaNBxDHJadLdV8hJc5JnZ5MQZICVkz8ShUH5aE5xRzQOPdQhc
kePXjBb6hstMzv/NWbecuL0O6ZkxWFtUqZqp/FeMctGja8KxgRuodsg24mJp/r2NlEawTv/uWV7G
uUb0A11ikMq7cTAw0eaxWc9yd6WZTf9a2G/wCiyefZLnIPbPG0ObS9Y83O55hvEzaV84XBcLPBDm
RmPmqjeAd5zAtj1aqcQHNQLEs1H8Cndg6aM/j646USi2dcHsxHWW2m0QFGKBmPAhOiQCf7SonuKF
i5X1XU0qdhGYDGCOuTqJWSOeSRHUEBQNEE2l4PwW+0s+m3k5kLVHf7avrnsLdKdm6KdYK6J2QO+9
T5lqjg8/NapXukKdg83Mbp5rJ3hZNQBsrKKzYVOtMqZx6pmkFiNsiQbsHLMj0sZ12TDLKpxPV9+U
Gw5BTSdgzNVxgTD87+IFpX3Req+Q2hLxLlHNESW5hIUuYZaLpCUuQFtSwSdG1t6bnfCliIYxpWKp
Wno76qf3aWJw1r5HklaEPgwH7wSNOMNFTEieEMIw8o7u+xcr60+cGnEno05xxCx5z1y2ro9TDtxi
xWs8TVzzRfFFPFvBtCJ7k1aZxu3Kv867avb9dLCr8ty7fU+1uqFqV88/S8bfOS9XeruWuRlawJ06
6mNQ1cvMj57P9C89RadIuw+Ja6cTccQf8B+ExVrMZ8b61+bDUI4n6q3f1PZw2gpfowp8Mjf1pWY3
UG6Jgpt3Rxn0R2qauMsHUXeWezrqesSpjxnSeifiFeVSVrJu4TZpWpADz1W7xitWil+Kev6sO8He
w3b9J39LPIq7Zzfq14z82Znpl2bjtMT47KJ9TkG26CCYeSvJz5Ev5z0P5XAxcE5Mamb0Nh6P+T0t
+dLGgAswxo7PKTjpHKgLFOHpDGsGHPxTRcqghZx+L1EZdwseI6iwBD7tzfSkQhfXYaV5C2Tyn7/y
NMZ+8esnIdqSxjUONAArP+s681wXNA824WyVJaMPTneyJ54LstOmwi3hku65bsuEppxbnGhxhBTO
ck3jfR3eTgfAC1af/su6FPHlQIOeYDWrnCFXzlSJqEGjmBhRUtLPSQ6S3V623ug9uV+NllwuLyHr
W/ZtQO+jSTmOkT8q17TmSHi/pglsXKAFZLkeE3borsNGgq1SgutTl1F/JNwKVFrGx8mebn7OZhoV
+v/DSP3ljjobPwf5haUJo+HYZeX4pkVVs2pAkEHZW0L/USRFgMTdbgrKUVAFYgDpBatsEpBkNtay
bxTyhUOYZSpQwTzFD4b9bP7iP+ooZZnGfxL3JFYmaQ8i9BviL/G/zLgfvm5TK/voyZO7/BZyAzy4
ixUe2x2SonSlzTf3cEJpAkbjo0CdFoKxGWqKNtmoLlGYPuj9YA60kNzBvo1dW7Panm+sh3U2cq/y
XzcCkMbPCExDfgC1FiCo18vPk1Y4bdz6AUB1Rn7H0Lp5H19CCUGJsd18ckiNsnKLV+c/0NcCold6
N4QMD2QvGwseK1v4Tm5z6BQZM0d9Z2AJDQPGsOxKsPMZP1j8i88RWTHAfQF4gZYA5zTSDub2QDia
/ELfWilsMbThi1zVFVsKsZh/C5ff95etrI47BkNvhkMC12/rcuRNTRCleyiln4fkfa+5R9NgxLtd
tBtKTyQaj/56XRocecnhD9Yovt5+TSJe6tV/DA+wfpnpKcEpOKCQCaMyBGj252Thd9LZbJ3O+JrJ
kdtZAqhNqAQGhVpP4qBXW3eieIHxJZkiS/SVbGdZMZTIvIBJVKDLjB77C3dHnrTINIazxjr1SZBW
QOoyB4kNbk92D/oE90kLW/R3Q4IdaLc7cW6lY1wzigesv4p7tPEnrTZ+bE1406vDp24PrL+sVwdO
T6AWt1tC0kiTSl3Ju80awA3P8FU3QxznP9hlSd+9Q/uvGZz4g1wZOpiJvtsFkKGky6S/n+6yL1Rt
qRlwalnbIvt4+lLyFxr1Ju0+qE+tSFlgGY/43VcVhHUtY7N3FMwAyeY/+42BkmgfOThCeWfzRJTQ
1ctBG78WeIKICrVg0b0e8Wfnv2vFQPX80jB2LaXGwyoqisRGewfK1JNAzqnm24sB05Nmq1cslEpi
HkJu9U8T+w8r1EfCG11S/LxTbkDW2XzyhVq2NcghHRKaiaT3Gxe1JlQP2WL+X9Z4cOwTuDhSasG/
yUkOEdC/9bEJd/YH96UKWBelTjxdA6MQ8N7RnJDJaDWJmnFST1x8W1qrq9zzOqiUu7MQVwV9eOX3
f3LPskVFIicF8BtQ2chh9iaqR2b00UfPQNyJEciNCCXUejSsFhUjXlrg6V0XktBZgyJlAOL1rFgq
RYJcVv25wwBTtqBzNZMP1WMGuVOV+4zj1HKYmdUH/4SBAF7nemH4rCQI+lh2dBSAmwvu64nqs8yk
DjD1qIgGfwyinkrHKUJjl1TLtFyOeT4s7493S7lBwOJ2Ns+FfkaOyiorfhA9Jm8gmcC7PuIXtcHu
LP+73m7Qw/Er/ZYutvPbOI1QdPruDJtt2crYBeTz6xu90dwmqmiAiUjZ0tE5Hi1185RFMZZh5QMl
t6MiFxlBGftWpTO6kOYwYoQx+DfwyoiCpGP4VnoLTAOAx7ItZ3P0wLJNaj9F4nL3BvKtEINUxy76
Xp2jqNur+Zk5NCNAnjTSlq535zIp0wFJCZaS/VyhFp68DyAmk8fCT0pXs/cBPHW7+ACOopvT3yxS
6iJX+uYo8lCT8YNAS9yA3Iva5ZYGnGYHy80uYl4WMXYX6WJFAtwcQ33zIie0G1BbDrU65hGXGlWL
VFJf79pahQbAalUr2lD6Ai5Pks7pZ4StMr1LamV4q+1BofALsIVFAcf+Oc8dXtYleUKF97Glf2pX
wb/8wXgY/5EdbmIMAmzqM7QX0K0ZcHjmh4y6QGLETkhHy+ipffBV2LIrC2CK1ERf0in8g8fX+N8j
QZWx0ozU0mJrEa0Km2dSRCk8Oan8m3CMNVIU8g3kUGJZ8ktw04CtbaJ+y4VVExyHSrvYO5adyo//
29SyGlHxyfGGU2ESHcZwBEfodghrLWE/rTIbFlch8iBRK/gYogzttvCfhTLpjiXre6Kw/wCMYdyo
/ro/8IgOxuICJpQxLFWY+Zj57MlUr6OCoqtDjx3HT2GHfTHshoKtoNvPUxDNma/M28kt4D7VfT5s
+cmOoMD1AbDIsmAcSjtIqKANUjXLE04P2Vzb8YeNLYMYyyNhPwPI+UJ5EOaRbtZ8k6xGvy4wet20
ukeIhhZT+xtiwgZ0YjhnLW8aF4nHLU0eLpVciziCmaou3axwJeNYdsWQXazU/f3PHLLfJWSm+jQW
K32DdLKpFYiupwWDnBZVGQ0UqeQAQQNWXGElbh+/uKsCqkBrSEaPENX/FlX4oZQNvaL3+sTXO78x
t+yomt/dronwtTnWHk4daTOf+kHMfIZFvkFmyd+xldR+rz7FtMZSTQpEgAnX8WWNVaOmWYDnAhPC
dSMG83H0DuP7SWZPrF23+lYclnLKqlfXKiw/xovhd+WF2uyIlnWJNY9+69/mA17Aj5wyZ+jrVIzR
sBrsylSqmh4KHc+ZpKXE6pYH1Q1sS3hEzKrmjCRPFXaU0jPeyCHNbWuZMxSij9yESJR76TzUX/se
UD+mJgMVj35Mw6W5lTnwTVvIJFOlKqGRBg4EbvavxgecLtCYgvpB9wygDhNHh77HUSUmRSoD2iv2
F4nY6mXjXfHKq5C1iQqP9b4dQL7HHtlUbDIbzv0IGIJCZ81fZTsvmy3vWkDdztdYcLWzGoLtl1rf
REeCrP2DbMeit4cZuLULI5LNQYo9rGcKWzpRVFat6rjzl5vT7VKoq4IUjHKo6PWSeK1eeybJZs6Z
P4zImM0ZuuWxRtpXWJcwWzH32rr5fxBVrhu6FEcmiGw2kgG1/Uas6DwA0ae37ceSbgBkNkvnUu7m
+2KYhN1Wvu0DSV1XYPuvt2dF5bkiveRQL/y8/46911LgGN2XvGbjJwFzhu6X6SQdWBraH1GINrK6
3zJcSRY9jpPBayN1rmnX3BQ8gr4ljtr30tyBwgVSJ6kCgFaQHB04HGzooJ8A5+MKYfN6yA/C92DN
+ldLyxaO49ZJv5IYcOiTvsXg4MY1r0QNn48Xh1ZxQXmSHOZeMNeJZyUKNIv9f+a8UIi9CjadOO8k
QSpOA2kC85YRjKBeQp8Pjn9P9veT3d2IDJwPleJr8TxcrJmuVZRlNx5zPwaZPHtpUaq9pQbdV8ZC
VQRQpcDROhABTR4hqMcfzgHBhWQ6fwpSr51Sx9da4gMKWMPnGCfdq+j7ziXpcBngS8VAcdM+KqWN
2nJXMYfWVuDUTH3jZ+tCCacewolEwxkuyQ8WeSxo6wbvuZxhVF3IkWT7ukb9MErvoBhxnCX70TD0
6PrrE3zB/6b51Q7HNiRLwmSMEaa0p4nXZhmHP74nAS9Q4yYHgoBPmatKZbRGYrbrzc/FFCBBw2VF
EdODEx6feAx7/0HMEmnms1RQ32P40rwTgoLOk933LWzLEqJqETMKKBrtH5KBydZ9gWwjsyd117vh
O+zo1USgnV5kVXK0Ph/vXDxIzalTozOAnfTI4hti92Rj9Eb6WVJMgkEvdXT17KHuyx3+BDmr+P6N
6O6xwbm41dfH452z4epv/RfsO+AKRKIm17LbnNN74EQWa8Eez5aDENw54R8KCQ5/bKMXngpGMfNy
r1aYVHki0GFalKowFtU/efVtenuez+qbZfgCDdYeSFAFLFAFswHYirny7xOPmrViLAfebaZXONTc
Nx2ZjCnL7I2TZRoErplWMQaGGWtmmG2aB7nxDY7YNs3nir+qipXCkd6X7aXGqjjOHbGvWyG2qOS+
pTds3qRU1ekPgp6HhZnvHQRvUD8DSjW8qrWvf9B9Q1CBLagjTlD46inypIBrANCmMS/mwP663Seq
h1WWS4TFBQYq6f7zHFu6VWWFuGDNd4nW1fHxCxG8c7TZNJvwfiG1ozHNhLeMC42QUjcRaBkwNtEE
EE/uMhlVDxDsiV4AF4Pvo8xMRk5EQoUW1mkDAah+phVFuOk3s4fgWM8PWgvrGqqk8Dkc0aDhtMaO
rPloQMeF7CCz+sFQCwRlK9JKV4mecTAAEC9Cw9mtxhubEFwUwBF7eE2kfEnDEtcycYKNPfJC+nOs
18Xf3CJqk07kPKTvOuj6mhnjU10JGAm2ntPU/u6LmTSj4jgpl6YoVVSZShJ5z97pdDFNSYs7uKDH
Duq6SCcDX4ZiViclMtDMolNAMVlkvTopsKkiVv0rvzJeHxFQCWMsTTbD/iqxo+zrgPPhXQtQQNRu
YOyq5xRarMf9yqMjQGRa9iItfP+s/Zk+PA/cDyCnSVj0m9qekMGAedXALf7rPwYkvV6Sg/hxjxE4
XMeHtuer9JS97cjf8lzmD9snzKFcgkZLf7cJte2lTrK67kW83cppUvqRcprmN2A0SsLt8eV4ti0S
jE5k7+MKCCt95cMVt4r3O7Rp49Utx6yyF+KF9luZAtNLQvBjovFoDQbr5UzvIBsJRwMBo0m9Q8kK
PGG5TC48HMC44xNXBJ0mzAEw4dDAsWJBhodvi+X9LaYN6hUI1+Kol9Yt/yhE+K23mzJjDJOkOyo4
rDvqQTptrTNxfqTTPGqw3MWTwIpAOeCiKbZgi1GLR87ouXj/lsBF4E4FpA9MBge8Xb4FNdp7AbKc
Sf0s+QZQd82ZPA7LsAo1PmDjbZYada/+EMNfW0C3w4xbi7x5F/Vbgzk991hbVZwwT29+7Pj56h0N
0cN6Vmkow6sd6i5ETgQProBz4qJHY/mBvU/2f3zGPgL0D9kPZFIe/T7YLObJp4Xa0Aths5hPoduP
udDNYJT2qgdfbfwVSYngr4OgKZSuslvCpsv81CYBR8s/5Xsa6TKIrLtzr5JFg77ZS29TAoHghmGU
oOR2cuNoFEQXufiHzLtp68nv+e/nS5l9uSt/c/rZDmRTVICu1hG393nrrSLnHixARqfU+E1S+VYc
S5FHYyiACSeTscywAmr4r9waoDh7hAsonRFAhqlxyHQB8psFFYS/bM7ksAZNKBayHVVcTMbtMn9D
0wA6fgwVd1wUY+OzyJ+qWUY0ufi/JcpSlFdfgexyEHSY7uT4H9a1ij1pSC9x5Tuk9DIDdsfToIC/
l1y+BuJtOMKVq07Lk8cyOMY7M5+Kj2JdFkVhbLMDcsfP2k1F0Jh0ONAieaYSAgGD+cbioYAAiHgk
LtKNBM0Ub1r1uM5scMdwR9G83aXhapJxr9hUB6JdvnZ40iw+aywjoiXj0RRh1Bn21dIytaCnEA8s
b6Q+k/lLxPmuLuqSYsFUBur3+uHLMzIMmlopT6N5l31RfiSXtP3w2lUBf+FZVl2sWViOEROM/1sV
Uo2TX2YxQtBxbUdhBOAsXffvKLGOfw9dbF/8JNsPfcQC2A9HSJymE+ADKzceJ+xrEPBxaW05QL2v
qCsRZ+avBjqVt94YufwkGyyYmvVZD5xZ5lI4P6e4BhCnM71zZIDiHaffx7XZ9C4LQizCv6oJKtRQ
AS8Wn1YmYwadm452axVbI45shKWY49KYr90EfiPKZOXfBQ580k3Hr9ZBjCwP3+XlHhpPCioKRTAp
V8MTHqDlgbdlqxItZLvvfuGjCV0WyKdjs6YJgL7u3Eg/7nm8sXKgsK/lEDtuuFFt7V2qs1zjUTta
+664p4RCnST6KVczHlpCeHujenQ0bV3O6+E5lIRm3+E5Cr0Y40/9g4Fzn/HUabl0m6dDrSXXtBue
3HlbEbGHsUOFLohpTDpJgoCr90pCzJtFrvUnyVe73zeAMpT1eB5vsJlF1HWgcWHD82eEXft0imQb
eevEbvS/yiUd/mMEwFiRm+3Sw2BxsJqsDMwZGn4ql6Jl1iNNaHGGuxxGrBE/QZEjMbZoYqHu4kg2
7ndxd8+fpSzs4xqnYGg5poQQJ15FQLZXe4rl80eklYid8UTPAnaYXrhwp1lm+162GeNqQM2Wvpwi
E7s+1Qf8ChucKezn8XEUXFuloWC9jRdq3ZOKE7JKypaZ+b/E/qP2LxnjtvowTQFUXlU7Wf8yfSjW
nzz8nIueNCV85CLJFYi40TvJ203T9KWm71kJRHHLunOjcMl/VpHwC7LmWTVgmA0cWhfgcw7iCE/0
XWS+kg8iDe5fZ4JJG255H59+3AwpgXmhUHKuhA2wGdEQISW+CFq/ULs4+RMq5IQiOWU8Si8mUCnm
skDhdcfIZL1OAZ5Clx/7DTBpMftOcrG0C3Gjo/1SHaNRPNvWbea6C3IgTCKJXYSfCjOeaRdMp2/I
F12Qnn2+jSwJHUoPGXo7pqO/qYkGhU19mOvsEy1s4E/A8+Zot7TKF9bqOQrNSZB25kzzirl6cLD2
S+EXlkCG0oKhQILJwty/fy5JwXFAf3HqwH3+Hpz75igN1DvvHzzDjqpumvozAk2IkGM3A2pvK2Wc
ohvssoCj/mPuZL3Lqqno6xdH7AtKzg+mZ7GC6WslXwx9fAoo6IjBtI95e4ss3pObH9NEU4SkAzA3
XphDp3AdKqLXqRW5d98xXjzn/DTLDDzfyy9254COZgxioVXBLl/uyO17GhwMP3rZ44k1Xqn6bzaS
K3EdVpr90uoTj3xr/2PHDEPPaoF0xc9u2R0N373nJaz8uUca03VJvl2DRiOKTpLQfthLw80o1S/P
78lwUpECvGXzQa3zX70H0uUPpbVUam8P8o4Tm9SFdGGwYpvUJKX32Os6T0XlFlYc719k/n/R3FSm
h5DmKrj7KXzOgjcY2Dgwj3uApuqRuLsh8zKy8ocdVDbqDXC+UMMavQ5BQme+pYzuhKdb0vsW8Rzj
Lqncsyvd612090qSgG7kibym2aaGP/T1/g653wx612bGWhPCe9AWMJvEGrmYFz1BvBwrqqq/SZhd
B1f6x7p0HkY135OjY0xU+b0H1X5KinxfRz1smy2aDIuiNZ/RR2PoUVvHTr35slnZZ27wfPHiYhuB
aUe5FDOwcuKEUtHNWRrQ+VDR+cgMxRMjtFE5lL44pQ4Hrfkymh5B0OgDO/FDJS4kggFETWWmkrBG
7f1oSKZrRakUo66nu+VWSb70+RLKH5RXbAB7p4AuL4kjNtDG15QmtqHjoQl+/hM3H9J0s47F5vqU
EYlrSBvmKAzkowf93tIfVbhadhK0jAOY/y+XZRT6cI6F9BH1UDIjRLdMUz4gdU2P5aSVrM3TfAK5
kr9i2F8h+hBjsXasdtxb5A8TiX66NdqitPK7tLo6D7uvxdO4DCehPCLm3ua9FYEAxhi3V+H0IRwA
/ttWvEEh+wrPC86pljdjh8LvPUxp8c8szP4Ft6t7nTLyjPffwl7H3lfhjOClGBDO7j4e6MLx9hYa
mft5H0bQGf5TsKrqt88qB6+SF1eyYl7XC0XG2U/xC+ov0TKrHKiaFX9GF1sBOewv0ImRNGUjCyaK
uus6Hwjrg69a6fHI3SFH70z97h5PEwvxOaqK5eC2qjU3f4i+qs3TEFAkfh14YHy44SbXajr8MsPq
LK2s6UcZboaA3zPnMn/XA38wwl23AaU0QnEXV4wpKOSTjKcfhFpt5OiEtMMwZjbbGF/bWs1o8RZl
DNbHkjCG0SdO7+9s8iXDSPyx8rECR3gHnaB4fjQlvzm3TX7V/sVVjAO7AE2xPtMZp3CEMUHV86mR
2X2la5WESOW84mAQuG1JPgVhtLFEX4XXT+ycHh9kmmI9hc6vPCbWlrx4FdJev6C0iVavYPYR9aZu
tf5iTI4n+Mq8ttlwAbne/fo/7Nm5Z0YWOReSkce4d9WwKR1SqbvHTliS0gwPJHTVRrPIyZ3bK6yA
lpyoBiTFb6fQpzV9Bo4U845uaVlinjFDUyU6nrpX9032HsTsppGx11JoB8mua6JEZotdMyVcK9oV
ff3hZD1ZXIELmjjv/WGTaYpORBA2dZSPzC121HhiNXfwCHfRD0V8n2s4VnlXbjGIUYgkYjTUcUBa
xkcccXIdb5D5gYXHbx0xjkodmJifGI+so67hnJughpeY92yAzdqzzB+I8KhvlmkRFpRgZKdiw0M5
ir+XjTglee9uiVUkPCpLZDVGsnihprFc3DvvbIWmJJzXz82g5YNK468JC3739h6+26n0y7BYIDYN
s40I6JMePfgniihr0tsgm87jZzDuGXxeJCuIR+NiUxMyCrJPxZ4KD97/gsiJtFdDgwmE2zyPbUxY
a5rA3bQVEzeWpez9OV22gBVstbZq80lQxYb8cXXzKgpbeFLnQzKmGvnu4G3/1he+Vu/TKHiBgmfz
qVd6X+0ifjIOo/4tquzNWeo31Ou1ZcO3Dc5WQJYOp9J1kMn9AoPhO1YQwoKxaOy5hFwjifKNf/7Q
XmL0vJ2u0mfM3qO0Wv2P6bcfTGj0VZxQxBKYNGaIPoxbTpkmFUXTxSR+gXNeJ9S7WvCECwhdW0mV
zAP2Wqh5eOAu8cGoIivQrXxREfI9AnniVEBqOk5Nznw+deASLxrHtI8XKwY4wN9vohqeT+5C2m5e
H+8k9NkIeGyN3Trrtu+YUb895hvitRi2eBquptqcIdc/hbXG+HxwjCXz3H5TjhbfVAUA4CA31KEd
euZN5MwVZmpyVGaQqM/48h2PXfkUABsCZUbJjrwVRRUJAiMyxnEzv5Mbguhyq5AvEreg65Gt1VMW
o3E10pfuCMn0mTV0irtzzm6ANiqf4h3U7UwnesYXTYJS5UmsgiTLr6OAqFyQ5cmTQVRk70BCoKeH
aTQaK8Pa1i7hyouWnwJ18BdMj/wT8dsZ4EyTIM/+WTAYABiTYDrBQfuG6WV6lnGap6SrflJBQ8eJ
6sG80/DCPiSyITKIppQgYUIJq2WVYbrsMBIvWVtWu6mKmCO2BofyCcrGOQR/c6UuXnyX2CQjEIvF
sBfAirAN91JPTK2NM1WIwGt6fLq9Fs8rUonyZAZGsLkMMSxnxbHC0PncHVcnOHQ58WWGTljXGMjY
ykGS9Bvw7HNyhfCDNFeKovYYSZpnltqJ8DyuuYNDUujmWTSWihwGYqGHji6ZY1j6KcgBvnwQd0L2
RvTAsnARolLv3clGyd9TZPgkT9TBFiJu1KG3EZtuCvsqVk5rfCy8KMsVx/3qs2G/e7cBqeZRqIF6
dsiWFijAnnEb9ZC2H8sbmVSyZqOjgBRyO0hCT0NPFczPP1EOoiIC13zmEHGs5rsU21P4m7EemS3a
l3r+hUp4m0uMFOR+IMLsJtVStG5D1hldz5AU7hyz/LuUSxDfQ+EqJdWBZkhI27zrHVqYXJ5UK/PZ
3LZgSognSXfmODROXWkFBLXKDs7hIMt89kqMTg0FSqHeK+/6hZQibX2LgwqBJMoYju3QxUk6LvKG
RVJO1FuVyD0KEsu6+yIA/E0Wz2WCFTpbKYpZIM+x/SGiUkpp8XxHeLVlwJfXDQ2Y7aJE0Rq+cnrc
5yLvwdVTMz24TdERa+k2jKvhP2MNJcsgSL//2hFZu32Hwy6mHcueSAEHXf+1PLgWtGQMj63aYCOr
jbNIPfMyLQKEN0GlHL5MvL0W0XqaR7JS3DlePRPZbcGslnfZDgZgb19rqrivKvmXBFNnAAnk5wZU
mM8axddQHaKAG+fFMC1N4Bd1PbrgDsToBwTwUctkxdGmWfWXLDAPbvJbO0Q/ekbvWgWfcrus8ol2
YR8C10LbM/d4BWDqIYpwQ1KjjEcyIOGJmDcJDDk+BUyrT3DWavr6dTx+J7yr8/RIxI1e7W7xlGCs
c1cTE4Mledco4vaE7PCVgzqminUnY+CLMw/irLjQEdvCYgiMBKvdqcSPGshVKJ1OXfED89cvMBdx
foHWWianxY5iw3gBhvOYoTFfQO2ac2KUXkw6aINbPCpQHDGAOtoa8U9OF7EOPi5qIXDd3jXGKxA1
mCmpM3rvHK5YS38Py7vCv6NDCcyLxk0SH3atujVOq24+ZKVv/3YOvHLmcFN8ugEVT7R+E1fLX7Ar
qbKzNs/ql+V6SVd82U67F/i7hE/pq/pWkwBQxOJwqRqBQ67FgYERMHHx5AoP57SGmVvBydZQodaV
QTl+k1+CU/4jLdV7fWuL8u8MbvAt4hJepWBxmLXq/6CqNurpq5F4E4vWKLJVVqRqDq9oMx6SfThy
+5fjr5A4F3ylSfIICKpOBBn91rbhZjVjrOPTpue5yG+hwm93BvknbGcUaJ/ak1/LQohbRBfmlVFH
/08KSRXwA0UX0e4IUTUQ1pVb8Zkfoh9fspXFFoTaJ8sOpo1BahpNSXoYcgJpvURqFdosBYNzW7sU
Ppjrk+7F40TW+77+KlxGUu0I2tLopoDkjeloSmPqFbH9ligy2T4emSeyTuzo6htT9fSS/jABgi1b
yzp36OPQNOJzNRA5nWSMsineJhyrnyfHPZuZTupQc49ZFgBjcRCztBPH+AD2Fq3GPa3qQkLEnfX6
W0Ckvo1Ov2wWXsSZ0qwdJBo4UEQTyoepVBliMQYj+xZxo+b2ZOOL6jJUaG8sek4ajMgwhef0/YcK
SVBs9GhJBgv6mUN6s7Y31NQkMgtg2X+ggvtvBlbqNKC1KoZb3qACwmzqSu12Yalpz3Ctf36xge++
sGh3d7hj6b8wACvotLQ5el5okBVV2DQVsoW7g2Hx8fe/vSyY/Thfgaw5ba4IEO8uyjkgbVCdNc/d
V6LE90IZFBF4SNtSWT3VOoqD8CGpc611rC37DPN3l3pFgSfmOGy9lM0aP7w/n7EJ4lgPu+4/WF1J
yjMhha23Kv1V4rdCP/KX0XNbKg3bGKcoyL/a8wX38k+h3fvdKY+ynJC3/dyTUWrJZEFza1mQe/iY
PG5DivgDqabINrOGOp4IV7t0qbDMuePybZH2osa9JJLKUpRO4dJwhHTNXt+lOlwnmA2x13750k0r
kVPxiEIb9gakjevhnNUwO5Ls95Ex1o3sRCDLMUnbk9bcb5p+/eALXHPQSeYfiPwirF5XFnSBSDdD
J87AABsfCdovB7xQ4tH7M0BqMLAbPw6Q0n/5Q93lKNMRCFKNin20mpm1fUN2V/FxfJi1yq87Wjm5
nE92csh8W3XaFB4CUr/M4hlmLjwCHcLqk4apO+LcPovPCecIc227kdlbf0wlHHrA4zaR28QIgnx6
AWv1cD324u/umm5o2tYwuQ7686UDf5mMVfpg+WdPtUrU582o7FrabowAweW2d9Z7z4IfOji5NjKh
AmKItH0x2uRwkBrrRaMhMgC2LDgYWzGijWVms1BCAiggRR26l5ZJZ0oQd4U0m2p7toaWCxS9//VY
JgrQP/3VOMEZ7Si1s+faK+Bra9Nda3aNf8G9hPpFz35c9Z9S2WX3k+RJwWIVHQs7Y/em5/YVfZHL
/qsCKmEqXqj0azCf2uKr2SsEPA5kcJE045mKobvFZtK4zxKvYMSdPh7mZu5OWJsIoJuq8QriZyDp
xUXMm1mJmAhrnNY24Vamp1dQgMxsyNdv8lfdMwLmQcmeullt6pLU4CAWqsxrtPLROQWFi4K0WQhP
QmyyuCYtYPV2HwzCoGNK4fCdU0uTjhbrwBSXN6DebEsF1CchtNd189mKvVXYPB0Uy5B/UyF6FV8p
z07aJHCVN5BosRgSlRVuFWu7/qNgSOApEvBnA5B95e7rgo+MSBuqYizLOmajaEM4birvLpv3/jz+
fI/qG29ENeLPu33pazAPCz/4sWFlBqBdpI0e23dlEHsM0zzWMVthYpO49/ZpKw27UxFBYONVn2sP
7CCYO2J/RRe11Ovj+K6o1RCHpS6FSBBCRM8iccM9mSp7GkNdTHIr59t8xXC5gHQOa6F/aZk+xIWr
daLaXztN/0s4+5rcOo34uGLatWjovdp8pVhyKN0b/sZeYH6c0z2bNjVDThf7/puBcxEYScgLb4Th
cf6tBkCQzcThCiCwbKcEy8dZmSceLJjmrPms4pG9GvLAnkbtRtMgYVLrj9qY2BaDSdvAA/1a0J4q
c/A06GeaLDcMBEGiqCFJDg3/hvuXSyxGAxiJh9cQ9g+DUeSn2L92nSiPAFANE3B12awD0etNkNVN
+nqNYEP9bwGqYG0Jm1DBcnEaE7rnQGRs/pbzZKhROPGGQYDps/BcMCPYWI9L6XCHXemBOv92SrkA
BmlWWFr4R+uRKHrjDkyGnKaux25f/bWWjVdiwB2weEF8dktSkwTQGU1aw7uhYWG1oKUFTxZ+wzsM
LEL+0pS6dqMCCZ6TU2LIa5G/bCh+u6keuEqLs6taicYNjrl+zwzeKfjOorWgPiiU4EnwTXTGrtSm
DWSylX3VaRRQ68mKSBYKzRMnXmdX0KakpMz84W0fZuyybnIJTREWhToXry2vsGcnjaWQhceodCrw
yvRgQDT+mZpEQMGMz42dK65ibzk8o8xNd+hQDSSeTPjoIDOUqcGrIvKEZtjbPKEzTPaPP4Vw4SYM
keQQbd04pbEGMTZzzfERbWgK/R5p2b4jw8/vbACEPPwVekutX8DfK6kk45IbTXMrBr9HYp80K1+5
JxYcjosmCnIEzZOTPtFKmLRXkpEvekUNEqcAZKN2efcGgCNh19juN1g6WDzG7O8HhQhOgxHsmd68
iPtlk6sCRt2vZyt4sCkd1eCXawvq1wBRLCZbg0lreYFosfb95dcMPwJZUd/bH1tNMdd6XxAiKLSO
+Rp58UEdk6BtW2pkr9+MRBhCtlLpdL68ACLaPbUo4Tyi0OGo6rTYIalfNyOVo0zPS6zwNVXQc9pK
ZErOGeIIV6UrOOTa4OgJvmoBP3b/S7nmVAS66TbtAHCcuep64bjqQitzbaGD2kF0anWiwApVTCGq
a/tPrhIB/FCDp+0jfqepvcC2z8+YqZarVscaxirPYRjwfOMd3Hi9y6He7HPHpTdOY93NLloz5yFF
S24rkguyUGkyH6JvQ1xVaTk/t6O6UhCKz6o+Pe79jKtjfzSkIrUZTTkUzJr83JPCtZkEOTrpFVj7
A7Df15y4LKew/0kh/uL8ID4o6JYcar6xIvB3W4MwpsSY6NyIUmH4TolF7tdPnZBeyp2t7JAHo9st
ES9/7Pzpt6Y1kgoJaB7RT1KSKTS0QO9/ndpm1x+AVpcqRAstB9+m6C02NDnAyqXtlczefwA/blay
HmwcnPeEp9YqIENyoSyyiIi7WLH0w9OMh1kq9bxPaBx8IhWNKexbTYqKrqaGYIhVPDkaon5jhPqb
jc8GaUl1/9fclwX6loY8COC0QfW7wO0qxowEMwib0MogkttHZ3qXJyeMlu6bhrhcH8KpzrNeeDcW
/KSeQxEG58fnfYS2jANaiJaOnuTyPfDNHvbx8ERnMTNPKJFQru5NKdofwIOduu9MzcZVv3m8KiPH
vfDXXHN8H5tqAZ4h0SA6ohrt4tZGCUfG4sFKwpgWNQKrl7c051v2s0FoI9mvZ1DJXcY1z65mHhwz
VV16ZbP+bLnswtv+xmM0Mf2y+xVHgKr+lQSbr7q4MeZY+mJGB7DbZMJEb+37Onpf4Elp7LgWq2pJ
FWdJ9hgV2Z4EBgKCs/ovxPf3HTnfFOZ5qmN3wHLnUVIX7Z0QMU7jl3+5PNJ0mZIDGzWa2TbLIrUJ
P+/RWT1Cdtv0usFsDS0vjMW2Sco/VJupR+rD8YvlbbRfHlgc+as6myb9uXP1fi/9ap1VukwUL8Si
PkE+QykaWVNVlbs0vXJClY1gfOElNrz+wFVNmkz23UNJfeY1IARRmM/WH+O6uqexiUhwB1CrzBmK
nPSYidWNMebh+juumnN9DiX2BG0kRYi699/UkjaD1YnZ2j1uTJZwSA5yTh0Idyu6YjjQISDA7rkp
jHETXR61ZlxGilYzxFDhnaay0BdeZjkT55Fe3rWOM+WF6qLPqjRnVj+jmjme302KjffN4G14E+0K
3MaU8GtddnpFcoE0qzlKXPEtOLxBP6+B8qZEl+r7GuRIzeCtVCUqWCc3FmSVVMN9Ov5LqrjTpvyY
NDBI2Sec9BqvC4aHhOSnKfJotGY28w00hGhHvweTcH+hDEq1TzQBupLuPqY9xjEjKIkG3ADgHbXo
Iyihr2uqk4Dqj3cGmWwpZ65AO2So9ihhZQw0I5Mf2wgB15mUM/sg/yj00gz8lspY5txYoeJFlLys
tXjJQpEwATcUpNmzv6TpP3Gi2q23yi8sYPQhAE3co+ABy9V5Wvo0/ldt+8YOLJPfzF2iNEuXQipD
fw8wJn2UThhfiZA0ymVMXMd7JMNzl19kYmIyjSULXrwHe2Arb54go6fRrnFLBMyvcxljBa/xJSRk
4RZAyMXB/RaFB/262K8v+lPYxb9zDSLT1HuV7ba5q4MR1lOGREnjLL1NO8e5Ej/zudyb1tJG71+1
XKjk1YQC+ZanW8eZoEyoqLBJZmnErMFUli9P7Hb9KDRMqaGkq4yDuq5tVRDZDwHornCFcRgD4Ugu
QdgHV2lKZKQyhM9WyN2iaFYpplGdsVZDucdzEzpGkIqN+E+1bAtnqukCXObqS5k6CUWcycoz08fY
j/GRTmSC5gVXTpIZiyyWf8ZaCyVfNC1xJ1JptChB8oEPi8qm9fZcB/223lfL3UAUcSZPwBtKhWxu
8BA1Zo5l7wojZi/wN59XhBNObUg8rhZ63Q+Jnlin5WO88hViJypP6VXOaIHZ4xS9JFsWdZqFF3cT
nOmRDBm2CZQGA/rx355I7T1ZHJP6qxbV/q8/hbCbqr+W9Tfx1VmNTStSB5i7vPxiAU6hLqqtcJto
aQI2YUQyVzJ4Ou1uOdcRhTMOfcN3W1mirP2rvelkTBMyZGL17q6HuwdEn6XSBV4RkJtpMnCpES2l
3crUmAG6TxrlaU/PgCjBJIpWlCFmLyweADELYVhPBAZUIMxwSnTQq244PLqweAlyWLB2J5tyTDCn
qt5mRvDHCjmSw3ClvNmILQDa2OWt+C49eV7IZ+NguvOmdgoSGp6XZLU+DEbT2BQBODupDZ3vgzvQ
mifpxBlks3ThOE++lF1B0UA0t0hC6yst2RG5l9hFo/3X/sNNZupQYJUdJVikNjRFpbZzSwdlPiFu
w57mdLAnPqXeqLpX0pSDClx0uanauQqnR2y5P12BCFeDboFSDdqy0g4wl7s9cAmENUl0pAitqlpZ
rYre9FVKkEVkQGGdic8G2qHY7vEsQxbQNEK6Zp+oikrcOnB6M+QESxnHTs4g6auJFzBlRyY6b+t2
0LlAioGftYsd+ot53HpXO71IjiISGK2nCVv1iRpYOCtSrd2Jvgvkqe2gEYq3m2meN0uW8OwR3gIw
EEONLSKNE/T59pZTuyYvB+1JjsHRQfA1uB4E7owlJ3hfW/9qONwk8AJ0xCQqu36pQ5/gGmFHlNtF
bm6WZulnM4mTn0J+ssEw7D2IajsQI6wRnzTqbCn3vmcOfQHRb3EUGYtY+5VpTfq3/24mb89yDRjs
rfe0Gz/V2jQ6CN3zriaq5RtbPITfhLbBTKOFgaqrqqED5RDvC1b3ac+fgheDZlIxybmRTMUIDHFk
riY2czgT9cEHvFYUTpub/ySrUgC2n2osqxHwAYLsI+NXkn7g8X7JZcCgl7L6bVMmIWn0xKxPLThq
RbXPgmkB8xC1pWMoefVGKVXBNaqPm0B2NNd/0XpXjDSZCJQvVIuZZq4eILl19AsT2s/6ywhDFHBA
kYtmQ2sZqH43XdukpepGk5qaGJvQ0Yl7+gIX4VWxK64entgqNv6gODk50gFVhY7PhjsIwcJ2BjPn
9Aa6vmt5l8ZuJFlVzS+aZM6hkZtcJRAufB+Xr/1rldiS+JVXc3FbmnQOiookzMInLsTnOOc5MtaS
lp9nVG/8Q48RqgQNJ9WGFXxu5ImHofJqfIEtW0D589O2YLknaWNJVajFwn+KQTVf+a+vv7wSm6Wg
+yeEt372fTijF1P+QNR82sPGpPfNn7MULK0c2ILc2ljtzqB2JFsIqyGPTwdxbackW6XLGK0pJ3yE
sv5uzLan71pIFdBKkTAaqSfSDXIqwiXQwOt+baNcUgkRNp28p34wx6Oh1ig+F5rf4e++CkVmy/Rt
795bab+4HKM2xJA+QVPgVqTEckZIhPV8LsSiN7+rUc7zCLr8D71ceuHwCapVhClt93Ry/MAA2CPv
mZtMJS36wAG+Tz71DEQ0SBiOz/1CVf9etJ45l0dS+Fl9egHDFSYtIBSiXmTND1j8bFtSzuan9Nec
/5AHuw7Hmab1V4r1TWKnoRsDYgnB+vKnQ21Rh2w0npuqhoYDn8jGkcEzNHYKAPN/iU/cSpv6ULah
O1f+z55hMkc0teew5Piif5H5g4Cm9HvBJfQs7/lrkEun95mh52cTBlB4QMHEmtWes6ysh6uJh3V5
g92Nurl8Qz9UktPraSqKTHdx0AM9X6lEX6KHs2TqNK17305rr4Gvbj8iUB+0aE4IWTfNvAnsNWqY
fiLlZdioPrGmP+AodJxQhBm3IM5AWmH6wSFYKrg5lXdUy6AyqRzxU1nbhWWqFD59CbL9Fn+bXOmy
LGDq9sglhyHMaZoloJNAST6TKzTamRZ1bES/ayXitSsIVbPaoR2b8LMclJDOup3gU/jDo/8B3CdB
bXw2/s9GSeIzr8wy+rlmqm1XsguifYjBjPnbijSVVMZd7wvGqTyMO2MQukwXUP979pqzWg3tZiCY
Wmg1qlmvgTmlIVoPnIdaPiCMoMpv/eMBp0EdHdxuxoxWohjAg8Fcpvf0CR9kZUuvu5GEZbNX09+6
jxCGx/fOG6CHV/kae2b2txyU7O3cIo1ntWelKdfm1tMJZTQLZGdGixuAVsmVWFeotz5vtgW/L7Ad
3weWVPMeHnPwzv5o+3KdRVL1VoFBv7lealsrcn/obY7eBdBhqjfmFZqpZlzpG1aLL7Im7+XcbnvJ
GtjN726revNSy5mmHO7eyOwv9Zj8VoJqjb3FwVWI0mtGIhCcR37pdt/1kPrS5vHs8OQWqvsb6x9n
UYWrRr5lftjKy1j1bKytrkVUSAziv/JGpXUsm/D20TAbkIGdzYkipRj+dZObZyN6zesP2hfzAFgC
d4Q6Df3S16kmilDxKLDJIER9FjrXPapRLyLUtVUbRxTc9KEoGQuOqn4KP2/Tg/Wbot7iEvmoRM3n
xWbLe2vEp5Jb3cTtm28auVsR8ixdWFlc5pa+KnhT70PwDaXeoYcnOi3BediNvRCq8VDjusRd13+6
ko1jqaYPZmviPUZW5omaH+IjKNo971JDCiD9IIKuId/k173FGsDyQ1Nh+qOjL8fxy0Uqih9AcHNw
Wvq7ABbAV/j3g5JnyHJ+JDwnamV1/8t+0PUnOHDMo6Op4gH3XSGq21HS1you34p1+gko7BoudLCf
lZjcgdiobdOgIIQBMLz1HaPdlq3r+oYd6KvT0iCoLILWSSR7f6mQKIJq675Kn1a8hv8rem4vf2Xc
DUu4H8jJZbK14AH+/5dU9LwHXiqdegk1ngI6np8QZ5PfuNtJS9m0rLfKqTAG3mjwlwtfE9NKhC0n
6khmHVHZ+UO+ShZykIuf+DmFkFYUEL7A0zLEvT1Zoyf+YPMYF7wpZJYkQsV4BdsD/p23+z7gkeAP
2aZ5P8fmhI92pgWNH95UloFCEnY7ucb74n6qz9x3W/NNwfcRJkk9aqGEKHPxReFMDo77On/PHRUa
fMFSWrKiPuHz40C+OG7gatik0Oy8KeOk1LeBQphCG9/UEqInyYClxmMKokWIA/t8cPNjvlnq8boi
YPsmYrjhnrDT0PSHEILtzG4uhUpjrOwrFxuUTnmJbvKGN2SV5YE3eNpZ/NbUbfo+zU4ixjFo+oCl
5nuub4PINslWTxXFoQYg0SQePouvXBXPiz2pkOpmv2rIXynEcuK8PvVWvK9YON7wQHKjJrqNDXVu
YzW+IK/ocXuQ8JKlS5B0WZHJNhP9vIdMCTyy6KF/v6OnjQqAGmA2DC80i5R0vNbNNa3hH1eOFSle
plHKlI9q5U4dHnFnYO5CyJVfCXU/c+ehwQ6qLjYhyvdO5JiY6tbNwAx6UdBeKwdsVMibrGhNZqC5
uRA0oEuBZi/nYcl2DiMl6GZPnRKvB5VtvA8MfooAKRRsun5DRmJWEgJUlAM5nxzR/VduArSziRDb
SNMXFJVpiwPYDZNwPCMcXMh4+RM+5kjruSmVb+O5OcTUXoGN0ZUGDkz+STV8L47NTq/JE1Z1DGCF
3s/TgMVhszEKTv0bfJLTwq9nyDWMIBWvzDBuSoKUs6xL0dgQrgpzObKmdsXXxxp62X5NAN3eTAnh
emEI/eRYj6qp+9hf7NqdxztaZoG3YX0nNAhL0rT8wBRSCP5u6Ec6xF6BJkSZETirJpH8g7nKtudj
OoC5H2ZSVIIYcQ6MI4mFZC6mZcsWmWNRHn7QslGeG9Pc2uUOsgmhrA1BAcqwSml3F0W86AbdGZIf
RHW5odOlcLIJ1cLSBG3Vrz4jb4y5CDFvEwoO57mHPm7vOJGj/hmrJ4qJXro0u23n0IYWDQgSyVxN
RyV0J0uAbNjCguFK8Gj+x8YKeAsB9WbD6voXHb4dNu4pAoLlHPkR9NSSJ97ZmpO0rWevJPyWszbq
pw9DhlGBzop6lT+6OOtO34396mAFOplqN2fXq9hf0Mq/EocM0ZzPqNcezQC/oC7QI9K7ZzGEtWTp
TE4rX5HzUUjGLj5kY5vJh/dS1FXIBwRzOvFXxhFuuoxUNO2Gz05oipSLE4VJUHFpTSv0M7IxVlSm
6n5zVLcUO569Mkzi/i2E4pOJZQkuqeWooz/S2KBa8KijtaxlAixG6NxnJSO6aR5bPBQ3gNazx1ZQ
t1aAeVzsdotjp9B2m1/eEUwlWnfMHqI0lcRESj2tlqea1PK6A+/c8DlNaO3hvI7Qi+OH6QzaLHNL
fd9YVOhoIyyE2QvqjWpT3CgV9ofHuaIkqF9vDCZ1CKRQ3PdT2fJwp1NbIkXbMY7/tUeEpvPI4h2T
Z2rtmL2UEMtMfJMurQOSNRPETNtNeXdIJxCzYTfpK8ZTwmAg85NqCxOECwYaN8fbp6pDWUJHLepO
JcoIh21WtlGlxjgHqU1mvY3y1+JmkdgvmqT9Q7UbfmAw2ALtEkcQylT0LWGG+r5n+DXLlYbfFOKp
LnXKWD70h/OYS6jld9v5oUpkV6gfqnLiO12v6SllsDjGMgA3J/OzC9EgzQGlsn80olL7MWBI2nrR
1Y6++htDLA0wz4iioNkBy1Zwz30AchFcJIjV5u8Z0HibuLJxrzMwevfmHV+8R4gG0w8gCnRWOHY1
ETwc6Qqb0s/qoUBzQC8SVdV3u0H7zwXhKZl150oBBC9XslWQI1/vssAngL+S36QwpPuSFMyD9DF8
+eqTUyQtCRThdyHzSfzdQiOpV/ecePh6prrJHD1R2dY8v81toVtCWJ2fJQGtIGDVR7cI40YmCF33
7t0GXhCSDbClvxd8qA2YRqU1x6KCHYZ5pNplfJR21f/mHt80moCcWOT/V/NHycov3RmBB4hrqZmv
S2Zaa5Yi6i3tpcMoNwLPIl78v+r8zqpnB+bjLuMJ0yqy3p+gshnOvnDiRMdeF9ek7dEfESl3Enbd
VxvrFOqeFRTIm8HJ8SEYSbaJVdaty6gXrQOKWIibLKL6AvlcKRMdEPydy3gEsPE1mTuEmcMcixxw
yIK13IdLng/xMlyKveiR+OVFcrQH7cgXs1s1BGrgARnhCndmEZpDu2Qfz1ICrRktrRu8ubV/RRYK
Rrk5inWIVcbT7WqCYsFPbta2v9w/NtG/grOpniK10pjLNjdLf+dtMcOli+V0ugy6fjrMBs8s2E/+
PYIAg3mxqDMBrwerPAtmX0E2q+V0433YyEB9IHCNkPrJOxLxIvlbYl7KAp6fNZSyo/O8gHu9Cb5H
pJObmIjUHHLVS8hvyVv4+/6+I6qFh0+K2kG0puk58jZEBDHisKdjSRuhRw512m2rU6WBPqAwvgT0
kSmbL28VrS68OPKaUEQBjNxrk5/fCDXAnwVqDC3L6mOS6bV1EKmiWbDGuJnk5iRILOsTJn89xO8D
dJ1YiT5YvyABEqA9Ln3c/PSdDvb3ywS9v8KmrrOZ8DLRVQmcOzvUJubm0VU109pL3pypjBLdWC8p
TKd/mQ6GtQvvpewBSccUPK0Z3EH36M0Vx9g8VkrUWvFMRBq18bimf9qBbX8SKFrEH+XmcbF/9Efw
45yN6K8/eCAvUpNiJsdsGTQ131Wcn+TZy4GSrB7V09xD+TPdFJvhrCFz4BHg3E3a7xsaQcak157S
MN2/QPYAltLWtiodSmMEF9Tdmg2PVZq1vkDX5+aRhWbdO1PZctNYzDfc74WAgYg8MJOI4IhXREiE
YNVbP4IUlXvK3sFgs8IV+mtY+gBp3pFpU2MiKwpcrFJAhNZLf1m/X9XmWM8gVydhnj5eGPy5uYaV
XC+WrNumXaXXKRu58BRjgsjEAh2INLgApz8k4G6w9Exp6N2Ah95InBvBMtgYLk1+K7Uc4zxvvWTg
t48zW1MmHxnZVEntzTGnhgJE/9lfO0ng91bUEGmtzZ7Ycf+M4ufXe15pekWuirHW2sprIB5s/A+S
FwDvpIJ++Sq+Bx3KvAWXgvzcfuwLk6vZX1EEM/OuVb7fIoYSDvvbS8hDJrLeXoLvnybJecWw2srz
vAu0nrMGYOV97/JLylyvxZQefHkqtPG8LZoWvtgKlppTJDaseUQnKA/8yBAmkHsmzq8mh+q0+7lk
JYZzmjOhQSUcwIwqSdp/OD7WxbY03zHajnCJY6WBpD7GGK855uicLlE/0PPJYNZ0PXwTkqPe6aW9
Vl32JQ8y4Yd964/0S6fwwMVM/PlES0Rj6xKZX/vX9DW64SmcpaICpxEssaxkefftsg14HKeFDMhd
+zrx+3IqNkMC5/Kx36dAYv8VRn2cSxwbli4GB4fxa95AlchL8wID/0ctUP2oIb2jK4kMREU0xk9x
dC8yYIcr09DrrAxGBWtL18mdkjIdLVNN85oJFYnc3HTCexrzRMGTwMigxTs9JhXKzQLTYmqbkTdU
NtN6OuoYk3luJn6JRYLJwPZf/CgY/hSPCUu9gPe69Pr4FumvFRqi0ejj0TyVRq3GFjj+ar4dELUN
rnBtmBfsrUbDXQlo729fifv3c9IHOndYpvMAOKsKDffJkBedq1F80spNmCKLJoOmTLGsn+fKRfne
nGBzeJ5aw4UFy9mmAvvVzqSTr5tV/k2Q+kpjIaTgW74suSTWCNzcZA09rpc0SW0QhRH8mIPCgdr1
LKZAg9/oSABuTVsbO5ufF+gDaLQJ2sltXqw6lyU0I9ikazt9+Vj1ckeLf8MDcTr56IuxhFa1iwRJ
1mlIPanh7xNbcoL/WKsZtSfVFj+QW3pJd43aZGwyHpNTCBhnPD1ZZ+icbGygaIxluhv6evAdJkzv
YyJWYVWXB2V0/tlpb/PTa9TVSiTcQ6XTkQ8J0xZlgfwIPVUiqcBS7NIm28cxdsyNEYvxfS/WKiXe
Q+qEBcGEBQK4WdHuH0YnsZTws67EmxSbEo3zLsL5CHoGpMsv5A5Jaepr45YjQ1RVlcLaiefE1ugA
BH5qkCqt08lk3Qkq9Ha0EoRy0l4mXVb5Uh9EQBXM2bmyYVgTT5J7dli6ZGLXf49wmN06KoVJOna/
EmlJ23EEH80TABV9aQGyg9ycHpW+f1QV2RPwVkxVz2BjVpQxW/isdTTcyWHfjRAPRWWkj4Nafe1Y
9FCmEGVpI+w5t73L/0eaV2x/qrcWE1oWyiMhLsEbg1Sq7NXUlGtOOCskUswgqqCF0FqETMmCrYnl
1cD0dw91fMmPwLBMcEI8eNxjuXgXFlP+Cc75vJ3FYifqCmwkVZN4jigB/xMFytCv92MB+9976w8w
q4QWqjGoy6A/XRc3fVH84qS1TNYM/cXvUT4R3ICQuUqAPw5B+trcqDwyMLCIuFLcTyXA6uimrpfB
6sIh1rYaRwy2svzVANU7rbIt6s6mqEZc5WI+mpW/YihanV9Bt1aWMCDnlWqNcqIrpUmh0a4Monyk
uDKhmqISkH8J0A7nojWNeMyLq9FMNW+UVALKkcdZ6S7lvYezv8nD2Umh2i4wpcjp8Hnk+XiBrkZ6
bKFve76pmPTZ6He5isgVuwyQoUsQQcJV9wYEccSETcQTjctsFY+9C3AD8yKEC7ki73oTC/m9BQrK
Lrb9rpuuHficgd+XIl0H+dzIeP+08QtZ0bg6g4xHHTQaWxehZ69E2ER8Ha3OKpqVQfdXshvejpjH
sfdpR/BA7OeAlDMEMn5xBZpOSuBHmv+X4Xi4uUDiGZuScebxqVNYYfT98z+P4YaoCQV7NwruesBR
l1gxlikAimnGVQj55aDtmwX+Q5HEZMuBQdEdPl5SG+asPukgCvALYDO0YG3w7yKk70QH0wfGTL2l
FGwHvLsBXNKUtJf9suQY4ZUpw9AiwTh7vroYw28Im257bBAzkzCAv2qxgQBpi7uHrqcXdUbpG34X
2LypKM8pd/bxv9Dmhc3tEI6AiOmtVdeN1/uC+Ja4idblM5PChUggMdkAy6idB0KjWn7YYMyp1fwL
D9vQEYwJp8wHKbp+gJHnYSfiit933AkNECmADcN54K8aHFCMmf0vMQCieu8HkL7joxuG7Q70UYT5
vZv3r7XRproH5RRE3wuD9TolDiSCJJrn6vbJwv9foQqiA/F8Hv2TADqmniiumFI6HvxJcsK7swua
GqBcW8EUuPkQcHYLCaGqv9fl1YW9r2hGpCe46gBctxbclKfT2hykORZsnr9xV0XPK4Tg7V/FHd1U
kvfhAbvaD6MRaZgsmfY5PnvP7gFNgHitJEBYYiTJBmUHkfaO5VguQwczsWj86JnCZalt/Y55naB7
4xKKM+BptT4ejXtDyYXa00l2mmQpUlVDdxaFaokN0Gsy9+a4Ovardi5NaRNuFCX8sxBAkgEKCObZ
QS7Ggf+0HjL5cQxD5oeJ72Q7MfH0GdgUDbCbk4IZf1CfZh/FKQzZIvZ/KNZF1sqvVUTmZhO4vQYv
WLbxVjtP3L9oUlTIVapIo/gQ4GH6DW9kY7hMkw7UnRBj3KG/Q3ru4yjRoT68YVQb4P+fqSrlv7+j
mSTowOxwAakYe4WRApMlwUyn6A9NnfvSNAh1d+EjxNk8Iurd0R+lrtkTsn9xJOHPQi/lo8CsyEuF
Xk+RVNYcfnLfGhFjLTJGYJitecBSx7GD72e0GHbqpE372wERDvzowVdvuSa03bohT3nysOP0KAoJ
RI8Q0RlWQ+ooEWvEHCfgUh8auQihx7/0k5cWOYsN8ZZstE07ZPwI9yCT8aYG8d8xdc7WSrcvYghc
nMyJ0b6mEZPscUzjuMHXJyZCCcWJZCaObYaOz6lu1Dqtc9X5nuy7HgFvwEsIxFcNMTYBrQvuqjpb
reWxShbjqgCwHWAPuP29nUxOqfF99Dw00CbY2OoJQD3C4ZpFBRUw49TbNBa/rcsI38upRw5IGikw
JJzLP2HMpgmFIWY1yTOnjk/y3pPSRB27z0G1hHPdT6JuIOi40k9Z224KcWeWoHnd9OccMa4BwkGT
Q66o2JwBxhqt+gtZTDSqws+/zEpxb+R9+crF9MBDwFhS1DCFvSNmyO7dL4ExuSFbgavQ21ZZddQP
g94rb37ZdoGEG70ZONNNfIFDM6de6K7lqPQWl8DnxxsBtQ89z9OC0TjsnPERUsBtjgz5uW+up5nf
teiMDFvyefjQAkc5lR5lLXrF6z75sQ+xGL4uD2xhbx3OxunQQch24YKO/m1WW746AMskqMk5FO9C
QuqHOR/ObiMBlDe5Rj0qwgLOjniOif6CwEe4jiyulDvQbFUtUQ3azjKACui9o/ssZLcLNs0QLy2i
YVGeD50QEHf5cZYF29at3TMhsZ5ZYToCl/oDOkICb5wNm1qVlFdICzIEeCYR0ILsgGmrh8H3zZFE
pEC5ZmqJrutxIzwIgW3QXJh1Z/72k2aLVG6qqp5H35i9JI/XhQYWdUFsNo0NUpEBl1C+FLQwZ2kK
WLVnCtbQE7hU3D6/FFP4dcqZZmPi1r/R3wh0tjk3NH32EjWFhEjXBkgMsvmLolf8mUPEO4GXt1lD
vPs6Cm56wUp1wxXzfZ8qZMRMKl1u5nq4LEXcvFLb+PhyzCPr0bsKiSqQzhZn/hKoHXnZqu9oqnPr
ZCQYVDESowNauOgb+sQ/8jR0IEoU8G3EajQSTQMzJr3wKWUjolPYhowmzhVHM5wOhFx42JhuJXwq
7DMmgRheLqgwhE4wa9lwvtyoOx5vFi9UIfuQFoUHi5IDQYqI4DHwXops/y61IsG2/vaWx5Uk4H4p
ldju8rAQ2vN6bnt44/XWeBLreF/Xzs219AeR2//HnxxQzXAFl4vQUNYJBfC5GSSyfI1DeTA6Rxth
3rioMaPd2JPILPuzJy2iu/be1P2Tz4dI6CPtYYwNzKmrJK8Q3x4iNbApgQshbuC4E3eI2SPNViZB
OCoyJOSmCztoOt2jIv0Lpkp5Bt6ivU9GSlVxyn3dBArJZ68BmAqtFbRuTkjjgCrqeNhE9UrzjqNV
XcWrQNSCaAl2RRMxv6WpSa/RmOJeTY/PtL0R5VkVvhno9uCUoAQ/YiqAZT7QOgEUYkQ0gWia2/FS
cXHwGWmtH6gJysVYLtzzrXTM+yZvDuXGm+st1bJhEvsU7t8OL6fl0XBwunQXpQaeoYaSckY1sFF5
sTa9ifyZ5Dg89SRcELhePDE+xO8SaeuoTf/fqd3URVnzF/eXHWOQ2yKhO0Ok0+KdLhZE2MskrKxn
SyjTWMef89FZUHmjBOAR3cizPSNm7scfrPvLIQtxwBM6ML8seZBHIiE7SGzP6eJl/pZR+XlibKxr
A15cbePG9OY/RzfDGUk+6J6ZQldJJHxLj8OIPYQv+coFfRMw5gJ3eCJiwCk/b8SRxKHYMn5Du+w/
G/yevEJZ3Ey+DH0Km/Sico9HOmN7bQHTkw/pzCMHC4npYCcfUYEkIYiSjIqfAIfArlpzQcvrxNXX
QxWQX3elHG/w7Msvg8HTAfhhs92mcb25mlcK/GvkwSWXb9JydJTR1O/MPmluONVIKlAEoeHryESf
jC6kezxcWyduT/VTTJiE1ng8DAPXMXwBWRcTlgnsXVLrlkQbHYM91TdYXL5cLQvbka7GfQlbHgCe
u9zfMBJbuEv7lJOkSz0kyQlMpfy5tR/dIA7SZTbs61iCdzZ1OXvRPLhk38Oc2x6qAbwV3ZCugtsM
VNDlGZgjE70/AjuAl/SC9UrE/VizZjvgiw3EPBo9t1KUhEZBzRa/BhA8lZyGnLcDrM1UBxz7YoJ3
FLPHzFQgUGFFK7quUsyhzHWbzigsRGKAgD1nbXg6z0dcV9JXDtwcSae1SDwN4FbG6+26JUzMT/B8
zKkq6JNK6dc3PqCMaTYnDXnAQCYbPwDlqcnnxHfE2KMjBTs7FFrPzius+ExpLrwHxXtpBTGJyWWt
jWKTQlRXVGh2qw83Bg0h68MZZMLdR8HT/vBpo8VT7QR4h+gr2pD8NcehdwmEC2D7wmcl/XDCZ/+M
xqlO9fDCWi92V1CywWRizVIC6GeH5ddcLx9tmxeYVY168m/0FcOKyaEVdYDwSPXUInrvaGci18Jb
FlXysm5U9y6UXRs5FE4oTKHc1UYCYIeLHesOzZVr7g5npH/qVwReteStFJF6+D2TskFbAuUI1wQT
TZVfHxKXxMWtM3IzabAAW0Ll+/iJkMP7V33FxKtvl13XTqb5f4u2XAXEKPhueWy97JLJL3tDMPyu
FD6BNexzI7K9RxKkE05/szfVcr+9c/UjA+wAb34Ew6VF7ZieIYtGsA0usNggWHsAhFSTza+txTaJ
apoWxZ6aj4LWywOT9CsAh61hHdlLPgueQhPCeVizi24UmngHQBMb7uO/jaou4UsuKjdeW9jMKXkE
wJUp+aQcNV0vKjU6G1sBYsMIPvyVcONVjZbyd8O2GjylTP1/xSid0V9WgoRZKLH3T1KiutrsJaAy
0u9tPKj3nPf73LHHWqR2agozxD6tbBCFztP3n2L6FwDLS2BL6ax6AhhfztpXkQwO+wBxxnX2rvJS
ass5fnppIHqLOb2tfMlP0vrOdhks/e1udBYoOs9POlctE1cQVq4o3buYXfM7OaDKFLfHySLvab+u
BaBxE35DjoVDP+g+zha3eZoIXHh71ka27ijjbCLeC/IC3RT/Ju91T0WVjdCUBIg0BfFN21iE9xli
KLfxYmcgwKonk62x5pQmX2Wfis5844BpqTegzAaCqmuO8IK73MQ/gofBb2qqcBq3C7iA41iZM4d9
s8ORF8qWsHVXkB0Fjw4l3MOgp6MBVKrqNFFHlYcggXKBSsJoEznhqkPFk02eulxHVpBs6OIqx1Ny
C+anoqMXwGb/PdrJdf4RS5Y/hWiVPsmicCdYzV9yOStNxNu9MKZIAwIOA97StAXfblOdXjolWBbI
a78jK3+j9l+C625a8u21qwvA3l6QHCSw4GngyoTbpX1+jC+UZSp+tTFkQ24BrRttkn5qMpSKKkrd
IKMHmz2nR6w/tpkQ3d07MM/LtkqaMwP3fWY4DlbIkgMf/FQDXRcKJV0JVi66bd0uWRRr+PnQWwgk
At0ZMHhO+PzphSSaLZERrfJEWipAAjShGJI0UIFVd7+ZzsCUw9GTCz33eIRUCqIo3P643FOAiFKI
Tjz5UhvmDTIuRe0Dp1pb7Akkz7i3ergLelSIqZJrqs6DUoDNY/XKolGphse1w7Hrje++Tr3lQhFg
uQgFl1hJ4c3mpNW5QjXAZ0JhTwtwJLAKhXJ9eOuVO68HLqoxzO8b+yg4Ng1Pw1LcIWJrOonp1yfQ
94s53rgdpfa/+vlDV41G1Yu1oOwfWpO/wsawVVLTdxzHZE29JaGTBF85gVyU0MV+pwE9YRCvyEuH
uoSI/nPYNMxnNVZ+PezW9CZSUJmvba7emoSDEBhXNkEVhzzTtl8E5YB7mwAzXRNAWTeraUYdLd0I
vurEHQt8TrYHqOZrCNYkX9f8/9OLdjUT6OkpU6w6rPTaiH22yXjLeAxR0XAGWghQqHIwF4jQrUzL
n/fXH2Gh4nU0k5ZW+wVramgUBY3drWAfj5+wdClLPhzrZs8p6PsxyHStFyCbJiUCY8XoltCau+Er
KDxQM1a8/t4VC9HZMGazV6ffUpyu7OsSfiyQZHVMGTHyRbKK7dusor4GxE/+F4iCREMXnLMlsFK2
evzcI7QSKQ2c+UVaJREzZPB/OS/3GyYD8ABROogdnG19t9hOmnW0ClOw2p9mzsAHxWYRJH3OW57h
FTmxs5BsKxf1MyYP/tFMLWbBAcZA0tHz5dipbXQkA7RjZOqhP22N7sFPjUPHa/LJIW+YvWT76AQ5
fbvdHf8oSRB8YLx8T2hUj8qjle5ZZ1nr98iwmTRE8pl5ATn+so7p74uCgZ/6mJBs1Umpw0ekvXEi
HoGLEm55qr/8oXPiB9EJdSzo5ksSzFwKRFkokNsRKXcAneCg+aPAtoIOOR67azCHOyBG3b2HL4/L
yb8NvIuwQwxdHwGOk5dz40huBunfsc1gYd1wboiCW8fPqdeFjjYS7qob8xjz1ZBwdsnMjVR1eDCY
gMto4OaqMZygqo9BBoP/FA/jP6WV1tov0MeVYhdgTMdysowzZcTXp0TvNRESDUs0WFj3b0kgZ3Zh
AP10U1gkFriFSLIRoDNW6rQBP/pbuzwmdUF6JCKBZMWsvqvrM2X/FTvJLozaTYOVpc22mMHOtTpO
qeX4QLbX+4DaIcOXByP5RUEC+EJ/wxRaHBw1baTHEsxKS+Xmbim00KuMKXSiTqOsSX07IMXnL1yJ
OElyXqm/QqQExUs2c+/qvPxzrbm6jFPCQmQ7lbTVvveOog6RbjcsjNOSdwUCTTZh9H0u+mKSHstP
IMUFDIhvuxqokXhcScaG9IfSvxAcit604PlVABhozbvLBxzW06WGOi5zmUrYeSk2quQDGAay36HX
0WLwgF0T+CBMdmGKhxJ04gkL7Jb6V9IHblMgm1Yimch3+BizULnVIS7o6/ElrNEPTxKZVHx5WZnf
gdsspkpqSjPy8PQJf6feuTcqoN1TEfMAIOHDzTODUwyLoAdkf/ZG/74gUdV1Hmefkl1WNPax56UM
q8eQ/g05WLRiAZrekGg4aK/uLZ3Hh5C0/8V8J3SFny5+BkUY8O8t0eUhPfzu+FP6Uck8Icak2VCh
vfLwogFJgVo2QQZ2knQ4cxhDjP/+5xMKndIrR7gAyZv07u81oriItiMZZ8G/5NyCa4rvNmaU5D93
P55HHHuKMq4r2T+AUV3qmOMeS0abp3aoXHcX9OXRAO67ETsfaw2hE57SsS3l9p5O09WLQ5K58aqF
4CpAdFnvAC3Quay3ZGiEf3AqhTEnNkQ+M/b1UugBm3gITkrf+qbSwWZSFIjQsIZuV0O+T+4Grga8
+0dEbcdv5W+9HNpEA+S8BPweyTVwxff/z+tBR12kliUVFm3Rh0swWCOH7zpBBavZnmefkNmqBWHG
YExQ7nq+d6aTHIP4UevP3Tju08ZOqvcooQV1fVgUy3K880P6Dh98TAIiFHR3UtPwHzoEcSDn/wgS
iP+vPcQaTBrvP53SBzjOqmuRWf2xPMEzJCtNzHbBEbUqWGiQpyZJ5JythiPpmYRzR+OAJl2kbHdh
ARBVofo0KmXTggfijQgduQEi3iN3j7d0qZ9z3tE7HOX8IL8wlyQrpdATVmg9XQ2F0xMqZ1NcA9y+
U7EcweuGLj2d+c2pIAXJgh7mYFL11zBIlGLXN3xq+FOUY9kkss7TvU5sjceHNhEIwfCqmsrzx4Qb
Jq6+Ru2WRoVqaUBtpftvsc3uidBlyvMvECZeYGxQ5qOfY8Dxxw0rmO2hgC/GywEm3d/oFSBhsCvG
eERXD8wghtAzURXkodDlI8y1LhgTQmxsER2J/KISQ/9A8RFKQ4opgINcjLdB/5tLtW7tVtj8DLLl
VdQ56KfBKjvqbnw4+TAzBb9j+uBhVvJOxioHAH1GlN+RJK2uTqfwmpkzQBxUWMs7Fix99Z5rmme8
JKafLDhYE0s882Zzb4Mw4SIihVQJzEVWMI9ciBokZohHXGeSTE6FCowDlTLpTD1uuQQ8cQpl5e/V
0mN45/fq5VTNEPp5ysEROXR1MdPo7bGmnAaHnmT/FhSkwSpkZ/gA7GoX6DBOx9kkHx/rNFowrFim
6Dg/wSYgGtJcHNa2hqTEJ8FWBTTOA7yw/heoHJJcam2qm5FEMGcMfYP2M/dR53Nk0qpzkX2Ny/qj
0BDGtOhGzDJB9SySntPT4OJMwnNC29WOhygce4FlvRqcYImJGDpjU/iQ7q9Qf1NOL/mViG5NVtPZ
ADX8U7DNkGopkwofpPLqDt8G76Z8ItzZt8f6+BCwYjimBqXwRCJogimU0K4FlWOkwbs4m4EOLm0s
NSAVK/3nKlOy72aBXEnFSq6exiqCrV/pv38mbJOw7iXA9FItJsm89WBRhwAe4+EfkYMojN2au7DE
o03i0iBJlI44YEmXXU6ecPB0srTilj3qLfYZXS8yIeLdAeahqAt/nE54qTEE6uKWGE7HolX53KGt
jDDUkT+1xrdHGqLIstvFgl4EIUUcycei72xbB86uBAber7QcwWiPdSrViBRZERTZ1RGURHsGytAW
anSbJLABbvouDFcN7GD4P7YV5vXsZUgKm+uJC77bflgfxOfbkpHXseVYIKvw2hmcQ4/t/hKJWaCL
xYRPdOfUpQE77lx/ITEJwQ79aX7+E0pROAiEe7gidTfhdZpZErkhdzVQX1higjxq0+W+1QMiuvdn
w1CeXL4tK9K+1JklB9c4SN3EOXstRbx27hRNcdgJqRdowpGn+0IBfMCv+2pTaNQn70gMqblYy+Aa
SogsBuOcuybJUSayl/FSaVVUJR+HgZ18I66UdSM2/dmdx6ZfWjlBVO/IeEbB68/eOeumx8Ul2dgQ
sTslt+wMW8+HOZjF/1XUxkQpyiFl2sp790U+8KmLbgC52J+FGAh0qgfaGk+7y2A56pM5/Gpyqoxc
BHxrwwOX4A+LwZFaU7b2o5VU7y3Hff3u1UKYFDYbASJqqCZVyEakzKD2UQ3AlPc0TSthD4IuzImz
GEDgc2EZ6DU598mX+cOWzOajGvU4xx9cYYfaxrEqRnHOg6v9KZ9QdfgUx6wyzxO4G9vzciGuwGMC
+yeQ4fV9/EmOXl1bkB2TXaXGePOLZSnIwwmhlJbs6B1/Zi95f+vmevgeHOp7WLzRgS/q4pYg/5lh
n5g16ULa24ZKQvzPnEQGfbAvjm5om604TTvRA6EGq6IF9kffkJuH3S7evZId8TvbOEGMOeRHSRHR
tdpWUvJvXARSry10bcyqCp/XwAhzwADTzaRk8pmQHkmdXKc0r7laSp7Vq489JzaVyafOW1hl56eY
lSXsTQgT+6Q8XTGdm2JuIea7iZxbwG1PLcHzNvFd2gXkwkK2vXAz8KLggurYdtVtFURKDZL2jTT1
X9M/n994BjgtUQexi0YijX3gCWUUaAU6mtirVBl6ytXb4Q/c12Z7GXrkXOVN5b8SizGldaU5uzCO
V8fao+gXAdP6JZNAm3wHwZIQzDrSE9HNbA+QBe4F4D0JSNDsZ4oEGH4yKw/qgINCecyHf730eozE
2ApHLtydckFx0eF/Zjd2IN/HTdEQPx9ChnCChCdMIBYSmwGCS3YEFptZwbhQQfTSqEmjSr3nnMFS
1lYYiNA0lPBv+lo2mxpkqUnpXZwA6po5l6A802thsQBAOdN3tkt0Z66ENVLkg2l8b/KIMxK/lyHE
4mYK/dOqNmg+yjypPBUq34k9mHqDROEPo69RycoQIwOCRkkYF8e4DlsPw4hb7pDKOxSL0pPo57iR
W68n0O6MLHRuyCx+eL9SRrH+9Lt47/EEzEnXVbZLfHPKo6dwuls8nuQYBXPXU3gaBr/gSA7xyJPG
AMvnrZfjY7GLaqykjdozN9+CmEx1AC4mhN8qmydVyNxSWyo0fTRYrqxfU4y3TG+0x1inkLZM/mCM
Zf/GiobcL36PqAG5YyCVlDAeNyZVwMxgHa0AmQN3Qe91sNKvKoNkTuUvxUGBZaiHOJMNL/IeXjr3
rPLhr/XjTuVjyMRZ+oBlpncmg+gjjpa7U2pEDBK9Dh3H4Es3GK9RcNFCLZRui+AaXoRp+KHcqVt7
qnRyqnynJHp9WMpiUy9umlDLZTo7ePdsymhFImteE6H941aD7JUn/cSkDvB2iGO2iAe3kqqSj1qV
j8SrgYQxJ3R6N6qpOjDtwS/mKntifebhiuc0usnRXdqcSLNBU2Z4u8XHlJI4qBjcBSBXjbrQGOPb
tsq1KbkrdgeGtCgFPWws1t+HfoJDbg4Tr215Kyy5ZJlQX2lX3+T6nKPAJ9g6JPLTrWnmISthxOj0
GhgqBBMppP1MxrZjZ3LAKysRg1pMvV+wQ8MG1Qr0PaxBKNByh8ujbM8FfOMGltHMPl4tfA6LRjF6
o++JfUrkdst4grBu5qU69OXyzTYUmQojxEQl0CHhGc6ZsPhjOxayuoB5VjghDsMiYOF+GITeqAf8
C3sLngrb4hJOQWtcFMklTkXAJynpktdMKhe3VVNAr8cK0x3aE2QRLAJH87hMzJWQBm/dp8apYT/d
yWLXNzgAE2LZP0wVW+L46bQpfq1EYvXiiw3D+BrPuBgtLzzn0G1lEfAaJYzWLak2AyIQYpzRRmkc
5UPAgIphg3i4ycMgXj3Xw1rHsaY+lbpvBdcWJ1hkGZQoDkETdoP8Cwypen4p53BjTVhCAVfno4fk
oxFAz1+94E51RURuW+VVcUMgcoebVzt1khFZ3fB16wn6vwYoaU4L57R6og53mLjnCLEHA922BU46
jdq6yWYKNgdT1tfXQuukR2jyALxnOaujniMaf5DmD3TZXLzkNhqQk1ajKbChGOWIy+gm8P1iB0d8
6N9W8daaYBgrelNvNT8BMVD2r8EPiWZTd+uoyO9p9cU32NHTerD75wfMRhQl3cM2qyAVPUIOeP2b
rQr8ODyKF9bvdnRZSz1AwZ1AAgSgg2HHGo9GyTLZF+LePD/8CMcEJwhPYIB8Ok2Q46AzSca0KfYr
qr88CHKwxMn1XXaSpi0fbKQiuYCiRWi+1guPFyYESkBBT3gMt9H02U9IuhNgBm0PIX7vga8Ee7gR
BVuLhCm13WDb2zRiWfvGXrP40hYJb8Mq9MyZtVcXdXvQZgBKmmJrOOs2fzffPZtVqifEyFQ8tKie
k83yvbSujKmzWlkahblMm6gT4PWcUe03Ah8E3LF7crSfodNxFNUzW3/taYtxT0wM9MyQAvDmt+Xs
x6gFTKWIvge3rWKExt/gC4lJtdiSYirX8+3WQHjUfk+2cJ1PE8USnLGE21gwT4wKsZrcvTx58pQ5
CLUNDB3XcHMbPjKV3QOzzjhT8/x2MCeD6kA+9HtJqWKikb9oplE2AXj6ZQ+RJl9THrnCdq7ZlT7f
jGZRmwk4oK4PtrNiW+Rdz6VTMLlhcVQnm66MtJrduEBtEvOcoCL2EX8MfZWk0DeObZ9xYRc1VwTZ
8/GXH+hT+hdomB+A3w1X/Ar6deodnFDn1f6GIOWZrY5Gj/4WJcltRWmA5Gj1RgWoOEhzqeDuEPaV
FRk1is88EtksbHt1w1Z0EimH/GZgItyl92xw6UR4rtCJi4TOmnYef5RSmcdearylruX3z4pXWmY2
NpC8crFX7gAEABdi2tPhsM0lXNKfSTGXnNXoGXLe3yaMUIG9NiXoii4hI/wcQRuDHaaycwQYeySD
QeWUy53ol8DHoqgMYCxFuNmdaygutqKmwuzR8ldd4cTMmM8KcvkrB2LIpDKokmrrx0WBNBVy4wtW
XzxWlBdigyqPRbt7s0PkzKtCMXt8uznJ1a5Wiy2VZ9oNGyLSHdDRNkr6qFRi8QgWgnSmfOLayfFp
rLBDMTUpVhYtulJGHA8b/Cg5vdb/+LNazrmZWcOl2RqH3OKtDbewgkaQq7MsbAue9dVQN50c00tY
uXKINH1+u9PsTa5BmnFSQRV1KsU+J16OZxjUjbWIgyPUr7smSEPAl6YgVhTQx+Sm4OBBwpePAM90
8H+GWLY/hggeVqT5EvHRDb7jhY686xqPyPEyDpycLyo8pme6B1wB372wHkR22yzrrDVeFIPB1oX8
2gzwzC+PmL784134mUBw1OslLUuISli1Ld+hTXclmSHX+Sw4aontqKAi7tjYjhd3HEtvLfAqvVt4
taspdukeFHD9wqkDn2quortgUox9yxwAKS8lRmp501nPE1CvVA4s987qil+jdMNLwDSqIEXqmlB5
vmX6Wzy3Vpk1pyBIFIfqphHIaQH6+a+AEnEzYVnHksO8jVXu/fnkmFa3LplseVAARPy8f4kBdQgw
c8M4okc6t+7y67X4zSVTpxHaWPFMrwGranblddKqLeq23OD5tNGSrxiezWVSAgJ3SZ24S0gcrxhc
FlA2XcPJan68L60DGJVGPfkp8Rowe1lVlvFmecAv+jtIsrTenar4ft79/CUNbJ7noJxATm92ieE0
YmgO8/qKdOqlsvvzsRzdA9FKtwlWt0eFfKUGletWTz/sE7ypbgOJOzPJjJRZwhKAfsmjE949Joya
dx+YVyJZLhDFhouG1b2O53SQaCvtNJW8SWDbY2t9hT5nbaCd9CIFFh8mXOHV56KquGyg+fTVFM7s
zIyv+9RVWYYf35UnEJUkOzhX18tEk/3Z01ODJW8ygXBZtxZuQZWb7a8r52nsIWQvBKNA/FeecmWs
cKVTXotUKIDTHy1nAQILhdabAqBZN4tJz8ocDptNEl+/j1hPqxsNnAZYLGVwNaMn4dIz4noGo4dp
d2YuN8fD3gIwjHjmxR0aJpbBb9VMLpWPvw908r5Lfz0tTdevLGQnbkNd46rKVO6XCd6KkOGqSZJN
E9OStNzkamE/U2gAYF9PQYGJTJ8yFESs/f6T7tAvNrHEO309EijihzoMHhhGhoN9v+B/dYDSCzyv
/pIYTuT+PtgzOYv0FjmvffkVRBdsCxnRqs0icSJUjdoHEh9hSXexHozGGuBl85i2aJdbJB8gJJuH
IusDc6Fef1Rkp8xE4/c6bLtL/uI68naxeQRhV79/o1mYdWUaYAsWznn/5OOSRcTKqrJBKsfXd0Xc
jiVqvIHyq77NWhqqvenFp2+7//N5qot6KDe4t9jlpZ7DP/UBY+NlW4NoIhHmHzqUQYrUf/zPQsEJ
OhqrF6nEQfdF9R1WsNoFG4yWWRP7MwfknOvkYVoOyVGaHWpTqDGJfAJtQrWkxKlDW9DyZ+9vmAF4
Hx7M+Dpo1uEZWJvacEYkHbsa9zlywnhO9sCeWdBW5dlJzcL/guPlJcpdk9ieFWkVk0XhjKqUZI0T
dbJl2/BL2DNCQr4ApXZB9GQ8j+erGNlZVK3umDJk3cL82qsGowP9/wCKp2mm+geAF9o623rEpbby
y/GAmbq33bujWJWJb+IndQHyRgxjNlbrSt3WTFbscdqg6kdcYhwdfFq1pKB/SIVOC71xEP+OEcmF
M9Cj9H6ub1EmRgh498558AylYJW9tWwQ/tT/wc38QU6PjeDqPdkVnuoq/rvzGOjqnyyJifEY0gtV
ZVoMerwrVzFRYAqq0kK9+OZALa6sFQXVy0gJGUs+s61TAhelSCyd5yKuxYt4/uvIGTNA8POY1k5y
0YaGL9qn5oH5WQxoIZTeFwgBZhbCD2J9/cZybh/7uhembHvCAAt+XjEtjSG4RdEQv6992ZlzIkeI
S/JG2GN7+E3lM0O2xSwAN7kza1yjizpXkdbhnWcLXqmTlptEpuzdxY04ZV2XqCRko5j8NL6eH2EP
Zw6frhcJI0kQnPEJhy66M8+Yp1L5URrCCdWzevCKJnEXRrEnXUqLONFVTzpvgXg+3o/tg36zGE3C
nBBcYYl5Dz6Ve0fAfWE7+hutagWNi2TXo5eMUTRj3Uj8PgCqMg7IWHQwHwdmtMA+fM5AH6x0Cw4n
IWTxbvdMI+GF1gBMdnqynq2CDgjHLn5K0Tv1N6Q52CK+W5p2z0Qpg3iPIjeZvcajKhSWQzYzDEL6
ODUrr0GeCKhr5tn2a+YMszZdkEznMa0IrhwMJDEv0QzwEPJAXVWlCm64hOpTD9NygksqwoPbBP6x
2JzFgg34HzWkSwNt38cmE98JgFiSAh+SSInLhZ2GXWAlmqKonz38jLq2VFvUUXVOoYzOxl1MF333
22/8MExEKFpE4E4c9eL/DYw2lgMH7xJv4kGodp+l7KdhFN5eYPhF/udTctrPZdrPtrRb8Ix6+8qF
rjx66eO8T3Y4UhAZqH5j33qFUTaRnkrTe2o4TGO+vMq1OmagwNmn3T2MiUALv2jXuFZ3lCjJhwJ7
nzyDh6wCN1tr1lQwLB31DoEXCOGBxR45/rT55ctk5Nk2hNmtz+v29CnxN92w8kSp5zoc/AibbbFz
UwfNbu3iE4ihXGAKrHKvMQ6A1iDfPIjUOFWYDMIOkx6Hr86rscSJH1H8RRKAXg1aN+8cljVGO9ff
lGmAlqaOLQOWvk/3Zl9dFxCsXruNDJjpCJ6kHLAqsLYTWIBEhZXTZp+7decYC3Zy81aBI6haZ7N6
eXho4niAjZHkgf4nODoyM1lpmsYWCfzbWR3oYRABxtR59pc3pXzGIMns2HDnlgNqHZIuPN4WxZT2
lJAXTChPHsWCTMsHW2/sIU8FsGVUXgR4AI3/1hxRE9/WNcV7bcx+32MoInuRYvitHdPqtl21nZ9p
/C9O0HbPRkAHDBsVb4/9oXSkIm84eDynohuRsuad0AWtvJmqP3P3W4dBQfkBAShoDg2uYcu4JHxl
tnl6EzSJOafVq8NJ1Rky4UtdzkgFpVlMXIOTkfbtEq/1NeX1TLS7w5fj7XcE2ptVB/hnxAWtEL5E
eVfXpIyKNpHJKTWQjNB4oVChywHjc2xHLwnjx/PllTmdrdzDEvG7RPsn6M8I8JEeEFfs8nsOJJ+c
nPqpbppD5HVRlxMdLjKdODO9a/V7Yxqfnm+KSrFRxmqSQZVfTpQ9KrGzWW3UCTf0n/zkVIpwrT2q
8RbpI6flCJdp7POQBS2NEsXzv3LMwKvV+m0u9X/VPXmIiWGFPcQ6FQ2hYx2xNuOzI/4FMf8mpVpg
AcdDVJesxeUAJG5iDsCXdJ1YdwAiCG8pCqG6wKvjIjWTgbYrCna5wpSYN9ykBOJuRsHxAltbD/+u
vSEMKJrMPzutoCYb1i2yU3fTMckG6jzi23alTnFq6dJenr7pMqFUzDtGRm147hKPlVOlwLv1k6bp
A/ytlKSstlFBL1q/iQP6QUJRm9sX4J88BJRG5+Ann1JsRY2elBgBvbSmDEH7JLxXgvBWE11bI3L/
djdCKoKgiv8/NS2F2b0l6axuboO9g+dYAMTL+j2dGXVbH8IgAe57gxIc9NMtmaAg3Ay8aamVmykO
utk7zRFSZZYXmogIbbeSSk5BuXrpE/9izjc7xgTghXiKuK/lxch5smozKT8JHsRT52LZAWuLSDOi
ZAcVSJMVcsPCAqS4vKWbdWsln8IdPZLWqtZ6j1rH+2b1Ie46VSsiLa6jgDPYZ76B2mI57lo0o0ak
XCmtmY+QFjk+vlsno5K35C4Jp4TGK73YBrsgmNUCGxzscw7GN0UtvTm29RgW9nrzsU42svSnVZpr
UiKcMUjhHDPndqPnLk4DEx4XQsWtOnBQLpXR2KeI7f4Njq68D7OQpiCCeP/M62C/mXBCx0WWD0Ht
EDNYk3fohSG5BiHCwjpVhltYxBqXL9x6KQc2q2iKh38zHFOR/irw3DoaNvoAxIAwFb/VUZ3OTgPs
xU2nqTDejl4yooxwr+wBqwmlyRhTufZ3iG7koJtxFLJCNvWJScv5zgdizw47Ne4J48/dZFf2UiAy
7GAoe4vPZBHYlTgvPq51N0d7t/TPO9tjw4cWjzIAgdBvZZfgyXH48GOi9oAsTgAi9W7PKFEml1fQ
hBqhjH6E5kgDtD3koYquqMepUjgdR7ugFMoDttQEAdS/DqQrhFiVIbhkC0VWJtGmuaZ3Mu8pNXhP
bwIPzAeCvS8vGpeHBZnEDUiLrrP4Fx9exGqLE+DCeh3wcuIOAv53XJ0w4kcw3DI0UEyfPVs+YguY
+KvpuhJJeexxqQkRCtODssDcnJpqH/myJ5NpXDp5fefwE9gh5n32eT2jGqIbOWv3xmy8A/xKj/m/
TS+UJ2BOhE8gjIPFnodQfVBhfAupHgdtVSNzh3r307M1smEkulzQ2wnMV0LAa6xW3tXuchZ7t55G
wIcUVqK9RNx/76O8cZWQgOLH6wjg9NDefsi88SuzaQO5fMNEgcB5sLC9RvqsjDAoLj+sswoYEwjF
Pw2IiDokjvQrL3kO3QBw9smDOT5qNO9W6Yps7lTUjxKBM6z9022rkNq4wkrd2P7bfvpbUuDkUtBi
BLtY00lBMCcu4iJOAK8AFEtBph7RM2sSqcKS4b8kZdm93tDkhvComuU/6cSpzCNDUK+ljI+nsvRk
8ya0HkFvBNYx1PR9EJBwkpL8KuSxden/EUvC1eAqSrrNX4jjw06+TfCM8wsmlo2I0hSDQoJohTHP
ZBx7ZJSAwxLRV+wLdonxSPTGVkZlQSjGgrLBH59e2p7lQPHXRYv1jVR01vHFASxID/28LEZQ1m3i
zYmFYEjTDwPC6ry/Db/FVVTd6GbJUiFnaVH05KVmPo/hSX0weCQBOu9iH47cdrT+r61e5PeU8FRS
VPvrwj+gFv2unUCm2wn/uLybi+YuHUIbtXYVEKDxIC/DqcRcRrQJ7yryQGnS+25SrlCuwh9F3d+7
aPQgiXqgtgXQ/rQamFCm87Nw/tqhq6PX/YyD5ci0OMdOUn9MuFwbyHaCdLLN4L3NwLlRpTV8tywp
q8IauXRghO0vxY0x5FGgcBCeHTxmhEZL8BHDSbX6Oq86ba7rsH2JrhJeXqt3tjMeaLlBgGT3mUgx
sHkCh9PkzKZtBQCBx4hRUgu1PgprDnFbY7PVgt5bEXJaaF1ahge9MZaQyuhUPw9vY834+z1ss4Qt
F2n7aQh77jwCxAzOMq51HSzw/elYgmXCuzgumMHbwTOBHWc1kAcliIgNiHf0fKv9aEBu/trzVFCB
wHSBxu7a9OCJPNg1sSN1Ar8TDCPxJK5tsBAMLb8FWIAQ/2yFJA9YMXufkc2TUaTs6JqOfVrTt5HV
4r+TcgCvo5ZWAUQAvWGQ0NC6la0Ual9fh/qz79A0be56AzSErDVx4lvdJAXO1eDiLCt2/cbQSDEs
FxaHUIiGPWInVZ944JvwnhZmswfORZk6hstZ0NRWKk//cECjbxHKWWVsJen4B+ZqO4F0x7PCK0dp
hinq0HZB4PsskhDAEmRNR8C8ro+YclExyugdY/I4ZP4z9WreCcanXNrZfKn/xgEtObA0PVw//uyJ
BsZrVElOgZP/bE0rxthAOg6iJstzDtzgBTJlOAsw6zPpBj+pWoWBpTmhl4t4b+cfpS9nwtROsvAS
0DELUyYrhFqkIFIqe4Qly+ohwAaT/Nd79j3sjbnxNd9y7VHZRFt2/555knoVUh5CIEWYS6VFN3a2
HkwY0Wc9yVqeLwngFkm33dgFO2vjEs4HlAUMGra9nKo2R/qOoFcNb/msyfpfInhTNH2tQIQqv335
atnJiSjPzjWoIgFS+AwNQ3hxcBaHZMOpN6qndRaCAwaKQwkgf19TpygLgZd1UPI6sANjwgVU3z9U
X9QiPT7HpkINQn+GgU7fYjaT1tTmOK3XUoLaE03bAD8fW97X7FUyrqiGhaYPIhwmB7fk1og5Eln0
kkzGpVLvWjYAQFb7hA2Y5+BF0PtK41B7pd8klOocIOWRF33sUoFV0wK9s7ulUcVqXehy98H/paQL
oaeKv49GxXTzfx76bxH9LsioQF8vK/EpV1X4YwyV6pks8UZ8KZzHp5HUH0RrSKI/kohJXlZHWOCL
YLM86Ami9pIbaC5JUZvr9AN0Hg2A6ZMiGm1qCAL+fCIiFhHniBiSOGkYRzMWM2uQR2pYhIjXyJcf
WdDg8aU2p0D11/uu0EIuQZ9OgXISoxUfehYr5WmfpDFc+pwV7UlnsH7YWvOIJfkOf+EnyB9tvRCY
hhWiiVBiNgs3/P29RBITljlIPks3mPXKRXeUmbm+sp8kC/Qk+JT/kTWoywxj/rWniRzMzpyvK3qG
J5OuW4fzaosu796psfqQi8ur4h1o7TjZFgK3yF9b+Twh8XCp+vEiFmTco8KqaZRnAKOslDs9htHP
PwIGKp/U4Plme6mGzRAuMITrFEnrsMgKwxq7oCpk4tQuJd/suWv8RBfrURGT8AFjlM6vJrTndTVL
70JaQWI/ralCFDGwp0R4DtrSS+8Mcvc3RqDwhen8Jk4JmPLAnzyqTiiHCSIn7feYhMZvtP7bN91p
qCX0bfESUmgABv5h+cWhM6kJs+e2gW0cZeHCNYb66By6iRRYbpcB9HnmF4wKtsIHl5Ps4KZ9cKHY
/wdVkxVlz4bxSGG1udn0ivJPZQDhjd69tSgfEBG93bKq51rqr9FNejBsmXE0yh/GNCv0MMOV2YX0
Sk1/uTVNCq8vUZWdH30HtbKJwEu63KcUeJpbqkEGgGL823m/koRyq0gMmuH9WC/cqpV5vKDc8IPy
J/vxKk+l7atGXlIe5FA5E/AXHFMZTVTpa4b4Vb6rlw7iSNSowiezae0v34LnoW6UTXxmXk5nTEOH
csG/AzOA2WU7k28p8eSIoaTHE6BtMokkiQzcrDsJpuq21aqejPp0W8ijwqtyC1ngwoJKOPDSHcBz
g9lIWPApI6VJvYwBlUgws991mG796TbGlWCx5kNNkNoOePYGtIZbb1IlfA2CfXcI2i7rR0jaf+on
0B7q99L1H4sxUtjASlQY1022yideWE7GFEB7rRGJMV0Q8jg/y7Yw3ACHLcBgR5hKrlRqiAzknEOx
huqajVjW0hquxBwoi1XkDvzO1QxtjeUfQQcv+3wWI7o22f9tweDeoJ2y8PlG9459hGaksV2znz5g
Mz4d6ZDPd1LI0HqW8sAFJHepM4vUeVDi8lZXqI58nxXJFOsXaMc/kf8g3m2HgaUQ60tNkILlk3Vv
4wUWjGXPWLYrpEFUpCUEKHb4sPaGvfuXD+b2tOziIosJrfiRRK/Hr6dQS5xXXYhYSrzywvyRTIR4
uFwQeaGdfxfFOJodVSO3xfKe33uyge+wgk1Q+y8xoEESdjxM3IINm7w801wyWuCLOS4f1D+P8nqa
4aIg7wle36ihUyoMJMXQXkfyAkJCH0sT3rqd3W4C5L9luoIdaDAJcdIGaVbnX02zwAZpVZKaJ1De
U2/lXd/yir/ataBuGm1xZVGJYT4goT2ZCkzVgxrPzdZH9qS28jrUqQ8JXxlp8XP+tByTdAoi11bG
H/vlp26WAO7cZZ3AbMgdYVm+3hKC46zrI0v9gQUqyHamfMY/MV6UFEbnNSu0z6KCN/b1CnJ6HWtb
E0+a59Gk1Hfu+IbEcJ5kQjVpBdZtzmXjdxJ/Bz5uH1/CmYytv8hveX5K1NM0JGgAb/zKS9N2TWuS
hW40Bz13zC5yGKF+VpMyq5zzrSMjaM8ffDYo9z9+RBUxDO3S1DZf0jnz79svcgVP8SKPXeAmwKKV
GmYp1eCTTfTdxSlpj/TveJJeNhACHgMMDkQ56s6GKFiQUCEX2uBz2iK1+Oc6qw8F0YyKNQCoPNfP
52g+e1+7gqYBmuO9Veuvml8YKHXhGp4G+Zk662Qri2v75F2ZZADrAEeTCfmaSC6hW/9LooxnNdY6
e0Dj0uMHS0HJuc5sG3T4pBHgpnMNdRQwA8y9I+QdYwqYE1Ze7YnPApB4zFGOA3l/YfpZashJUZQq
167vEKtDPfYuhzW6/blKS6zY1yVmqHlBYL7/UzSZetObME3Xvnly4meoaMreaF51Mky0gUpoIAFU
g4r5ZFFNuBBw4FPjCDHiBdwDOL9EUa/HX87Nr5eSeDBILPZlQbw32HrxjdHq/PVADHX74RczZVeR
zA7HhN6YpXwZ5mTyVSUNzKBmQ25S+zA7UI4lIxa8CuUTFhKtx/z5hr6m+ymy/IItEvSNTnWcakhh
hbVUz5jImEyIj9GxQ8PijEw7wjCYyfst4UtYEBHq9PSgqcvWWpu32jQW514FLeA2PYjG+M5uSL7x
tr0aZCdL0YDG69gij15AbNaiLrXov4pwAAtgd5JsW8ZRBBw6r9CMigJxcrohrgPYQgzp0SOVgKxJ
fVenEOxWv3rjgRw5ZLFsfDftNOMuoYUbf4Gg8kTrYaa7rqkYWgpvWdMGCp/VN+b+3J03QhIXEfBb
1ewCPVjG/TNy+OtCG8F4rHDq8v4lTyk0+JdJzZxz9+ijnYLZygp+xbek2nN4I5U9ogJqA1Td969A
vWu2fcPWKx9DkUnQdcF/Yv4w/Iz5van5xT3Hs6pgsl0pLw0QpcXztXoecmKiY0RImxHpHJ0x+2/H
xnQpXtZwz/hoSNaqy0VV9JShWx9o/YiGZ6x+9ZIaMjqPM8NAznWp8pwyVuomKg2QKFZU7fldLDCy
+2g+tkbpQAn5ipMbG8fiRlIrkC4HVCsfA3ss7QQHMnKm2u4SvD/MENERTUFxQU1VnR2TKafQGslK
Fl+hH7KJW6bUETgcPKQuSn1wOpiRlxcgPLktgRStp9jY5ketouAVHoR8E2UANfJ0+0a4tFL7UrUe
aD5qnapi3oUIGaUAmc1chPnajgH/vnSdJ6lwY+EzYK5LrKFOHdADVNlxaiPB9dCSrvk3CDbIeGri
p6+NAxApveQdQDiuFz8RUHv/RPl8YaSZwjhXl0Sd4oHIyBPcw4i0SW7smxrgMg/ELyxSCo7KlpEv
MbzNaY0e8GEV2xL71wBVGwV1A1lt9wPd1E+RQSFV2SW82xpel1b9pu0yaQ7DnGK/MbTcN1PrPmAz
vV8ScaF3NNxlHNBcXQJs+2iJONpfT0eNKqkEgLzTQeuL78DZXjQm7amapq7tYWq/1P3N1OeX/fkU
gFt7yqx8eb/zxkveD3T93F7yWg1VaLjdRob3/8+a+s3gyTVXO54AvGTVrdXnWaM3k4rIdbQop2sc
ZH8fDGch0QxgUf2FPEdxkgY/1dyHrnH+j+mcyV+JNaJgAxbiLnhgz62xBLXG6F1JyzlqjakVH8IR
1MLtIbgi6wUyobhHNsuQw4EGO8Qci74miHA6zytQdeRgfhVzeWoHoHYSV6azsxtjYpUcX5TKOZvJ
nAxYuI48TRuzCMw7cKCgeBGFP/agBPalRAgE9xa7h5qoiKPuH4TJiR5X4htGvLgUCOyWSIxvy0tX
2DSY5ck+QFUtuEEesuBpisTdTU0TQA4SXZIB07OLAOFMbixCsdBWF2lbyE6+bgRM5bLU0kjiQl0l
ioI0i19bM2P1tTZcpUhD2sPJSDP53K67TpkA0p6LJr+WbTqNKsT6D8yo0/2v5ikY2B1TKDJ5BjKB
LezxYwBQgO2tmrHGnIYJ99K0L7omhy8CUaa8ijH6do/bQRB5EHtRXdOrdK1eCn/lBrul35NSKNiS
u6uHGdusCmA4naW83mX0DLXXRZWrvygbqueT2o3BDg2lN8uNOLDRodVuXxcvAMUsUeZ7CyhYo63Q
ci0AIKjGRH+q8dIivFpGQFTB8IYqSyMPr3QL4vE788XFllsocpIjmP8TrYnFk9VVtnVL5Pfk7pqh
QSXXk78DqXsZb9dji+WtXkBgVAHnWGKAdUsMTAESJWQlAouaDHoAsviAJ5Ei/6GxV0GqoG5yjT+9
JJyT2aU5QLmOphB7ZuDDLAnwOZr1K/A/YolIJzW8X7KhQ6AZgPzHmkABAXxc6nXMMsdCFstKqSTi
NHf3o6fDZfZPAeY+XLCPBu5ImTIUlz2rWsRqlougO9lH8pJFd/aHEi3ksj/zOtI4gKlSQBnp/nCm
RiiaYf0Dj2pPU97JY4LnUz2M1PcWTqjWmfFnvV2c9vwuuZKb8DNcp8bqnvzRXTpKIboZucjZ1sK2
a3lbFhBkW9jy6sj6LEKH88ReQPiIsWRGpdq21eHhRQ2ZXwfs8KpDH2ti2v88ieCpmiNW34SWEfVD
l51zufJv6V5G5EERIWfC69vUayjjNMqf72wJ0FaZFN1Lv2pBALBQnRvJ4M9IyrxXZiO8G/D/sPqa
C24DMzZethi/UTzd9cMSPiorfOmNwTaHRy5yPgBppHw1zctH+P4QMiDMaQtMrq0emd0ksm9hLLba
h71n/YSETmip8MhJD9t3b6L3JTx/Ul95ErVB5Lc7x6EJ4gfhh4TIu1qnlvfC5prgcnuzJaZPmibB
30MRDtNAMwzRKTjtBlQWZFN7PDuZU8qw3aZrh/yclc7qoc3EFzKhPCicvZJAScxIIpStct5cpGZ3
QSqdk5ug6f7qd5Ji9RnrDGtZlIvUvWPesoxa2uwF6FJTAsGOZE00QomcWITREiG/jbD6ndiLPLnV
hiML2GCI86y/YppAX/zGz8yJfFn+9abVPKbCuxux9n+AVEmYBIspsyO6V9xnFUbF11DOhsT+uZYl
j95zWzWFx99H0YkcSZp9rVD2vhv1SycIbXzFPYuAU57WRdxM5xbLKmujLdISqIBr7XtsgTu2F3nV
h1bc+jhPpxg3OC2pVvRt2fcDjpk43Kr5t8X9maReAdIEY+AL2I5a95qc7Gxc9cgcSjKNDFL/ocIN
xt2bYt2FLAkf2F9vc12ToA2yPkabed3Wrah9p7WnkLAZHCRX/syZ+pgSOBZ4mkYejO0Ih7rV0uh+
2Pp5qzw6tBbX32Z2ozPt89EikX5B0ETVxCltc1BVji5QbmUU/I85qwyU7MBAC9E73u4lC03knp/p
+vY7EXxlEPkmFVf9r76rRcIN0lNIXrycWz3CciiQXLG+08z0a1bn9AJ9YUyslziUwTbTUp3sGhBB
ceY1XxKvBB02v0982V/W00cZX54UyJyR90ybjGhDiNTL+aGaiUrbMBjWCg4uAx5Z5hyCThLc/NzX
762L7CJlUvWD+CoqI6iyTru3ehHRUvKXK7KpoIuoMGOsvU073smh47IC/RELV+Ysu9qPZ1w0l6o6
U+BoZxE9Mu+qSKsMC2Xq3etr+U0MaduCaXpp2ezRc3YG1GeJs+BZQX4OT+A9zCWqmMBApSmsyUWb
7Lj2oKTzJ0kFzmaXNmnBub3LFCA9cXC2PmFBBrf/7HV3Zw0a63zakHbDIebcLXSLEhY5/YJxgge5
lj2hmoAcR8/kH2JSgAP3ssNpMQti5dRGcBRBujcWCCX/KMVHTsuovvkz208/r6Qy6rPsZMQSL8tO
f4gihz3tWcJY+YFSsg4T+rMnqHCvzNM8r98bITNugX29sM2V3alZoXqjYzUOjv8UdPp+7nRsmORv
c9oW0+h3urpXUiH8kA0FQcrKWwAk+5G161Ai3Gk0qFmK7cLkaMZ6LnD1XzDIv8UWSkTy6mKXdhcz
QRFsfFn9ruKqHLIwaVEEzKQGgXG/iF39XBA9Fnv8Tujoeitfp6hL6RgCASmGF+/xThlD8j+1Hx+w
KQ7pwY2tXIp/8fVM4ZlCJk82YPVK6v3YF55BYPejDRD/+/EAT2nSg78vSph9q+RPnJ/kzipvoYsX
9LCnSsl+w9tG6IOkl0YceeukwHXXcHxC997MQCOGh7AmItCFOvl7FM0GHoO4Nwf+TomlH2mCXy5l
QWHfthoG4lAibtD0aSLKxseASpD6OMkXmRxziInTA/Bb2ltCTwesYP58hrKtLqmS/8gyizil3qyn
1jgOZbt8bzhKes5i59Pfj/WHJ6EpFrGhI9TdXoywLH6uqaU1x4KRlanXTa8eIXv93xYsSHesY1n8
3nR7vWRvWuwJaCDCKFe8mk/2O33AtOh63L2rA67N7nKCSRwSp0aZBmPmHFrMYYgwlP3TgQokw2sB
jVVUVjHaw/pdMHYzJWaSQi4Byw0qy5RBlGqgHhAtlAiFJ02AecIHLy+JpiP6X1UoM2MCSB8v5zyA
r22wfrSGqYopubKAf91EVED1/fNOT1/Vv5jb+ssNyHxw0IxPRjsBtdpgiDwkfH1fmP1wbyuDM2AG
XnvbyrTMG29iFjajWa2ZHtiwEMR4fXkT6lhkCICqrUFO44zclL8RcblDZ+o8T6awGAQG+0ury/8d
dM30r3OzMWOwSdDjLs232gH01mO64KE/bTC6vrpY2F04fyabpFkavBdc4VovDGvxoYmZFkFL4bn8
7o6DZ6fwtIAbVWT3/v4a38ck4iFRLQHl7kfiKBl9vAu2U0MAKXCzX+6rzohsZQtJlR1UYyXb/p5s
VlXujlksfBCEfzTenCY3yT1NIZ6ADdlZsyklJ+rR3PTIH9pJaKMrpmmzLw5tBkaOUYFK40rnrZru
mxeVBsWwuYXoJT+gnUvX7an5aZo9DLyy4W3OjDxdmHbwEz4v5rEaIb9xZPtJozMlWyUYeFLYKVr2
0cnRW1flrDFtn1TuVl01fRmjwNfpVQJdM+8prnakUNechfs5Lj/LnmHjzRxcMyK9GvexnZ/PiKGn
1Wwh36fpN7B2cb6f16lORdjbA/Z/lC+qVhtFKWtzpua7RDAAIZ36ftrnfYeZC8SfLv/tS/xccQwQ
kEeEZPmBHw6TEO8vpm0EnErfHatLeF7DVmGPTn60Ver3cA4wDL5/WTQzlPjXWSvGjFwxdkDSoxIl
+p0OviIWfTvS8P0qRUpduKrSAciVSr06UydvHoz7UWyNdSlAqZavp1Aao/g2peaeGn7RkeIF+y5x
GQjViMrh5zUJYeDAUCL5rC93YjIWUESRpniPYVgsHdviFQhi58I5YD18GIjALgWqInM04jvu+gYZ
IclE8m6UxuuC5WEgkz/Muh4CH16Mpr5rYHU2yw07/0Yo80037IYeCZsfTotjmrApjw5vxHbKyFoc
n1h6e/H+QtMelJnE+0dHq/7lanodaNUE27+lEGxgv0iERIRkj3UAs1yjYhar8tC/8Pt30BtQiZWO
b5duiQMl6Zj8l4UG9thfperhfexbbdvJwgJaaiDnBhnU4SxS3RYgz9zlebfZ7m4g5xEXQ8ldX0wj
2Gyr7AecRlSBdIANQwCVqF1WFTtddTlhq9gxzIR9KWm2bofO0y5kkS28sAVGoqn2ftdn9qpBrSzc
zGk4jugSKMTFAAepCLBcWzQWouYb/k4Fz5XxU1D8vMu4qEqTk+DBXKYumc+FUtrCWc+tvd3OciWR
KVIAaB6bicosOH9xPEDGIwAhiXLUOOhhTowUU9IQKbUqwR+IIiD9XIIOKjhdZPGrm0okygfA3AaG
P++Ik1RJ9J1FYyg1KK1wm/Y60VdEFHNpVaBjJzcmXn6HHL0isA770XivBFbHYi7DUkgUnLflCfYP
wEoIpW3SMnL1yCC4c04KncdmiwPW0TDeEXd0lZlXecBi8pyNJbiFWV08zFwI4ZIhXRsUZLzZGJgz
P7FGFxnNpWkZUdr89TwUSNLC4AhBGMc6QFdSqwb4ZZr5QRjXg41A9NqOxhL3kHTt+64eMVWMBKJy
iT6XChYkZZKVImc66dh/Db2CI9MetDCt7Vsi3DfXB2+/Y74xFu6y6ojVwcapfzpa7LVaEuD/0QLD
rR9hcig9qVs/y8pCCoMpCl6g1nnwkExLaBvft+E1HT3dn01MMrx75ykDmOilNDB57Me0kM+CSw7M
Lbsn0c9jd4SNEaKq1X3t6LJi5JlDEbUyIg33tfihhRq0pFKZb9c0iXgWu9X7/c9TzgVr/Nh8loQF
RZn+/m4Fk8ig4CkwiOrCcf8SvpVRoDhJtE31SVHoevann3rX+//OfIibG/GXryZ88yJnY5JWVmop
FOeDwLZkc2Thzvz5G6S+7AloES2owQSY6/UyFxolS/78QRkvUkBJl/TRIhB5Mnck3caeppcHb1EY
rPunyQ+jCKhYk0PbDplp0eExHQRMkuh+NPveVKr/irhtX1T/vjfY6fmFN/4hFSI+TPqc8XxVpY41
YPrbxnRjm4/Z+NB4SQx7q+HvIMgcQ0vLgtLDIOskXEKOYfeLm2cmURLpGp59kVESjkTZqEW9LOJR
FM10xIHDXWX3a4S9SqewFZAgtyu/apQ7+Jt0Xj3hYpUoVdEdbPCmhue0q2vpsCv+Z3Qb4btiOx/J
KYzTX/2SdTr45b82fl7TJ5UdAvPUGNHipKXSbB/viZvcyLKkYYtiVn1d5TH0bGjjWmVtWJIXhGAL
NZTSSo3SNwxtbf91ogxGAzMIxTaFcrOMmAX0dDa3rjYW64NBlsbeEx7PbgsGMu+bM+EBbviJ2E6Y
c5xH0I2Ndt8ouich8iy51BhbOVNlABA1WAaeiw9arDe65tUDcqCl9Dgux2QqbvntYHWAnA5UWKIW
xPQ0mmhD50uZ9HtwYiMvprEs470cxkHQ1Gdpg4ekhVP7lE+Ia8SBnIuhmk8PnunSQIyKx0eQG7fn
u3r4ZjuBvddaHQVkzuSad01X85f8QbJzQ5pyVCm6kXPI+74GPALQNAGy9RwZxLgD7b98FYhNd/0F
fSTWwF1kxCbG/E/BYI/Rnry+o7YZeXxS4gj2dcl/PZdN35ezsV22PWlNFXRa6ncegp8SVnixrkNE
uAOgYEL5CfiKSiIbnqj/ja9geMs62i8NdB/fUjtxipjiS0kmBdvJzFp45mt0R/e0U7BnQX/poPOQ
FriUKdt0nTvri5bxqBGXyJUMNs2F9pXr0uUo3DctuLPsLjOP9lYNDk6mYC7wOFptSHrXWI/Awsux
8gyB8vd95ztOzpC9DvDy0AjEZZeY9PXm8thjpYmB4dBzHzfg2XgLXQbXU/PqDo9PFu5Csv/i5NZ7
hrtzl01cmYjp70JsrXAJiqc9Hch31hdmYH1jjo4GeoJfpd0RLVwuJWjbnnCuoNxvo9D62lhXYhKl
oaImNAyOYGaHPQ91UHlSZj5xyAn/CqBmAWHmV+6p8EsCxAjH3HxUpfHdV1SiLPZQUlU1umR6/FUT
8ZronetXvgx3RN3fvm04oJsyaynRTLvLHDgdWMTBkFlTbjSZTu5feinOu/K8nlJ8hWMnYtY9DWeM
8IKBhNIE0O9p7iOC3VYzIryuNIVhzN2HkxiKb4mnm86bNlJeAjcqMLNiWxFTD2JLO9ApzXegNJY0
1nLbhiKjJTav2iaD1JlZFCXsMsxuHScHLxAWtDd5yXmbM1vL/rMSWSKT14ZVggwEY0qqOy3hHYCH
ZOsP5ikodUjjPtwLw7MB/58q/MIUbEGzumsLj8ghOTQWluDTuwvi7p0idmR9WVMuRYwyDGq8dzWC
YchJl1W8V838p+PROgmiRQCf7xffQIweUScl6AHjmog7HHgcAC3HpNvRyw8wcqTrv0giw+vdz4bp
zD7J0DGZUmE62Xxqbfx0Cbc/D8jb/HsFIhcZKmAa7pSMBRNi3BBHycn8nPNwHus1rJ/wFrFlg65B
0BrkfXA49wW01+98LgbCGUVLWv7yOTIdQ+a9tnpxTfZOhMLE/MBUdYDGI4q8l7rUnONuK9fa/JxG
msz11VdUzv2RmV1uBzmp5pn5/UvK0+afTAGt0D2+SEVvifi3GcdlEOb2khLwg1iRD+GIg+0IdDaq
Lsc4JxP/BA8FDrQeo1mb4VsMNHujX4NJZPn0j6gSXBePJ0iaFHzAMz3ceLj39RmR1v5U6gfD2awv
ZznaVvRIvmEfx6MDTLsWVOAXy3SjK0KLMDdGT31m8VhKfLQBSR7aNuRxbPmZgOlY1bjNSuK98QoD
QSxpl3gnKNgFfx1uM/Vqmg8jOoQ6rRg81as3v+3hWwXTc0faT3HvIjF/WOoS4QWu5bjLqMCwMat8
ioWTsIWXivMG71r44l/5G6OpdFIIZBS28n/C5/WICMOQ7FlU1DTLgoihs+01tyZ50EOfN+HmBT6F
3XvJsUTbtL+hlFfR9Ce97vQ/skwdriqGh6kAMUsgsXuMMxcqRtVLnL+/m7VLXslV90MJJsiZFb7x
PU0DxmKI+996U/erLt8tF6THoW8JrLsfXYVXqs7pKioZjKAGBKioWZZZt6BUg6yI2sTDtvopimVc
VHC9hYe4/UUj4MwKVU2dREHpR40fW7O9b/00VK+iRUYXlb0JMjKna4u5h8Z7bGGvBQyy6+iMRI6L
DQwZycS8YWvVuyYjbe4AzzvuXfQa0K8n412DYRxgkzXPD2EY6VdHS42g/DZe3b+BGUz4kCwXeJrl
JWXRV2y/PRFF5ny8YWUJXFdGr2mq/fRyhxyt4vpe1keTlIOjAJxccANoGFYXOzWlHZDrppSBrQuO
rbczl0b/p8m8igRw8FGMZUikrewzwaW/Mah47Bj3N4Tpj2A9Jhx/O7H7YoVp4Yq13BHUWJ1RdFDZ
xjVWvK/6cPaTKAg5OSkOIbDNowXpstB8OfF7MiFrIa7WAMmQ9kwOV4Q2/PTdJJw2fNWaK1FO7QzO
Vdn0ztJ1H5DRy8jXoUp10NXHFiW/D6PCYbBcTmN5QeWLnrOyzOAdpYC/AOHItznitJ5MYIlbLB8d
pSAE5qEko6v2Xomf3nC8+72FhB5LJYfbGbSSmf8sInGmmbn38C0Rx80cLmOWiA0jMyR41zX/oR2L
5jXL0chAeZifJmVPSyp41A9phUqRedKnDZdIBid0H8yAEwnl9yNxIQDF4jedIVixPzQc5ItdVoqO
afaDBICAoaQq1K1Iu3ZmBuWZEZRT7CSBmc/Pmq3SHUwiLfI+grNljUd8EIOpctrpYVcilqlBTd9N
sW7Pb3BT2gsFE8BhamHAeUl232y49hdfProeUZuiZVH61irDiWQYuDDNiWZpquMMwKFsd2oDZx/b
8z1PM0whShtes+BX8pkq+JshnHz0JYDM85dMB+7zYeDU4uoSeObVO8zIL4hJLFGGUsBevNXSY98y
e2DY1chmM0V+KLqRRUBwaMKga5wa5zNAq3Dl1egpiI8Kr6f6s05LrCttDOQFL7d/tsTf9a3cQqNJ
jQRwnyXKC3aZBBOldtB6Z70e0ap2bkSfSHT0vc18TP+p5Qcu7wOivfVdjDBniOvGtpO6SJ3cQJuL
eFhej50kKBAIYMnGCWYfxqFbF2gNBrYgdjxQkp6/+W0S21h31/+gd5rfZmFixVudI1tq9GwnzSRq
cLi3sqd60IeiIQMXPckW+1qacnfqKYnT4yy6CPtQAiyVl1HkaJeZpOILl28Ncz8m3Vzhf6XluuAH
2TpjIy/rOayXH8MJkfhhh9XF5u0B5yAneZ195JhnnyJU3M3dIT36b14zlQlzGkSgZ1W8BLP9pQN+
7f6ZEym2vZV9CkTiw7NqeVay2URcZVTXZhKkgAbPTzekCcZa6LS57gm2eVWoiVxFrncHBtpKNDe2
K1i8//RkPoDDRviVuEa1eBhlkDRiOB7vT1kyxeJb1JKpJZR6PmzCYRygRaGVXNOKSxSiaIqAUsXa
iKzuyB/9XlA28MTzyBQ1LYWovk+iVqSso6Q5cP+S/HBtMDVmP1J5HREwJ90+V8jzzypFJzwvKHo+
YwyOdIek+tnPFCebfxFiGI9+icOp1uLsPc7QGSrnraBEOBGTgw7mQB1hyNM7mCRJe5sGGz5wO3NN
+NcgkLzZbZuIB3jBH3YfMlAyJ/w60a3PXrC0BgxSLhNbMzfZN20LiT6JpB3qzvo5FqTspbTZKR5J
w7QgSp48SEWrJA/LvD0IdZJEzirCRb+vGBiTzNZLF1PRh5xpg2lKI4fwbijVPtgBrMKSTmt3ojsT
FXV+LmS2asM1rY4uKJv/mvb4fRqJtsBYcjD/NYDEAxaOsGsDcsVLDP7aHwgvvETrWqDD5BsMvE/e
E1dO6YtXcpLblONfhXiuox/83O04HIKzHvzHO2uWAOEc+EdxZEiFPAi3jJiLupb0eYCoYPrO12hx
0p/yfvdNAZtXpD5LibDG5aXH3JeIxx+jLh1wUpOmsuUoHH6Stg0HAma0Qm7p9LhktRFEI+sY0Vbe
84bnRpPXcAPWLWqtzV9WiYqjFVggdGojxC2+401TtZsa2FZCM+BFOHvBJzJtzmKYas9ZJRphMlOf
XJzfaDJFxDMP+euNxB1YQw67jF1xb79+fMrRAJh3zRzUghyvu0JuPSUVNx6piec73dwsF8atSKF3
TmDJjtY3wTcyHyqGdbUf7vKKCuXYTXhYo5VresMRo4qWqDeRk7PLzKHLk03hjtNKPefw/SVdUq0n
6YiAyvr4lxggaX2qRpbBq29nwM0JZvFcsKMzmXVcDcGmvWEcKZCOiWFm8Q4m6sfS80pQWYVx2oUE
YQH0dpbD1fmgTWY/qT9cXAI+1kS4dUukPStmMC8fxKj4NyLEnNuU1r20F1uYllE8ju2y3LZtExzz
eJOoBEaQ9J/uMGC7eBjcSxEwnQDU8mQj4KgD5pIDAwGimnmmgmJ2lF3W13loG/BETHCMLVkHfTDz
i5pcK1XuUCV6EtdmkG2/OuJydtokHw9IBf0jwROJmUZFhezyomeKPhrRWNhK7fb2BgeUxl63sar3
WsJep5xGBJY+8Jnj5mSS8HmrlFtNb6y3DiMDaDxW6siyocEM7rOCSG4x0MBjME96DWajLPP8d5Qa
M3j9BVFRy+w/IdYNhw+xDLNpY4A9P5hiP7RlNNlg0/1MFPUs6/qdmVbYfbY/L580No1PZxj1uTVB
GR2T/t8K8tuo/2PT4eH30jV6HndvTkuh7wFiZZBOWcfsPbMm5EwizeKJR6cpq1F6CwGyIitnmayo
A6RGbZ5HmW/ydhjGEJZ/Gs905/S/q3/OJ1ohw37bPosPe3H3KLW8eoVMLrpTWdcixUpIqheMVWMw
94Ia5tGrqS6m6oBBrZ+672ZWDr7J9CsDuKynaPS0IJaBpCqCsFw6T5nBpoCgceRKv5SRgsNWwDVC
rCHmo0Fif8Z8cGFupqgysAlKYPXEylXk5VVJ0ETSJxBurzNqA6/fFa+/L4bCA9byR0HNtgPt0dzd
ku3nG2BCb8WDVuyQoyVSfpuPbjT17+2uoBim8uo0geYyP6LiN1ILJ5yRVDxxuSBstJq+HNjKZWhd
3jRlvoevCQA3WjpfNz5qbY84VfdTV+LEubUIIuAdvnmSXyHQP5NHug+0VfcMdX5kV1VSInZWvWxF
N+0UwIyi+FwMID59O9iKzTSWv8Ai2qzKSKbls7urt6MkuJLWrM6MjTQw+hCk9LrIzQ2sUMSyai1p
5p05gP32VtLO+lyEqoZyhlOS/QlYXz85P5SwsfKZ58+dpvtFLPI8m6BBZ8IizB6YYiqa84aZjDp3
RVPixBTC0PXp9Ek91OBJuyegbJQ9QYnaW15juyUZofBt0NfIO8+tDCkY5g6gylwG1g+niWwciOSo
0m2pVcFUrr3qwOwRjMHEcLcJ6MsoYbbAG+oRfYzZ9MVcc6GZv2I9A3BzR9bTD10+Rx9dPQT1mNAi
6hmrsXq3Tptn/GnTVdWVcPhmQiLqeVT2F81Yjklde7biQ4ueMzbfh3b9yDMG62quOzUiexVklCZo
Wo/GepBP4AULGaWd7X5vlcYChvDB1KPQvcBqtVX4SfIf0Uov8s29ER4v+OVrlDw0YDClxaax6GHU
vwIg3SQFIxiKuMIORu6ZqGKGFfqyVhsOxx2dr++d+MnSgTq7s0wLRqkwSNQK7VvRQJkYOM3ySYdD
UpjEVAkkLTa/522YLoMKPgg1xR8jEyB3aiJHm/i2HIvXymUcEyLITSfNphIufUa45XeLAf+YyrOH
m8FHO8D4k4AzOvOC3VIFvQTLxUPNmKjfCfILaW+6lmPwG57HtZvXHT75nYZ6Cu0nymi4TEQY7bAc
ysrJfozdPezUpCH/ysx4se0gI73DNZcTtnuNtCnGQTV9Itg6j/cza4Wa2OoCJOeBPHsLAI9eq1ym
NHfx3efaHBC0+oHe2Uel2bq942q/JQMQ+OEh2ztCivKj8OE8rW4zScg9ALNJ1kYdWAx8bf55YEED
Duup/+BRzVDdc3Ytbdr23aq7vAtC1R+oKSICgBlUTdAjl7fPfiQZD/NtTTaXMLRugLlTheIOz1nd
ptcx/gQ3BaSVubdYKUEJRXn6a7SSIcuhL7nr5gve4Z+P7XLVhfFsbS6OuT5RLE7ceqLJ/whSdZug
fe+GJlsaHJFyqH5rZLid7Fu/6yA72qsDCVRz6nbpjYo0Od9IJ0d1hR4uBKT3G4h/HpR23AvshV+F
DMIj/+b3QuNBs96BFE8jqu/x3pcr0sIgjljYy0NkHRlDBQmUF7YXU5m+aEHjbOkCLrjDFr+sDria
6PqFJ7znMK9DFsSTbVRUOjkBWfUtOcYy5gXYPyKs26avYD/tWhCGkOnU+1w0YYwOdRqtO+S2YJlu
SoDIlWiudft1u11BoCslBgqLVQTxc0RmCRcIzSeMn4dcFjlo8x9sFrH0sOQT60wyP0AmBToolPvK
6+iM3ibEs5DbNEQcI8jAAAlRyeB0xP/lq3pk2CxrUbrRvr931NqtiLZY97grskmbQqXfm08gm14z
WQfRc/6+N8fYu3zQrIyuWZwuQVDMLla/DWkd6eBJAzygBzXfgEY4xVZzRdktA8oCSWYHh1TkYJZ9
KHhBgNS2LqZ2McFFFHb3NqD11Px/3jW2x8awgA4iA/+E/ZtNUC6GmQJwXKAGVSEf6Ac9BDCf5VuE
TeAyorkYqOA0I90ebcFX2BXm9vSnseSZuAWu2Pn9G9Cnton3OaiQV+z1xqBiyFFMG/IfpSaOb9oH
3AYetTqUfWazMYUYhcV0H5VDuieNRoezY8/0Sq5h5mCdzEAgWmsytNIaRAs1n6UwH7Xg0gOgz/0N
m71M5cWO4QAgTvIeQH0eNhMKdQwnyask2SEXr3up1sNtQyM6GuXEohtantKDcD3tsmMi45oW3MO3
VxQvM8s6uPFVGxe6yUzx0EImjt5y7Sqp0TftCh9eCE9fn9k96izVr57yCR4FrmsLY9i3joXbONYe
5VQKdw2xt+FyB9yUgNNx94qyvaEe/sza5qtFYsREVkq7rFR2S14Lh0+GciKGHB4T/oEuS9mg663I
5/yL1PLxufHoSD8hcDxeG5rNyTYySnp8d4W0Zk3Uvp6o4xfIoHk97qf0HC2eRJFwAU7V/cswAibA
dFXldQmC02VmX3S5hV35fYF1kz7K6P7IKICufG/fP53vMPooJuO57Bes/D2J7NjHnUUD8gYjreqU
/dLulNojgJnO/BFQC12Zgu4n9zrm0GIlEwVXtgZgrlFOQqaRWzjiLIL6wzY0tbfNXvgRsj4zdop7
MtufIk2BkjOjIJiSJIE3zj1PLu1ntzI/cFagLMeC9HhcXTPashlHqUZGN6pGQc5Z0s0QAM+KeI7u
1RGYzNq+eIxZSJkDu2WrxcMhJgc5+H6gRZ2qekAj1bU8J92MM5QWH6ASaFeCNOctnnf2KIAaRO1m
b0loOtBB8U+gMt9tE2ZITqagZYPjuW/VXZeaCqjL79R8+KU91Oq/CNY5PfO4BCSHs1vsGJN5vBoL
6gr0AzP0XSj54XVv/E/bJCxC32EKFGjSI8oAHXYFTfKjuU+1GJgNowYpXp4OodJEH4Q45DkAqTNL
HRIsfNWklpLcbemM3tEwFp2Vo8qQoj6DLfX6j5CA6asrfIZLujQR+0bB4WB3fdWNS7giNf/tiNiQ
2dWZdoTEbVTaWO4y+y2NDHJf2BS+BMqktfqJliw0FYiV2fGjBNlmNPG1ZLMnKn8YYiEiRVowimzo
mZWNDCEoWjhNA/hLduJsTDItlXNCQJ7t5LI1VgcETinUdEDlcuA2r6PKL0VjNPMmOkF0Ozu1wvCI
D3IgJ3sbyjRis87+XDHP23ByFZYBIfIij6TzUMSLod++QHp0e5ad5LBWsdVnHopHlM0OI1ByiPbK
GRn6Ii3o3L9tI9HMu1FBb1Sx9RY8N0Yfo/HIpk/KGnJS8R/0jrNQz6+n5CEv389SyXMbXRDT2810
2KZJg7T1Dx4SpEXBGHKKWgTtzRphbnCJp/D0uErLnrCIcwxrYkbRzHIG5mF5BuoOyQouKqkf8DPG
cIvDsKQ8ZcMBtQmBMPbCwMripbaTHXzHxd4xkhLgpepSSw7WGvvX/nORG7uAHYq6Vax8VwifuSGU
i/mRutL4LfgFQAmoIAWTTxV/Afhv531Jiswdqruc5NtuwJWZ/HJY0E5D6e/46tIviwFd14RAglmy
7YPnzHwXHauGm06dqjOGsel6bgS3BAMlOKHqs6tus2bdHnTq1ErCkMD7wdYFbk6kS9IFwtzo+E5I
vNCDE93FkPBM0A352WGWYFZSO920hh16XMy3iV1Sz2zP/RBTo1NAQyzVljtCFR1YyWKSvHf76Tmc
+tVHNVpy1BB+Bo3qDEGAVWHBLgERJX+MT0bbsbFHr0DiTxqK6BZNjucE29dAPtToevMtbA7rrUdd
GDyAUVh2qgsoto11rgyuXnsc7wR5jQiD+gzDElqcZZtfGMRm3a3Jrgd4yKYBfJcqxaUJd3sIjDFE
JnR88vQiu9xW97v9kpOLtF9ewqzkCFW5xShiXzATE0wOgPk1x5sGpOtIae0n+CPXXPALBZPfpFSI
7wzv2h9QPtjSal2XaXTgLssoXRRuQHwixQ1pEyeCZek3VkEGNoJzvifoehTNlqeLShLuiJ0loEat
dXaW1SbKw7lO7lk/8zUsOvCeOeLbWWCYmB3oCat+nZKvJ3UAh5WYLhiLpBYlOl70e1eDIGnDZ6z7
CSLSXFtZ38ny2tC33XVz2Q2mwIfT3JcnL6oJLYn1HmxvybupqFGpHCPK+D/trXE6ZmVcvJuFHZb1
D1kvgOO7W0/Qlf9wsNghzwU/52biXYpMlMG5+5ukyu+8jfHWY8uTaAoVLw0mD8DOrW4pIR5c6CqN
7pG4N5xkilkbQU45xt7DxBNk+iCN06rJAQVjzKntOq1VPsiVW41qML6ibOfL09IIB3hvkgIdlx9G
joN9rQdWqCSB1lCPPxe6iUjBFr/zSnYbGB2eyLQhgu99Q6dP4w1sG0USeWBOsVIsLfODqtaNIJYj
QQQVzS8U0TsSUaFNnc9oe/09/hNFjc/ic1bG4NKB6vcyQ/AcN9NK8Dw/SE6lAsdAw/FkT4InD4eR
nyM73KHXLS9jaWdDxc5ekbNBvlfUTz+mMXw8BQjlSbM9XKFznjK+c0F2eCm42jgyIIcX9jtWtWlO
ifHlzBAazME0TPT2Ob7MwfzKypjOohuBdAZN/Df5sl5CMc12MJn+amBlktLKnzPg8hu58DS0P2Ed
WVczbw6iUQlg38r1u1/hRPTz3tSNkqSFiUh41flmoTO/0udjHiC1+9tve3SluBET0hrtFYyKNNTi
WP1p5VMtsbJnwMG9j8ZDpM7262MdQ5oX/NkSbaEI3kaE4Obh3xXLMS7M661UVD7Vp41VhBN/C3nR
WYwKRwc8X+z7jyH49H9dkva49lPKG4bvRHxjbbZOUSLnkbmOhRRj9U739ls005fyLDFVhErQmX4S
lqaVOGJ20ERJmTOaXV/vOGHWIqamedPcUgaawd31RGGXbFsTqOlr6qnpu637lbSAa+qYya/47DRs
k8r7XmnsokkeSnRtQqlofl9oBGbaTHemIKBJcQ6pE8DxuFzgdQ5scBdkpfw1uGg61t3uNT+BOC88
VL7kZ0tyCeLCdfTIMefUNUEuHXGwH9AtRa7O1Mu4kI177LFxra+6wViKxhfQwl9Q8nuQko0luXmf
XcbVk0l+PaEYtEEd3ZnarcYITbyS2qTqJQ6kvehcqVszduFOt2pVg0B+5jokbjZPPWKE79Y1/j0p
bET1BUNnR5O9JdS+tCgJTnoMqvygcwNw+DHyS/FD7AopzntEAKYcCgkOoUQvJaXGntCaOXq4CM1N
cRxdpKDUOO6nf2yqZTxnSamG24O08ruThXmcb+hb2kvIn3wuOW5prVuBv2LHedp3IW/xlzhM70y2
+MSh8nzJEuYfqzYT1ry2cSpkRIfeEZ81wQr520Lo/pPVShedMztIARiu2PgKEo70u1GcEdb4QONK
/8X4yyrqM42kRg2wOxDfsSK2sc1FUhNZwhXzWJhmrIKl8z7v5hzjE4ekE4LYpljCXuY6SJP8dTDJ
6M8eBFwKeZNTADS4056H/zGw84CecfMxFH1TVC/+r6LW0MO6UWW7tnLCPDhQCCcjfrmOgKMI1YDu
JtlpjYst4XqmkAdZhZX9zRxONcXfJot5sZl8lLrTEgbHq5rXmGEXxvBR1MY+CFFipW8cOdZoehfz
LTmmUOCqkoUnYB4S8C3kLyWDzna0K6IdotZWqJ54jlz+Lzh07FeXpqjwfmEz7prhdqJZ0DeBsubu
unYiHHhDJNx5rLr0piET2cNswdCBxAYx/Zs2cfWYS1HM9M6nrJG+TyRkH9MYnUeESFEesaU36I4f
YAmd8BzUcxD8ZoJ/qsgKSgYu0JOMlKhA7NlDCrFFNWyzReAYLPDms/cyOXmXJh2bH1obBw8PDyiz
EUQmCwnKe6/nbmXji4pxP0x00P6YPZSdjw94k85F0vCM+CtDaIGqqRoM9Ih7StF2oU4Xxq23qxFg
kUlu9vLtaTZvvmb38M2Jh/P5v7Q4798veIBzQ67CCL7LlXteSZcBCD0Ix32b3yfp/AJnjyVqIz7K
nI1MwVkL/zaiCGjrWXJwloLMJFXbRQLHtsMVHbc/voRjJMQN2AGvTy8U5Yac1LFJIGHq5twqqXWR
krJHqUsBng6QL2ToEJcAvmiYfeWnCVN16EjoII1bZNHvgxIUXhE/hr9HEhWWwe3UpXgHF+eMwr1c
sTpO7dQMSnuyrd1xldLj5cSr2x9s+VBoIR1aIChU81+K/ORwd8yU6OvcJca9Ow8AI77qbKtT9FCm
X9TrUEs4gpsUAYN+x81FXnHu3pSSWlfmYwETeb+mqOaaBs25A0hlKa4xnJKE7MrXckS8MEl/F+BN
TIgaXSQCJIvsTIGs5UQ2zBtFDrnY/GpnjtluD6grsAJEUxtOrosmktRYpJxbmI4tl0XCTdHXLpR1
yYpfyYIU+HzuoPm/B8f0HCYhTt4DgmUYbqfRKlfg3ZCa+hln9Eb3TAuw8t/ot2DV7E1JDHmcS1yP
ILj/jW0tjdxcV4hx2GerWTBUqIu1WWVdx0pMg9BMy6GR5Ox8magfhAyGKz7mbn/wtw0oSgXu+D8y
spCJisGPArU8N60ieBIojBA7lAf7CtbY6WIf0I08UqwOxJm7R9QncR4BH4YqftbHohK2Plh2OSZz
yU0wUE2abgm/XEGqdvrIH49HKnydHXoW6po8QcyjrEPSU0Z03K7sSNyudgd8d57CwV800hs54NRX
WASvDOnmdD+1DTy4EeO8CfHP80Cu6n1i1i+HznkrOv0DcQT/Aj6KMuV/UOD1cPatktYyKQxJGwV3
OptOGVGwW3cL1fD7IsrUY8a5O4jUYqbFgAbuvWceEdhWFAOjr1aeROnPoBNa8cHXmQbNkQ6rSurb
FNqZPWtKnwrJrMMSmDK2SQX28w+2xZ4+DH0OPpoqNRQcN/uB1j98fR8Zsv0+OinYscr1kEKPE+ZN
VDPX+zBICdQCnlOE6ESsCR7uHelsqJ0jfJZb2tCdHLMhEyS7YM6tGKEuQnHAMnSEcxCeLaKawQGJ
aPEMGKqZSam3rk77Og2kk1QgZfP6TURVlbk2lUidtk33qEu0X0mYKNCu7LKoTOAIZJm3L34/HvRw
MP0kG0NiKbBEve3jNcKje6iJYYP7vpXNSQ4Ti6ZZdLS6UojzJzglOK6k+zzBL48vLsNwxPMZZo62
eCSw/RmZYn6qQRhjWTTaUo0FZu2X/VSeh8XLjzQyzaJ9haL9Jpnltlim4dy7VpEqa3SSGOnBM4D0
vi431D0/k5BapGH9O1Ks/tF0RZCmn7DDJSG+TkP+FOjF+4KjtrFt3yS0n3tVW/p23w3S8tGxwstk
sI1LyBClO301SLQzwxEJ8gV+o/6nyYEhHgEJmMBLaDP1l3sGjVsI7dsjydfCjUqMo6Iujps+H4ql
bebie5JLPe3WmuKucEe60H19FuIUg+B0ehX776QYBY0P6o5CV/wVirooL2H+x+Yhc43TIXVyl0Jk
dfnMHIlH2h8KlN1sX3CUPkIPSY6DSctJxjCZEu/2Hqpa9lRJPVCDZUcPn1qx/ZI3svVm0ONMDqgI
Lw3ybwR4TCeb3UPNQTpKsM0gdMxNVQ5qQy8m7r11wlbte8fjeiP/mK6bI94d8CQFYmo4bduxC8hf
jYFNJsA8rwRU4qGHrYIkH/Y/4l6CHMzr2mHu4pjhTtMEKpSueLrV/qJn9rkjPvDTrx01aAcssvK0
SZheh8FdmXnSckw2iRlXUk6n/MyhNXhc8g1F8rCvIhtplwDGzHl6JkW4B91B6Eq72ncteuS4PcM8
RB3KJV1l55OTv1HJt9iAcwA7QjFJ3okU/gFI7wXFVsHzv3TZ+v9Fyn2jvMFc0RaAIvnkiEn0hcp7
oPqhMBTPwzu8JSWOXcoD/e4RjtTYkqYZxnEEj2AcQaoXnZwZH0+YC8R1VePpHRq1v0Ql2PALxNtp
dGyXiDfclWEEESWvKlp07IWB7dDnBW86OXViKKuMWbkjtO/AtVAOyyGQXuxDl2G+eS2mOmKSsGtX
wn4Gs10KoIUIHPXCMle2vpMGqiTQa9UR37LMcYTAM1WJ1IZFXy6FweQjQd55YwxGOLaALGhZSwrN
9Fn4ojiX10w/HE47LZQPqSgEzNT+F2QU6+gGS4JMNSlcVjgvbkP1OAEHjn8nzSt4WS8AxHozB4v8
0VajUgkYZSI+z8gwTF5n6Nldjs7TQLHUmkHDxCxxPYSr6XxgOG3F8TNuFZONcm3fDfu17S0G1XJy
hwu0firsDgvrXnpIw/YTOTQczJaeQ1bRINoTg+KMIKLY1yrGXrTF++cCLmKHnGsUhAe++inD78/d
+ZJXNFMJaUc73e1GQU6aNEWlERgH0NAFOgG77FFJIhcudFcmPqBlKhZHrMacyVJjxn1I+zp0YBx5
UI5tqg+K4L42e1+BdG8G6eNQfG6VR7oYW+KAhzGtanrG0ZRXYAWIPc6gFRmBOazQ0x8Pl6Yhn8My
bPNvX3FQkcWGH+lHp5MkCsBahg8QAR4wOTWIuxTT9H2ESuXmGsORpk/mbb/fwTqBKUkDYwMCN1R4
ilkqJ1db1jvYHNPSFMuvDi2rqd0pmcw0wp4p34HhDbUZ4I7WaLsnGqvOVVRYDAI42nCCmeTyWjAf
QkH/BHa6V26K+39wA1ecLUtFtGJcuQY9dJnUWMfl9go4n1P5gCabIf7KDt4Ij+M2xsoUFPh3V9jm
eXDvZa3m4C4EzOsW0dPwVSKvCfFwB171siSaMD0j8dG/wIVMC+/8XSFiLCFfOiSsEd1fT7DScZXa
m8wSTpqGm3mOQBGN9QWuCiNwIgbvGG9MOIiTb1bwiUtn9yxODfmkSI8zENZQUABFlkhK3u/R2v6g
yZ5J70YYedd7pAUnz2+wcSYhKQzIkFkzDI/oVYgquHa2v4rAhjr7kMssXkuBGXRLDY8LaqsWDWN/
DlJ9bajxcAtcg1ErsUbjW4lAwn8CzFX+LUSKpIRRJvnmOpwcQs/r43+0dGDYJBAnepYWxPMfjJal
AAfbfRX8wADc9oBU9b+AfSqFagc622vYYmdjot1xflUJ3UgdMBTGtIHBXzInQJy5C21gZoFrjPtv
ygMTyWskX3cPNarbgb54GVbVDm7kNwigDZg8lt8NhvgYR+3QuTOWoTH2kQK5jK31Rh3T/rnplzJW
qC8oQ5tzFxmjRXAiCgMy8GvTJ2ll2qxJd7T0mTuT4eaE5fQ9LrFLBDQUnnhiyxgdJnDYBXLBoyf/
yG4aiE5FgrqLVzPed3xW+aoOc8vg8ky25i/Q2zy4MQ9kw87BGmTLEXE1BcICgmv27UJ4reTVuN+a
ERln8eAtU7FTniTWoTt0x+YjxphHHRlFlFb4y0zOpp3pjOa3pSwGQcNIU8gZw4uvrYdzOgu0uJBJ
IVg6xwBw1TllfcgNnliCsw30fkbUNBv8UbdGrief5vmvtSPuWV2/NUlBrSqv2MKtD9HMiD6Epra9
cUB1BbmTD5Q9zhM7lAc0ncpFM4M87OPWziIbL2qUNSl+NuJgHzOdikMOXzrUXRTf55HpJz48nAiv
gdTMe1uuv1wejlllW6FSuMJl9TaIDDT8g4vOIyyAsRGcGPmYyWpEiwllwHgdVQ+kyauACeoR66yA
8odVIo7NgMVN7tmhMoF23LHCG9lkuU6py9SHM4ljRLjikxuNoWwJ//r1C+uuBMmXQ3CdfDgjw721
iKSpdAfYtynifN9Pioztmaq1Nqp+twiTKQ5311lMSBQ2wtRxyJJkUNyVw3IUvXpRw/UIhtkZtVgZ
jrlZZjCSNSzCVVzokkocrNvaVNZPuRdGAsFVBgvazd2aNp1qxuMN/ZZIFJDBZqpyRGoMJd+Se3Kq
b6xWvfvcb5k9ImEEzAc9q2qGgjccxEQTbhPkvuuk/nUMkPwpc3uxbSX+aizNXf/h03kCnelKb7cv
An9KMA52z75oIzPQpK75PBjfiHWx8a4nUlfZjyM5JtOeZkkOdH6e1WFzp/NO2Hea7Dy6xrZ2lfxu
ogHSDeJDoBNaQ5xcX0juSqiuNViFjLNsFxhSycgqU2e8mwtDKGJNlCTyMhxkvzGWIzsfRKVSZZS2
QJ64hee5a/MlxVi/sK7yUjTUJPLLPevLwEfB9d9xlXkK4aVdSFtsKIz0yjB5acidAZaU56IlnwcN
2OP/N+gBDzekCogr9helYarZ082fLMuhjJl0UPGXHvmZO5fhr54qHTAAHG3tJge1qgkZQgx8jb6C
AuU9wrF1ynS4gbchCLVqhlU42VAE1AUnUWVJg8eMS2hI0kSvbHlj2Dh0YrT2EZh1t35to2PTixiK
BuPsiQAmK5oukw5zrQVVLppMUbsPN6dCCGLFk29yKBNhMoOZfr3wu65vqoNY/OQn4uL1Xi3NkbN2
FVTOnFXy+U8XrpLwcKYkwjxZJQ29njnDiaEgT5HcPyCWSRDd1UsizYrAhp8B43V4yCxWHzNWlD+z
6OkpGi2ARsnFI1A7OfwZXjfbRFROan1u+dKIsouW3h9kR6wGFxa2Uf3injyBLPznJ8gYr8wISk5r
nqovpNYoqUDflSVi/Mnjn33WWLx4oR5d0MY75KeQIMgi6khbDBdJlrol8lXOUwARrOsSL7h03hL8
TpdH1WsR1tSMNHeYrTUfsP4Rs7azYQVmlj/umHLDOvQwNvnPaNwewV85/k/V/ap3UneJaBDmwFcj
jiBq38HOqxl3uka3VbNK44mWRfDtDMMkLQIN9xkMqOs4Ov41689msb43qLkHKuz2rZWnVBVGfAmc
pE3Y6HgxZneoPYunH/FB0iZYDdDYNHrD5yPG43nebWwu/ODojb//M9VYRElLG5qdJFcrjZSIcH1P
OezZKzgZIlG41e7Inqv2dwKauUoautHgXxJ7EFfQUiTYQw+yljAINCDA7WJ+RWfAYAEZXWtnychp
QxYEHT4r/6BQd3GrEbg1y/RNoU6m7qOVLvuimAJDFfAJ1EV9JJcoEAWorKTb3h/UUdTD9qPuDwYh
BeuEP3piHt1SBpB7fU2Yjbk8GzsheLhsBEvgd9L6Q6/YJalvqZ63bwIC4nPl6hfEllwLZhKoUOaA
5l6W5f+nnzv3NHfuBiIahSgxa4PcMlOUFYVLui1g/ccBQZd8ZIdp8eiA1kUYOgHz7CAuBRfAHu9W
rhVCw9G6kLIopXmnFhAG+XUHyDfpHlSQj+o0Q3K5qjDkyLsLMH4kL77kL1ometjq5fK3BnspT/nm
wpAwYaRyPxyHzIlWCf1k8yWo+cbQLd51l8ujvbIRUJUiryDagJuJ2DgHeYRJSVksBqTA61gY7w91
IF+a59PIqixS21KhDuiArEW64iyc3Dd3p1JODBIrDaUJh51+QLpVn/4HEB9SZg5vKaEtWuYXlsZ4
dyYYOaqhg1gcpkPLAwq4j1IzIVkQZa7m0LH0Ta61kGkF5wBj+RGuflAYfU3E9Mda3hRaFzk+go/l
g9vrWmTmmNP+eLLHTe47Ahj5a5lfMKlvcf8Y64/7G9WMh//RGo7EpXkh9/gO+u/3Z0h5veq/VHYI
aldQ9GnyPAV6Umr9oxsu8DM0ZdlsaaoBqb3oOJbMAQF+KXset7NWxXtAo/gWK3LKbJ5OsPWVaf1X
TD83G3ee5HZJGMWWgDL2FWl8L1loOPC4vpMPbCUWU0se1EaFbA+8cJOhXJ5qULCgFJeMoekW/dNs
YgW5EBkOrwFOlA2FR58KzCTczyWlzGWl+UcvtuhDDaTnOeT6PYyphRxgkOMzj8aAPKnLNsuez+M0
ykPeVT5emWKAp+YEAlNjZKnMuZGs8iVP9753UgWUGlr/jV1FnFRZZ3nrCvEePG+LrKYriC7Oj5O0
yAo6CJqVN2id0Yf4h1p4UkmGMDEqp+gUaNVq2uYE9yyzWtC51Bv0L/JTKgdOXjd9LEjS7d/Yz8iR
7CSuXc4S3WIXxasH3aMaTYqHgfxJ9xHa+KeDMGwfgw/9guspw+wU7gL4Z01Lzy7xVmFKpxiCRQoM
hkREI9fQWc0P3KwQkHNDkBp4zAAToVOWGKX1zM77CY2CbaYdI1oleqZX0stgmMQ9x0sgmHQDeYG/
IwcAHih113gtWM/xbUXOcAIyCxxyPQXQ0QXK0/3XZe4jZKcCgFmQmxmbddQDLxvkcPSd42uB7QNE
X8cXVa23tUAYOmUxlTU31j3ab01cG+qjU8qFBL2bDyctjKr2NMDdsZBJpbag+MyofkW1/Bj3izxR
asZbx2LPErzx53ATCL3+wVuExkoYvTGJ10L8XWPuKU9J3YpmbhQCLKn+vpPxIxT6dVfLuG2IzKpC
M/nvseQ0YgIAuVTL3+r3PZBpsPV0T6t5zY/F4+vvVdqQHwjPa6M4naPvrhb4VXFhqsH3z/eEhE/g
tB5DItpyiyxE/+jwRqWz8cxuBjjJRW1N4jx56mpBiovRqmtyl6i05/0A45ACdgcEx7PHh3J0RD0f
493fq3dnEphg1YzT7UuNIaAqYJe9JlUWwxm3fBYhBhfhgtfuztNG+DC8ydHPG/EQZ99FcL0SLX/6
77EEDLLSHRu4ZrP54w5+hqYfAaQlflBiiWmcSjq0q6vqvejC1saOFmJL+OQpsY+YcrmRRjIXjyD0
DNbTacxjrUdkvQKZLYr/OM4Rhn1QwO5/5JTGURpcYoUawBw8m4F1QIDnyBa/yfOG5ZvlI+Uni9Qy
E2WEaKKifDuCgV/0g2g2GJn8yLZxNWNLGe0AWVcr7CMeLG3d/6zvOBTeLxfXtUVYAyG7KHQu/Ll6
4B+fky9oOwOj1dJ9J/0Xo4eAtKJd1ve14eupeDqmNKwPMyzuc7jB0QZ9LgE7h/swpUW8/SxtHM9O
DU84lz1RG05IeLkv4sfkBHkMctaYXjT3RUsOIruNtdpkzEX1sANVNpahUATVa6JsDudCnmhebJoN
cqLSPT3dldhZOkFl7+Is2aYvOqsS5EtWn3kQZh1SZycpACCE3wEIGtbMh5F7wCQ/X8FhzSJJPNTN
5ubIs1Nh0SMHSfhhujV/lTH77x1Fy7Ghe0QgcVYb1Dbp6zwd4puK7GBFqCdmMCGpXNnMNW1F6oLo
ecbGB0d33My7ZD9xHgwB9aCPO/4lbH9Sr3It3+yi3EQhLXs4PyB4qpyeKLtj0kJ/57GkCXyueQ1A
E9BpHgyL8rtI5ngz4Osr7FS34fQHiiI69xdcSUxvtviyG6F/mo+WYEzg5s0/mt3TtPWOa/vN4eUm
3TbKLcKBt+fxzCEV27o4Lt+eI0GHmZzuXnNdkbzEgz6VCYZwRfnIbP2bUcm8e6fk4eOkMHvVIeOC
kEUdAf+hqYf7mQE3IDXoxFrwtwEOrv1mLKMAWVZ+a9vMH7hVf+78PGVqxUZajp/oOeKQ4VZauiIY
fzwWejkHbGGrpUAi2qQNnhTMPZxOBJMuRgLmJIa2KF0456GKoaKZ7TeEmr+cza3aHy2ecu1Zaivd
UQJZn+XwTAh/WfswrG30SQxrMVyM7PNJV+R1mb+rW7kxp0PluUkhQDfT3zC/ZUn1R3r8wg+1uX5K
Pz5xu8ixskaSW6v5pjD673bho5T9+VHkzlQkBW7Atzc+/jys+vijjdiAXlg9iTeK33hD0ZDqUmhq
8JLfSBejDc+HN//Hn+CH6/dxVrdgUpB+oo38i9OkfTwPZPJ+zDxlLFy0/MJ4TgX1hACV0Kn1uaNQ
kU8AhgPG1D5bui4BXC8bZH1c+xgztS49DdRJirCIQSEwHyYSZ4Ftq5+FROEH15IME7q+IKgVpiAz
xO0oL23jRFp8MxRArYM5BQ+pucCa4iqOAA77QufFJcvPhzSArQH1GRPkXn9t/Z+Ncxk8YVX/oGCm
J2u2uwvNNmhaF9ltBidzfhkbi/G2/u2WzEmJer7YskQhf+7muWzJfAdV8k822Fcahr2v/oiFtv3T
LI4J71zTzvXlht6FVmprDphFPFaF+ZIFXfV9fV+zCL/0RQed9rKP6KzDqH5D0g3fLRszFjzVU+V4
7xapVT6IMBYrlVyBqnmKQraPRQ6SDmujNYq5+7mBs//tVPW6lSuXUrWLLEDCKzQfIpwUkeqUOTMj
1JrzFPauj+vZ1FCaDboEC/kamu8pIGGhjNN0vZ7gTZl1aYZ2KuLcUZwMs9ifvYNG+vwEEJAf1m7n
SMKj4W7smEPV9iP0/gNVB8j3AGtOzm5m6q9iAftRa6dkxUab5d2/V0CKkozzzRZ13ktMg2p12/bW
do7Y0SGNFwyHLI4Qy26nNhBO+5zFk/rW4zes9y++Y132biCWoP2S3oSjHO8UXBgS/YknMJ4xZocJ
iVb6SMocE3Ai1bvwE5Y4vc9KDpIrwD1JQ+j8TX+Shjs25vvVdBz0CKF686pVNdVNO8UpLTMOct/X
2dHHjRIxFX9GUPGDHv9tELpT+A7/8R6mNbxrzMO2+8TIVQBIokfffKrQuo5CVWVxfTkqxn52PHwo
vyLpOaohhDK4pPRB/lV9VvIjlj/aHFqp1v47SjvmN5TYtOcb8ILsTmPwEhlY9/nsdELMxEYn44k3
77Tjpw3pm+IpT3OlHsWcFTGTK3OILaAKo0Zgl7nOPodI2AvVa2r4Z0FKiE3HjPrNTE4l62c5T4M4
sMY0AB7kGkyLJwBNC80AjiTRC9Pbzex7wnJmzjqMBgIuG50wNtnpZXYzhPFRxllI2xx3PgMwLRDS
jHRu2ALdj72Y57dtWlF4g1owAyzwa0+1xoomolegk5jHp2FKdlWi23q3SfCJoCaMxuvUKYb2TclU
CmwdDe+3TCaqLGL6BcgXQWVvZGEN4t2QROtxq9bRXusmQryoiRuDG3rwk6wYWGXI4eJ78SL9d2Y8
ps1UbtNUTB1UnLSBHYBfpOrhJXjHXuL1zxJupU4A8MveSc98ukrqifhXEEWvRCKzUWiSYCB2pTtE
uJQSY0TfnB/n0CCoE15gPZewkN+mOi6/QQJpfuqNsaXnMhUS/g7e4+/iNt4bpiBlRYYXDYkMZv1b
OiXorCqxlnL/51Y1yvZxjzsJrCyzcEf12eMPA7jEW25yCKyG1DecVAA6vIm1rn8aDHRk12tj9LIN
ehi09PeZbZobQGOfs/84GWHLvVKmg+f0hmPQ5oTcahRjCPZcQIMP0BpO1dMWNkooVwQ4G93bLmDj
6Ware7hres6YKZd4raUUgsrSZsSR0C9peDvSP0kEmWQw2Yh1RI/4QkFVZLmqtvU6pAhWYqfcrcAL
OHRI7BLrCopgBHOjeU+kkBREsTy5WNIWVLlPzi/ovx4s7pRyCXQIS4qiKWh6NlOGiTa7p0uMvDrL
t6zOn+hP0GT7oT5hcta+ez8ejTKX6k0iQcw+Z/9SLLVihAlt1GQT6fVCtqamiioVtfSXHU5hqqlM
1GI3hbuO51e2mDdJI0X0vKCTOWXLMwPw9MdSaR9Pmpv7R12r7nc11hlvGVtJ9tRA1X3lWTbvK1GQ
whRwk+mFH9dRCwtwimnn6WKBWwcVXkSW+HBrH72bXKhqgk60BFWvzIPIigi3wwXVfFIVhoVQHQbJ
bQNLKhZExAE1ZNbLdcSraJB9ucx/lfxj0U6c9dgfiwyM+IkVDDqI4nHxsTk2KVJ+LKC7QDDdLz3K
1knTdTeeG36gx+NdTm8Ut6CqQTXf2n00rM2Lcyytk66KTVrkh7o6j5zqRk/kXD/P+3FNoAsBJbi2
ssfzBLWXR+XeOvtCK9lD60XMMZQVRCXJk448HATdVCYLglD+X/RdBQ5tL2qeKACe2u5OLKqKvemG
v7tWdQsVeJUHN+GKkcbjXWFMRLnOjHY7E9n+d0xT+vUxriPb1z8nazHsb4muk8VybWuPREYT0KKM
trE0NO31J/TORVXefB8UMcu7aK+sr2YshwGEaXAWLDEF8XOvec/xub8podWL+BAHxp/lePIri5Cb
paYHccZe94mgr2EfmKf5BtZmB3499Vb7CXyvmlMuTRAxSF8Dqh327dDBWcZD/gw3GqjZIzWCnGHX
I2cy7zgiTxpTezGYUE99/oLSg7Nt43wdlvW9E+R8get6c15aMx64UuVLuM/R3i/TzYeIXXF+J4Zq
6jLX/b6nvZ49CPMhjgjmqyW2TZ7seSxOfEsH8O864YuUM35soGweL0L7dgy6f3X6C+hkX8POKnq1
cg3NLE+AtIOqOVIRS3jvc3GOiRD5df5s4ckVJtyz1ZIYuKThOe/8fogk9RlU5pPwoAWgSbnM2Eoc
Y1Z9m/lV/adxjzG75mj316tvLQxOGcRiUFw7oj5aAJ9AqQUcsrVz6m2HDrqz+a6oMS0i5hyxhqQI
fXHZJ/atp90uLMmmUmVyG+StsIchW1frRNFqbfQXlacmzy/6DP/pPWMDX+2w2kNpTctHac5gWXQN
Y6D6M1NP5DfuJuu0mNLZs3bVg79T4lcasQi6O8ff4aZlwI+YyaBClHlCLinFF/QHD4ZE+NzF2Gi8
ZpSeymU+sygPyjqWrGJ2pPgpk5jg/NbO9Xz4Mx8hDWE6K+0fi9mzUHiEcjuIztUxqYksNMOk0wXC
Gw+AsrOUID7XAegz0Fj5bkPtH6xe3k82KBqD7lYRsjrF06sf/V3PRh8hlm+XmWcZOYEzNtu/OAJu
zgHdHqtbQbsYwgRTndFUipKCfnNCgGmZFbuxZqtCe9QGiVHwzHcXEMwPRc+JYQmwn3Gj7wQVflxh
TJpAy4hJB4Df6Vh0WezMYeYlFhThCyFiqblW11cywzUWRzL5R8lDL4KhfFTJBOGFXdpknpOfW4H8
NSSsw+MdvoQ04A1OVDmvlKR17i92B/B6Q67liQ4VrWs9MsfbUViu7q79ulLPtRJIWO2x9+rQePwB
9gJPRMrFBaV6qVv9KUbN8lmN+rEMBjpQ9AsK+f1IdFg2QBXuoZMk310rvwghOcOoDlotcXoqiimU
tUknIt9D1oFcN+MtQOuC5eTcAIIQBpFZQvZuRmY/gc/EPXSzxqYNWYWU3jgxQLVKSfwmRs9zIFL7
j4acc1+ZOoHwYJIYSN6LmNjGa54zUjQ+tdwxHGJFbCJrw4puOTayV7aN+f2BHfCTTR5s24wkm8qC
8m1Lfl2f56KnSypEUJue1yoROAG0j+wme14L8jYx2ajh7tP/3RXkFl3kO2fYfxLgC25DpAnZLpFo
k3bXcSXsZdWdGhsrUEJi3dXQ3f8ow6iUjke3ubQ6dXgyXmSCZPFDm+rbFVKJ/sOB40z4Pfi/acSX
wg3efYSLyXsYaBs8hgKMZpr+YMzpBq11mKKaKEp5QXrwFxms2LfCnPBt/dTNqazfwBaG9xqCx5cp
6n4OfPiC1VZyu6loae3hlExUdzBhuT/m8V0nDWvewQC1YC2BNqX3eHdV71zvhE8dL33teQoLpX5X
tHLcqKgDFBjc/OgFCeh5TC71f0wzhOZOw/pF4wN4vGEM3KP2VXBwSRiP9vwDGTop63h3fh/x9JbX
s/ou3yLrdlJOmfsiiT4T4VCZA4NKhFFdCktHTQ5S/xEEm+l5XxrjaAraEC04qPrbrm07DxglHLW2
T30ty7df4Zf0qwr+rlWRVz+Miz5K2l2Ud2DAEY1qXCNYTNEjDubRnSu4MkpVe3rickRJv6ADQfKS
eObIZ5JWKP28gxzSIu8ub1UYqScfToT+p0buFO/91JiS9/CFiUsfkVTU2o3cpszu2QEePE5UDb5V
8Ai7LxvTiCXlblmwJ0aYsd3BbpqX9po5Mww+Hi1aFyASmP4QiPC/KUyIfTh694Q9HVt0F6BQAFGZ
OMEjSkp+TgmOxjmuec1GVn6kUErxhHCMb9y07SadHc+YXoplSN0slr0+1c/elvrjeXqGHOCpkEm+
Mtznwl8+vtO/zYj1KUSuU+3gS8/r0VPktcn+iVrPW4aMVOZpZz6flta+BDvjnaTnshuhoR7bPSeJ
kKf4pdGRM+2spBScUAB83dzl6tHQarwbrcqOeauR7TLz1pXh1KuHZv97KJCsCULAT3spZrTK41pW
Pna2160mAcwjjJkRZ5pBbqfaiMLfdVp3NO+e/psz6f4t6W03vnGJnD5Njr45snipzCjmhk0FndZy
lk1PW3xI82iTATgDLK4dRJxXP73nO2I5oV5CgTAt+kKO8jev8TN+bwgvd+LXNeS+nfI19MJYYf8q
6gUrWyVApENtI9yWca78rWp53KbtQE74u1W7ZWJ49+t7NQtUsVFvMn+aiVLcp88FJeLryG4fqsmZ
mhWkj+GtKECAmzzXZtk1NhXTX0vF4PQZewMJBvnb7ciJdWVvJA9VCESwRZ+vX5dlC51VA1LV0SRl
Tn9Ld2Nz4aIUtb0BiXlaAROzov33dixnJ8XGAPRoS3oyrFyz30GROrMDC64S/f6uRXQsfqKJY+/n
0x4N5+ysqHzoJ8lcR1plaEQMKlk+Ue5AfpOKYVjl53xj2mYsDZboF5rClK1TfhbGBih88ZaoqVFJ
UbKwIn+cJ6sdINn/0WLJBlU2ecJmJ00W9UMAeX7q2X9WVDngZnYVzGRIxI7kzZCBEt+hghxHzd/s
oc4zCBu2IwkY9EcWAcSIDNPRANrQlJCP+xciiE9IMpLcRzLY5WiwzotUJ44D4EN7PZxdxlRNF2U6
dI5dQ2PItcx1Zn70FfPDv/h8MFhuwwv9txwrRFzbx2IFCRuBMvsmuGAMj7zleBnjHlQIf/qxOo7E
MHnhnwiwqHU1+wba+Il8naVFNCVbWyWpX2tq5me/ufspsAzmNWDyVA8HNlIcERPxOX/K3NSImjkr
OYNrY9+G7JttvP2l0ypw64LdXNcO+mxwRUTn6ULwzoc1RCKpLGzQ6/Me2ukYJiwDvROh5/hd6Uma
VYavr+X0FQv8HKAmLI7WjsO+brJGN0Ca3/4lLXjba9EEU3dsJsOyRpPCoxRN6ESZsdXk9mqUKFTl
rVyZ2u3VQ2tYGsu0g6GLs2OjV+2KJMHU2xghKGuo0CUlFH9se4MfzKk4imp8TlLuqtEDgjnWthP9
ErIeM7XCptmqsjXxNDBrA7Ovv4uD0XhEW4iWR19rnWa/cVlEVyo80zqJfXNU05tF1qez0hnuB+Rk
eFYEP6zGMxe7ahNPJMwghJWdjnUoy996PM+GZQTcp0nqX9balEoZAk20XY79Jlq6vJxiaLYoO/ko
b/SYbWQC60JHbdLzAc5FwJsSGMBFpJnLei/Kh6IUCIkoJM0qb1Jqpt38CjW+d3YkTO0QbRrm0lVI
uLhHmV499/JjA/dSuWu6eTnqxf0dlI8sEPThZm729WySpQw2V0lDkDJpZ2ahuSDSRIxQBDo1ONtT
Kt1p9T0gjeuN+uleaII+CIsZGViIwvyx8ytwpOgOTyLfOJbgE079GlB0rKT5vmKoiTHkfmMoEwa2
fbUqv6qIl3ZdUFuYDgpiyLZu7UZtLmFXOWT78YjHc38yNoBWjeKAmTIDFTubs4n6r5A+EdzQU5gx
Kwdxsw10rLOZDNyVr+HH71tSEKJXYtERoxcycaEPFoM4Mpl0sI3z57lYuru2pre1RQBk1NVhWOCH
RcqWHdGSimNj7Jo/jOq3xo2+ozwtj80G47/8HB0TL7QcRfI5wEj+jRsGxIpNe0BKv5bOF1wv295a
bXg6hgVcS9tSIbTzkb/PGdrKmrvItogXCd7UqfHTCA4am1ckqQshnNmwZqXV728kDSXxHzv0vR6y
d5nVOJfdZBqaFlMraLmO6SeGtk2lYHJ4DinsvHvmVDYRlNAOwWDhp4Vcqk0LkaaCcfvBSlpv/8Fv
HjEqX9s/S3jiu8kYcb0hfFWYmRr3a2d5M3wmOLpu2+IfP50Pp7vQ5uC3Oxo7rxRStX0IvvVOMU2f
AnzrYVccPdOoepJ5UTAk+23Bq5zlhyiMnwkpcv0uMkkJqt5KgcrECJ4co8f8FL3W2F6EELUjsKVf
7hd0QZA5fJWANKbYFgUJJquCV0sexQQIx8WJjPYTL3hQq79Ganz6KwG4RlukJOb5esFsZu+ERsDP
1CU2EkeSZHpDLfGA1aJTWF4P5piNiZ9IheKeyvik4eEn/AXC1FtkirgIQ4cyi7bwrR3ly/e4D16Y
d4DeJvlcVKRQ+CuNdhVFn8Gpc3jzS8kRcvV5+4/vR1EPWahf/oWqXtUHghRndNBdFFjhflAgh7G6
PhmGjNh4eaYR7ohDjGahLF7SANOZCHax7I/ItllBSIWnQwWCMMUzJ69OtKIL2e7b79jGL+fBbvsa
Z72tapIkoHAMbn0igv5OX7UNNThmpb8MLdKcP9GAYyUtpExCNJEJZWxl9hxhFkmRz/Ysy6Rc5eGO
rW9uwbdHlxG2283GN/cW6l84vNCoxOtcKMqmP+FTAjIcdxZEpKNg//EbT0lExJwmdjHjTLlqWVVq
eYvVxMBtnyaSFIm8l3ZX3CPq1KyLW7Vc/ovZBeJ3PpWzXQNcOmJzVFpeS6eSMehPvElL9LGVRur9
ZFwyLNysIVI769m4tItoKNx/ddphtzsFyqYdSRDIylKubGJNsf7BrQw+RANbndosdrZ6Wkn7mebP
nvYNgbNTXJQ5pfOtU177PX1CPpWhnhdttp8luFqlG08bp3b94HtGEiXFAKZM4Tfdgjw4pCNXPnkF
Hx2Pf4Cxi5aXceBrGouChorDbfswj+jBe3mN3ChDnqOGQfhDeUjhbrcyGZkaZJqMnzAIdc8UoMCS
qmV4tni49LT51LIGBSQeRGZZ0caZjWdXRZr4LYyDy7lkugoOBPlQ0lqvwnCWo4UwGWvhiFiNl6Tz
WX2yRC25TdmYzeuQacOgs2+/GUFNnYNFM6ce1jlXxodtDukZ/QSK6/cN7TeznsgYy/uVoUPry8e7
Lm4xEKOuULMJ+9KCoMwj2ADSjXT+SJubG6beG0JIQA4x9iMSoUL/6pGl9E1LRnQIV2ClcJQEobzm
MdrFGTvVufg4/TCJDAmFgN3VxdzhszyqRj4UYXVrp9FtHJVNVnI9KUu+L8GPh+tmnApwv3KUgETI
APW72cAWj4TeQ50dpHInr0QTCRmAIyDGSDDbZFux7OSqKGt8m4IYVjQvpRBdRnij0O9404cdbmy1
vNwz3rVuVJ1b3QIBLp69Q0FuQ63uUPd047zLnbkhy1NHFtd5DMa0VBX9IIo6ZTyfNp6NR52CVGsW
y2F2z7AfAcubimjoqLmapHOVgr5jaWg10MUvY2mgiIlVrFiy1xOQIziRea59B62hKvff9DaekR63
rI1OxrZBTjGzAlX7UB7RPlrbIth55+wNnQuI0dWRvEblKGshnoqFhft1ttqD+NKBl+lIcg/gOAnV
OWTOTzNO7LFTTmNZPmOw0NAMFHGXDoHNfFhgW9pOciHcnzVRoSkIQB8ghIvHFNn2mVmDEIQYOnlF
rp1WEbzB8cuVLlbaSr1z45O3kj2UUyGAzLvpaVc4m80pwHFBVqtMQWlAdEEbNUWLAaUjchE1Fv9Z
+v/Ky3OrIHRx4/BDp8gNDec10ERxBpCE8pIyd4FzBQYb20ddFAOaqOwEazGIkHUF733YSmTE83Oz
rn4BOEmyOmLlyp1qUtjJI226T5n5TqRtouxREtXdBeWZYODof7+6N9TY7nS3Gzlv76uW/tgkC6x8
9Ukpwj+wuVynpno8gvVHxhNoGD26uT9/RynHAxV8HbX9TOGi4xk7luOCg5LnAFEhzvoX2bg/q1SR
yX/5MXtrcSClYc4LvO986N3fVqiZLmc3YmurEROFx+6fzZjLjt6Ee3PCx8K79LmAGlnmg64a2cm/
Za+HB2lJwRjq3NfgIMweKixVPhzfs4EN31jNRLKsBW19i/snsMcrsVwQDzBRjk26pvqPaUL1RNag
JthbDH8RWIJU1VjErajm2821PiwgWIiP8VTzouiczuCjopyhaDJRcz38Bogr/yMQ0YO8qbcxU0bk
lHuiOifVTZhGxjvgAKVLHtFkTSApJX8ZA7qJravXRj9rQw1O31YhiYtPcBOjMkX//EO/Ac15W196
jN3PFrDFbGOaW28W58KjULQ4XYBbaYPLg4nP/M35i3TBvcu5tWsgjMeWjsR3yYSQkiOL2lv6Yy7j
Syq42d+uxWG57HOzoO4IKgCSk+CigC7kCrTHZnGsUHziJClOdzIis9owdInkDvLdw+jaeVAMV9n5
ADdCr4VD9/M9yZdHuBBbvP0FPWd7nBXTUznPSYtxkHTTznwX+KYCK44qWgOCViIIyUGqJpvNxAZ5
P3N0kXNg0QguEpb1hDLJKqOJkAQ9jZWN5TUdpBcV9dicmLntc+GkduuSfmRM+2r5e1yynxSkIjsm
orGvrK+dVhBUdX6K7knDwt0IUih+gHMQ1d9X/BMX3eNd1dl9RilQXtjTdc6K+gEexskPKNKHuPoq
O9ddcjiHvmFJS3uVtzLEtK4xNuOmmPtiD/dNYtDuziQz2+piI4CM1xcMad48QWnmG/gbmLWvdd/C
t5fSmOu9lN1n8zmgW+/5NeWUiKOLKKOHsCKPH1tV+rOFR2ceNCtBXUBB+Q5uVt4bI64I2CZ596cM
duRXFh80HjLdAoco0iDQJ9Hnp7xb6TUwJbWplTjp3/wT7SGrdrll5qZT3JbIMaoQ3aDdon+i8PhL
xxip2M+VY8j9as4b9COQDTa1IvOSJL/9fy+UrItfIy1bPvneU+EqavJ8LksEcdQl+cdWVQR9fxnf
s86fnlg3oc9vPehChTM3tsiAreLemK2J0wnvLiqBpOZFAfHypMhX54GQVgBxHt4Z5HkoDomqdjlf
/O+5w50Z35auvRiugI89/iUYUUXW7y4l14Ubu3aW/4xHHvGs8th1vKlNDPglX1Mf4fr2awP01smF
n0Wj44PIp2kdP3+o0kz+2/VUVn5pyqkPpK2qvN76yj1jyxBMiU/O9Fy1Y3ANT4tBAtkRHagGDcXt
+Tsk4VaRZxiMRJt4SS+IgcC0o5Mak6bLBgZluES7kmYSCAROPL9NhSn8o44M4N/YmLfi6ojou/5D
CIDSZrJWaK1iDTvksm0mgYWYY2rjV19zUmFItkef1bUPO5EDFbElIxxkZdmY43glxHNIw5mTVGWZ
BSSmblzlV6v//I/c7o/dhJ/TjLFEhYSALfrf0Vf+cff+PFd+IkWDnS+qpZ9riIA7jEVhoKCh2ZWf
vSYNv93AuBxzVFhqYV5fVV2Z9yt6INks7GKzI9UYyorf8e4/N5kVA51Jw25YzoftPKsga1Wb+xzq
H8Loz8UElvddGstPDqn8Rja6eVUPzBaDGbMO51j0SsvcbTUCo/GeA4WTjnFEBAi0c324Qw4gawQf
a/oszCvqrNjkKAI/LyAhZvQlNEH2DhDe8Eb5m5VfygxuC8xXTzHqVi6VOkGuUK5EMGXg6tDnnJyp
gU7BsRbMj61JkYLkVUC13JzJ7Wy3Hq6mV34pBlK9jPxSipsMiWXJ3LJA2xKKvWyE6tG4PZJUKbS1
bvkzqfGpe4W21F/OesY1z5WGxuGsl3BvWzTbsggyam+XhCTIVgyow6U3qH2Uox/r3aooeJBYwWcj
0/m1HwO+73VGWe903tfqXks4244Bie+KT+ccR0PMsod0gModNBScg6l+a9HNADa/aSKjnY7TAwrB
K7QyQaBlZzP/FvVBfK3XHNxGeBGoddM2VXpMNrhyRtrQTkfg/7frnkxSwSWx5COh3bpiUTATvz2L
Em2XkcfmIATLQKI+Andkbt6Jr8VrIJR9NpZ6OIlREbI3v75UNbRiYmOCu51LVqUaf2NnquljzoEi
ydu7HFORi7G1OTE6SIyz3DU4XERcbjnP1iR7pWnV0+IbtZNoF0gqzWhq7CG4RHPTjNxRr3XbKxoJ
zOlk2UHW8N+Gu7GhXPwRzwe/uySi1MvRLLk0cFh4zWUe9GgtFYd8HBE8sygSY0K4jMUjZkb9M0z3
uQL2HRCl7z1aT8tEAcz4RmC4D0UWc+5NrT72hZJE7Y2VE+kl3J/Q9L1C1G6aih+R2sbP9HBhdEz1
Wg/5knk9YTJ2f1dSVbTIK6Kzsw7mvc2DxvofpAZ919ZBFrt3Aw3ydZOlEl/9RMFG3F2Hh/HuWFEI
HWa5IonE6KTrgYkxKCq5bB6C0POinGJ9g0qvCKuXnTIteYH68w1yhxA4tlKlF0dfcYPdFXvAiQv5
B8kWo6rNhmm4MtGsbPAEwJgix16PRPUdowoY7lOcxx43YPAvqdChjyadzmEa9cmqxUm497CfbhYY
fC4eGfivlANE1oMex0crKFylXPi1guwH7EvFgZCRVGFFUgdqRY06/7dd30UVJLpFEXVU2oR79BR9
bouxtxmuzHA0muSDFj9RSmzQrK+O1kBSgXd7Pp7S+nnwzBtrUCbsVMD7VV852Zkc7HisGm/h9aWx
EAaj4kK+lzaCMTk6WjK5WUOnAPkmStpY+vduXlfzKexpaoFPBaVwPJBDT0+b+PqnqxUabLh2AF4a
U2OOjS0vuVrZvK7jeJStPfqxknPtoc34FjFLXws3j9BWgsGPDBUoJb09UyhMXYevvBX+PLfdWGrI
3lwr8CatALTPORNpmSPLY0Xj+xgHTU+n5POhMGAaiE7ejLw7yWcIZDJDsMiyZLJPolsKyHtwLw57
BntaGTsRlLvTpi3iHtS2+m4lDrUygfkBS7OSZcyqRGotu4gP7miq1skgjlV7V0/cvKHibzkHdBBw
VCuRdGfWIHDSUAhhAUxcYtdfkyz/lxJMdDaVR2s7d2dQy68sHJzMg1q08jKABBPg3lGtm1Qcro7U
fEnhOEJrbTDiXbDG1gg+qM9SlDb21jnoA84ESkTP4UonDIOWA/ArcxR6j5LmJK9qCsmeoqLo3g/f
eY2YvJ428Y6EyiQrYlTgPu8Te3lz9Hu0I/nfhDAv5FA8sWZmhB1/0LyAhEbxXed1IPgPCOBWpTC7
LDP5l55M6MAxJIb5PgtCOL2kfKdqLp3X7MYU66TwsYMcIPX3Z6hiCVC+05PMwX/c1HL/LDm7I35k
Yj0IymYcEF1S/5eWIf3kSplN0ZSUBG6UvCIHmSmIM1EBJ4YGJXjuUy8HDFloPvL225wCaXTmFQtq
Jbpz6fw38U/l8uBoQAMtzRN1XJa+oyI6PdYxQmOpy+cq8lV5KD7EBzlNYfYghZCxFTNZHjpl9zz0
R0BE4nPbQca6dc7RevhbFMRg4h9rlcTQnrXxU9fvOkswRD0JD4YrnT5YcZuoqodfYsi6gCs5nOMb
Ho/GV6z6Jki8v2r/L16+uXYm60D/GKYig02Vm1CmuMuLlrCL4JrhwaE0YUbqgCgYlNGV72M7dWKf
Qi21Vjr+DigGRDK259hQKfOLOeqJl1D62Q9RQpe5SNvQch1fsAf/ppQs+jjJxDwWP5zXCK9qkk35
d2xNHQd56nVQ3YAa1ZabqoM7nWNEwt+5UzQeZR+U6MWBFO+IAEbHRDlOtS7UqYFyjtKkkNwVoLug
Nt4rhGgy9zeU85k0L95bSAvic7wZIsox737E4TxH+svknClbx2Ha4xxxLFRcRBLG/VJ+84p0xnIB
JSdQeBDW8tBkn4+iw09UvZXcBxWxyB7y4rCxizQjer/qgqOG5rhtpk2QTl+xGVB5fLGnnMwyrdob
uuLp0BCqo1JLOk3wZ1bQt9hXlsX6qOl4wpRJoeGKLCGlPbYuNbRcAV5yIQ4msGzjKy7PTv/xgsfZ
bBWD8sbPAjjy+U7Yr7HJVVbFz6oljF33X7TPjH3KCU8wipOZvE/GzQf9nP/baoOFuqTZ4LNVbDiX
qSVgKC2b1R/XnMZ95VjGnOwQH9HDOD9HsanKiljaSScf5FoJpMhHAJpU/XUJ9fEUercSBrqNJ78c
NkwprX0HImGSnCX6ax8CUGCDHhHiopePkIryU5vqI/Aj3eacEViTVb18e3vKpe6Me3rKs57ILvtw
mnvvuyje8O0wPblxtd1hPvZF4DWlbIg9rkZaAgR7IYq34fFallTj9tOoXfcini/Kb6sE3oyniXQg
1CR7FeAX9/KntdSgGUru4djJW7sm1QS7MKL2+20CsuydjAIgSG62Gw/gpEuyuHat0rR/TqyOKo8o
K+5b5y59HTJyvDPu1ztMoBWphFQ6SbRqgM+cGlH3IUWowORA1osYbO5J/7GZy/KiFvfuoJf1im2U
yJ3ThPqIyAuukBEkYOxiVPdj8MBVSMhqOlldohCmy9oPUEWYQmIrINwFMMKaEi7mYWxfH6rjqg3A
hvjE2bt01Wv6YJLIZs2C91O9uVBVYkjcgLgbjPwiduVx4Lm72YxthxqFO0HLVd/vyZIY4ycSxisO
2cU0VQnJEnTqhpoS6igBoTxftj0eY3XMkrsPxbzWtGbF/iTk05mxAEE+ert8MmBUZ+JoK9onB1u5
S1vB4fsFwzNG11OmCAxjw9Zq48iSJCmhwY5khBIjiX9IX7Wt6X3iYQgVHAqkvkRKa/hq7pmKAzQN
1qtQHwRn7wB2iQPs3vnHNTUILTsbrBmEOimIlvm2VC6PbpS+Opu8omik9kRQXmMwiXJrWulQFItk
KGk3gdsIEyDL2K0pEPc3MHhg2I8ElURmlYp3K4ulJcDhlvYjnRheS8LPH3m8/sATLiew2oq3jBgC
A7eKdvJMtEz2oQiG9vuNzrvm0ZgcsPz8MwGUDHAQeCiCxC0K7opA92OqJUq+uqxGkzkdNUHUi0BK
HuBPDoBUnUTgbRdAdc2O1TQFr7gikdgQs+oQ4BKksOPWgXjDbOMen6h8pzxwtTjPyDnMvhCyS/RR
L5Ce6rpXaHcUNqPvrScJYZw0YHuRtsPtZ69ISDAWHRasLT57pu8lubyB6V8/2GgDGTDO4da6OMoZ
RtQefy2vmqxnluVU4J6Kt4u5plLaqzBUBSCMHQkwuWGNhEGG1ArgzArmuCWFIFfolf/JNPpG92JW
R8x0rkiUZPvcPwrcD4DQYHHg5FZFL+7YCR/gi7G3jRp/5cRlOGnQmMGrSjosEBWY82KnYp5ZcAiM
iIvzU1iUpK/GFx6UU98v6ooKarWDe+TWh0U2A6HaadqPqOxPbAETAEnxG8czRDA3U3fr/jAXZmOh
Yerw0wIrJA5zAB5TE0ATpYv08R6SKIlXJO4fknP/4zemNO7QXXzNuNcWoij+JYHwsUY6/0GK1BI3
ii1bDk07mX6VJlG2FunCOHjQuiRdYjud25oNAIuXgh0nBtPkhnVkry6eOvKf2Du2kKBz4B5KXK7P
/9+NDW2MphTvTMvIShS27MrLVs3w8aXJ2HEyRqEGwStszNhS661cv5RC1FjNN1hIHUYfrtWblhop
PC/crbWzo5wS7wnQDip2tdgYj9tORmKGbGucYLE2wg3aD3HcaPl6uerh7pQEGVL9qAmoKDJqKNMd
R1gtJYeDkWtM3nKx4fhWQhtTJWqKsF3ocUVcpYvhbHIttiupNH20w0NeWjz3fycLZxRhZ0Lav/1X
GzkxJ6gutZUtbmJNUqO8/3Aets0JgaQaffIQ6ci2HJ/c1SJQ3fgmPyc2MrAKuzg+T8VC7c+JZtMB
B/5a0oW7J/AbTgy/zCxFCP94g5s2p9S/rzbr9ifBaImnRrTsa9mpnJI++EmW0EKrtZ+HwUYt7KOD
bygT35WNPbTgbmPev5S08fKb/IY/bQ4+YMVs6HL+paiKHATzChke42a32rqVqWEip4BuW5U5u5FJ
muXdRq0zEOt3/HR1ZRWIE0jvCWN5P34ojKrPCJZEqm/4HuHZLspUVugoeLCCtCLUGql9b7aqsj2N
Mwr1QpE3zN6AGpRC7yzkj5Od0Qn/sYXP9Agz6ZP3tjZJAK5DL121Ku1hVWzVMKTzNIFzocQ5gFzV
8lMp7jZw8pC3TfOMmA1foJJ0R1Ezt3XR+TpeoDAwGLoufb2+XNTMCz40kyj9ZR3QY3AzEqn7cHsL
aAuaIbLgzV0WKR+D1RqOaGLYNuq89Hop+w1tXXH5OyHBNXgyA6mMJIvnPDpmEM/FfjzkI2KxEicb
GGTKazKG7YCBmhvgZScqwUR0zjHR9BVhGpGEZI72Uvgj0EgJydharyF3Ky/sRG7UgCbgDYjYNIdd
ysK41FjnLRNa8z/uyrwnxEDZ+ovwwra0hREFMB5q6yKfwRXAnHqyP+KCwDkHnCMoAFwHJDSe+u7n
PPFfLovqUuBxDgN4nWay26+YuvYfO8K/PpNv3K5FXORBy1Pm1UkQvTADd8Y3oioDEsI1ToZHVx9J
89ryjaP21Z2TM/XFKZM8zXmf9c2xR5tb0nSDUttoPRBSOx+M7AwchlQbY0CHhYh55n4FrsGGDWP8
uhLYabd3l9+1vMtwbl1zHVxJn7akN7aA67dVvlvwEtbOOeTbMJlhn2HfYfcNQ1Tgoiegc/OpR9D3
rXaPB21vyiNYWogDzWgN6BxpZh/PJt8F7Q0VEfzSeOhtp6/2mP+EccMVCc+Rg0nuNAQV/HdR/Kkb
/PaakTY5uGm2ajF0WwyLDsiJrQDyEn+KA6Cwc/PggVw4mAC/SPDRn4LylpMr0Iy/ELC14fJQ6EZu
l8vuHTB1l6IwOw73YeMKwQz3QrNHmGm4vypmqyNlacaLaGvYt6VUNsey7EiruioapQxDclgC4n72
+Uti3xrk98GR0eY/SxDfDAhOYWwpZLjzeJQL8hLm+aZh9jM3Q4brGsEOdzQe6XC+/S9iXDo6nka7
K9E396BQHpfEnuvBq5ilmUmRa5mfC/hrvuj2qVvk1quMPFiCvbCgHyPL1Weh62HM4HLCTAg+/vTf
DussoNTrynHCwiTgJZTZF3Dv80Hq9lxDxtCOVggeKCP2cD/Ya+aWiYD3I+s1BU5EAKEbdCp0E4cz
GFZl8z2jUhzekQelsp2svcC44hlm3oJ1B1GIgdeJA3V383hVYE8wG/gJ1rQ+XpVyRboJPfMd6kLO
pPieUW8Yy3vJRmon8gDDN8TTMG3ltE8WuSusEKSYNeHrVXv2TL1SHhDC+p88KIVrVpsm+kdUfWkK
E96bBWw7Fm3kh0S38W1t59BQ8G/JplH25nSiBD6iQhjaGt6ZKIBQzdaCRjTS9xzmpCK5uZu/5UwO
fqEJB0daB79h7gBJvq5dSgItx949jNbYbB1E93S5jTvMIByAiPFGWSZAxQ6nbdUdSu0rRj3YF1Vx
x3d0nocPLmqFoPTIaT3m43tQPeHRdUjlqqn03Fw4GnbfDCI82mxe1p0yNRkvSiKclz8bbjpY7H82
8DviTIvuK8I4ahf7WvrNwAj9IKWgMlMTNYMzmtOOHZXPqybQpkq4WyWGAiSAzD//a1bdSIPfOYSh
g/HduP+JeXOedMUK3teAHDjJ81t9u5Z7l5Sb5jOk4i1i7HjNVjQhzfonCz3UiC/b3Wb7E930R2l6
8W0NXNNZJHKwO019Hrhuakv3sy3rMLTsiFstE/v3NcsE5OmzJoYsXbmo2elI7I1lKPo2YEE+qhhh
gz0eI9J6qPdKPjuPumDLgtoZ3xKegkB/dkpBTOWR8zQxRnB8MdXKChPAOLHjB6T17szIsVId0WiX
V7ppwlbnEiEdCbfz0uKqbtJ98sttgb8Lb49tlcPgCPbGDQS3JkgUfZf5HRcpdZ+qkdJ5PG0rsuN6
dfGIo4bVFTO0MLCvF1K/8pSSCHMB3zJRxM7ODg6HhEoNEGJUjcYSml1rmPi/qJp4o71RpD7uWd77
gPv7EvUKYt9saqM5xbsXmzTuTofj3YpsjtalfU7J9WZmKtRjPWXWcMYYVu3tMn80aNteDmANvaFp
dMbjpc3xybTF+HHAw4B4zHwseVBgJFyIkxy6PB35nOfulGMYJtYPzdbGbr1zJvybps+g8k2a/0Ul
6ZjE5PrcxU1KJycx1uIbz+5S+4X+hXHWzPptjrvLB3EqcAUehfRkz3AMfYecdnR/jzHuhHMOekJy
q0qj/gYHCM1HYI0wSCKWeWxuu5I5T6uCc5Cs3n7pZa2Nb+gv3ikPM34lUSxrPn+0LxTe4NEhPblX
0g0xV0zgjCbYIXxhzyIR4AYqisLWNLpEWu6vuoqn8bFOCxTQjTXVlL3/72ZElzTgufl185iDb0CB
Cnp0HMauh4hhsZKdYX74V6pysBzw91QhsdqBJZn9HBogWArmA7TkUJR1emzJ2PVWS4fO6/a0yhv2
PQL5tNWUeac8HZPrhisC+i68qEYShJSspsBUlBmh/8YZdUP8mMdqjLYMBmogu0Ykxqn1DWbCNULp
3ynpmf9Py441UbuuyRakxMZe1s4OtObYG9Id/ZEF03dSIWE6mMRz45+9cajvKm0RBRlsCxkloy2J
DvV9UeWT96xvuJGSBEdC6/faH/sgFp//1VjrMzeA5uP9qc6gQpprBUIh7rZMN+cY3++rKiho4rKO
cfQYisAeKCD1zzJdlyAtSi1M1jxRa1lDKsJpJZoCemfEAqo6vIPdfF6N0ahQ//cvKfxr7la6s8Oz
XsFHb7U2l5ohoaoYoWfpvhoCGdJWbXfRtad8K2KI+6fYoBWrfvz3fvkJ/Yyhk+ktnT2r102yLMbp
dsrC/S27w8JCLMwK7QMS5eAyAJ57CHPl5T2NeVQhCHOJk3yx0BuH0xTC+DPWf7EWcI9KRJMe5K4m
/FXljxA6S0lk1Yi6CZrHDU5HeeIkHBNiaWeCgXMLAoeXq8VW+/s3uEINl2quvRQ9GFlZhz/YRNXJ
jPwLX2CFAVvMeepq/nZt8Ypr1t0iCcJX3ZyRnIxzjvC/RCwOibjkILYOIB5XV/PhPUbxSzKGzuy/
Luvcgun+lxRoadWPHR9pOHclSixNb9a2h8+xXvOHBlAoJoQh1XNgL11uLMJUe1VWks/mOH4MnIld
Giv7TOp4gSBpWd4t0KRhmUrKmUD9+Ig5yryqO/N4SIOGvW3G7/rZWYL2BBe1Ix68AdYvY0x7lHCo
HxGE1M7FhT1/KIetRiZhbrRTYsiX0cJaKpkoSqAhzXY7u7Wc4SkiMEEoG5oemp9hF87iw3Acgd88
yZAianHjhZbRWfZ27tz36d1MDy8PNKzOJ1n4tEomZn5CsjhsfnDJ3ulocMRyIDccFVol8nLZCUEy
RZ5elq3W2YiN68j+hRrxkg4nb7i4sJh2m5bcTOlXJC08RhHx3zWnuLVuI8z66YjpDb33d6TtAyPy
riva3MkMusIaZxaoAxn3t1D0f51URFx/vDwyzt91HrE5ASkFayfa4brQFkPoeyNDUl0Lyi4MMDkF
QopNxxNqo69ecVVrs18RkEosontGva5Tq5SoFnx/DtIclDYIS5wDzqRFnDLuFk6+749DtuuoNkZm
MhJOcpppDLGXxQXpZvptftIKpQYrl3FpQ/WHaph3KNHJbgeUGN4r653mi2HdrK5Bpzoyi8d5Bb/c
JofEKe+vtn8cR+xRbSmBGx3EIn+ZBf54CHnEEJYgdUWh/62k/NTGf8Lf2z/yk51ZZsJ3ceKmh0R8
TO5J4eUqRrvDtCTYtT4eI89vM71EUsw1JKJZb3+I23M+k5d1add9ft+lEYEowkHPDTR7KfeDXnsl
a+3H2ecuNZedBCqdmnSHLIWgkUsmyQE8L1fBmRuEwBy3Y8s+ZA9Ep8XpSun6yhypiiub5MHbwaei
qMxwa9H6qXCcsEndvSWOz++HbEnPJg7pqMdGFUap6IbGu/ONLliM5vU2FNEj6U5HPCeQ14dJ7D2n
AfWA8WuqkyBNHWXoqaAUQ/S3DRs8x0/VKONKfVJj7JY7tFKgY6c9DaHE3mwMYtFPon/lbnAJ3N5m
xunDOKQi9zP20IEoGHJblVriHrPLpzgMiRB0g23A+o0THwAuk3EcqPFx6eB8kDLfKkVsZaTBZjkX
fq1PMRYIyvLjB6LtYFKKH7Bqjcb1Q7CNkoNGYgIm+Egz9U4NKkpIX+SMU09mpkOkRw7e6ABhmunE
ELEp3oIR/vzuggP3zs63JuPkijGnYuWSQLF5VxTJ37URd3WE0xxGAt5VGEpHrW7lhQuIaNV4IFCe
qabItuCiL+tbFAFC9qcau2Vl9M80qujhH3uOGJHv/62qok62CCsmMd5ySvckw0SEuagQ9NR6csMq
yyiZ7b8H/pjMBsOVO18a/cJxg4LHFAdq/EwWnPCWf3Zkqw/EvvQvLofr9BIVtMTs0/jmT+ce00R3
bXoSgKXx7/Wcg77vZ7ePutG+7c2Cu2TIUw8WKhHuAEgQ92fqsy/BVQt7rIBF3GtyjDeyUW6+FSyz
fgRc3bljHiI3bG1Q4sp5pCrsoUCiZG3H7ZyrVVECgFSFFfdSey5WDWtXfk4glrSEESJqjSaErGEs
yiwvL+6H7Nt8E3EYiYKr4a7yONdWlqUfFPWdzuUWZX6d19iH3N0pWwfWuPmaJQbeVrN+hThwOUqy
7nN4SRcycRKm7qZkZoo35tF7U2r5UGDqOuK22rwWWWV0mMI+7bM8MPWGa+NDgeAuN3v4LxKScSDU
Fc0d+nGuJoZseMLIP0J9zsmTO0amZCoFO2wdPgpOfGY2j8vS4fcJmqSlzMCnuqO0igUUKUZr/Zh3
ptEQzYDBx/Ea2uzg38yk7Kd6m8GGxVcGVL8EwvFEmd0/2oOhTd7apKlROALyHhY5UVcZyuur9B60
8jLEBTxqW+eISNntOZgPkKGiR+QP9k/pz0J037an2L45eMNcRhXhuQmMECFsTGCmwUc5WW4t2R2G
LDbH54ZoRAX8ybPSfMazzRVxnYO3DiBcWgDM4IL04TKo0W40J0gO7XjGLf7MfsfuUj31hCheKNvg
vL3gZe+615ByEMIr4XefqUVaot3ClSD0zPavaDoCefvJgC8EtjUbJ9S4JeDbvULlX/H7FGByDOX4
0xNCZ43fjoi8lcDf48SSCRhTWU2E2h/DqNf+Fe5bFZnVwrF+bvsnK2yTY0zeOHhoYM1q+gFmxmO5
RjCqfzyi1tCKcI/SwbJRkMANV/3qKUGy3vOx/TowpQl2WVerKIdVfiO8qVj9nrVm9H1AMPq9b44D
fbRPh2NAY2HJLHowkj5y5PYMr8UUuWMHdeQuvM6AP66Rfsi6WmOccBFSqc2/jna68RN/1oHzA0Ek
cB/JBf0oFYKjw8dtTpwaWOZ+uTenslGcqfvo0HJLMvCz9hMLbpmWnCk80clTLM74KOZSRGVSMH5q
RWfkZbMEPIR586HZ3goyLV3MiiVHNeXsEjUxM303x6HzeZnYWpEWvH8ir57TM248M5lZQAsh3GtH
amp8KzEAUXYIgqhUsEwHQB5S8QeWHfLZN1hrZiZ79q90sGez49BLLOmXZwcW5gsHefc8UURYyNo7
3aFbEB4cQgayKTClLCgIBqj1COwfLtsegvS0ehq4S5pRQlEWu3lKaztwF6ZsrWHeWeVtyk7A19jH
AsRMnkAAoSewisdNZ1PCCRQuWXAv1Lq1/kkmuY/PXQZLZ3et4qt1zU+0YMNqA6EhQb4x+wyr/exd
JvnDedLgWTbncL5lnCyGmlrz2K3itBFQMvK+TB4B9RdcGuk8adUuJGuecDCOkK46UV/T87bGPmBG
twJgI+nYaBf5jzTh2PRglRl5B5NoSNDJzHb3UecebTowiqzNRAb6shj/xiKMgO9sU8p5hf5802xJ
uaMnKcPCsRubP877QcH5//GIqm+3Y2vmsRWw9vN5Dn2/O3NVBJMbuHxXTaLJTXT9/dPnuMF2Pob4
gDihkTYnOhmut3S4ov/vf7QvFOrKyHaPGuAJIBoPjNOab/zfYby6DNltGr5D+qwCyL9/DG8wnTMD
Mf0fXFkqzLfJf/XJSXONg6wAhLXUxhm963glqnmK9+jeSdgzb1WBYXtyfl88/Ip39Rtm5v4IihuU
KNde+q0IeydWwmXVvtQTkUnsS5ouqnk1luDFSr0fsicBbwsQXQiM4zxgtOFG9667YLthu+/JPQrv
KteLf06AXSF3qqsAQkfSjeL50jJ68dYpk0zWO8c/rFXoQ3GZIhQiROwNd8MVqZ8S1/8CYMnfL888
qZnanQZ8K5wff5YFclRgXBrXUV2dk4weWuOAXGItJM8dY5aaLoq6ee37bqjVAW4bABE2CuHfinLf
Ppcx1kEHzCkOe73xBSMMN4zE1zR6mLIT5hAgkvxuLrjGaYDOzc7FJP2xRUDoC5PJ8H+IJbvBTNnR
hBvdlq9VtwsqcSsVyIiwFYxGJPnZRiG1bhbs8hiIaKUOxONM9429AFAkpCljR/KAc9ZISx+HV0DL
XdSzrKUsNaUFvsOeFcB5o9kUo8B8HYvh1anEAH10YLWBqsGQ4kgXEzv0RJA/dzrHn6RDcMacAuoc
HK248/Mk95vt4tBS+0D8w35RQn4CNW/57nDzM5kgCJCutH3KDgHqCAfjfHj+tbeWNc/ivIrPbbrE
DdpTwANK7PdrdXjsdxGG+brDvYD8+AszU3zlHOk8yDZw4oSGXoOoWkocU9BY2KSUxtpjPPn8UMjV
zMCA87AaB7n0mFzyQz4snj9ypDWGLwkQVBBYrTR8kALHTAoIurF3QY8fKtsdyZN9ATGAHr0c2vGE
WaU+EoJxZO5ex5GnD7kEVmFdKVbbPsp4MjPv5bxo5F94L81wpF4sGIwABbuGrPMkK1kf36K5DfN+
IZBxuwN9GdpGjvcxkxc6nAfwDJ9R5/q7do1wQXEHjhbqwml/8zx2fuh3a9sla1UEPhQUcYQ27MSA
bbNqMYlHTejmvPgGbcYn5R7sC0KcI6KXk1ggdOKQwKyWZKbjQGj7gz+li8vLm3hlas9sWMWkaBmF
9WIajelN4steJBLRCW0QyNVWQd5adHJB1zQE2X2C6HjMiezdsgA7VQJW/l3Jo/qaHY95ZhifsYBa
WT4vWTrpxJ1pI/4CChRZa9i9/CtL0U94mnRJAI93qbbZoXcG9cAclXgGxZj1WDpPEbjsGCzheydM
ZI+P5Mbz4fETEPbbZRLm+5SUYdB2JOiA1YjID7U/R1XoAfHUoBdT3+Duh0ltjWqt97xNm4WumupF
IsRn0bjW6aUsZGGT2N8Rwbzf+hZUFIyj/H0XU9F2ggNyWE1sOVrREZYK9kjB3Jk+hfGMpoEdDajV
LXZpAt9P9CcFKo75QfFZd7BKNDi/GPdHUh/pmm7Jz+OfB+lk7YgPwwlZwJ5yHMdjQCVkOGpuJR/q
a6icOuj//Jhzj6HYEBM470u82kTq5k9sGJ4e97+MFVIAr1Ezg9mjsn9jOf1dZTf7D5nAqEelpDev
DL4glIj0IlluTo1bdHt8s4AdabRFRXhhZ+Bg1e+h94qGA47BfT8PauAMnDBZTjoIIzFeidZgRdmc
DMHLq6lzuWP04pyp682rFjbmGfYl171WSOQfyDWzjgkm4TdpN+zoT22JVVMFpHfeYfaqB47T9YUe
+4Mk21EHsa8cI4LMnETMkEcZ3NoGctu99SaFGRTgsgt7IkKNMNuIhIwjLmLGpQpEjfs/qGcby7tG
CDrH8bnHoi+CCnX7utvpj8qKlaE/P4RnWRZn/scJQna/KuRubl2KA8t2sZK3V3LYT5ghZfJnX78q
uvetJAAJE/YLNVWqa9iWcAMontsHV7scCy/PVkE/bTlRkwSbrvvUA1blpV+EPr4dw4M6jICUZjXA
JrK0LztuzRm+k1GdPoHszWg9J3TerIuGjCIwf+585t+jl2dpQFNFhqhDfDKFUmKQKQQNGjQWaJIu
qr2qSFJhqXKLBNhqCvZcPaZTUWhh+sB58atOZxx/RDZcOsyznSq2mABLMfUBYeKzH7+WxpTYYpnk
093STKupDDhdcXDkj1kASCBC2bineKeptJJRtl7EaKK+3yJiTWsXHA5o5AqvN/YAf9L/VpdqJ3aR
xqALB3ezUsdzhFDtLGt7g2cLsp36BZxNKMwM6RRbNHnKMC9T7cTNLoRRsSI86CCDQNEUaSJuFKAW
OGZ9JNCyAdiJTUxy9Gd+EOHsfE1weOxPJQz6cm24zOHEknJ/63Pt6YtInv5Ie255Rjb4cwKyY9/6
0uR1e71P5A9bjUkZDZGiH8THzD4rcfV0ls+ygAkg87Z1K5TPGjS8m4rsOAkWfRcubmjkyVaffprd
PLCuvML07RPrj9u321v0hzWBjiJpLPxeYfcXTexMH4/7PsbDNdu8+ZHhvRLEZOf4J9MYYdzcy+oJ
3QCnTUa76qjj+6EIwigst7+jIbtal6rzxnkof5+4dJ0sou40V33rwo0ZfpFrSsJKp4X8HNakgxF4
/Aw8KEoj/0p5iRk5+JQs6NgaCEm5BneMu0BFECdmP3C9aeY0hvRDUk2wQSFotuRHpXZO8rM1Ev6p
1/g3eBj01BkXN4Oy0nV9v1vijseygUX0XGMrhhrFyPZnlr5WNzZfzsgDMoqd6qJKXGPlWCPz2Y0c
XDf/jZPycKWZKafT9FgqKmpd2oWvI3ahSm80rmS57rYoNWCADnahK5rjiYXi/MWkPwkcRua3y0Xu
kSdVSDW28yqCtJKzC71WNdQfEKNazpy/HTMiQJgnZpokytLHmEr6AUk33qJxjAkwU/cDejibs+3k
N69XvXsqqFEmC5bnOY/UDlFHjABsWKRLi9z+M92qtzW/aMHh9n7m7mt4Rn7ORnFfCdIGcAkw5Ife
vdTIH2jaDoPbvGM85PzDPvBW9yYKD0ztR8BF6a6Ds9rMRCeq3MkImP4x2Vby080ebaJpPi2k1YLv
L42SkjSXc7fgXfs4e/komZwvt/3Fmeal/hMFSBwxYJXvko3dnnklC6dMnEm8kEeJ3RJwNFDr/to+
TknCEE0ooZaMeFyVkszpcM4vrs9Af48MMzPpOV5WQh6VvRU1w7pLsRmeZ4nT2tJEwkBY2336InJJ
NNyDewpsOC3NJOOUMSLt0HM7QF7UkGAhyZVWh0+oRZVf/1MvB+E7PF298bmLSzveBY1jyBQhDItJ
eZY8WxdXa2aXTI1S8XSMzqsSbh6ligVLiombvd8NETGtSjTApKBHaqZaYjhgYbSqNGvu7IYVYrnB
s305x890JS02RaRJo9kS46pte++Q1Igl18B29/UdF58jH/7ikjCNdZX8C4LKk5MlASUNMqHeOVja
KcPbwxuU0/z0cSQ6VkLOzROg8dR67QzOEUt8Ju5mp7u+uYPPlveOcqM7q7FnQXSB+qTDzkwtRFhQ
Vh7mpNMZlCuKmwsXHwNUMoh/So3KEPwFQbaAU59CqAx0YvAsIVJbmATxjbhQALd+sKaf57SCIAwy
GrIkSr0j/8kACVbAs/vRAXsJibS62K2nlMH3BJ2PKF2a0zU/mOrkcIFQl9t0veDUzhgN9pHIHv1u
VuuZng8JjWMsrfjbHjPs66gu8QO8EF5mCJEGStU/d7PYCsOLPb4+ftotIQ9Rp0xfwRxTlyEuZPGj
YPoNOwZZr0T1TQSYSNTAxpr3uA/rkwHk84jcW85GCJGWZ0KontcUn6HtGvHre25YH6dylHAhfW/R
XDau3ZB7aYEQfcaF2Z3BUxJXoXXHeG83aGV7XeFgOBL6ywsp23YeHWx4DrZJF0Wu3NXhOkdpGw4F
h7rFfCpxpk7f430UgxIzgmdTygRD6+NNmYZVVex2FUvzocDQKWQVeYh333yYicSeg45E8AKvOHgy
srvEUXdULqJqGDpXgE5Ke+X3h4nZ9otZJsQTpy3yvdG8n3wxi/F3co8Y+K5S3r3TTN1XEyaKxLH9
swrFrEeLA8XypAqtxsxVorPc57/COpUehOaMtorDPpGaWReKBw+9OD4T0ilPNG3peqwHA1e847pK
HAqOzgEXVSvWU+SX5wEgTu+q/Pgg/RTixeLuc0C/laUGDBcgBLpuRv76nEuS/4JogXuqR4jb/dAZ
Qm0oBg5cbr4/6fdQFr4dVBzSIsXN45WWQ9qxIUahtB3Ery2o0yUFRs9wfGVYN+W+xG1QZvxTsVD7
Fx0gMoiXXgEhS9/UyhxDNXrir7LlQ3UlKuM3DzQKOewHrfS+/8u1noMSDCNzqQP8O0qJxl9D13wb
ETdqN47yfevhGgI8Jx88UBSu1hIgjqg50N5MDoqNqRxRxj0227ogTwU1aB9tWZ7j3ASx2GjGvGf1
YHWOCidE323t1C96kkys7hyha21pywIDwbYGiLC8WTAKF4FI9nEnbZPrubLFezZ4zvrOX3b2Noz8
eHqS5jFAZhCodA6BDh2e8aNVSFlyWKSJ3a98Sbl/wpTi7jIRNZgyeQldGQumSb4aCTEs/dyH/PYA
mR4RmkQRr52ruYSPVxjGvTHz4VI9v3KQsqIsfAO43usgGo8Nl8Tr0Nh3las5OrirSQVY5AL2o4S4
Am5mUU6agQXLuSfJPEXOSoC6Awsjp+mE4Gx0DShKLhLyf/xsnqnqtDan9W/bcMxazRX3hDUCbPLN
dKuc9Dkq36r6q4uuL+qQYhZ9FcC3OmSjjaKuNNf9HFxuesWE6wvd3+NyPCZQU8hcNijjalf/uv8t
+cI1iAKoOKgX9eF7yM9JVqM48TM6YO8qakIBF1HLyxJXBVwGxEVS+reBu1mmpY9jaF80iW+bYOYp
D2mgwYtH4n64goECLXlmBfZCSLUlU+68SWCWGybH2V/h5EUFsiY3A66EDJAlITCwtikEttczsH9H
dbNFQYcPeYMRC0NeumtgiCsLr+ffPw+BtgvUiXtx9Sz0koX6E/TMAxfwUF5RY6oQfl/JOrEv3XPm
u0tKrLlOQLmagpYEVUfSr41cuu2foflMtQv7EAvPHX9qZUITEc2kav9UhdjFbqt1kPZ3PIAP144Y
UvTy2cejdvxeSWtxR0YEZqQahEv4RvF0di72NDlVsbEFsSekKOXb153SxSgTlTTY5nP3VEfWMNGC
xvgsOIobs5iakT0T7w1d8+yAgvBNNCs5erfrSa5k4JzhNrtzteOM2A3um5G16vUU7tUavltqawr4
veHAlUMoJiB5cIbFvzLEYWmLVDhbg4n5+MjXnAm8aR8WvfAmsMlvJKKN9ZFLIQ3Y3GO2RtZ4Q6be
AIrJnvnDf2fN9EXfYCPkv1lcd+L5QbQccWeyHIX0wJV78S8uE0zswPNG2wAqi7CX+dGoshZfd2vF
J7SwlCIs5dKh2p1y3FMgdlL3JNjXzgsOgrfUkofIVD6JhLV04Sh8kmHqPR1vI5EPb8OXc9amWZZY
LKNyfTtooSifOV9j+X+LpxWdKAlXE+7PhVvt6y82mrpFud7/Rh6Ec+BkgT2uDuRpYs3uEcse2cIs
GTZca39IIkgbxTTqm73pHDDNmpozuqUCjpzggBGilU5mgF38Xr46xMZ/mM8jgOyTONeK8PsMTruN
QIlWBGuoJSxRkGEMimnlTk/EES2Qe1Fsp3OOQjgh3GGVJ7WuKaElGOu08kW3vrcI0gBqnqSJIUVk
imwrK67jnYmzdILN2FksJc3eLOn9rOqposOHlxlOLUwn1Wo7yNMhRUkm0Jjif64liRy/AM/tk/38
T7p92O1tbsBCiNGl2vdiTmuY+5NNEhOTsSqVqW4lLu+L+mJgHFdEmSn9C+oLGQFHsSomhuPjYtGx
n2/n34OIOnT5t0+V/rIIfqwbISQO/Kefm34LsbhfNhpvq1O1N3Vv/DDiESdJMvPtxh74JD9GlJFf
93rIIRJ34e3hVwo3qBGY/It8PS4g8KD68/NFZViJJ97lZjXNSF93JpS6eArFPUDq7X0LgPy0baTT
ny1VnS6Vs4V8VahBOxiINf71ZHyb908u6Bu1RZfQZZqdAW+P1kjEh7tRoRyrzikUnB0AQJcs1zrJ
31O2kCdJLiKAxg9qH8140Hk+Gd4d1/QiisZELi6+QyFCLwd+M10CVpY51+81sweav2KawJzuXIXd
sVp8xXOHdFA+7q8gFdVux+ZgbyqAd4WympaC0aFe3Unq+MSmH5+mjY1OMajwJjQhWKe+hqcgc2Lw
yy8BElTDrDHGaAiCWS1GGHa4QHGxl+OaKY1CuCHB4PpA6k4veNScKucqNmvHwu9lbt9cv60uZVgh
jWpc0NGxK+OcifNeaI541XwePYuTyGxU3F4zOFCObHBXQQTIswff4RoY8aAg+qs5RA2tuO+ne0jy
5rzd0Z/E+foK4IX4zYFCTP0GAcviK3tkI1SxRDSUWJu0MNHcnYbDbXAsztGCe0gYoIH36eTx9rkc
dg+65xyfki7KzKJqA5k6STzNu4I+3WHeUbAaLUm4AQdVvnKaGW3h/1mBhvJ8+bRXKLIAoqgqmAuA
mjFSdH4/RnmLPlD263PLktKZXx40la8Qh9YFSsIuxBcUtE9aIjJnOpIv1TOaXFhE/Mjgy2uqL3If
6Z8ZAfABuAYWfQUM9Egg4FKnNm2PdehEJhRKJwZCoEu34GPeuvLDqtbUiiDepvDlKkQYg1Y1lqyw
vQnAzsgM/J+p1anrpJbfTIDJYktSOuiV/gAdtj8QWW7mAxR++CTuY8zwbF8mYEJcOUqEI2fcwiKh
MYcjDwafdN8ZvKZqWJ1SDhtpAzLnRIPr3K4udhv+ioqSrZgLklGPwMx++AB/VGSJb2SkE7EThkDG
KfCMUo0PIOcRb5CgFMRrofGz+tcoMO0ocG9xt3zeJbVRsAsc22KRGA17eq/1PrCWmYCoDvyvaFgj
7booPrGwmKfPOLVIQp/0RdV1Xin0YBgllTNHpUKCRgOTh0BRbS3fF2ctwNjxqvxPcJeEdfxbpF7p
DzkSDee2KPK73xP+g0bg4Q/c+JsPhJgWnY+5mkvsqJ0WLGlHjjhjWi4RAygMm/Q3mCWXfMyLBVNe
L5PWsRTKaV5Y2/ih3Zk4XxXZyoFuQ1m8mwTglU5RbvwZrR/DXfiEHT6z8p6kxaKv4PMrE608ofBn
WQyocfqiUAq+0l3SNzhGkLZlDI5InXSwyIgxFDQmyO8cKLazlar1r2k39HF2HDlt+kDqXu2W0+Dw
pndbMsGmOtPVyZtJfS9TaH+U9kLIpnUgaEPY/IhBI5FdgcISbQSBgqQku402g/WoutYOURtuQyuA
h9OyU5AGYOpFl4Mqt/eDdo2GKwygi8CWcpJt4+iJJbWptSVTIwX6SxeMSYoXNWhxupUtz1r9OdO3
nKadhHsk9GkaRNBn6vRjidtXIeUYPkbLqRr43eh6b7lrXo9P1gd8G7QsH5zYKzYnkTlueQOq8tOB
K6kRcwGirFI64NE6j6hseA1NkBPcfvmVTUUjoygdvwz31niQ2kkOUH86n9hvvBoA6SRXrmRmi7xH
HJAPLqQ1W5UHkchJ72JD1Ke0gZbjM6R5/CaM8k4CrJ3SjT56JqAZeIffYCJiefATlA3biVS5ay/c
Tn9grLHCqiexudx0mDRxpjlK0+67ASJFUtSoVs1uQufzOLxz9bMo+kAy16DRacG50L0b/pVX7Lob
zRBQmw56qh7yf8U0YGTzeuFiCYXI4ozqiHNBNue+7DzSzk5lPAObyIzFkUr+x4t8j+SRVmcavPsN
GfeGTioBrZaIcgvXVjDAc5QaR7jIHRRo175CFNYa05M6jPi2iGHbdoRBsYwDJVthzJ0HGjgxWEtg
53jmu2kGGJCNEw/hvcKR5ot/Qxtvq1I0ZCBeyddPwIlKMgoaB7H0gffvlDIJuhRbgIH7LFARXV0x
iuPzx6olcB22epj0Xj26zO15nZu4QZfJUERQu4i8RJmTwLCexeaB/qm6qecCmfYI5qGtzoPMKHss
K/nlNlRWRz2/XBTQIh+n/EPZpmr7wQ9wj8zIV1pGWnvtR9AJ5ElAq8Styxw/9R+5fXnfu0P/pqqF
avdz2WF211TZ9UPj23OXzHKjzs6HiIe0Q46F8ZD/TGZFrNQiZoAWByg6RLuYDH3o3FFXsvvCkn9I
SY/1TJLwwB2cBHQJGO5UxNDxqBBz7pIWglhy7SNotybOnKLGJfVhLZNck6r2rWr02NW/OOu6/0ZA
27LPdP9b8ldfpjQOIDXsu4gq3EonBP5DL3HH76v1jz8ev8WbZj0XlrOS4Y1NBfYGoygWaipg8xEC
4/Q7pXD1AxRSBE1OIs9e+k/WeXF8UTgJxUoVdz4O4q1Ci9yHGxC3Ac+CKa5y4n38qi9k1zyu6exZ
/o8/fOu+V23G624jhCiv7GFHw7awyv2DRccLUUF8uXooU1R43TMx9Ft4Wq5gqIXHbJekmEiba3Oh
+kJR54q8wGkaedDX6lqmTCkAl9nfx+gZnCqhtL4zJQupC7Xc3DmvwljMClGCbu/nKmqBf88BiRr3
ccSsXRI8ufX7JNOa9/IPKmf2T4ckhUtvObEWWqrT/26yFD2KbnHTMtRSY2pOwdk3Yrw0uYeKYsLs
cyNgsi6Z1BKVa1bLesXKwHh8+VckyRDXL0mVopbm4AqYL9d8ChgIyWtJcv55fKrEGozL6uveU9U2
ABka+xt85eTE/w5zscwdJGj6RoFzmKIRCgkTBDZ8X7GE7sm+AwMq+5yBSRHuMshqEzYTF2MXnddi
XajOpztGyI07fBBCCqiUWjDymZ22GqdTEvYCpJD807C8lwSSNw/CJOEaly4028TA3iZ4UJlTO/d/
C0Qzbsz5NvOpMJyGFsKYfuFs/eQhojAUMfBVpgsWouCoFoo/6Qs+tSgfhMi4856psyvYF3fGtvZ/
9CkNJ6lIIGUVzaOaWa5bVhnkbxWynigXuHFCh8bGnv1a/LXg24yQ0fEzyYfsqn6pLc7zrU8jBWBF
XvD6+8fy8fzzVgdddIfSHzvfmrYw1YOdmttV2IeH6zWXb/PatuoXWp2kTaqxzFO5G59dfqZ5D2NX
gQRuC+ELG0fD1sEOL9yRyJ1k5036XVq+qEf1Fr4zNfqYM+CWTGU27FB9UIyYjD1G9oNLbdqOL21B
zXP7veTD9k9kPW2RKGIXUoHjmFmpiHZujafpqVXCliC8CCWu1imYNFV3V9N4eKbkFbrv3YqFZ/uP
e2Si340VQSr0iu8jPYPzyhTUIexxzyZvOpfC/uu1yQp/qQmUBNgFsVBWJ9f/JtiHoPb+RZY4W6bi
PqOSCi1TpVP7MJ2bhBqqGK78Q+M347qNwl63fKeUekHxF+KPwjqalIkU+fY0Yxpmz8QSmVGhnkP2
emZf0yBeW/8ZGhVD8oiyiqDy5h04tabuJETiFi8j7B5y3vQtau4sL3oRg70WZSVKrxgiklFoEvwP
lhOpWf4Yclo/y+tfXEk8IGAxFm31xoVg6hXEPjYmsXXaZioTan5ffFdkw55YmSTWDO42v6lxQZx5
pSztsTX3y3DZGtOzT3m+XUhIuQ/el/lNIzW07p3ks5qqiHNAvI+v1PXD+PuVOKOymjbOf47VB7/d
Rkgalwy2CK5WYNw8bmIwejS6vTaeCl8PkUuBgeN514mc5kcAiCZFnyJvTtThaMhDoTiT3xlH3XzG
yoaY6Z6zea2MsBeF+5ncOCdSfoEuj/VK38dAtHYiP+RcT01Cg8gmag23NXn2CkwvdAvF10J6+zA2
IuiyGRWrmFPGMmxk+d4Cc5y5gjo7MwanSPmh7HCEMAaXRa2wxZ/CzZm9TlUY3AduyAGhIkKnCgaf
iMoxqQRkUfFKzC0Sv6VWxTDWW5005xaMYFDqVDHJUI4ESPrdXBIj8TEg0fM43X/DGdZdM2XnNxYr
X0LDtTMvYtLe8ihmEs+jgKYIRDtthA/Zch6XEKbyZwlR3cU7b+u23s8Gyaqg5plIOilaEQ29NBNQ
EecAKUh3jEUNdLRbVowtLFnVRpcLxLXIgaMKG6rRlHEyOrcnI1zHR5PPx7gPeOqyz6ChFnVpOw4P
nP24A0USFmJM83l7uv20iDhrpkOUSroiXRoPoO0eo2WafHFOZaX8BCZYb/harcLKU6as4F7EzVCv
M0jBQ3GqOHPrP4RKgEoBtftIICVo9/eACAvD1QIh/uFMu+DM5kwjORwvUef0tYAFhDCsBcfv2/Wd
K6s1gYeKn6zOSHyrledMXh4UgDgdEOYLspSGVUUJDfEScuN8LVzGnYdL4UYxixq96ATL9p7DxMk0
T6W8qTZOpUTTDROh4h/0nDk9gwxTcKe+BEgytPlJdnln6FtLLdEaT3crABwRDnwIX21or6G/NOLy
L02ejxoDrCfLphvgdLcXzYMMkVm41HjbDc1dkVg6iQTS3ZM+wo9jQ7CLPz2fFcV679twegIGE8YK
5mLvgOjs9Qx876ai0OIaoDv7C9TdfHh+olizXKT3LlGxZPCzGKPW97K6Tm0Qphtbc4IXynUUM1ij
P6zq8b/XBkuKmMnc7SJ1uB2QCFfr2R255ljNv9J6G8zQGBQnCdYDdmSAtQPDKc5AwRser09zjs81
QQvhwtlv4/iAiIt6zL2bJhLL5IyMGuAO01qeKfYV7LDcUjpAXof4LJPbk8N8yaorALQpZES1isVh
OUg3v7R5f9x1VJ5zaZx2Z+YUaA5nAioXznFuBXpAx+rt2iqDr9MNwD+djUZSk65s0PkmNR48dJw+
n9pKcy/Vof31tYd8en58pLuH8VfH+r/m/WCV90BiAs1PYLisP+wuyyW7BJf3U0U4GxFKZ2TpXMSZ
MJFqn/D9TC6rv9YxnJjBS8/KAproMoAoxp9clh6XjwVYFv44+M13eyQi055v1o1iENV+t/wnB8rh
02TaF5rWSY2Dz+if+hpdxmW7HQAmrqrCZz+BLuXmDOKzOHY8bccFROnz0eSI+R2VXE6eoI4JLmwH
y1MjM1405L+LRGy+ARuZJ0e1Zp56mf/pH04LFr9ynaSQOyYX4vl10L9wamQjOJB4d8T2SQMDxaqw
XVkk7u4CfgXt/q3wvEa42lUQBTBEapH1f4/G5EBdxkXrxr/IM4Aj1miXp1X1dzSfAqcqW4WHfsww
RFUNytHg5ssGYxgGFiiBRs31Vtug9O+6P0RpfFNZYMnCHtqZug2XSFpDiOOfVj7BCuZ1VxSzjfvF
ZK9UUu1QtMtBzk956CQjuNozg49BQ5A0ED0J84Ji/sAYON7ka4RQRDGHMUAxXDsP3g3oMAYywu3q
0gmhKcSn8p44oYRhxXEeiNix/7epw080vl6cr+tryLOASSBEeIuJWhxMe/1u+2nrZm9OSIogR2D1
wt11auT7lyXuVZqCYf13eH9RHO5jew1nSmQQXs/v4R+BZ2NulKZMHyqW6TaNJLBETEDDIl2X8OLh
2fAP7KfetIIvsTQIliKYFRwU0oddw1ynCb1zGZj5eCCdHjm3Xqg5UUYvOhqUWvNQi2Utz+d5WAL8
jrSBI3nDnEwa4j7QrDs12w1XT5MCrSG2w1L0zIiLhvowBhYjbNVR9wHMSWrTHas6txGpUyN+6q+O
ChS/XzM9bYREUFqbKRtH4Oz8KrJ0wx9oxekY9PnjtJtSggfdSbqSmqLYjrnJh3pzOthO2NjygmQ7
9Al4aUwARSlgNFZ4ROGSsH+Lv7CNJ5tT2Q0CuJaUYspW1chAxmHCwQzIEybj3nGjEJSihlSstrSn
YNsdYKrG+G4S/Lf/w//ZQu4hpzMDFWTs+eLBiBhxEN1eK71L16jslZivfvBl8LzhobBkKA4uzXGC
R5E+C5L9nsukhj5axHV6zGro/jdKhc8ZsxtL44aSW3itgBVhgoOlxr4zYqEStQdwOTHOJiTNK6CX
jjwI81JI4iQIAFtEmQExloB9bpBEKo7eXWFjVszvKY8I9oOI39uNEKpcvXmqAtU2CeMwJPHpQzjT
K+g+q66ofCI+3oQbB9WtFJwJFOtAzDvFkoK8z9f0zS6gORN4Xwu5ttuI+6xiulIbpemzg2Gh6Vd+
+TN96x34xo7Ub1/KbivrcLQL9M/hwns+34qWw+EzNRJCQYYQTweYn4Pg3fz/Q+LiPmwSUDFwhGuc
/2duQahM9oq2jbfLHfKTILxRHiSmqJ/ERdfMzyw972xK1s1G8IFC2Ebl6oIHYfj7rEQRMZztuoBh
lKtUWktQDarn7HEd8Ky3BDKBaVCZc4M5h+nmsyAUIuRpG0q11ngtdI5OC68XTTqrV+JHA0tHAgjI
fe6AX8WkMWV2ndWRcHmtUIpAKol3JfEsHWZ/Hyy/exVwom5yO6dKs5tn2dCqUgpWrrecyfxuO0RM
3/mriq6ZKjiGAbeEmZKfIWTTsNIi1JiWLnB3e/EMRuuPN0Jb/r0LUdlb5VuoJVVE2UoB9N4x2oA5
3dpoviIjwjmUNU36quYIHbcHE1f2O052L59LbkJVm7BBtOebn903z1Dz4Th00a6GUiQCu8YvmBf0
YNAuM+HLOWF/hBwjtV9hIo3xoXEegmOpfOEwxwTe1SwuinndLYG5uLPwf5p5glBJ8dlK82IJm9om
lNYuTmf+M5xW6/S38qIsC6+Yz2GaitCtBaFJ0kVYOFce+oToqavYYd478U10W19gEx9RxDuqtMoS
bOmcas+nd9bR5uuW2p6Pt36jzD8FRyESnsqyfKpw1MSU5B9ugGwiaQ4hxaOYL/HDw2FYCY8pg8uE
OmuR7/dF1ix7+KQT2veIZkVKRh6Oibgol6lPE+Ne9PjydS9SzRJ3TWQHexO/FUwWjfnxYccuyH4V
QT7Uszq8Eag9ySbFFw+3mG3QHtLf+LyfbLKnJsi2oXfGpgKfindIkF5v/ld8gBd/tyLrPuSji5Ex
f4wFUIQLTkBmXKsSS9HYPrVrAzQnMNa5SY65T7+tw44mi04kuMRp3RSPh9vKhUMfvrOnskwGbABl
XFIhSbXryVWl5tFrBtbOcGAxgxoiVvqqmKYEHe9JiBRbHrBuN+YSMoMl2rj46iVHQVFH7Tt1to/L
TG1BCBpZc9NfjnryCnOrRMJj9HkdETLbv3mLiQektKV70l29hhG3jSDddbEAPZkIyxNl0kLbsXw1
uUortLnRWM+GDPZx0kLNMcrocUlahp5IADxJh4FLSyUvQ9a6IeHKPZ0eKLCYbFPKtlILh8mJS7lB
Q/QmZXWznRJxzXBkB2YQhMcSJMEry3eaL8teIkmzaGFmJhDpOaCP1NWAXkgKJ/K+87buRK6kZKtl
ewbmiVfdyfYvxKtzH+n4Q/5qGr0frJMbFI4647wj+Ytk1QaVSd1fI2PIag/r7Os6TFIGYFHq0esR
ZEk6XVJeksOqKuam9vvPPag1xUCTWxg7Ct0slqoSiSSBRwnBfahGl6OONAdZDsO8C/YyocQckaez
uHNjoGngoyhb7attu8EV+uF2mYtmoHzhSUz0crAD0bNVQFIesVyhK4uriJ58911iNSwe/8ySDqZR
dxkYsJhJ3tSBCkU6NU3nNiGyVm2NENgBisspeNKA40fllXEhT3khM0TWZY9OOdS1G6JRde7XDv/i
A3SNV7MBK8VccAAM91L63tj3kwCetSk4AMjia0o05+uBHFiuxza4EZAr1JejqG5BCtd9hf0eJSLj
CgMQUx1PRNDVm+6SKbWPrKSV7nnWy2+OxgmMDRbZIOoD8ZkwApwACKWB07Xej+NJgf3qroqmSvjD
ZBPj7dzNJB9FD/BL5whSEW6QeFKSIestTWcIQ84dwjcA6RKT3rfAmVnDRJvmKcoL2z3uV+4LaXhN
tolO6JCChu/I/oPQfnmSsBzFnv3BTh4gCKBFJXSd6ttL6b3B+TFA4IrmiD6r6sivvNAcPMjSx1Yr
qyQeaOgJQ9Qa0yKPIZqM2NtJKBnu301LqaLR6O+4kQO4aXSCx8CRx//XBivmNt6ynHpAVu049/1J
0qce7YHO9TwypitdvzI96/X4n9pzAwMLhpf9e5bbkB7BWPUnCVrBdrMj5yEQT9fNITU95r9UrfvP
hitYWh9lMQhLC5HxnoiD0zJSuMe3oUEJe587nJug5t+peQcRJBep9L7LBYlY8GEPbzIrNUgn3Ipc
A3u3YQVA+zCZ4CfVEQJyAYdVUKfUgJdE/U/EeH5R5oTJwazS5/Zl/GJMyYa3vhFXixTiLZl+RdOG
7e1EAPIhcKEUraFSktXy3zqWkTnH27NIbljkR+tq3PGnT6M9fgEmkcJCtWOiqYvzHNEmog3VJUck
yN6Jt+m5XFss0fp2S+Tl96eWNUU67JdQGw4d82yWg1klo69F0L5aJzqnZ+tdoPQeYKeBtbQrv/d+
q70Ks+OMvPYLDc3PLTDrngmmfKXMCsPZF20UWQ50ahc3waubAtxzAuti5q2TsWACH8K65TBLOVhU
ugf1OTZPPn0eb71Usk3whxUl8HbYmtlgldK9RW+X89Fvvq8jBKoc84D9Spb0kvIWBCZbVi1VNzOd
A9to5RSkWNDYipaCVlYX+vfiskgMz8qgP7gLWiD7kGTOSVf2CYeITEKbWOsIySm2Fp7UAVh/RDs+
T8GI0G5u2SUtY+Uz1mMKLjVQ6zkRZotOgNyR3AW3px3au8PlNBYJkIspr0TaTlC92vdK0Kbrw2aF
33QEFIcb628fWw2zB96FNO7LkIisfPp4L6niNxan7Ro043hb9RD7DyqhYlz0g8737sAmvKxiDNsV
Khqh7ZFEsqHbin+Ji8MQhHDDRKlNt2iF3A5FJWEeVYmI1zGhZIs1bIomz2ltULXuHFpbsRg4EtBW
FEtWD/TFXLG+o5T7KDdKucHmOKVofO8p9ObFxAIsvG1AR/IDQNpHBwrF3t3W60pYsx2pDHehDDXj
3hFaPNjtiJWy9ZBy+O7+I32NtSlsY6MoFM81OVttD7r4lZVCccF0mdSeUy/PhXJYgqd/Rj7L0KSC
HBOllpWxpzkzDk/VsRG6tLwuFJyJAVQ/37x+gl9LciTcKsu4rw7e25dIYr3TDgL8ds8nfmWeOEcB
OEURWhJqAxz8MxlIx99O6NTankyhDt8U2np3/L17t3EZvVMpZdzFYSmkGPSNTA1sXHU92nlZNaVh
QEycsT4UwLZct8hac9KSMqgMLu4mkPA+M7tQLSCT3h63FWZw754JhUNJqrCYI/OLpIw0OBpop7DX
OpxL5oC+q6ZjJCGDf74Q2PLQaocKodujtiU9Fls6zxMxQ7w5/PHaLjXt4gW/CNBuyNcOFdOeVnIn
kHlctXfFBEo/zFgmHDL4fgDlhlo9WOji6dE1wADSf7LNh42dKEMmlFSZ9MlOFC5z5LXykgdsSrNj
NjdDUtI2k/mcl4zntzQULDPrHlb9eZh73Q4raijeuJhIul17diaNOCNK6ZT15CSTqPwhVCuRmEE5
nFsAeE4WVY6vlotOSkmwT1vcijADpc4+jYMpb0MJH3X0fnueBz+X++5AoSZCL5PZcNkCbJksye7/
2YAp+zF/7S+sTt2LLetBoS1z7z8HAEoeDc6ezIqr9AxeO3yLgPp3q1fqEjtj3973+gTclbz+AJ7E
a3BYtTviXS5fdnjjP5B61Iue8MQM1/g7ldTerz+4YXpIhhJaQ6o4tGo+cCOKPWS7wX/sUCNXaCj2
f8pvdlmulBpuM+0HE1pOyptNjWxbPZhSbd1Lzqez3gRGU85kCWIFc37V455nX6CghctBl++uc1tA
SbENAW3yM36FK2OJvZUQcuM3dW824OxzbHRkannHs3lX1Fkc1a83FGI4UZtPQO5lFmh9svGY7jUg
cLSIa6xbB/qCIch1UUsfzrGHScAGfJIGQqJX9Cfg7ZYgRNDolRZOdirWfapBUO9Xw3ffkjY9WaWw
a2Ef17mjQ44HsPX0vHxuytqMZIgtA8rrpcttcTboNcuWqHv+qC0MbRFWZunEFt2iyAx45bNo1NFu
6kCampb6OXmxQH21dEhR6vKUYP/M1oMqiMgUtngINV8BlPTvtu0TNQ/ik2zTnzGfZQlfB3IwJOfh
eISAP99J2pWyrWPLmSIBKfpGaVNP9pgThImFNFV597Wn9h6oPT4KwVM7wDca0E9hRkp0oKoNcp7U
IgGfe3J7EVOIGmQWqhe6qGHQq1fYf+uA6hRKm78kh/1JtGibQQsSQWNYEh+jO+LcvQpFfb5+m5uV
z11XZtjhIG/9UWaj5Qg4ZDFamtuyoLezqQ8V7vGwJPF9TqFKyKsUXfm4BfYYd7Qh2KilwmkCSah4
ikfZ6d8tjNnKIOR50nseSZsoUtS+ht4J2N7BA5+O6e6jgDOtEFY/l0l8qb9jrBsSpWI4RihRHmLe
Ieu9e+Phl1dpUcmpbx7VyKciD2k1SP6lnc3MDwB1lwLvnGqiftZeqVS8F/j4XkEftbqsdfsRVij9
1oo5SGRWfvhXg7vMH3EaudJzpZIn/xFWKc5An6dm3rFQxxNzXMPfPEdLue4NsCHxEDU4Tjlr007f
e4EacZLFvz4wNgDe34rtcFvlH1bmoJg9WO1ghKg7M6E3apDxMb1neqLDbi4WeJWTIl3ME2p9jMbh
aTvi1MtHxr1Mqlalh/ubafSitigeZ6gLcxgq+HFRJwxyVC3WoPyR7aDSmpomUlJlMFEn6tdx4jGb
khea/1S7FMlmNxpZRAgqZniqzrhiGDkHBEhQ3PY8+XI7bRZvTGVTlzjxAw8pNUrvSd8jEzyGuTLT
5XBwI0Kyshj4pbrQbwg9uXOcswwTWp5GPtvv4r8yU1B6klF5X3f94GsULYLMxPTz1+0p842f4lEj
Q8fRaq/gglUFYk+erf/Xn7NiQsGDi8oUu/qReif0zwBMZvqStli2gZJs2M8j51dhqgMHTsbNi3hj
85kjp7X2nnEH3myYS/2pc/gEgbKeuZl64LwkChsOw2tZfe0Zfh6OYGLLbJAsSQJGECFVsjbFuw2X
LkzYO40i+y8aWO58lJvi4UOpVIgm970daDhRbTbbjs8vuPyejQX6+ggkiqDymfW4u9FuWU5zHG/n
POXP8VKFdgPhD3ZC2tTTvesaYD5iClaoxOa0b0vIHZ3hDlTvKpYpdw+rgjaCQEQK99B9Bzp2wIgy
zuAdDZDyAjCF6z/g5LX9W7LyvswL8tBYgpyHV9/v6AOJmmNBLfFvX1FyUr0ixD0SuZgSYD0jRn8p
dZvP9pdXN8uUG0+wTsivlxafpyz04mpcbvTAIbOUNOvNR7pL3mSiKbXynLE8PDlQgoyPnqOPnncw
JiF3hWJrjI+gpNcPJqqaikEhaV3YTQBP0/xRdqLwmoA11aQzqXqzupeXHSPaW98nY1hCk/8O57SK
EisimDKpyzNMrXUWCZ4H1aNNbAFxOw8kYwMwYS9yDSjRFfQrZ/CcBJ7o5cPd+Sboxy/YMAqaSbH8
fWt0krl2Id3n8D0nBVDf6z6UWSlrZP0mxCK+p1HJbPAReRBKfi+8tk623LxMWQg0L1kHQ3faQdRm
Fa2GkKdr7BJ+V49LSXI9PhQGdTZey+gi62gnNYheZ6riwmPWoMkiOYMhbeWm/IDK3M6S+h4CJSD/
ufrv2L8wILJC2aZtgKWSrdEv2EOXU2EmsiUG3lG2vLB5jp83gTnQA/pBzJ6NdZ3cp7Iiqe5KEwWo
zS0A5VdiPh8rx8W63pIZHf2ecTKBw4h5GYErzm1jsJ7taIDV734DNUz7og23hUEHhaLYka6TMu2y
D9lw2PmJSOBBeDTXZn5FA7afC0ZN7XkNDX80J4Aoxue7T1Y4IEWNrABO+W2++H/ca44N+NWJJR/P
Afu2jgy4TtK9OcOBRfptRzAoAkFNn7sJHuO7n4M+iTQOb2MSF76iFoxeNLuJ6UGDsAhMDRGncw9N
N9mawX8TH5A9NWxpWpbdWBlnqiAKUiUFvnJKboUWPdaAPwAlLDjR22svLvQPt03RMngO/OmPTt+y
xVdDZoMbwD1tsqBBUxDsw0QuFxSf1MGvzV30UUqaAVcAUqUH/ZU3mlkgwKyGQTPfhOckTFJCIfIg
hx5K0F8Rib4oOjSQpSjWlZoYszjs9h/gPI2xUDuxf/frU7uPJgmi7uxRlO2vOo+L3Jhjtogm7fgo
ILcGDhsmk/0UEFg484KA/5tTNNaP/iZaWT6eFGT6g6BLrZc1oTJB26IYzXKxRYr/uBoNxsBsj1pp
2XDZgQpzwNGgVnGwaDQ75CLu4wvMZ81urCA0YwwS2GtE2vAZIVpVVlUv4Qfb+ZjNDbLSpbF94LmH
kAquwto5qy4u872KRRP6uCMIIJw0bmnD45F05KfiImj8iRtiTyZZVLfqUsxsZaop8CYXR+eh3G1f
QqE6y4SU3K0SJCpKX06U5MoIaxHp+qOHY++FWyV5JfpRUvICqtQ+mKamvwi/ZUjumn4Ftt6usltg
N1/Qkfd15OYHCzUPCYY5xC7XSK4fQdrQULJp6Lg9wSnxtWoPyIWIMFl4yBsT2J8dUSlLDMwFUo96
xx6HlT3X73BwMJ0Qd+XkFfIhwEvzz10zgFy9/FbXAqWgGYKL2ezmK6dawS6pKehZ2D6uOLQT1ILu
Bfn+OcBTsRks3XmD/XZAnGDyTAmg1I3O+U85PixCiuHRK2UtQuySSVt0QjZvyGrtpp3THAQg8Hpd
iDu3+e3l6eviQ0iwSybpmTj+5BC4ZAKQVcqUVoJ6bzAZsDwV5Zq4LS26SF0W9wRQHflNbCAM4yVB
PIk2CgE1Po3J2FheQHMLbhiWSwEzOQln9OgyMQBRgf8k2c2+5EVDVZMDQJgnltQxZ3QJAtNuZ6f2
zU6RQgcrP9WFbp3+UqwbfmUmfLxOSwq+Zj1bMAa5YiwOt6SM/fv8/68fydHPnyclX7em5gh+kog+
BzMBJiy5TArtm5bNndG2sd/Jelaq3A70lQ2MAt7pQapRa0ONFqXZxY/e+rUNm/1dZSg63mlw+8hw
4J03b+hvrFL6JUzQFT/lezLps/5BaPq5Rt/pF6Yy9UdMB1Tj3n3Kxz4CXCJKSGibaVd1NUf5x+th
8E3tJTVAjdhy7T8EuhzCNIPe0p6TkJdn2iIDu2H5mOQ7GSDEaOvxkl86SkY0GY2fzJuUPpK/sroc
77Wg1JD28flPLgFy6JDleOtDefqpkIX8tzqKUY5JJyC4b87TocUZOMLYN0kR4lsC20k/w9It6MbQ
q+vXccj3LT6W1q0blQOkYLGXugAAl8Cal+kOhRe2Xq6Cy+NExVQ0l+jseh3OMAqbYYt2UYxlkjw9
ym2Dl9vw2T3nPV/tqmVGdlavN15K2ispxbRlRED7v0arwdMlNb9z0G+NnCPxnLsaCBvWxm/WMiR0
KgVi458wS2N5x7GXC+nXXTM/6+d99806VoxWApu/NGQRwdYKzVtN1K4pb5izE+kLz7WToYJTZohv
5sOHK02wnOFMd1YyU7KJ9WePQKK/e1BhspQP26DaU+Oo/J1TAD/cq5FAkuBSe/QL3/obHbVYHo5b
hwPONVW4SKjHJVt6Ve7oc+Jd4TOzHLb7YfQVtCMsj+8RDj4s9PLecnAFArwhLKnLM8BFXX2WA0k4
8ynwddTS7Egt7W+u97tua9xES9E8eU6OJsnpC1YUIViwT/hG3I1DOWj8c/OBoSyoY1Lp904W6n1I
geBSPdQZ1aDZA7Lp2bJHRoImBxK9yRkq8jIBzCKw4UcgJLeYbSk7xqFOdsK2TH0IpBMOxiUKw88P
5M9O55X1miLGCOaGZD83ov7AOIERM0qpqRmhTWfg7JC6gqMy5FXTjr2e3qjafLttYpbJakI3ShLC
CrKZuAr7D0SBNkiviNVy85xn6Wz576F2XFP9Ya9Alhsm1MB8GXYe5KaTq02ZySNqzo//hGJ5OC/l
9nOPVm46C1ytXwKGevLRqquowsEAtMYk5mInW+ejmAbC5qj/igHNSUEU+wqpfMaD9SMFagYicMi4
9D4B4ATsSmhycLFuS+O3i22QhLzfh8YyX3ysr9wxPxvBLQjxZMtjneOODFRxbGcRyZiyyFm48PN+
FQmZTteK31F1e/ImkovHBJsRSGajSinBX2Kl+KKkf6zlSmvv8KasoJBDK7USsNDCq3q4fipppq1U
6Bx7GHyCtPDbEUfv5yra+Lhuv9pgEWdKfwtKXuuai/4y2v9K/hb6XFkymCPznXCV6mSuy31KkiTX
V9Kl+eb1vVLb5SxUBInKPubjwKxIj4s8KcpfHnx0Wr5SPwZKx5PBx1VCo/BlR9Ldo3oVyo3QsdI7
AGTfgcLUSn7iZbxiGRDerNBF+edXgEqVIOW4y6Lw88mAbbDsh10Mracxy4v+FwLt0maLhnGVlW6X
SsjBxM0YZtikBB2YWTVMBGYJwXIYlRFNOrxaXO168RUipatEH8AgRFkH1BHGVR/vY5ZWnrykJHcg
G9rqa8mI15REcfM2Mnc/6t8qtGvWmSDL5UH3xDZ1fQYAnh4RzBTU9vDPSNOS2rA6CLFdR6wxc70l
NvyL2q3PZaEX6xzqpJckO/WxbmyPRQAdwd6E1dMuNtXhkCGyqKgOt51uwK6mf9HHu5PhEYvNo6ws
JAMuYsWFhgWNkNg2sv6LuSL2slPswNiCM7lQysu58fuEiQdJwgnZdwOxzrmKQGc9z+MEfSRidPTj
eWCTKlH8xGp67+0i2eAXcmEM7cKawUxWjP06gdW9q1pkRZr4GmMVpCmLTevTFjY0XBBpO73chzgj
2DfFD5Jwn82ocQydaD/ekuqYOLFu5xeMutR4ITLxxlwJv7/Qrw1gjm5cINHyrhbD7/beiazR2SXp
v6533V1+zzvmOp8+/aXe5tHZRpEw8mgtkLt4R8Dbl7Y9qTvhd1cWHQSUu6Pa2jSTlGtxUKl/m1aa
JmXBV04ts87RfZDQ+qZXCQaP+IvIEgj9XOvn7itrw5Z4OhfzR/E72I8ZN97fyfnHIYI10Y46RUyN
k+gMGUfu+ZqQnK+s4PRwSlOKG/W9DvqATLNH3oLJJjT2jkdrlpfLf4UIxJTcPmP7cDHEtr5bezGl
qNJL7VkIkxqg5MjpBxscQqPtAYapVz3hcLzIk/M0YiWOnH0DfO0Upxs4Hz+2BXP6OS7+5hlsGvQ6
ScHKoChgVQZe1wmlIqNpIMYgLc9MSEdVwEzAxUnStbDopR6E44zT5nikkQU/8OYjObypiNH6I7Ld
QR21CBFK7qtifuYaHf01FmjtZtR3SEDRyJ9RaPWLU8z+RHvt4Lf2LyRm78zB3ZOPxgmThIdNASj9
i1k6frZVFIUs7qAuXs2OJdKp6RQbLf2weofiiQ5WKMTkQhkA0ieZXJF4G11k0GU1auON9w/Ks8Ae
pjV322/jLeRiwbwhmMhrjRSIvgesEXsqUYImA+1gIfOYTavDdGLtsR9KLM5QM4zIb6k5decgbB9U
GhTwoeYLu/On4MCHczx68bfvQc/g1GD6SfG3NisgIecEye64kXlpP5tQex8KlxMOCGj3v6H84HCG
xtS1+JCq6blTCCSTgg0MC9fa5aB7CeNm0714WpCzMEPJyoRfh+s4WLs39zeUIjFy5UrSwGRWTIwj
lFNB24pOJARSzOacaqRlg0KzXD85xBkS6fqiA+8sGWQA+RSvDxP1hV0grKnD5UZ6P3eGO27sOTW/
CbvvM0o+qKmME6dF0oDhrkz7kEbbwF2E61WK0D3evwzu/3A2bt0EXW/U77Xb21RcmeXRlkuvQ1NU
LOpMhnJVaAmMKa6YqLtBCpRsAdgbstHyRIIFdZqpxzCGgDMj38XN1rl6L4xtNJwnhcGBV66oIjDU
rvcrPc8gXtjBsMWnSeqEx7JBZ7H4eRHkU86aAS4oqZt2QyVVyxRqCkFxU4+3L5Egb55uwTPCRvpq
jCjlm79bTI4I3DR505ugzsTfzGPCblCjlptxJ/SKoxLTbQJXqdaetsvJ3GM/cDgBftHMW8dx6IJB
laieLU16Ken02tFonvW7hsAvsdN6cuQdkIhn0G2i3XFuR5XantIEQumpA0fT5wExAPUHqD9RZjXC
R760VUCtJhtqfklP+htJT5aIm/gR7p9EAomHvilX4UnDTW92g6bcb5IwE+ggU7mScRJVSYRxPo3C
8yxjUIGPdZdLBip4BKStyXVBbUIe3LJRCIADeN8bra5JCgRVd1wbGrJhiJlEInMZclaGgtZjIgsR
JydbHKukL4FrMwEWjY1UF/nC0/myJRf2gHpJ7K/EeMckt5eH9ahV1CQdmdKwJJJ7cNFEYyQaBqPF
avB9GqrxMtdL3ZCkoSUEmQR7UMHBpcmCvJy5KhY5CqXuzLWKGNkeKBtidpBvIvz+IhWvR5OH4Ze6
8kbHTOp23/jc3i41mdXiYzwi1Zf7FdnmAyQGtedE8Si3fSO4yN73ElIGR4q+wKOLG5g8Ocnx2HLg
kpj0l4388Zguzk4GeAbgiQQoaNFBHWTfu+9f1heNc1vSY8kuMVOB8D3O4aR6FVdF1Cm7ZuOef8uz
D/kB99esleJ451giLsmrZZJLAYPah1L0ziGNDRwLv95SNlvQHjdd3BGmGhKPi0jSMW1qGz8CHTTn
yIss1HJQYjSOgyrh96KUrEQOrFc0G96FuYJVGEuD90y7AARU3iiTHSMLWyz96Q2G0kF8LycGAg8o
Mun/SZBllMZEPSKjMKOlav3cC4zhKcalFphuV/Oq7/V8o5Wo42OOekbb2/oF0k337wOtK5w1B2iE
85G3oYfHA+ooBlFrek7VmLeDfm6O9LK4x9ktIhpIWeE68PE9lEpO8p/sg4IdrmqZWq2Xp/dHLvZC
5ocz9KyjPn/aD60DjezbuEA+X4eh+kxmNCiBQgJlSQXP4Op37SKHvRhVFK95Zf9TZ++GgLfNgeNF
lQaCTaUPdu5hOxEKYV5l2y/2UytLen/TAMke31eo3Y63KYJ5yUzYrkJg4ZUUPCDfy2SjMUSASxs7
Nlbcpdpft9QpoFN+LU6lpZIxfSBkUdpi10whN0UX/WfqzU/FLYQMrY7jdqq80OvqvzPUh2BSq927
WLmnlNzVTSEgdmmzcWqdzKA1qkKRpVymsHpF7tJY1HpnKjctZ319/KVwqQc73apMEbrzNr/H4yC+
///RAheju2FPQHebp0Xgax2eXIFtGr0H3YeqNhQJdLC1OfhR5Hb8aCbnfoiZCP7cZ+CfjNlcQhiE
oCf3Y45uRiwlGCWEV/yTBo1/xaqEY9UBAqPDNMPCyUUbdU3Hp+wWMVk60kBWqF3HkmJtHnSHxoLj
2dF/Cxw5AS/nppoqeK7h/XxuL4dGbNJWkq6YIE5AwGkweFVftcMLwqHQM57XoqpTHSvTztWW7u7a
g220ttvKQmpztMDlHE8E8ktntJURLd1o+f+VrekuxDxyW8nvUFqzH3lexaaXxYCoDYxI+gfNTOM+
Hk2P03FFUxRMjQl/moWfr3ma/SnxG26TZqnJ6eLG872eEN7e+zKPV0mg2yYxWhUNRjtI2IgRYmnU
B/pwaPlnv5kycw6yzQo+H6dGFt+uFgmG29fs9VlVFKolrsJB++ogYnFhgqglLd5PlZ8IG3pB8GUy
XR62nYnZpIMXzLKBlcpXqG503KIisPX+7Mdu2Y32b9PuLFssgO2891vWnWGaWcV1W9fYc9wPJewU
2FNWG/ofmdNJRZJzR4z+A1lgfGJKLdu9U+V0V82UQdPo3O4Py5Rx9NG10Tx0JT4hgPr15LMhPSOQ
pzFndsmkouCfdLTNzvnP/udBFMYztHweJsUiS+StmKpKzewUwTC57TelVyoVmw58h5Q1wJ8MuaDo
/DMBUhVcbl/KhRPc1nQZZ/IQuMLcjYpkCfC/1H0BQzwV9XkdnmiB0lN0roR1RyKnNHkHG1HEMGjE
DLdG8ZrJi5dvu2xBDCvCVDzgUf3agkP2XD0IyFfa6m9U5CGv6E7FLxmuw7v7/yRZihukQc7a3gBS
xBB5YJCQzZg7MhXgz0I72Pc6oeCQFhMJd6Aue19DkEVpZzMC8hLqyM8+lF7LRZyjWJNGuqCPhk6k
0/RwO8JirIHNw6mS+aOCp+UrywL614fnIC1yXVewSx+DDFPSt2fNzYY2ptdqshNT3lDc6kz0y+3A
c4jIebEfMKb1eiRcN8sdOi9u2qXsnt+CKGFkVR7mdB+1UwDHnrKkXf4byGDGwLNeRolE0EVrln0n
E6ttO0pGCFV4u/OUkGuS5d0y9K5qOJK5E1IKKup62LVxWX5lcPeQSxb+ikGAcLkyNju6HzJvL10E
J/tFnsaWpmDJ571FyM5/mxMGiawo5NeYMvCoBwZ/6we+5FkMq79jAkLwARJlHZwHdIMz9ZxJBx72
EmalJC/muKikYLpEMI5LaQETM50hD88YpEQzY5+omYixgyK/5LUyk40nBUXNhr1vstSkvrpgm8Nd
mM26f3cNTnAchDQqrWb6HhVRyX2IZclN6liGMnbHppVyPZdhn/276QxL4lfbAhK3MyEnGUrZRaz7
i2V9GPon30H1LaeFtIfhpFUiCLq2loI1EQ7fA71xUmWaXPFRJbQSo58xfNF1SiDX1s4WH9l5rm+t
aIr/g38/s3z3VBSFffb4Ur2VE6+7rsuHrQBa8fZkyDMkMN5xaLyAipLMZR1XN32GXwzbm8xzcPtS
ZFb9sySCzSjG01LceV8KCTRYf2PCSNLG14kKXtomcxyzDwHme+ihfxCI8TTAqUshqMKQ2pF5x0XL
/yvyXjn53Eyvfki3vRGrc3B+sL2yGeysRH63Iwt5WHJj/Xf9IG5U6X0VOKMPXyF2W9Y1Jflsl33e
NPLEVBM3cGXt+xwovc5ygMk5uknZS3qHJymYTVXjJtEutdVgKlGTX+Pkp8CL9ap5vbOQkrbWaPKj
/wJX91/82me0diJlMsXdC9uMQX4vfi+NF1cOv4oSwxNek0eM8RJ06+63AjgW6GtufV4Lo1GBfym5
DZaxWDUNs1NQPAVvdHxTlTYccD6xqxEu6gH1aCi3RQaCzxpoPRlY/cLydAQaT6NN6anj+4v8ZDKc
20m3wQzKL12+8zy3YtrWvRqjwgeOrORZFsCEMNO0G6MMzv6bywdY3wMNujC9Ezs1f8oi8UuS+NbA
r+uqaMseOkuuyvITfXxosY0f6iVU+mtnlJui67eE7J5rP6emC+g86UByb55ICVg3Gro9Rhg0xYDu
53IwiIxL086Wu6m7T/pkRfD1KaOz3CDqwdRQOV5NsJK2lQFTTcLJd4ks7w8Dh9rH/X7h5Xq2V7Gl
xse4miDHT89v5nj/WfQtx2dUHqzUs5UiEyI+BAMT+H6nAe4J4siXy40kmB2L2NnwUUumBQhdUXip
PnJyjxydUlVnEHdtuKnL+A6sK6LpjlgTKReINokmOHaBDCteYzXc5NBVi1Ga5EV/CIZsS20aRxxq
uyyWzRVPEP7wqAEazILJIY9AvKJd/IhvVeyYirhLovQ1b0upi/idSabh0tXlI3vDtLSZBOLInowj
dYgKEz0piedl6rzADYc+viNC9CQ1UdKNjmeHLdlyrN/KNC0hwFCKC7YZRPl321ukD6CyV0nxO8cx
UXIJxwnrP2vPboVSv5+OzOg4qvdVH0p+vL9CbNVGfaKsBTPK6jK3I//pY5IbjLH0N1ymgyXhxElP
GnM928zALgX3pKBoNQgRxav6o2bBeSGEKDvxJOkHfMnK/3802a65OIvSpXDGrsx97te0KAXYdciu
e7K9B78mUFF6UkZhwM8LAy0DW56rVgFMQa0CMYmE8EDle+NNa6AdelpppWl/8ZwZ/uzBGylOq0SE
ABKtNPXLyVCJ3KXxcla44GdpC3+71dHbeGa2GaFOqxL3nvKOi+Gy4WJaXcRfuXcEIVQbIciNv6H/
M5/cmiUiJvEfu7xfKONY3HnEfQroSI247U8Xn6Xh8rYbgr2RMQODYK+7vXNIzavfU1HobqlWSHdU
kZNZvN+rIGjBD3mYiqh1HPtqNAq+1pgrvEc0B7gztUjYjYtdITazIsHnMCq69TEizoRwvnfIELzd
PdxydRwoPay2qyr5jpPZCqfKqBXby5NSVyhyU58QnmxSWNaLqyo27FNMzQu21ufpRXSF7YYocjl0
yzY06BT3tJFEqPSE+NyrmqEKcTrdEF2G3Q5Y/vAm844hZsIrRV5jy0jvNRvVMfeuMVG1sWFPKPwo
rf/UzgiAFkbrXlg7sntXI2ifwxKGk1WrfMkUJzcaoqn8EwfnY1f/N9lmW/d8WHweq/mRave2Ql3F
2EHNLoQknnaByABbn9nnI6KclxAaD4wZiyabE9awS/By3mtnk/Q6Gbi2SuaV0vEM3sUcYnba9rOE
4KG6eKbQxWFGwK2rugVHnk6F9DaGO8R0yOmmqqiqVIrmumS3IaVPTZtyrJgDhpmntpDypbNFPBQT
GecDb97Gn9WvvWfIii9YtQqR1PKGWdZjoNEANUYlohLQq+i0VGfg5A1Ot+aTI40g53QaPlGqUwOA
ns5HI8VWG3aaaawhInKUtwvjMTngqh/90e8o1GYkCyErpE3mFqXF7qPD5GgFbJEqQwHtZdpxOYYX
9KEQLKWB7A0t2JB6G8nL1Cz25Z1x12CCGQy38YSeVa4+ReBR2L3fh6cDbYkwfGkgK8hTaIVlh+o1
C5wgkcBCF9vsc1A3b0h4U5PvM45eYAlQ6F6OYwonsGdQ6b9tGomwVT0J1U+vG5i040Yj7LG6j/fa
F5N9kswdjBVyCeE3kGaM2w6iBFWmvKJelesJIzkzrof52y8X0zuu92KfSBBROgiIbC6fLqsDJZ+y
y9Q+XRt1PnFHnzXLTSGAl8sAPUhyoQcQDzlT6Meg6B/5vcD0zFe4VxWomYxNEUiETa083SX4zHYa
N2bowVZHmSmc8QHloePXbIdZ10Ajr+aM8R95kGBT3ecIIkmOm/rxycsWV4yVFSPaeyO2/Bqw/raw
zh4Ui0VSY/oF0ibBOkcfeo3R/2oTHhCgxGha0JJo2EdVz1JmyxwDhcn32HVDX0RWH97jqf6+Yo6H
DA832aakoTenbUZSW6QC6tlVhYyOELwydVZ+/CZYr2lQ47770mETs25p5Ri9vwlHCPXYuurEAAfd
eysJVnIE4NM3ZMU6W0/jhKtY8gtUE3SdSMECR1o0Z/WL6mqjj4BhhysF1U2dKyd+7XkttlYuSRWK
NPoigO/HdqEUaNvr2G4AaQFqNilLR2o5XbDF1C0HtjTH7JvFpzgAlkeaZSNJ4poBZsERgLXMpHFk
BudBCwUULdmFLigHFCKMd1M5dTTt14IYSaO5Olk8MPXFgUzR4q4v3jFjP4EJFF43fPmH1WHhCW7c
np4Pbb2qeW68NheVhxbCUOo+GRaPJZmBTlC8AznntsFpwqNDQNNB1Xg7pPP3W3F9sh8VxmSFccRR
MjFwALJR38Gts6uiWet+BPHeRHze+EPEjHQmeuDJi6P9XsGBRnyPDSZ2JXjmttWMDjCTxmhGDeQD
JbRBJeYTSnxnAESNZYxe913AizHS1q1Y3lZkMcRm+WoVEwjdHf51opRempi1oBg4GDgImeJ3uPhe
IkdeE4W9NMOZhi8VpirB5+5Zw64j+tCAXmnnX7wyl0fq3c4Dnnv35pXy6hSWgmuzv3kUyeH7y+k6
H8gHT8ribfGc6WNlEVr4yJBpXckRtqMauXFQWOu4U9m6u/y6pOXveWDSJ9SC2bn1u26NnIpecxUd
iEt7L5MiAFfztVV+r8e/H0WQ/jawecuK0aS4TWh/Uc3wu+RCm0y8TqYznepqMIW1aJAOSVuMRSd4
UTmTeXSi6OKiWaqDZyCI8t0Kyg+lVSJwNsPLXT5U9+oNZ2AahIENKW+qF6Hm/y3Op8GkO0JSe1V2
hIWzXRKY0AE04nI1+6Lra95I0PC2epdQ4ZBaqcC5aU3D6QIsBTU4s8C+EoobB9JDnDjtDXlHUs53
KXuX4f2UK/GGNAqKEpvxWEilbK38L/k8I8KR+YA9D1/CmeiYKf2rOmEpAHQ5KMLvtTXcCb+W2rlg
Oi1iUKAsZQ9gm+tZjIgqTF2ZkSqucgN51Ao4qPpjCw7sFjDcya1dZaQcYkn+yDsDyV1wk2H4HQhZ
w+/+X0gdnuW7GqAYO02p3FiYqzVWo7eCLJvIm8wnivTio3fMxBfd8aTkCcvYmzavJSUZmNwgGhRt
wI9Bje9oyBDdHQLPh21Gg15meqh02EE9Q/coUfyu5Ru++5YtlqOrQJ6ZLfHFF2riWWZuzC202sjV
prZPWMNUo99Z3xK6H8odGAfkd7NQ6mfFibb+p/1vvhZek9nW/lhemNEGcArwWqpZNfKzuGyCVhYF
d+iAF8c9goLruxUbeIDK+qQtYIBCVfCID9zo+mMbGTCkjMEDaOU8lz4cO3zyD5lc/XfJ+rqXfbod
IVH7OpbietSQ1hJ59Fk9HxqZb9kmPJGI4C9aumwDEPSHtRB+3/WHrbWmGuSlaHg/JgfL9v11x79M
vN5Nbm+nUfaPKmoLDGBszPhpYccfELVoNy0mwGYIxYfWBFxAVTbt/gEpQu7sVZqqw535pmIPBFVB
bGZkxmpGzs3xIPGSyKBYGTWuOAEgTGWg/S6bhaFzDFA3HXuLR10lI3zXcn71f43R/6ifqNzjs9Xl
VOy4BdI3EabRppIEE3RMye5fbMMBRP95AfNgrmd2Y/UKBWvwFio/lNxfL+P5yfsoALKQs803J2Eu
ZBTsRC0q+GoOBEkil/nMn2RanSjLzFE9R5KBNDJLs6oEnC5/SuoZeaWDJtdy9hvZBrpv4VLxwnhL
N0Xyfc3YNYysULyKY7q5TcwvW6aeHQO9msoapjFyQ0fQhx4TDC2y8OsDAal+BVFUMf1QqonMSkL2
XTJus32d8YrWxaMaDk6fgP+TWfSklFsTpwQgtaV+7jNiIOY6iit/othrwkPMI49QpMtfAEQk3TFt
qVzVWvMbDsdEEvRaJfPSMP9xcav5NEc74PYqeX+MSFhSwWsVdV9ZkeJI7hAzXsbu+3vJr01c3yjb
8OTU8sxHor8ICaiURgSVrZTcOXN+lXwFjjhQvhbXyvh+RbV0Legqma2We/LJq5wDpxzj21Zl+kyh
CSBV3TcGjom4q0kNcZBWE/FtYxvGyzBNmqQhJbOW92gpgZrey/Wd8VJcNlmUJiifZXFJ/F6Tt5X9
AhlhNa8v41eWmql4prsSww+yYCN95MGlLbrEz79kbTUmghm3J1fp7ZAQChAsKPvKqqiMY4Yv3T0m
/ZbBVWDTZaJRC9//MGkyTSWKTKj8rpfyz1ps3k2/6+7lGHgNeBNm5km2ocQdGaykzR8Xm7RE2n0b
FouoHaW5V3O1YLrs7W1Gp31M14PrcK5J/jDpxCT89m/B4t6hRz/aZP0UcvDlC4n8mYZ2UyI8nwTR
lPw/mWJ5CPJcE/TFMQ11zjEywL5WbEveT4lLv4ALXf4jZx7TYR1GCdiYftVWuTWiZhmUT6AM6GwL
+VS5KYgwWF+1wkr7B4HZiDf4LOCDmgmIKFE9n/AG6YO81N8n+YrLa+W0ObZky+0oaWKHh6nBphb9
uVilPf5FndX/p00VF8AraLsmCPX6oSteXQppcYzGpc7ps63GndXOEW9tn4qsOwZtXWmGNITAW3rx
vVzRa5TbmC//MyxUgyAtPvEtMcuPP9aH4H6xBfZobXJdTdTVkQQb3fuljpnhjFXFM/5hAGQYh/Md
FRxIN164qVdi1WE5XGXhFKH021raHurHlCg0TJl+0IwJoMK93BA6keN3TeQSOOaji+7TU/F+MsJX
TqO+31W8sROXU9fE9S/07dxZ9/dsAzuExT4FKFAO9bHLx5Je7e4hxjOsGiZwHB9stDZjWijhNIoQ
Qh4q3Zk+g7aE5bB76WHwBQvs9J5NLcNjxUZNhOImcfsZvynIrgxO6br94ptBAf03Kud8DOa6ln3h
mzgt1V0L3flCfeUVjU6t31Rx5m5OMKcnAiKO0kDRKjIhPkBkCRdcmqGhBG6jsIpe6p1BN+t/a0oG
q1t3BwOyhsHKgMEvPxkFr9e3edksMyBmjgcUsxFqBfS040JWV4um2oiVz7XevVzCbQlFNnTx9sKj
brkTZjY4CqMki2YegIIEOQXtlZKJl91wfNlyGiINP+FI0r7P4yYyLGbF1uCSfAdsTG+mWuuOzyML
bK8xNCvWOxh4qhnMIQd4OyWgbL/4bdWh9EikuH+os6TlAL4mT0eBUzne2Y4DSffUb4h3x/Hg3lzM
X0waklSWEOfWMpbuUa9I4jSemDOUo//Y8Q4UrjYVQYBIl89fSaouPwabuEF58UEgTXrcqpS3qV6J
FhQ6n87j09gCkANMt5x7JSob+B8JgTWpAlYe3fDlqc3CQQ36dLGa8KAx8Xwj3FlbNZI5MAFCgycH
U70mGrtQBvd6X4tTYn/QVzs1ODFQ6YSEFrc4bMWgYQs8ojI30YJRqZBuG2oQKcYN5JPlKyPFxDrU
ToOXIUV8W4yhKl/2timnUxzj+xhfoNQjkzwZZCDhVUKvZKF3dEGRJaJHXHvq6n3KKe9zBQb7Slnv
sNd3Bf2nQuX7L2wxFlOeV9VunSnR0zqijba1EnZDKBKogEqLBFjW+47TFZaW8vTjw6RIeV+v4nSs
5f9wpXO5VKqAJNolbk+kh39yNcHDe4mUwn5dRKuWMK/1CFKsYm7tlTlLi3AMwCcL5a25mVVxUGAD
j8fS4lzidJdBEFlSHXzjIwIkVgaqowLviqCAc/FTs9fbGfffs5+aGHxrP/6hmzGMTxSZc2V2NY5j
R7AGCAV5HrX9Y2ozerNXHC6GQxetJAP7kKS7O48RNNQsGWggd8mO/f+9FNbUChEWTmdGFpB/srcy
cbvZFTi1WrgRzl1x//HxH7v16vpzUeUQx25P7P+uWXaunt4qry40SwY7Gr82yvkT+FNAg4d96rNq
M36BN+Dmo1DfScxSTmfI7Lt2ERdE3NDztraT9IBtapEcrX0FwPXaRhZ6Gj0X46TFL2mZhZbMHiFI
4JCLiS4BJ0D7J19ST7i4mYxhYXVzI5cYvRIyP8QvWqdj9eY/7I5kzeKbA+95VbeQtlRCzFBE4Z+Q
lJyUEdclvJlNkuAJSAvlmPMS3/UsX+XXoM3Y45rDhzkdsF/2Pht5KtPTjxotOKMPIGwMFIemmjEh
H/Q1S1uDQ+gvJswWTLnUGE8y8f7xZWVo7vQx6Mqoxw+g3PDtxM3pDMl7wj7L1AJ86/r7ZwzcCo1L
0rHh7gFg3Wl5QBiOO4GdWGT3PKPvkJFN2JyMjgXMtLCF1syrZL6itKcl9VKvbjulkdsc2+hPpbGR
V47QQG4KJGAjykChD00L9vb4sPGgI0XnkPIuDsqMFcd2XAfc3FLkwltKK+ZUBNPtWP+jM1iWPcXC
ErulkybsAbGc5rTNHM+48em1ZyZA71AT2/LYeln3tE3bCI7Oift1TUDlXS2wzckwoxc0nxvzAlkJ
S8sLxdekQwVWbviHNnvbZSq/IYxqEDY1eFmtvwa1n2XCz2x0E8Eu8JvnspT9fEd200Ze01+lJEBP
dOKDeKvxBXm8SNq3ObKMRUCpajX+3M+kx8zkTDytafuuVWdWRhrXGMvdMqPxA9ZUZAr4tSFvNCCZ
YbYHCvRdqMPMEvS0wF+DsflE77BA7dtHgp/IArcyrAsaX1GOfuRbl72ey58JKoD8QNot+i/b3dA2
VRyVB8qXGso4CpKptfOBAwOffYgzKjaxJCO8iQ3GwWf4ohDFkB3rSiNfIWS+1CxPL4n6/lhJep0E
6Czjxu+xDWem9yWWwzELSI1a8gJyELlaPm+8vjPx4JYk5P3qSox9cePPaNqQ2Nx3YN4t19SMxVLw
pduK9pjo/E3cKzM3fiaophZ5CCLUR3WWbX0JkIjiAK2veo/1VRNm6zoy6ZO4lWNF2u04uIcHvw+C
HlAbPaopfcau6AUSpeuNhD6dGb4/cNGizXletjZ1uYAmDAtBvHU2UuXP+mpddZfDBhj21Gk+/bhs
wSsHJT0WVI6JGNKq34xSqIL9xwDP4KtnceIkJm2IndBu8pBfBRYsX+BydIlGRZ1pAF7J4rijYxqm
wEvBs1L1eEAvtOtiGPziybgfxUHXUDRtLqgbvkNTvGg0LfSuwgIastvVVljx2NxFQ+Dxdx4WxUiK
rG8GSwZAwcDbeDkwO5lfULyi6xqpsHwL7DGeXTZWsimgIr3bRqyBvwFgdgcMv7xVsTAC5h3rWIwE
53iE3cZ8qMkJrt/IBYPLq73GDZnBo38Nz6LCRPDCnAzZic1t9EPAK7sKk5Qby+zANEbjDDI2EVGs
+Laop+wX5/7iDHgKWERhVuufCu4UqC8BwCm+gI9jrvH2qv8oLbkgfS6cjhqeibJp5LrWruCD9IO9
3lc7Gdy0PINf1cukH4avMYBTuyxOonn0M/+euJ7ttJZYbiL+V2h08yYnr7R93C06POCJOuf2bni/
XXVFGJ98F7u68dMma1WcpkQd0CBjakHm3WtxPj0PdUrfwT1CWAURqjWvFGvNzh+Q5OfSv0NB7bYE
0+7mhxtveZmOAG7bsiNtMmBjwKUq3CehU68i11QuOt+AJ9hHtY50t6BNkVc3rTjJHabNAWLC+2Hv
E//62g79EiwWYA5bIRgC62xRL/97ijHg6VBuP8zvc1gm9HXEgyaZSgAcxbuenTyPGAumNtER4cz5
7ZNThhb4o4Q3bZSfNPV7dYQggojZXeYQoKg2pi1+jkfFgg0LgcaQFbOfs83hFPaxNZGXBg87VB45
HeYdnkjtkz5hUXdKQkYDRu7k5mOnmtUUZNk09UypFkVn9y9GCIdF/LwhS+kaMTEhR3VrCJgtsRQl
Ma42aqthxJFFiuZsvHhkEVuuNhE97OTqQXQEpQkDqHLZS0zNMNx1aL49TS6V1Mts0HYvG7nYVnap
I6nLvm9EtVvswAeF5KnVI+jBDDMQLi9T0yZ/oL+Hi3qK8pRWjb8NOzRHcFlaSzw5rEAiAAXSbx2M
+y87hzk0ZJIQAYeGtiluNdH8PkaRfUbftNFKKv8NeZdOtan38ICe+kG+DEhqjoWSq2RlNwUPPJuV
Zx0JdcKh77RtJB3P8grzEa3Rb0Fbqsm9uCXsxJP0zJPUEm+FuJD6PFJxRGSufY7tQYqf1SBVEhSP
ZGojFZPFTVKOHQBE9+duhUKiPYwCYgPkBAg0ourhmeLrSw28pIlCSWxPorPoIQ0tLJPCQqrLe12e
HzSRV8/9jJnK9/OEImpusllstqdzFp0IzDlcYZbhXwH1QG1m2qmXjERa8CsckilLlP3j8QcSRtza
D18AyPKAVkpvXL5x+SAV0zaDeAsj9wb/pVi+yWiLXLsLdiR/udSnId8/usKskx5NRx9ccUfmAez4
yEHJ/xe3j730gGXhlIFoszdxRYjyrw/6rRD56df0WDxYmFODpy2rGvmyzj3iUaw1C5t9BazTqq1v
PelsjGej/xRmQ80CC+dB6ivbIr2Vd4lghNYzrfy5+Jb0sSP2CQBX/RBBO5gepbNso041lbKkQH4i
s4gbrmGWOfDjHuAY5uBD/rKRo0DtzrNMokyRW7NtXQ1lqEBvH5r/Oky9UoySxiIXnqwusupoh9wj
eOWMuRkB/2xAVhXRM7qr5NIdacqVKhG+6VrsFRgs00mV7PtVxywX3fmUWY7xCErOCIBh8mBjl6gU
o/7Fx9LXiwctC7HLbnnE862O5BmUMOeYLJX+8ardB3bfV/9NGLxl8hPlYVFphpXtS2u/GlXoM0+/
tNMmdslHMXUWyua5vnySQjAbtFDi3oswPUEhscA30/hWnKuBj/BtCgEWAjs1bgtY2/56RpjHZ+1s
DJcl1bofzcaYNZONuaZlI41Jfmnc6Pf3B4DPUyaY9TXgGVLgKZwWHJrT1yAZXD34BB8kOkqk4j7i
a3XPHWinx375Puh3QmjSBT0cr3HUREy95N+eKhPAs8SCAZg3uwP1Mz6RHQzw1aUwTzMjAN8b1bq+
Ao1u9K/5h96G89aZNLgY0+syO/c1E080UtHPE9ezjuZZxYNWHf81zx2hsVgOcIBB/ZfkLJ2Z7kX7
feKbMU80P+Osll89iz2CUQg/6ptgxecmryzT3mHvjRizGeJve/4GCv2BfeY0Z+uKH3ipTFVxUSVt
vv28EWJY52UlEpfe3Yxc4C5sARO2qS1uwwxpe+t3W5pYrhPB+OR+DodXy58f95xbpnEHfomqgWeB
jnuYteJB1Xo9FOfLI34fEQ9LtvIBlfn5HpVsqgBDWQ/KCOpCgSQBt2OPRt2mDAxAEBF3fPSsZp4X
wne8WbV3gXZW4nKIvGFbgVZsyzjZ5jM7CtLByV4EunCx4IDMQxxJRkUfHOtrdqDG6wKod9dyqG2f
Nm1I1kR9k6NV4Nha+9ua3GZWE+0yJAzTbIHXeRR8eezGdB07iBKXr7H734LHAcQLP1xelAEl29X6
O+Vmof8mMaOBrTQJmMo6swcDO2D33xLkpTAe+/Pt/+4IdKpfPA52h5v6d+AaOgMt5DQp9khpRDLR
RVLMy94fNKphvC6OGBblF7eDKm6YlGICdAUuOvEgS6298o2ozuwJv0CDgzdhs13YnbIKxF3cZogo
2XnLRBpDZnR891vt7On2oX9XKSu2n+XsnLV13J+v+Xl/VF+eXyd6GQuYZh4R1ya6DP01sST3lzAE
0WkGNomScL/7V5kpVRt2CzLDAyTUOyLfC6iLHVVCsYR59IA1Owo1JEjiZUUA48fogR29OmSVr15+
jOIfIJ3I4ASX9mSWVP+r1DZgeITpz6JJSiIxLfBKdtU7C1xHUPOdlgzUzpFo6rvPtOTLYiKRt06U
MpCtOkEQD6v3Md9GLstJejeBzoQzRFmKCccOcK0fgccY0FvNXBM2kAyPUTj+4qMICrGbOeTHbOBv
H2uh9qfhl+f065xvvPhB9BNzN6vr1rVzknfO4W3cFla3sRz0R/jAjSP8AjqtALRpYJO4l/v+pPt8
TdL6XX5Y0xKKlxylt/NeAcVSkzGBi2ef8nxcYJc9tbdiyxVraj1HpYdte8bxPIYmo1Su0jDuD9GA
5rt9eLwHVbWb7r1r/p1OxZnZmED5Kg8uQbhmhrNb0Nq98Yb7Qw9sLOdopgHv4B+eqX+WYbl0NASe
/264Z/9+tvlJcr79xHXx9SSvv/40AppF+KFx3R680ilAUA9gBzN8z/0Sudr/cDGxkqP03tnSKe81
itZd7c+cX8duqs//drh9iOtPbrRC+etDltSvWQzttbY2NnNkidsB87HIKcRHY8fSbYPsl0dBD2qq
vtgtCC/iSagKu0pqANsslRVjl+wMnak4ZN1u4j8hX+vH1sudJ96ZbqD9jGZL9l3Lmgk82oeeIbUE
Iq7DlhOjMtEv3wg/ltluQjXvsnP8mcAU6qc4HILelJkF5UsPEkZN1IafVr7RaBTbaQeYba6C2pZc
VPwUwzUZNrs/LACv7l1F/H98udRzMhUphFJuBkVWrIi4btk+Dgfjm3FNR5su03QVQXCr+yFipjw5
WIVTqtYJF716BAYV3z+rS7tmhZ3hjgBw11csOxlX4gAaUbmZe+JMHxmnm6XYmmuB0dG6Hr0kWkeR
caUQj47q88hqYoxfbANxY5yWM5zFYH0dQPQ5BtklYAjRm6GoZvzSdeaAeZAIJMI/vHBM2KLXqd/E
TXUBKf/90szJYRpku5TEHdeFRQuQCk8FqrIaVOx7ZK+eAGIawqgFm4C2l0FTC162n99nbqnNlGbP
A0VJPQsxX75aA0tgOM3g6xflyZ/ILW1cdoNiWodefbIuZmnn0zegSKkHvdIT8pFvzOL4iCqtVvpL
dqtuBsEEQGBKXIFBH3//sjtc5iJHRHytai6JTRkosyPW86fhkv2Tml62UkWHeaA0A9KKTgDoE8Td
oBOQfc1i6e25P67DU+QTgDjbPYyuobTPif746IqYUy/IvWQw41h8xPHw0QmKigDK93Fs3OWUlKtC
3oir6KJLKDv/ftLZdgU54WJbRXBTKONrGRj6oaY60EYtzNHLS4O32HtvKqZTYKSJib/uw4uwYMqZ
RkYddi/h8u2+cF1IAftLV1G37qTnudN4w8nagoW+zVx/zUFaWtWwGg9vrEuIQ+dpsNTUBHWTBBQM
gaE1XDurDydd+U61B82VUBYoRStB74vrTv3WOoLkOAr7Rtmpbmkco68vEIvceTjK1J5Y2oszNQ6q
mu6drIOsX/cD0jbZ7Mo5Pyel1gjj7MacXRS1ucSPVxp8mlwk4ljRkb5GPR+tzb5Vpvz/9fxVqkjP
MbaUGNkmS+WYgGcHylZINgYRWPfa6vtvcj6tzxLrjdbsbSCr0nHKMR5s4+LbQJAGRBSI88JC4mBe
/VmicbEjA9ImPjs6mLg9f5s39jvgxKn9AiLg9CAAXqyjv/JZolP0mvX1mCpXzoNTff8+lW/7Lo/g
ddOWlTfV6IgfMnlMcAMyA4T+JyXeflDx6rfzNUJ8HCxc2Gn7UmucnwG8crKQGzhro33b0vX8t5cB
ULX0DtFmnDOzCYLCvzh4f+4gAXHZGXiO/P5166BiV4uJWKeA57OKptWmPE37SMzCFNgSMa1Be+0b
ZKtiCvWvJI6B7C6EVvkWs7V2gWXgd+QmMy0bEypxxtfd4bj1rUNRimpJQqQWU8Bv62bGgYRGRaC3
PwdYKUD4muhbe6clwfTYHwOX9ZUqTnEbFFu0MUOxzM6n2K1BekupFYQ1tIb9EuwtSfVaxbg3v1a4
Idl+BhXoNxK/SQC6cUrDRX/8AfQQ+t1U9q4HsrSxJ8KSYad/hn4uFWqrV8bzEuyqp3LlXMQ9IRYv
wA9ilH6xrkzgJyI/5scGD8nLlLU1prQjbTOVDmTQn9ILhlMQ9jHk6YVasoBGFBCbCPIoeNrzBVgD
sZytVdpR4pvor7vzgKV2hSQFXwmPa0SbOi4OKLQCHtI20sQZHY8H5wXV8zFqr8A5PFee3Jm+LgAi
JLkvTSoUDeMalde5DnjuRTPBEZBmy+nor5HAQZ4NqUw4CJObW5X4wC+gi/6LpNtIHMKyIzvYCwDf
l/yoQwh29SBZAmbw9GZdzBWqDp2m/IBI7LK9wRwVpHMKZofsuoR8lA4juWBVozaX9yWt6FGqnew2
GeuXp0tnEEi5m7foRHYGCXSTD/VB8Bo3qg2pYwns/03ClhmIbLD9VtoHEDBryKRQT0eu29ZhvCHJ
FiEoA1bMQxZeQlrxnk21LEDDSX4naAIvpQ9jbY8YehjvsAJo77yipCSHPpuE4nJ0pIYz2CXui5Va
qstVLJO8XHL7MbievQtKpmcxmEGhaLSOhQoIfUaTyMn2HX8m/V1EooxluM/yFe+CpZ7f2+qGqERz
4jxP8+PlggtvMyhCcI5yHUXi1BHB86zp59+2+IsxDfOnJYyYm1vKdTAOBcwWWNq0c3HhX7ozaEmx
sKBVFZr209U0JSDxSUCE/fHplSa6fEsqOk8o7yrZ29oz6iR8V9jNVC74P81OUVWtSrxSp5gIL0R2
WE7AWEU9Ufo5hTLznHdhtTxsQwwJwtSFA2n45IvPU94fTpBY/vfg2RCXPkz4jFvoZ7akbsLIfuTM
yHHdXaTHV25RyNZDqVpFEkJ7s3fvhTaI9u27ehQK3MTzj+sLBe2lJTc++208yrKtTVXCHa8NqN2A
+i95EtHY04NTeRibw9gviqp/Uajh3u9UQwcD6P0A0JPvMCpnj/Rxt+eU7XtAPQXq4J/QWwEocKH+
7hv2dWZm8Uw7DQZyqXJMuNxyokfrQwZfBsOvbmRU5tZ548mUd5OoCrv2oz3k6aPNvMxAMQaYmD5e
1IBf+/CiwUhqeLtqNbzjgt1Vmu7oE8BGI7i5Y4MYVuu4Md1CHtFShN9lGGj6kKabmrjXz/RJRWxz
OpVJuXV9951dtegULdgLRbK8eP0lzkaRsAC763TgzyYAXmZnGcOOUBnPKUi3qtYazAQi1F4NQNIh
LhijEhky4+kWICpC7tSebca+c+ieTuooc6X/MAiPfvqvWg7GtY/vbrYgDtIO3b7iQDLLuYsoDUsI
t5BQNNVDV5fD3DrkQfUU+sTFS43kDLPaAO2ShmQk9VdFdseeBnr6ntetM63jqEi6DJFAHi1asYTE
6u1Ri8l3RU8rVAH+4jvvA1gUQN+bHCp/HDOH1PP3jnINKhI3yuYSEbAUk1m55/zj9DDIiwpj04Bo
AowPxz6AqQZ09DPyyAySYBd+aDHSbvARSMWIGpwUe2OBcCFHf2FGodSqWzZt1SFXxHZGuVCONuTa
B4rdjIw9CJA2y920OJK23eryCVU2GOkj46I0OLuPiqo20Z3ea9G3p0G3ZQ9D9U+gonOm6gRQSzec
VlLIGM+jRFc6U3h/kAlp3yva/9Mt+73ZXIgyG8JaIcyvTLDL+bAxOpv5pMBE3X2/9S5v8r6Pc+cM
hrWvavR6XEq/5LLU1Iq9rNzIv8w7mQIAJ5WCWXetJrv0YBNZHDHOSxRFueWxPryo5eNOHJtOzXcM
nW3ehFixG8aYUeDO1o/vTlhWBx0mQddzzFDoRIVY4Kt2LJHy16Zexa8vVUjxQkQ27NZ/nWxgaEWQ
Yq2JeULs3kTVSgVPpRYsZ2+QACs5J7t8E0Gh+6m6g7mfu/16RkO1s4Z7u8nBWY79TsMdkelD6WVX
bTeN9FZvpkUS/1yr+rDewrlJFdC10eBHXaWw851pnTRPxz6rSTPtT1ugdq6BpjbLIS3hlf093dVN
siShw2U+ls27IuwE7ihhjDo02Bsp3vuITQj7Ay4/ehRpV52utOXdidxyE+GPsQSVLWr5sFmrX5BH
wYydbdZcxdiZH2CKx7v0/KE+WdlxDoUC7lanQsMyQaIS9Gj8rhzAlKMwEzdGU6GgLNgnHdNfE9Dc
Kz59Q2IHlRNXftu8C0YsgZ4TpZb+9pT9tA5vpYRl2fWF3BxREni53Fvr4N34QW9JnXYtv8ezUmWN
gwDA7bNj01an7z0KDtTJJ+SdmBJgfJL2NMkdAusNdEfPZv4rvGnRMbsjiXJc521/PBtdrhx5LVoZ
CYFX4uRcZcqiGG1IlAdzQCQLSw+CXn3kEbICT/jXAtrGh8G5boN2uHEVXJe8V4T5n4TFOTqFDalP
32/8GC182RkNpHp9rxyfZPliUPADyCW0F05VkqcuJH2B2apxM8bv3iT/KkyaS3gS8l0AexPhCIFv
UvbaYwTe9zQ+tPcWk9wXXQ3HPmSgAbTepRQ9C29ymX/mWCgn2b0M5k77AVryLPjD/oDSP8p8d2f6
ZempaAmjxESeOr8XLrOdNoQrOAQWx1Dtie7353Ganarn49X5YOxUV6TVzwHxb7X2A1maGpPFknc8
AV0LC+K/+yaiDaiztazV+t3dZXnlPh/NiA70LeLK66m4sjIfqZWBQ42rd4f8jtHQfUwWMSJ4LfxJ
/GHo3aLdu/YCpTHDzE1BgH1TdK9KyLgo7LRcL5x3esKDzuTppMc7+kPe0zLgU+yZOroymO+XGTt0
ZHurJU4Op8VOWm/88qJ5SCWhW6wrBPsr6h3d0UjQy3/+kp0OxuqFyBrMZ6IkovEiux7GwhraPzKk
zldtriPTgCHDPO40FiTMgtkWvodTK5P95lNtG1OZAc1K3qYebNLYlfBqbF3oubSPibp9txYcfndR
o1cOMRLMBboTk3F3xkolQMO+s5tdy5QluOs5h/GDEZETkydL3N9H3dnXGJoy4BEFqwtvKVQs+9hF
eZDaCadqL+6B+rEHqZmKUK+2UqLcSVzUYClzzLLrJ2sTySfN/zRw8z9ZtTK/5UKTX+CvcJyjBWJa
rO1M4L2v2G6jshiMErsQofqsmRCx4/VHEkyesVr8OpNq2G61SGhqrg+5V5Y41XJyaYpeb84zClRG
FpNZPePNCavgkAygrdM5Q0YzRLxzTZvriAh8FMliDwnp5Do0UhJmwE/er+Whj1pinP8E9OZ8SJv4
XCJ9KGQ2kz+92BPsyZIX2mGpD1pu3RPeGG0sRPSBNZl2jvvOov6DZouVj3i9sEFshvXGU+SU+U94
tr0ksklP310Igd0py/jW1BMWYAjJtF98g0SfFF7UohJkvi0jrXn7zGgZwm4IM0D6e2JBS0f/hvD4
5ocJNdRVf8MakawG7D9yHAjlj/+5Yg3N5aJ4o9HdTOCH+ZiTzeQVQrzQ7Yx0up4KmG1fP9czWZ9z
fsYm5S4YxCRzYwxbXWa8DK1ICnrv+4HqywFJESH9cex4CvQrqO0DHyohxAefmathgLenIWvEFyL0
jjkf1VtJMfmOYYjjNv14J+ow8vAvAI5FhxjVtjs92MaKFCK0pQWWQJzQ5Ifw99eVogqLBhF+uygC
+sWM+FGWCpEewesTC42Yi+q9FFD1eAwvhIT+XV4YLLUzmdyYoRjvq8NnHLPFagyWRhKLg46zygD7
/X/tnMTnmn1zT4I+y+95pwe6WRZMoXa0rjjigrlA6k/mmtkoEogjKtcrD5SVGpQONATVC6oR1Cac
Cnzp6CaWhPhuERnQdoLC5Zc0WhRPbqkHhdJTnKQlN5M6AOa2cfGbIzPEjrd7q9n5ceBixCLfo7Td
l3GvATKT4LcFW35ZW43kRyTK3u7KXODIlORYnbDYJ6Rqi/zdmgQukGqgIqwL1Gzpt54QZKSNkq4U
unAtdjO+VRLs4dyxB0YW9jlyZI5d8LyTFIkBDLvVzyzogX3o0ZEsE+BeDU5eC1lw+YjLnLbkdmB+
j5d7c4SoNBr2RtU9Fk5aUhl0Y+Qf6rvTGRFvnyi8xqIQkhzsAsLASJUsCSHR57T+h0cTqPBGHC3X
yaHMRB7O3rz5mYXKFodO7Frv+jTpFs2YWRSLjwQCHouvY9OxVyRmIRNGPeQhD9beMvNYcIcRlLbv
5LgzZSESKKKuiWCUiyhhd7kG9mM18jPclHCLG5MJWpG0n2AxeFLAxKUgSL5UksbnoNh6QQiT/7Is
xOobspFudXbKAMpx/pJsQDDAR6++V53hVrY7xRQn4CDNbmz9/I8bLYsWwsU15jhV7I3ezLu9hhNp
2f3ayixLP/thOBfkL24+1IWtmwUyBUD2o05D+MLtfwOpeMgVWkRvX9aGtLGY21syh70OHl88wWbd
hAeM02ca9p7CFmWZGu7C5ftOfutPixp+CQV/YuhzHe2PlCx6RBVDaMzi+lRb8l9qaU86Yg13VWH8
qETG3yloUQyiCS/YDhFyX1IbxFUph7pHRgBHzLMaqM8P+IhJB/JHlZAeosQI+ogY+RcXvPII8nep
f0RhXoNEiB8lcGnqZ8b1pjd+JFplzBbhnsswNZo9dKiYIKks8ZKR62r6kLiUfmYJMHa+G+jkV1eC
cGrsQ8L+jAzJ79nHU5PfeeoS046WgyR5DNv9LkRIVyIjIqBqv3RzkEQdU1pUwWFByjTA35lqj82v
srB+mlG3yH3OenZwM/UMILNTxKWKMxyajk0jwFM1hCysmEaefuEeZjSOnAgRpf2mkMDYTbOpZx1R
OBgJfIRVb7wh7lw/6QqkiqiU/xDSQcmJ+e37qQyyem+HP0+H60LMykCIZRS/JD2BmizoN5BZvIZe
n27AwW1OfQ69f2ozQAuFAsrYPL+MlrE2lVhcAjLRAJgRrm97chbBLAJHbvP0w5+l2nLXACo/ZA46
pVERiOSCgTj8snCYPGJ12qXZXyDZDmnMONT7rOsdgSqPOgbRjmjzYnSpFpkcppGjGC+tnwTogLap
fJnqUXiH3K88MUUirqJvzq52TQHT5zxoaEYOslgfyU2e8aY4SNgPd9z9UXO35EuXodYFhXvg6mS7
RtUIoZlAScQyWPCf8+fjk3Ray/oiJZT0tRGOGmOQG4ii617h+siIoMM5CDN6Q7fxVEKgyZv6rFdS
CZdxbtl4ZgrWG2Afbyh9YxxE4Bl/y8iR5UDNihI7RvJZL1ae1tO3yzpgJXeb+9DgrDlLq0xWHNet
s2FOLeIffkh0jQMfXnVlGEWP//joQke83tTQRlmekDJk8g+q74sMpSjo+oPs98EH8+lIZ1Ec/UZ7
H9nSN1TMczlC3oMuQue+Lfh2U2TgLgQvH/QQHrElro3liSmEsqRKv+RdRfvBWOgOS6aC29+ivL/L
zXWJ3L4EbmZOl/OyDMsF1ip9+ewHHeNHE9vaIW4QDFqhrX4B7eV4zdHA+oU/ZXVYlCwoARhPC28x
pufrP977VVOoxLNyBvOc+fX0wlHGwKWFm7stE2TTKcxKn07erkTA2yLSXXXqgDKRdCbW3k99XsRh
U/Oa3qoc4/SHvzDI+SpncK3LDOCbwbvQe8BBwLqYf7Fl/xEAlf/vGVjcyzl2qCPSvyB4sfI0GtU+
EDbtwj/zN6dcJvxy89NkBpGy17Xrl7ohYB47GG9P57lskuNS7Qtubfxf2pPEyDu/lSQm6zkKQAKM
1w5iDpGqVEWPKVHufBFfHu3SboZn2PPm7Way7xxA2Qsiwe+reOwyUKpcmoKLItgd9FkKBNWDhHwX
p397s/53ZEE3O3qq8MC3kHWY3TzKCvKfZuXyb/AcPVRR8J4UWrH/ps5ecY72MacXewvpFAI91RLn
zkdmxohwct72NXM+ARbeNmkXnW0VsDbGU4n6p98cncA2T+/cr2KrUNGa4PlTTsp6UvtNmDB9bB4H
jaXk5ymvZUhSkzXSUNI7mAuRSLiAmvxPo7khPfJhl83DoP26UN91Ql/VrXzQgGHWWEmfPbl39hUn
prMMuqsr2e8z059Sq3LuMMcUvp2IW0R075g+D83hEOkm3n+3ofJDNjazUeyu62hCL6UBIdTNuX8S
2/f1abS+nDckzsU9lY0+c922VXNu6katAFtVlLRNLW6fkEx3jECrFmAC/XAeHoGBkfaFq8jUadil
Hi1eWI7FLndPw7oKV1Bp1/9/rIdZ3cfqgMkRI0Ci5jyLGFVmMH/U07BubFkcXINVcAM7yksXCW/G
EWvFAMIJWD9sXW0y1aPpxUJH0Igdfex8bDjosUZ7rZrRLQHlh9W6uOSwU9cRD4j3TS4zaKUWDY/w
dsmdUXYoDSgAz3wPUgtsIUoBi0tEEL9wcwOWuw90KHuSgzbLCP70JJqpQv/lA3qgUq1DM+O3y0Sc
RbYaXkMSs/8jB0ucHxWdryNFNuplDQGQaqdkxFBXz65DEVNmWgapOsQYh8SuhNu/R7RgvhHLPHVV
v4pKWJ3v++2v1VNCuCc9BWuZa4mr99ocIO7MRUm1dUIRbPtNfYirYgCRyH2kVSs3l/DjCjmj11ia
x1PXwCpoaJg2mccLKi8JNvbidmtXSIuhVkw6nQCzyXuzoThV9XJe6NUJW+Vut4erOkiqaUSEIvy5
9MZVGQL3jAmCCuKbBh8oVSPumOwORTBPuakd16XEZEyLxBSPySRJ7v1Zag4On9aBlvjo0ofk4BcX
ATV7a9Iuq8Gw7OboBR9iwGLBXNx2k7JANIMttbrYx/t+8HD57ZZn3SEjolMR2Lq8SxqtL3pARpNO
LXawi4OGYKJT2TP+AWEVpcNLeRBy50azb4Xgtgj4BdvUGY+UezTZwWrpXCLG0/L1qRje1sdCFgz4
xJNXWd91Lec4Rs8CuJYVl9+SFAVH6qJdIADG9vhB7zxksg7DHhEQu1D+BU73Ala8sySqDSKsgryc
Jni8kyiL+89ZqVGq0KYRCC/wsKFB+z/TDPyTxYt1egvHnCcRdiblfLnmUg5hliWNjWhL3U2IbfLP
9gVzvhKT0UK/soKaUE2zFjieeVL5EbWBGV+lnjXhQnCT7q7AWXBs5XHlRh/a1dJ//Lrn1yPmBuiS
dnBDeW4a04RleTEAFCrg4m1lKDtzoMIiNui2MdJY4zDNmclRD2a3kwA7aUxZRJOtJNCeLSrwhgZs
9g2Wt4ujUx3ytJ8GaDWFp7ddhK0Cq9r+lMXxhpDK0kaTOv6y5yGrl2tBGJF1w7gGzr4XOTr4aIaO
cX6TtY9mN7jUowcnkUgevWHngO4dzhYyIOt1qg4lcbqONygwAXKo5hlmdM/YeYKVsyTXOSTu2oCE
+zhcKrRhlwvA8nbPWBhCiutTsqhYuBi7C8z0oEvg4mUlKQzXkKWlX6t82FUKbMJovyh8tjVwfaui
NTTTLagPSoe3v2SK5mP0P1CD6LuO+DIPe62ypJaK35/MquPqROyuoFdFaAM2O2hAnKa39w9e1803
REPCqhdMauNi13jeAyki1s/tlvjA5jHgbTjffe6h+QbIcVcEGKPLrQEtKkR8TygVuYdLfFTbobJP
E7D8fe+aiukOzAPmVJi14KFIxPGW8I7h/QJYyIPRruQmV+WIJ94QQCTWbdTg1lltveF6RG8O3dif
PM3MWECmZ0CpnofevNUbRz5JpN0979LMn2ipjtcRh7dsNktEAX6aB+vyLkqSTVIeh3Af018w1Sp6
NgE3mIiErWhyOoyfDxkNL2C0A26IWU1HZ90Pq3OgMfbF95hEtNrD1xalmLh6qcBno/yL2T4OqPK+
UbUoi0E/F3DdKCmya1ARP5Y9L30vASocelCaDRN5M8II9QTsA6zOMxC8YDN1r2vlxMUiXo1KqGOT
PBPY9OVwWgW9HsoMkHdSU6sSnhZQdDkfarIr1Caa2Qo6fOFLTBrbmctonqUuZ6yxWzyCOHVVSLHE
IYLinfQnt+DhetAMiOXiEY7lIr1T2KpBG6i074k+fy+9ozXOnwCS7Ey5xy1MhNsRQeSIkuL9WlQU
7YL/r5LuI13A9EURHPAMgsf/NmJfciLre8XuuCg7m8AuNVWemh5k8mDWC6WK2qqfPKIUjCosekYV
gINohsELGbh98ttZLei7vBu+XjuamnNQlUF5ShcDhKLJ1hTAS/7it32MaFX4VEWthanYWa6B9RH5
0gyxrjzbgLrJkedSA6slpSWDuiapdpVx2r0fmozXLqoEpzLiO9aELm79RfqfEuUKn37R6rVZWeAv
GdsRaNpqp7R22a1yIomc6jeK+iH+p9ZkDv4wPcpgy8Zu3hHXWOzjGOSr0DLbA+RfboJmW2D2cOOL
f8z1MCdLW9ev+iT/AMlMFiEkf4/43+nY0u902AYlpqtp3tM3ZVEYR9k937jcB0E4m3GhO1u/JlNm
upXNNBu1b02Mvi8bPABVgWggruv8QxsP71AN2cGdtKQPNPtJTljyFsmCPSlNA0moGJ2BoilfrcRA
HtCprHdZmA2PF7t+Z/Rugb00fkjgU6EGoKL9xFq+4ez8CoNUr0nwS8F2G9tGVkWYRXQSjGYBd/4U
Nd0FtRzgb2x36MwdMAgcVDHK4BmoR+E3Zw7YzYGzeOsxlRQ7D7OHzhyvM4gsAzIK4H0BmGcm2gva
x0ARhvgItQ2WV5TmP4dhx5PdOGsmxFcIVroETGByIiVbBnZQHn06wrTT97px8T+lCJPUA6/ITqJL
HiHKmejwlQ0XihhJh0oQ7GMwcKGfr8KpEAjvl269yXWrlKTXfxoXszYcmK7Rn0D4cMzxhr7hNCKh
1LpLlsHWsIBdTO3v5KwLPzmwDalDQfkyWfAW3Nm41JhPnRLYcgjT6RIjsmwGkowivw/5p4PNaFbq
kveDvj3nlS3xDW9s3lk+4RhRruBDJ4oAlqLIziI60M5Lc7PNf2Gc9gpnO8mjOhg2Kg6gGw4oJ+81
lQSLsHSzYjQABEpoBvnXD/nngkAUZo1B+KpcfgsCxvylfOEwbPX+ZbobFWbNrRIpIHXFaPmiNYqt
BSnLaTZBU4iR/LZgrPBxAeN9xniOqXYw6qIfNQFR9Jlux0z+UlrJVe27jy5Qiq6RHwL7kyFyFLrY
OnnW09nho247ISq0l+7Y+uhulj7E6nZazGnlOEqEPeeHhjQwoa0fCRXs2BtVGTz2p3lqzFHzT9D4
dGk0h57Bc1rxqOvUo/0qaRBf4mer5H9XXhK65UN6we9qxpp+mflQYzApRD1M2ur5Van3JccwBfGH
W9KzWiLqxdALvP0xSfsBKx7o70H42OTDZZcM63qWy/ljSMM7t4VZmnmwlRTCeFkiOLSAJd3TtTIm
6DLWN3SYRzlI/8dUjTxyzFvLrukC+nDiF+b+/NYvMVVe2gaQuYS467fCQDcYgG918HQRMVMDe+Sn
SKKPl3JjNSpX3SphNdsDwqzImhzguSpX5fEw1NUhUrhBXPrkZqC9wmH2dCWVhAqc23e8Z7BoE4jq
6ir9t9cifw3leaUhg3wtxV0Yvx/rI0ND9AuMFF2YQYijdet8W2V3e9QABnnx8betSwjTfzL+A4+V
DPIHlAcdDZS1OPf0rHE6jzsNE3GaQauQr9XlSWkccDCiSf/mNyJcXh8Hvb7ESE4YAZKiCfvhSZ9N
4IiCxWyI9fZoOXQFwJeEi0J0SLZ/zg6kgKX5DitRRVLnuqHJ+kEupL49/4+hgySC3KhQLda311L0
sjT4in84wCtlQmOLP/JAjWP6PF6SIrituch54Io6JzstbHdquLmcw1PcF+B5sYVCQVDlRib+w0oM
MLEHqYG+3BsrjHrVWM4ivsnvqofmdDabXJwfffT/Bkh5/sNQJUgP/TqAVPED7BRII6GMFDQxpqXC
OpqhDn4Picx+D+X0Nuj7Qw2dWFEiSryJUKa/E0cKGn/1kaF8uJk0HEqH6Nr0vLf3nj9buZgToLsz
w9PFDMGEPrF200o0LRtIP1bD1N3ZLRndHy7d7iI7TIfRbUclQRvgULmTNa36m2P11J8cuf37IkE6
3I+xtGkB69OCglBkmdswboslABD0yQaFEdw+W7sX7og9Eofne8UZNI0+dhYgeEjSnHRh2MmRypP6
KPkjnqQBuxxUc4p1wmjYma9Qo4ifjWPalDVxOyVKITtlkmb9+BNFL9AdXo2tEV4/eZVpUaGOU2pn
qFWL4vYsjWH8dKZbGWXgl6j0U3Eq79VrsySd11l9BLlX6CfnSfamKB8kPIZMngKm58CMaduZ2nSp
szxQSkSksPppizRBMZqJ6At66gx/zZRAT/V891SK6yjPg7gY9m+izl8oZ0r4tXnYCopXOOkWZsu7
LRulvCCUvkQVazFPA1yOcmcX/cA/yqhaGJlxoAT9DQS16n+kHH0f30/60UGyi+nHiBkgQ97ixhVx
mXDZjcMRFO+qljI2D263U0r83ET9mYfCVUTA0CXfV8RTvwRYc3JdRgrUX7x9Kxl+3FGixJy8Dhbv
ml/RKU6wJgQLEgAmKyYLrtmnrJ2X0FBuBalDaNSVemFYM9yWPKF77lDjvNGKyKnQk13aIrgLqgC1
hIlCPL7rU1ALdqhVLk3zFWIQ8dz3+AasWCDb8sXCGM97wKYZAaQAoCbLGZn0dMXFU2u+ch+gatsv
I0SGqYOLYoNxWRlnlhbUXtWypj2Zn3hiDdtoU9MIZIWKzOfH/R5ghv5TjtTJQQyoAQ3raig/HAYx
E02hjGNGiMnnbP0jiFd0EJZzg9ic9TAcgz+oBiiMXmr8H6Pk7K5XpRs45RNWXy2A3egrNhDpM5IC
1NbYQkK9KElu0qDgjYWyltgvU4/knWchermSetkrI8ZSYjuq9jHtYR9r/0H93W3O6WpImk5EtA3C
qDP+xt6CpjpxxFbGjt+FOJEZWth4ArAl0NPscAokzeVp8kP0NbKLg8fS0WBe+poHBRycuddmVGJk
nXZ5wDUA0PD4NVfTdiSj2KPwjqbKgT6FJoWPY3yNHJliD/CfS9banPbgp5JaH0F1D1OjuI73T22p
ML06aEC6LnHypH+7FH1pZtVXEKL3Zz+bOedRcHvX+OXHl3y1UKT6xLvJhq2kApLdshee+0ArEAFe
xbuqbZhoRxZwR3JFsEu2kEJpuhuWEohe4vWj2QRYMAPI1YjFx4yjF9thwqAdEYXCn4iUXalP0/np
S9FzUeHYfVn5d5KbnA+TdyUFFTiOinQKayAHbgrl3E3b7hkQQuIFUU2pMy7MpcKNl+1mhgXtufzI
Jfl10whRp2DuUubcsAjT6u0uuWEbERqkDTucmIl9TGfmEbVRy33gG66biQQxhkE8KAk5a01ls5fg
t+2q17PDtl0Ba4mQlLZt8IRrT670j+a11fzI77spAJk+RSALGxbrn14HVAJxha+3KQZBR25D6rKJ
YAvBNhkVeWQ00pQ0MSxQceYgWyTvvU3xvdxeue5IhsD65nBeUFr3sRj+RIjRnf0pM2P+B0QG9o4F
xbf6O1v+g4M5kO/iWd69iur/PBoyFUxL51hzrAss/ZbmjVMDBhiCrBK8t7US//M7GhY0tD5JjhOP
1aiE6uwGsqwwbtp0wAui7Xbx/hGUE/B4Q23FmRGa2t8x7up8He8UlHkA5aXJBP6m/YTuQOpwFTfA
yfopw2WFMcGks6B9n8QLGApV1+dOot3kSZCfEwCHG7lmGb1kShC+D7G5oM6A1aT/27kfVq7pLZ4s
F9UcYK+sIPWFxaOemg01hBdzqSmbT3wo5C78t8oN+aQG0uspNKWJaCljrPQ69sRElDD/wcJGseB1
uNnkB7O5BpPmIYUuAxanWa/BSJCuOBUhCKJx8Dz23Ve2cmpmJyvTSTrskfaYDWINdWhMMKvRTTjl
AMLJnr2enK1WU+khMf08iEYhGR7uRgwQcY7wAj77ZyB5w6OukWBniKQAITDY8S+gpDpBCQMxeFQC
nlJNGRMkn8cJZB5UeUE+TCpU8eXYuYDNCrx4ANbDYEg/+RIhffIOhD7Ya2KsnUtxMgp5BaWhpedL
ls9uqxVqANoISz7qzWUgqVa4JUQduC981YH73FyYV7wHyHGxaNExXnO7/5//UE+URnd6Ssg5OnoL
kV4G8pTKnHuCA4qBWTPxtDZGCbqYuZXgSHKO8mCeXALyeFStH/ZM0kKKrNJPn7Yr36g1v9T926VC
SnL6D9TjQrkC7Mbtb67xS5UmmbzMJKJV+DwUDzLGQXEJV9ecViveTc2wqsfYjIx1tDbdkOgl0WmT
WjGogP+gqaM4bWSaYcmd7TAczadrPFcy56V+0Ips8XoVkqMao9Wff82hw1vNha/IXvzjWIIYr41V
nSFPXg6m4yUef9o0CPHpq6qKmloO1rD0IgkctfQdo9D28M/h/evgfE613H2XZFj08oAa68Lt8T4F
VIE+AMpMCWT6LvTWyj1I9F9tlD/89L4PB74tGi2iNZa0fDzfYtSRppSR1YR8wEoDTFTtMdisu3Hm
tEDeW7bFOLfWcA95fEDewhNHCdk1mMvCspH8NHYa4sKZAUIWOfyf/vSsxWhhw9SK8Yc/B5ZBx8Ny
HbOO4lVLle40/6QDexHl4SRReN/vkquxm+MFv7NpwTOgeNqRSqnYZk+IAsRRJcRESgqdgQOXFdvE
3guwftd4fUaJmbQazNU/GdqQQc03ukP+Hm5sjoLYzP845/bYIaP/n7N0eoTU9oaG/TTmz/XRPRnN
FMA8ler87HuSAh4p1vsXIjkdTxN4Lqy8Sa8MywCR6mYtErWUksed9nwRZWU97OOpQs3i4S0fMh5r
eaLlHNFtS20hW6+kvemgwjmrIhM1t9L6H+uFvU1kPBNo7UbyYBPSvXXIGEnB25Bmy7XipT1tNi9p
3BwwskMV7BQEAJSXLUthRhfEjjwjrx9guo1rEsOKTqS3Gk3bpWWElujX1xTqy61PpZq/LeEvKn2N
eRs8tETvpuz2BcLr1BT+gqqRGNeiEbHlRgmZADFkYRVIAz88RrN28mLNZJMneXllkyAIy/zv4Ft6
sEj2ihP4VDxH4+RoRU8vn1xEg8+jzuTCmtqPimynfbT0I2zC1X5LzG01+USn6uf4LdpXJRheMNzY
Q3vDBS5Ou5QxUG21OMiTjACsBt/m/XuLxcq61T6f8K+IxOuHKuuSPxYOD31qXMUudlFx/ChwdJK/
3eNkivCLvgtBG0zRhKDtv5BPFucu2YUX9q/kEtBaA843uli024cI535CmigTDOU/KlBsDxz4gVnf
/GJ8Y6KjV8v27KvdBP/cOTXkhBnC50MHPizTM5Jb/jonLwgwDcv3mkiLGbtHMkjkYKkyFFPpAZFl
W7QzIcO2J1as1B97NooafksnIbbza1RBJlrp2O6WIZBdRiMHrUgAmgGy5kSghZUToVgG9c0Sgf4l
lxJg795xmxgkPHtHw4pfbqyHiT8Fv9+SbNA9aA/r7mQOXXoZi6KADMmVDY+3Q+ttW6xe9/tc23oh
OBFVUBN2txBbHVLa3U7X4arEl9sd9a5yQQY2aEGQ7oapWBD7Lz/rn5V9/96rK5h6FEhFK5UjFeH/
koU0RGq7slEYHBFUB/EZcWHQS5yt1EuSoUNey4w5zbkXHPvo93OXn9hPpvfHPmrBUe54Pgac1wXy
+/dWdxNodUnk9Kzz92pQ0z9r7LVuSTccgdcZ8zh6sQwFhX13Q7w6yiKbJVm8QDoDC2vUzbpTLmHq
5vRzsPsKAILmxGxjgTjVgKce+3m83KD7pjRbM3jl2t5s4Czq/IfVXYiOmTZRN/l5F6hYGGP+d0hJ
FkLHwUQUekt6lQvleQr2YK48MbBWnW8OWvGr3+9FHq5LsH1PRrujDMSi3ZuvrgsANUXj5Ron1Obv
893eqStK/rvDdW0kmfCT0/c+xeKAk5QfAKqCJJnSTvlEDk/Z8xEwMK1PNzWcECytAvcHqYvry9dR
gYmI2YB1eBlAtrRrj3Lndc4JCFxYkaxtxCKTkrI6MLYLdBgHavo0jqLI7rZZ6UhefhxZCYsZKxyZ
kC/HfTTb1huxph+Yq2tTHzb3caDShVx8PBaDWkwL4Y8IdGs0YgWe6P176MwVDYA0hm21RBP0+jQY
qGsZkHG5FPI5TtLvwYm5LAD3LVE8jz7ysxlQ7gDWaJK6MUJpEowQsXLr+foTLzcKuSBnyx4d9hcT
Qc7tAbOEzit3Ij4z93lOVRAF5qip/tPNgKDftIpR8BMOE7nkQns88a/OjXgyyKbyUd75w+E5yWLR
EcqjaJdB2jBfw1fjc2OX024TkNbHTEtcYqnYpTvEEzyR+N6w5uFy7g+CJkPmCcfUmYasMa3W2Bai
qjJxbB9nKTmJSRg8gsG0Xt+klo+zMjxqHrVI4JrEwecJ+LWQfqnUk3E0kmYfjc51QmAryg8Bd6w/
aCxTpfdl8gb4jJh/jPtPq97njz+SVbQLQDsE30J6b0NBxTRSK/+3ibi4j5+e4O4esJiXzRC1Uu+D
yOdTOmPWCDWdzyE0IwKRvNK/EsI9HCg8Pp+cqNS9NNONw95qYRwPbzPlQruh/+3oOhWURwDSIiJa
PCXJrrzanRNwRbyjFnDR5XYQyb26K5f141lNpOgQMiHlWreuMBYNYbs1EBKd5e6qbOy5l6zpj5QC
EMfOKCqohJ4Fjrmrd0OPau0VhqMHKNfm3qtb8KOhGivZiabtUhZBs6A3u/cUC0pQUeh6lJRGmsWM
OcM/pCy2Cb/wJ4C9rt7QwLrd0QKoW9H5LStNgeA1quuZA38PJi8PwjvB17GpY/GRZpEvmt6Ifc9C
CaoRmmuwJGv8ItB7JMbjE/2+psmCPrCxiau9U7W0TEiPxz3J18EYy34WQATSZ8pgnR3asBhwzwnY
r9igx5cXIwHoyQPCFkq6NJnCjC8MdTx0Sfs8UFEvxBsekYjwax86buQoQ5bqwrSyY/QAg7DdnmuD
Ol/Y7QNQLNy3I+nCp8Gwsfzeq9Tm4+8qe95/AzE4nCVR3tfh3TTCUVmW++RHJNLDh5uW+gRMGWFH
8e+eHroz4AT1vs2D8Nt0+SFvyheLDDsb51VjdVj1F+K5b+PR06AEn0lihXgDezgi7IF/gvsN0JPV
iO1hPJXJ2qUksWV1oXrMiwyzyWcAkx1hxy5yRuKCUQELBTuf6EOmLGPB1Wr81sdxwz8JJPmSoP66
y8uk1V27PU0weAvZKHXylSKVpwmCYCgM3KvbLuEhKlxM8fg0V17UILAru5+wqkCyXFLvmzw+5lJ/
jDEsCkKpaFHxXk9AS2+Z31vdjMuR/NadDU0np8O+lOGfY/o4j+wvynVJMXF57gVwFas709lFH0VW
w2uhmHtS0RVF9cK8IZ5HWFYAwD8x7+/QbKVTZvsrTUqk1cpsG3MfebX/2iCvCwyHBX0KFEoxkMSO
wsotm+T0o8HsBCYRw47jgKW4HK6sLDD8zMm/2WjiGPzA8iktfTlfi89homCSLdCEy6ROeicIKfWQ
PURbQULw+okU4zBDC4iTRSAJqx/L0IhuHYzLVkTPIQOBCSltA8sVKy4iDfisCLYexY/XWSD+7ETn
vHpYEIDn8yU/X4Pzspq+adA+KeQrmQENIJ/btYYNgTLemZVijRXPvRCyA59VYiv4esiDJCDg7DLh
euWtZtI0Bq1wNp2em6HkC8SoMNYmpaK1QF0A7duGkmADG/48HxJ3jIRlJURS7fc2qtXOqXFgWh8p
H9F8dJFNq5N3tqfhKI3FPpuu+dcemJQ02X8QUlSFJ+MFhfhEqqSerAkXzMOgm13C+ZvRhENuEzZg
5IuvzLs43jbDzqVa34XAhIceFVM2lBgK4BN5mXnw2sarEjbMPHEpY3nWh/xM9XwF2A9coMs1gZHR
o3M5XzbvkyR+eprGxcFuz20H0lVdnT1X4QekhMDnsZ+L0oowapdRtLOHfwRkZKYTRlOqI70Y7rD3
W1LeopchFnJ1gAo/tC3qutj+eydgjRdAsRKb3bKLIhRhyyaQPN12xQvgaaHWJBbWAhWCUhUtqJJZ
C1IpcKwRW+BHEwpaImB1KHuh841rFVM/Skk3L6FOZyEQtDymIK8skjm29hRJ1X7ENd3IX5BOaNu/
vgfv3VyVZDuifSOnE7oJLT4ouYTNItrtnMtuzGr2SoNrnXtXudoWDU4LrVd/NLmSKFZiMjhFI8Qp
kWnPMmOZiAnq5tioLZKBDEdjFkzClZ0iJdgGbFBYP/NG/REgj2NNtgPF9tb5TYvwFREmiTCapFfR
c0HTnhGouLDRSYCFYnzcAcGnZskpgX1QUeYjwOkBvF7e4AIGeT60WkeODU4Hac2xgjk4rHLvC2+V
SEinuzdTyDDNhLFO5Pmo2K20Nm04eGq2K6Xz/qdwk0Egx43TFUvurwKHZKAX2F4G8jvgvPX5mu1w
7Uq3Judgcl03Vg5emS6I3GlRsM2FfEgNweP5KtxMdtJ7C7uGNG1z+pNQ4zWtmeGQr9AXZTjVjSOX
lytiyBSqn40G/xNfWIf45CNX97m5OAxXJmoqNUvK2QTJp3E8KbnSnqrYqib4aiCHr/3av/5Nj5ZL
jnvO2RBugZYThaO3/xJKS8RQKLLKXR1PmY4yujftKGRFLqEOgxcTWmTWtCpwoaFv+jztUMfFIaCd
to2Q/vqh9/V/Xeoz/E/9S13hzNLLabrCRSGV0f9G2WStXJJlrBn89kslN6YN3pnAP9D6MUTVWZkC
tZ8uSYun1Dk4/Z+dVvcTnUO2XwSz6PmsIZtrhQCWtkHp/Ojb2sfLY7dDbzlkyJ1VEPvGswpEikqJ
+x/GThes11fiStg4HYwzD4f4pfaxgvXjMtvlDkUDlFK9Z52Xmi1vgXL63aa6VKeRtGm+SFVA8Mr3
obgIkvxHuUBBdX+IW22Pc6NwOeuu3DvdcgcqPyzr2RGZ3gViWgyVqfuZE+6gX7PeA6oZgv0oLGZN
3EJ0JBrO7EDUVLWSOe4JfZUI8gqsmDuLNpVHAHrjeTMxJfhc6wmRf3P6V5uPkan8Jr3Vot+3vWRh
pWQlArLuDdOKJa6rfhSTV3T4amL+pLNIOND3+I/ZDYp7RbIL4oHfDDxQvy/loLXWCH53CnC68dQB
YDhmNjCFyvfwsSyvZAKNA9VPhAng0vNVfLQ/6ACUEStKPkvTdTceeMv1ZFFucfDKb9/V5G6BcgK6
Tupjc2Til6HPnefNi5oJwvC5Elp1ZRR2OiuLKFzCGEzet0p3zVPSXMhFDXdHLQxmKgNvFo9T/4hI
we5vzhXP1nCOYwyLYagyF1eGkquvUs3zcRfLGUBEwNkM7qgYWlGZMtXJnc684c1syxwvD+pqTbjq
87nMBd+xN9csfRCld3RPbr6dFG/lhTQqO9Kyvzgux0x5BpHBKQfkrEj8n6QqeAAFXUnjRmEMAel7
T2R16iD65KyuRrZuwPoco2epzrkrhCSxB35DzuLJgX/1ygPa4BOG1urOR4THQMspoinhFuyeYIJE
3Brz6AZDm818URPwcoiaYl8brylM0ZB9V3K2zUIL/tUv0N7zhY77wCRN7cbZg0MO0cFOn/BRCdNO
rS65GMZy7e6OifFdlX7QztmyEfjtBiMSdOr0q4o6UHMtSecvUbvqGt8Kb+1DzrrpusBl4gn+yf+N
EL5F/JoCcDVz24UDI/nu+3tlj/cAUyun9LAtxqc0O18yHaTIrMRhxpCtrsDRIW/G0iJUfvUTiV71
6GHWE6myfWLgGY2+GHj3n6P+1ft5pNCxBYCvHK/qBJV25QXziOF4ARCT8qP2YR5+g/0B0GFV0B9c
a3tSqKs0blguBEARCI4ZX2AniKASdO6800lVu7s/Qrgod6N45vW+LvGWGYtQk9+14YxoDQnGc9vY
A/FLA8XzJdqMjtj3/VAtlu1d1gYxhu7RdmVJSEGwL63dIRSyvRtIAJkQZmaGe4EGJdkoR5ENqBCk
/00OccDN48KJa+Q3U4cuGLEhlsYSULq0Ptnhlf7seZGLuBKgsN7em05hmhRk3YaGuN/WZ5zjRZRO
xbGS835fTFMq+TBD2v2pMmJ1/l4KN/I7WdV/15kJjE9V9JtXqLTKbFtzwd9le7ve3gH5dJWtYzBz
NV4LzdDQM1ip/baW9ELWDomaAl+kFnV03/RLGdy0DwxaHrNHpNUoAwC5QOcvxbN3zmL6YhrGXNZZ
xUfc/GUuB8yle4gQCremf8TzW8qwYWSk1LkshR3DFk/DLeXvnVxhS8JMDQ3pxSUaJZqllHTA/Zp7
ABzn7QuiG8P5dZZ5XeUmuYv9U5eimoT5n3mN4wXs87ikSrNyiJMZU1SF2hKPXcXrlt2tks3oyJ5I
MpIHz2p9nD3h+dvLaydFO4kMr0c3NNYiJ38/1Odzive0tlEZ3qsZ/h5emUZnHxNcnkkFi2hL+Br9
ZnM+52PPWE6JH+qpRH+WGm/6ijh54jsGChjSAB1TPOfSJU4fAptqC5bk2H5Yb7TndVURI6PWaJUa
WpG0iOdKE3df1kVOdpSKL+lwF6fY2c1q+7gLiojNNtawnXf1zTs232X6ZLCylNm5i0lxuzjK0DyN
w94xiH//VnoK/dbaHLF5L451Ox5QmVqBiU6A8X0eGSm5kYrW2YHgf4/meStb0mxtUqpBQ4bQg6Cm
LerXOH/ljLpT2fYcFvjVKZNW93DCAWrh55KKg/HaWPSBqaac88v2fZFmV/o20nZ23OjkGL/9PnU6
z1N1DXhYKhtylhZXkBSvkEP4HgPn5FynSm+PlVoZ3/zVt5O2747e7HEw/OY+8aYR/MoI4zyulQIy
sAN7FkrP0aAlchSrURJP1721kNgwRfF8b+4EDL7dzvFjsbUG18joRQpEdbekJccIVBF2jQT984C6
T+fdyKWLiWdaRixn1E8YsSRlni6Vkacavc1VuuKHm8vB0IWBvmI7r8oKexnuygOTK8FMVomcgo9A
lKjDPB/6QcecLlp687OL6jb1BwNWWitK7QO0u7wyqhi0DB0plHluV5bngu6AVJgQNHiBTuPVhJgF
kjndrxb9y1A0Vyf/FdhOm4O/8uJLD/JnzB7EE2QsMuBOocANjIWJBa2Szuw6uxFqYdIDpwKYfgv7
KmA8VWn2/RkcwPx4nRdSWAOy0jB2WWRlxjugY2vHSjQeU9fNbF4mb719y1GbFOrfIymoa4Wso+Us
6D6SmRrborNbM94fmVIu16glle+IF51Lj5lUg8l5Wa0hvY7q54MuVjnE78FUC458Wt+JhmCS7iNm
0q5GLAgxQnZJMvENgQIJIpFnOzg4+fkOUNtNtlZKvEHxaHOFtG7oqY7NPzhq3ZSVesPbe7fUYLn5
zWboqFVN/9vlwN6Uw/tws5/6E+8wZVNwssODW/hnwFWU1pTtmY/mnII481+/cRtyR+SRZNG5XY5F
nW84JKpBfFdwvVt7GGVGGh9Ob/H9UebRUjwAglCyv6Udcmc+ymQwYQ63qbGIGhd8oG+UEn+4uJKZ
XzAl0Aa5vdeCqFvCXZgwV+ss8jZZUNFQEzkE2I/5eC4LXfhgJijHN1VFQOZVbY+Kviknk8L6OO2l
gWq2VVE1SAC3khjZLBdHizyKf4gl9ROL5t375cPQtbn2Xc4Sc4LpkPnvy+HJaQZJxujMmVLQctlf
U7QAiPk39s9X4w6u6sc/94YNPWD5IKMJW0yuI+b0W3a57NT2WvLvzP2sEQS2tDmGFnafSDdgodcr
0BfH50+aRuCIIG0bO5LppnkfnuyN5FZh2ic+1R2lnyoxLIWufO3ZKTezY3BZxbDYO/SSDkFkOwr2
vp7ifb0Pj4E9Uuicv86UFWMMhIm9DfNidleUOvFFDDRE8hQqe5ZIrivfdPBiM5I26Ho8mb2JC2CS
NiTOIP3FAJgmGqZ6XnsCJWSdncpBjDobLaY0YqCn5vmjejbuvAyhyX7vro0PoJLW+0Dy7PVK+RcO
9EiqhPI59Pd1flc3inEPzi5pZKUsk810lFdQ/Hr2ZEf1vOCrZd+zJGTUwKT/v1Os7ZYxWJiq+oEn
BrZW9zTWyi84uU16hqh/JaDftYb06psnndaTrsFgWQMPFKupS6frdpT/693kYFPc+ZkAMr0IYi4C
+t6ZC/oYldj456+rQiFP30y5SM2fPBkhpOEBE8FF+kBccuN63ppMPHqiPjMUidSLChAzUBW9ovX/
AQO3iuTDXMHd8rNxxyWVPZlKwdyL5i7RH1+tUegiHS7xJ3y91+1v+Zm2Xf3FHSOp687OuJjoEOpb
eYTkJngZgAIqU6bAdLa5MEYCE6Iu6i0MCfhB6BZ/dcHEhkZO/GoDdlgynGRD7htvp9cH7xjcEziw
L6bjbDL50pNAyh2qlWuENt6Ad+71JXRjBsaxaM/Ua3dVeq+LDvGswX1YHh6iZmgz6SH3UHGZcd3D
Xngmz2y9b1aHHz+sQweusPP6LCuy+t91cYQ/0WVgMYKPdvLQMZT1PXKNuM8aJgfokEHIuy8JQ952
AFmdMlLqN1GLujlN+YRrqblPy8xnEdP8z+qZ1Xu10OsCjqYqaoqq6ru01daRvJQIDZshPR3Q5iIi
uSc85OE64v/wFTxJcXxFNHx9XukXxR2dl0BWHssyAOZ8xOI9oyB/iZali2LHl1UAsc0YKhCZrEHx
8xhsbh5F1p3gWVXaOsUjDDy6BkIV4l8+gAXUP10aXW6mYNbDQy04xXQlOMOmRVSXz8068O1rkyAM
msjnhimgNDrFebIEtbbVgnclYSvTSb5LgleTkxKTbLSy78PVU+0juciCvsuC8DUN1yxygEiNKCsK
6ogy+E1yv8lTYzqPZT6aUjrX5yn6AgjBkmVtOleL3YCPHuyUCk9SsieIm8themrhafI4XbXK/nFI
1dpdZjBbvgW7oQ2B33NRl8d5GKiB+YrJYMj5ubk2fvU7fefcUG/u+F3nNq/d58PHqzis8ScJYi3b
whuxZMWfdsxctM+vZwAGz0wwZ38cW0YKPilp6+16+UVU/rrzsSjYZ5PN3Ew6skfAnWEm0ErtS+O+
KSz1C962Kx8jChSCHOYjR0FmxkhAwpjN5HD0AFlD+vd3k0wBRlLeLcHDuPGTkhA3hOot+AC7CBXt
PbyrNl7JdeoIB/BmZO+/kQ0MFXmVIDPIrkHA3nz+9H4hjSdxOmI76MGLBdLd6SicsZbYedW6faMu
Ezbu2eJzQs273I952wZ+oH0COLDWY7ciaUJqpWkkm4gV+S0ZxeGCbdwtRHfOuFMh3upnp20RW9l6
mHQOaB85w/qDvX09Lb+QpOAywPmffea2MXhNOEgtltAzkb/hXI4sMtPgnuertfKF+O22Ko9RjtoA
tKTiWUgkq3QgGWAfsr4N2/Qf4VgDTREvWUi+vw74ZLCs7cmxuTKqSgm41Yy1OWi7avRMvo0nBFz3
Z7d9TcnyzHd4l1FrvPZQGhJts16nneCMvJiQ+b/9bv/asAL2a4hRoCtPs1rADrEuRxE0ov1fq6SB
Vd08jo0facg9l3CUz+QifQZ3676sjBF4Ycg2QY0PKmGJAZHapKBU8kiJBP54yj71Imls3/U0YgXf
PIZiphb7YSH/Pc4djowQ2TXoQKVR6DeIPgODP4LAbfaVY4QozuiBWjP3vvWvWRIsJGV26mqvjg/K
V4dMuSCRCxxM0CrU5hUrYLlid2CrSdZNzlJ47q7yjpr98AQwNsOMAY9ZYqh467kss+c5ndpFINWq
oe7otTEcR6nj7hX+jIzlVK3YQdP5iVzm6ogAQZMl4e5BztAYNFsVdCv+f9VWMeyWbCFvIkkKP7w8
hYpB2g15+1Z6ggCj+j0TWOMd3v7mxL1o/snhCqcsCugK5F5ekGMeWhMi13pepIZ0GQ6p61Sk2+Zt
vDe9O5Vemrh1T7abXZxzPxyZKLyn33qFms030ns6XQ7VnOHiW9regu2WPkzwP8IOIOs22n3gGmRW
X0RbCPULpDAMe8fyED98i/UeyVD4ZWzv4g0Apa25KyrGTbr/yrRBbRiGeo5nMEDUasfGyk4/N+A9
6jYKtuZWMp5K8wxt/CQZXuQcesPOMr1nBA9V2Am8kCq4idSZpwrL44gjKPOgnS86OWzlhZzoZNq1
2/LZzVlQYThKoYWZoTghUJGIwsOdtn3tCtgDctKWIFML+mcd+30B7vPNHR1Jr2ru6GXu3c7SVozx
sf7V7r0lrZgMKix8+LLcsJ4NUV0rm8Yd87mpn7/dnSLKi5sZ9L+FJXqijeQY3TXhBfqLeJCruFMw
qUCzrCrtU48OiMDoi7N5j5HZjFTcFHDRwRC6uxQmTzd91rtjJTpUW7paOfB+LDAPFgq64Qu8DzS9
z4NXGBN1qmLw5CLio6y/DhGKnRqH6+p14mcAXbbYs5FWqqyv69ZdDFBgHBozBB8PqzQ+xc4QM1/0
w2AZsvArWT4KLyPfSHQprjkqotl3KqoDLTgiq6fOXiY+KaYzbm7QVVg4s0hEBx7rryoLA/xeCamT
dozKYzgkoqAJkkESeMHpiZdtTFlFjEZdxiih97AfuHSrgtZsD8crMeAnjsuRreG0N/71OEwttRtZ
ScoO6hZbYXFdrE2v7CD9dzr5EROEaVrUcPqqVV+VefvLu3FeZJ+6Jk8OPj2WWFhX4NGbwoWt1z0s
aA3eJ2lm+NmygmIJRhuJYjKLu55jkTfVW2k85X2TItGNSWZvBVfzb+UeOeBtA4S1GKMNkkxfb4fR
tNAZmz0avI9lY8wthrZFN/2mPCvEZN4LhFOW7r4lNddnNbAQ+BDnb0G1euhiR5aesjrTW3Um8Ais
oT283H0hDztrYxLM8FNmEByjpnLyYMqNyic8xtxy41dL6g6DYJhm/AXhKsprMn+rHGJ+8jiwem4w
0u3TgDjp6S6jCKxgXtBNCqKIuwNiwUypH5yzaymHgofmPglDyQwXfNLqatfjZTaRZAjN3hSVPmye
98VMFphkKTmT7Lywn3B/PBvZiY0OJm+WecezI6tAobaiG1wtKMkANCDZeX1DPhvTtMlIeb93aS1r
YLtqC2yMpIVCd5pDC7R9ANmsbXTdbzZIoWCgXOved4+NiJqY1fDesQ9KCwO2zLZb5FOTX95DoQgA
aQytl7IgnVywRXcB/CPF8vCODDwY97s4rFAPhghIOw5qXDvAIzXgasaKc86YVoxUp5qbNl61Mjhg
N0zt+xS7qUlyO+kvx5+bHwi3WEDnGjtAxzKu8bAOwS+r9aNmtcRclDSOJ5VhahtXj+R4Y7DzAWTU
dlNoMkNIjnlMp5AHB6LxdIFDuMynCq/u4s8k2ipmTJVq+a1eE79F7O4xrhQWV5crVg+JuO/crn+C
RsvjK6SEiy1TaGTIxgXojQx4GjKGOdMIVy+O4CNU24aF5qmEauk7b8OLPSSBZnZ9kjy0fdoMIcHJ
fRxH9DqO9E/4charR/ls9CeFliRYK94OMERN4MAe3HHv2N6n0avXo2X0SnFlFQXQ3BnJ91QC8P4q
WDtA+79MInYpGByBu+ODsNRoGTQH4Ywcbw7WvCMynnA7buN3tfl/3HlbD/DfLDDpLMWRr573HISp
ZROaaWpu0fwnlw+rP0BqI4FrgP+dYfK6PkPwqduS/zlCy2IwlDeHDlRFZW13fDpF6Iv6u7Qws3/b
9Bo5S4hGyAPSMRRx96a/+xGrhIrpXnOhYmjSKABsxlrhLiGBJd2xaZEfghkOL7k3YY/vHVWuTZ7f
sg4dgefyq3CX8cpuXW+tcdCG0H3dYXbw73BjOjicS5y7h70V+I2rPvaqqwRd0bc3qFkCRiuVYBp7
kddplSCBOCTy7y1lOoQPSEbVqUcD8f07axF3eWpConiq79FqGge9N/xRJ+AxxIti9zy81Rp7OB3H
ZuO/0INqLVZ3gwK9vZWIOX6YuCANY8nhnTBcktWSw5G51ETbbwhWROXb9yPzgnR7k7V2oZSfd/Rm
b4tAMlNRiP+cxV0AgZdg0RapEgmj0fBvqvK8PH4o1bPA10uxZm/8U4MhTihbitTDKJZSno8WJXPF
aNd6STOSIhiwlQ9oILh8zwVmYgoxCACYpBQcijdfiiXqxM7cIuHuBMRx10BoVEKPpMuda/B5TryA
aL/nxeDUwscI2X6cRoV63ohRHZt8Eft7uSM5eiEHg4yKVYZjYJaF68j1gVl773LfOoi3GZ7X81Ay
8/G4zHjDSTCCXSVCxMpbbs7lhEJOA9lldv9X0PMgrnydow5PYNRmmxIANJ6nWgc26CIFiRr8MWZE
Q4VWR2+nA2o7FmTDmQQBTxj0jv5lNnjy/r2eJxYVdjehXQGSH4QT5krOtRuWdU9U+X/RSY/n8uo9
O+ih3i2GxQIk0EMv/Y/P3x9EfFlonA47aLK2XRb/CutmWUPC1Mkyxhfp1QASEB7Gg5QQWezGlZmH
rxxAKYbserz5E7lksMtrn6/7kSY8FpuHxgHvw2kBeZuR6JRtEQ6BiKsgXNjELNX6HqRXcn4MmRZ9
0cT9QbwBrkHJxkqdssnP9GuvC6WWX+foo7J9vdsZQzR1ZhZVVJ38lbswjAMabHqq1eTuwPxnZ4Lj
DR8/BhD8hE98h/yD/tOqrD9Ces2HmKx3f86+sITTGx5682a1ktbVl8nejdb534fSrgIyk8UQb0hH
jVy4Gzor8V9W446d6LXJzl2vHZDpRoQbpFcP1QBlkcxaMvEqLvg+PMsECp8/RZLdCWpKSli1p0n7
yRO0klnb8aEl/20ONnXw6CzFwDp2+XrSqJ/pz2xnrHw/j+jxJfFRD3o+MrjhAZijL62QjNK0BeKL
eTK+SGPgQlc/DVrvXyKRrS6noQ6Ft7pmmrqdcchyNltpK3MY8ZB2SpoEMRLXI4NGPFUvUq8Jtq6W
GfHhFyPsGtqY/l187dyoa/II/B68O0Bb50i5HJG7pb+nNjuXao03NymNmrcGozrZnOMYRs9jKLcf
ZOLK5MWLWGhOTqQEbl7tRQXw7MA7yIh4oeynI7cYiPmqAiuiAQTYQvfnpSrHlJYzanPJCLGOTEDA
G3unKUiVIfPmWqhVe2Xw99p845lh8dxh2KyK/TH1N99h9hEEuALIsLZpTQmDohw38h929crMLEsA
Sdkc8jxjH9287gnE7gP9oCxj6XXMV5AKGKvO4O7RQGWPzuDf7rZaMOGrFGRyD9ZlMOAUj0C1uNfl
BumuTaq7sWFIM1BwupYfmLKv5b9LKvL4vhTs6nXdpl3IhiSF8lrxlzpbFl3tNDXnZ+SrQVChTmcJ
O2KIhUDVJJot5rFl+HaTUxGSzMPkaW77gUXkmIfDiDO1fqIqR2GI4xOlAW+g/S3hAnHtNSmzqrsD
tk/i046hNw8swlFWlgRBKj3Cvkd4s5khq4Ep/nc/hZ9kiCe3mvBRi4DTGkhopawGM1lzLhq4u6ZT
8FHP6iqdxO/GQhIY9KkGawLhG7wyjNLg1nhHjZGn5LjNL3rHNXHYZ70mKFe70fLOzjz6jUGEbwBK
TaGO9LdEDUKDpGcERsxYmW8t6qhEasEocckwJsCvL/R0Ox1dUs4aObARfuBaEFtwt3Fe8kIYukkZ
WmmLtqry/Fjd2R4U/eF0SzJvRbijnk4zQgRpoEF5E42ULH08sHb4Ng5k6tR94KkMXQzXNTuS3ZFu
8+Q0S8W2PO0UEdzp7t74s7y9PuV5d2XKvK6z/Fo2ZQfP7asmh/Gn2qIdbamBxviw+2JGlLDzOLGr
t1zOcGeIE7f8lnj0bw0GpN1Vz5xAjiKFwcsZ7vtI2Z1i0DHheNUYANu+GwNg1ylvf9T7V9M818w8
ejnn1T6aGnxDc3X8El9/IEAb7cbLuChlxs5pRxUQr282ss8N/ucdtZhKB/YonDMh2+8WFHkDpglO
4Q+XZNe43PJSK61TwWgxRSsf/O5xQFPPUT2FbcxRmRVcdOrtRO3j3DMjVGuPB6IMzmBhwbCGCz2a
C21g6tphvyQzN229NaZS8fRM6M8kHvA1RS+fFsebCbldnLhYwG0povtsBKsXC4r1z2bchqzGkSZJ
AgsPkJh9epdQMGoRYXLr/DEDl0rqrSKY87L3TS7R2c5pBWzl6jLkfOE7oZe6j/5wvkmczO6YCCmf
8NCGaD2BHVXr4tVpkpggRnm0K6ZeKY92qqudwuWauVNiX/b8uxZic/ieK+S/v0BxnZM+wqNBwVhW
Q1AYaJ7WOMBX8V1hyPlbZlMyv8BjEyD2U60zbX8rKDqcG4HmN/nq3tB2hrNHep6rxxeIKJjkv2f+
Xm0o80JISOJF56fTlNRGaWl5iEhOASTFpJaabs8srvYXbTXKY+NE0RqODRSptAa6vpCge1oMQwa4
1um0HrSy/AY7m9xFq8Gt5qSZ/2emETNq380obvgU7sAHj5OsVyxDpiDurdehEDMC9OwNDa1AxWjK
NXpyVj2XCwI4rGvkzlA4bQc9QjoLlWAaozTwYX1dWks9RHJ3mrdHsQ1KBuW7yccqOz4jrzqrUlUo
Uq2X4jkZUQ6bl7jO6HwQcUGoORbfOjHYz4MLgDZzHNtW2q8MlkgpFWRgFZ1H5bOPA2RAU03KHib7
XLL+dLPGQ1eJKryq767D6NKskRJge2xm5Kfbzpzwn1q4tPe1F/XDQLJQcGA5WVYrBeDVA5C5EeAp
0toYJSOHAuufaDwQYO48CwzA0tiDgqSJpFOFR7wTgPvUzciOB9WywITmaXcSMqli9t+rVIvl3Tf1
inH2gYrvPGlCtSXZPypoutahQcFELZWdB8DNLigja3C6jrImQWFe/u83V1w2UGyxmRnMfqi1Qix8
pmOGf/hcVrxh72DxBObmi3NA6LQ1T5Ft5Zdfh8oXEGtbM1fhsB1iinzv/Eeper5xUYFy86gyFZdu
HTB/gwQQqjfhkvc5xCuK4jrBTCQdncW4s8z/9cY9J4MfRQRk+/VL17LFNGkOUEDFVuTqBhrBy9OM
7wnyc8GECYSq0uY/EY/e0+/4k/F+9nmOaI8arc/gHkrqjX3g9/hMlZ+XGDkbTk9qdjNgexLT8VdN
Nseaf8FePe1gNq/j5oBdW2L3rZiK965F8wA5L4vuQY79ac7mDYkBroxB7vAKjK4Gg73LuxcQ6ArW
e90qrky86ufT8mBscLYYM7h/F4o9K0wvhwVaoZDmedkjmk4JDafC42dTJdRNmbRUUkUbzf7N98Yh
SbrUc9DZmN0Z2FzmCyI+bwamAlYyUS2SPtyiiiNo7BcuXchqzfR1nDJz/EEUEAwn1piUiWc0xxG/
Z+wXJvICrFlfl9Q5MSI/FI8qwMrk/mCwY9MAzSf3JhGjbmdUk7zrDHs/nOQITVM8ZrmONFEDtVim
52H5d3rAXeZx/J/vWDE32qi0ddx4kDM+qyrW/9DPP0Oa80yatJrvTGFyQqPT6cfxnNoYqi8OhukX
Mv9jK+/HEOAI/HuyfMKYRCGDGBaoO3RzbYZSBuqIl0eYJogI0DUl6bAwrhf9QClATY6Q1J55Rdhb
5mgihKhzPQyP3vX3udhD1u3BUaUhfHXr8CYeze+QLnVd2Nq5FQFfHAZ/TN2GnSeKA1Ku9UxB+LSg
lzu+gsOMozwBj9RETdSiThFK0s7M2Q5bF2gZd7jn7//mDHHbTnRU7JgIolYisQ7ZGRafhyRFfVw7
Mpdz1WPChyU0c2a9spE+BN4WMWFkkyb9fG11OgJ5TTozWfwhVHIxbCGsfVnTp7XYPDuPekCUdGXc
l3p0SvljWOP7RNDf4vHPjq0QY+A19tn2SvIQO0QaZWCFMtQF4UkYAYAo5/SDntm4YK6Vgzhd/FCo
5uN9dqKcNSYT2adSfyeeKMtnj+3+vyHEe7PraR1rUp/Li3dAIZkFEPH2Sab2Ig/6GHkJY6iLB4cR
K3XI+JrPwoEMM5mnAQpIPHGRptCoJ2gaUcl5NCZlsXXBpnU+j7awf3/7jwNpVnrfp6wbfxGOXLdU
5uHPfmLYcZeCRJeN8ddZQ8rzVffCrDte09Lili0UqSQEt35Tmb3Jmugn17WL5aK5gqLeiZEgQQ9h
5jodvXXvCXL3/x2RsWvlWdrUWra88SnkJzP8Z2fSXJw2yq0lc3u26E1yQkqrSeSs6VMlHliNSkCv
Z+eyJl9koZvieeNjIjrKkqJjNYO/bHnt6p+WVSc9vAKln5s2miXWm1+yUcqAm3K8bJ/KzwhnBtcq
Lw0upnZ5CQCM4OCzU7Na0eKKHH9PRngrO2QEXsXQaKE9xfWOHK+TS1PyX75zyt2Os0YS7rFIdFuS
sL5RaNLAPb2jACBK+Xadu7TX96+PIiLTvq2Sa+up6ADrnXmMrt4DWIh/dcLzcaW8SG4XJ4R1pA12
OIrJACtTtpbuC24byhmBRXgkjY2ezKXT8C8xDV7JLIRSEhTPL8X5pz1FJSsLYTxHMyov58FNUa4Z
at3OND6vb+4B7Y97F752yiOjSJkmRUcqhzAU2O79w+9SgsoZsR7jkX4aNLcug840ErjaE+CEQYNN
HnZCsXYADLfxpgWZM1HknbvUxZWvvBwRLDl7zFXqrWwEoDEXUTMdrWI1A0tCsN8tD/GawYSIDhXE
HVcqWeSt8RK1isLeChj9aLbRp8Zi3ks0t/QBgA/XoWs9jOJVRDn1XUBk1M4U9geTuEgS450UZJNE
8fXWRo/HOoMtlMz8rQSK3Mq4Cz1W/v4GeuufQr16kgXALEhbgTyG9anEenzk8ioXbcfHjO+GpPqu
vFQy11cXEI4xj9RKz0IQNV2LQc6EVM0IuionEndZuVJ6ozNphFWk2fqAKakJzzxO8DhuuDJFfKa6
sm0yE/P4exdlVrOUA2vNDLPA1ti+26/tkb5ieqIzcn0kt+kjU2a2hFD0q+r0xmu2u4+qQx6TA8js
Armw1euXlHgFzjOpLpWaRmK6dbNX8NijcfxPaNeWC29KVlcjGeGRo/gehf8uLllXGFx6m5bJ6uIR
6sSyPh26iKwlT16fGZ+bpmC9cJRwRb5wV+7UGAliWp+D6xNBVXQSKkJKIxoflogxNCUTCYbTyq7M
uqnqXLTmKCRQUENPs6VyUN3rVU5sE+Dh4e6W43UCmg1UJ20UrgSRlOi70ZjNrzNDmRK7rVNjEKRQ
0187xWvukDKeaMzCYQs57KijYkYBuhC+0ZwwuZ7hsPzdipTf+1Y8LQ7lpswXLCaw5om1pDsu7uV2
NFE7lnIfybL04hECuy5nd270IM7go+cfqi2bdDb7ARqW5OU2V7rRH0OqtsegR2isOPEXP0RxRg48
2F9aMCYIwxEzXmwSlKJqwxtLte3MGvdJFCL8U2MRc547fwXBIvx5BH7bprYAuzsxJ3e3mZTgR4Su
q02WT2pQIy0L6S7qCQZUjbtZPyX6eE5yyXMxuhXyt4Q5n531kU5MIeVtHtKiZy76+dkEJZvuuCeW
NwUUsfffWMoxNfkfcTUVovWbHv34cYjCF6+wwRhprCOXiSuiQkwShngXOS4dfcoZ2MyjB2hDuh8c
xuqUCPF+e3gDMQhIFbhdo4YxioHxtusLwXBDT/b3mXMEvVFTDfvYlSje1qOEYhdOxmtt3sMlweES
x/53buU1484i0j0XxLWyPCmbcymeZ8SRUQ2kzaqhmKupUOT6e0YRji9iwcrgeF6RGM9OF4R6VZmg
yuOYZs8zBjtAvcUqcFoaA8A7e668dknQp/hk3czMCRMmNK6Clu7tAly7GUQkvPwlJKkE8rL846bQ
khdgaFn0YAl88BvFaTgDxSRhMXwRxm7Dz+F+CRdAYCzbvTdX0a0TFQxa1aZSArNCENeVPgupFUq3
1GAddkGK+nzHruv9T5JSMMI02D0/TRkdKKlyDR9+1VnYW6aglbpGeVUIbxNrhXj9wpfsbS5Pl/m4
PYV+clpSXoY/4ziaB+VPq3EDcWSbAp9AMIMNj+C+EN63mKUjnfxIW2+yJVNMsVzHNlu7/hKDHRst
HKtISGvlrqXfwWlDICclTu0zl7rj/KBs86VpI+vr/+70PhFN+asxxz2L8e5lN1ifHirxn3B2wKB2
bgHn6gTDbOm3ULbPpE9KYj8lSWR9wAOQzpgaqDF2BziqUiRZKf0AUCcjg4IBoHSN3vXA6zgamJ8G
6+QaISItRUUCQoyVh08n0faGcpnhoFL5lE9bRHRW0UgXIxzkvZU9gSdpGP2N3DeZvI63JJ/uSiNQ
7hcIKBEVjr1n6TDNOYZzSan19WkImwsDZC5NzKXy5ZLv+k9dhMxc4LaVr9vWNrmzD8iuzLsiPH1G
j0/atNtj1qRT5Jw1NvWb8Tn+iwVbaObADrvsXUSeHgAlGRNVKC+eeS2VS52ipvTOLfqBAN7LaC7c
5r/CGxeH3zEHP3lUvisQzlMWsWM+jCLikoMcgP2zQGS3UEbySxTYuYRqo3xD0xV/6uNUQA6TayfA
/voh7e1clJSi7Wpv9bN9EjjDW7g0Yfe58sNDkarduxUfXzfANLkxpiWWk6UTf69CwM0QjjBGpUtt
6yhWGiAsZEXl24XIVPMpo/PP/rZk7DAe2pj2y3TpASMuArr3xeVqaunHRC7rtWyRVvEFp8OLUrBY
vQTQg7wAyDlj0hCLge/YiM+zGAJR5ePNH03UYzb7O2bpRNGRECBr7sxzmxUyAEBpOZCT5ZUg8jTK
gvUW3UDllXrxTVoylVAmqyjiBUeb95NhkT+gUN0UGxkaYbI6kxPYw/0Bq2aQROGa7aEQBY/PLWeY
GEtUJ/yePUzQ1HMUPfW0O7v4bev1MF6PGEZgHeNV7IQk2j9l/qmfRXYFW3ySXLMmy82pnbR0oo5a
ejPn3YQk4eZVp1YIBi8jTDEoKjNuWt7MKi85U7vGciGD5+YoO1q7uEnSDGBmyoseH9PrZIT+ZIth
m4bEfsqunlCpV9CU62f9ohSXjGjdQ0gbEh3B7IxIrE3K6f1yv1BqjmB/WRBXs+NdnCpjtb58omU5
yrI5pCCxNKbhuri0N7ocUTBHo5x49U9ih2OkxQYAL89zyjnKveHSHto1L2oWGo2FTjKq2GUC89TG
CXpIbVStTMMSkISQZciq+Gaw0Vk4S77dnjbLslP3FwtQEj1Vny314S0D5Ql3ilxLGC2uD1WOe5dB
ITkbwbePcSBsgKHI6550FRvmrGQzw7rqXHdQumAcFNuWR66cvCWlts1gvKZCplzcS0LGSKNv9X0P
RqE4GyaCXRcII46SNu9OVfpfwQ1f+3IDat6j0TWa+5U74lkWzE3FfGEvSQq32C6gAXJKfJMQVkkw
oHwfjqUeZcsIsJeWyJwspzRDX3jkY4jCA5C47HcnE61XpsYdfvSx0JPpwEWaUGwvyaQomj/EK7lc
EvVFBkDpt7ur10thrjOic89xt8fKGlv0hojrQgf+ILZAVm6q7c7EAnudS0DEyKYZNzLbyqFfu57N
bAqNMhVr5pET4aXMUYYbuqKU/LxJSfNnW6DEHM1VV+ABZACGQPxbIh4oz7PKKA64m6Gt7edPCxGN
3TCjtYMCF1/stbcgqrA1pRvuF7c3zkiK62lmQDJWhCytIIMgiLB8RJcdFbZKz9lqE14KFOCPus4r
NIPpyQ4qqY1S29Nn/CGKKz0zwxgPAQuF4sPP1BdV98u5nUNxjlk9h2VjfGowi1l6F/sp76lfSCx1
4utf/cpApIsdZAdUvLY1SYZBWqjdWxMkD3gAJCJsvHIweyRUxCSVtGHgaGVG7pSq8UjlZI5d1QuH
ffojiNT5KO5wvsk1WmOaGTn5ao5gKdJmayIIYtID0V4TL0NIua9MC9kKC72my7RFcFO3htf9Lw00
jiLXjdi/0VWA/XM2VZ+WQayUcJXjIjb3H83n/Ar0PbQ5NOHPQBDIDIXXNUoReFxrU20V2PSW95hP
xNtlNSE/MK81VMRGEiJkXEKQx0koQRIOgNJ/E61tbj309FO9+dGg9NksZHSjHKxE/rHdhiYcW4Mn
fww1PNF6BETiNV1a0Ex/ajIB/E6VN+Z6CIDBIyq+31PBlRiJobKQ2EkLOdjXXvX6f+AnYaDhr0ve
aQEiGqlNuUVYRDKFjtUWHjVYxoFfL9Ri1abiQ3ciePKIAxvHruchwXU3/YuG/6xZQ6E8JLbDPPfw
HT1qvbVN5mPz5TvLF7S1s20OqYo8jglFuPCnZR4bMp2GQqz6dz6nX+E/g0Xec8n4KvLFxHDX7SNd
E34Cux6XENSprCCc65wjZJ7tsdGoHDdMZREpr1MoiwvC+4iveqZI5PAf/jqMb7LZjZqFuWMR2h87
dS81Uiy9tZvMDXJ2buyrSzt1nzn4+hCf4HmzmyCu+bGS35Hb92EPa2nFsQzABrE9QJkjsbjgZchr
e/T9sfEx2Jw0TzUKfykuQ0ioimJB0nluwVg5fn+5bb1oj/K+PjhxIM29tTPufSHYaeOJyaE3MnoE
4b5mfJO6jrJB6+hVDjYs/J7z5333yEECUSOpV+eVbfgVtQrDgiZT23r5F2ppA/nvVhEBAHR5BWcq
yexcsuHSJkPaI7ROC6IoC95YHnNEea/U605jALgyjVxnsQ08S0AvUKkN2hx68eEhFBKNZVffCBBA
se5FyDBehfKHpnmplcrJyPhvKQ8uklax2AHvo0FSsMAo6nO2g7ZLK8XqagTf/Wi3D8pQlr0gz168
ZnzYNBvMFzM5DfnPq08dqRExLnoPBufcZ1Kupwa1dHCHO2PmhtEnOvmnAXXlIYRYZ7SdNAz4dVkj
5zSVm1i4Kd8xyRoiLMEYKVHh1ehJBnA2yYYIb+DZXaAL0/9MWcOWWCpZyfyqN7hwO0lZhuoR2TOf
VW3Uby2V58puVg4pEzjOs8wxge/AVBd4L/Mx1VCRk18teIbwgCIHROVa+zGK7iS/vGCftxHoE0ro
UfYKRCvSf+U8I96P1dHsrM91DKj+ulL58C5UwxDbe75vGFc8wI3zNWIlYlxMS6UIe3Obgb8j9tKv
AWbGMjYhYpwBcHhkGVPBqmUAgqmxppHvCXsz7y4FVjnZreqIuqmULnDCFVBZnvnAwza25jTcKAsn
RZ87/vjxpoV+VpPWUVNgy7ABgoDiKQDDS28/VUxSux3FiJI6RSz0ul5dLNdqfh4G44c+x4ltjWeD
D4xxMbAbRTnYwiZdJc5qSSUwCxfC1vbiBokZRFAjnLjtZ0UnG7IuSp9rauE3NAmHqd8lltoRf9z4
76Zz+VkiwIN56ALme6PbUCOzJ55jOEjf/C6a+d0DzaYHX7YMnLdWyFbF8bKHI0PwDWDlBpFis2ZQ
kRS2RNVmltquUP/a2EckDSHttj88RJCu+M6/vbcw4JkzKXobHmTiG1xV4pd2SzPkbuunwedZdwMc
hCAoL/wCYQk4b3b8pKb/E5oKHhq+lrH1GYWeGJXv4nO3BFju/N2uDdniqHn0m/kJWMgcGM5mjuzM
XXGSxe8YxsfRGFBTeD1qrzHrzNTT/LWHSOzjm0eo8YPi5FyL82OaMcFI47HySENMCjtjvA1l+WCu
eb5Kycc5p9dZyJZt3zXGY2xzI84/lYEHkACB+CUFozjOKX6883HTzAi/w38oc12F7GWsf8yhmK0B
LrF5+JmAI+3yD1+tDcap3kmTSKifQaJvx3hVkZodLqiMMIG4PEdlbOhlb5jQ4UZ0YAkkKzq26Lov
pe8bIN/FW7quB5zxJp5aMTIU6WyV1HaNYRaOLNy3+f2tuGwkD0FMebXgOCti7CDeCvCAU/GUrBMo
8rodBQaSqFk7HPA9jTk8ftGLWwv3A67mUv8JNn2kbGLVvDiBtWL9ZGQsoXMsTiCaWSjCmelsuVoC
xhpQ76b/4jI8E783tJ5pPiYZDAA9YWLE/9tgRwZPqzPR6P9Lpy1q6IHWHX805hH4cixP/5tz0UL1
d762L/84HGGUHu/AaUTSQN2LY1GTnCU5aAL7blRx0mamFFKzdsZevIA79DoxSEr2KzPUtRSCsprH
SWA2Uj/+g5Didi3/WwtxiVKM8KYzUFVVZPD0NJSmBP5ALJC8VlL3hjqACoO/Ca828+d8z/DZpTfg
NOu+TWzOX7We/kWpA0OQ3llJy6Vrzjs/2PdYifB9srDBb7dV1557tCyS0XvKmkZNeQG+NdZyuJdd
YFxHStAoKs7UMq8muOKaFF71KPihiH4AAJibB3D6PXYa9JTY70P/1BwhKzbh1iG/bIzH0XdcH/Wv
3EBZd5IMfBVlkhGOSqtnVd+OO8bxCRjD9K5bSHCR5KsB2El4KSYCx2uS2UUORYNTaKN13PBKen57
iv50X7WXmCw0w6XVnN9/fTKIX3GeJg5+AE8zjgt8dU/k2mLZGJb+tfExzNV+8dVgZHg95A6oebjo
Je4KGfKZen6AzcePzbZgolJCMNMtSJTmGoZQ5aZPwFpaQtjFLKe9ZMoRRMix7vByPgDb9nlXSH2c
iqQoKexMOLf2KlsRAfDUUQ0+BnfPRMXUtz3ioVTLhdzR9xVzrf7tQPIkuF4mdp4DNgMcEPEknBod
6jyacni6b3v2HwSsU9Lcw3/x397lZMkViCfdnjus49AqBxvIHr0t7YALUwGjfRJXqMy6mNe8LieE
yjqupSc3Cu98aMGDmY4cHKKvfUsvvcIpUJ4nbWgCeWtlBRyE+JSgHIkoxvTg2nRDLezqvjZnm2Hk
A4THD/+ONHvQug9nksvyw7NkMRiElbVd0WXnZ/CiF1kKLkLcdIrUk4qGskpw5R+rpxx5K80js9wp
z920B9Z6PwEcChxC0+L1u1rL9OO7XOwQGNOle6fDXop2FWkkamn9WgN1cejbjBPeawPCjMOyT0lL
2AY5v5J2B5q+0Wax9OX++9Dl8ddmvOq12F4WfUdWawimxGwKKlE5iGZvk3GDKrIwKTDHeX71hsVp
DKQbJGNQ9KWbj4qJinnKvgnZO0o+T7mtrSe5eTLY92Ywzb6LzVccqUN2+qAvBDyg7E+oReWbdIIA
Ukj2e2zbfxJwYw3KSnxPPqcZIvTwPCdmE6A9zbZ6SF43t2MrQD/cPSsnTksEVtIOuEveZdlxTU+t
X8iGfnOpsfMLUp15FEiG+Hdw8hujR4kU46eBJeS3SsZEtSRyV39z4mJss3RktItCmQ4aw6HKx0VZ
Ce3XkdvfLtc20wApr+B6mVnaSAinQQ9BFTQN2Fn8bCwbQs2cg5ZlZvKssDMDasVjZUYXl3g2uEsZ
Ssi5GuF7TQW9Ctyp8xopdkivi/fOlkS4HQ2wq6hB7eFsyYe+3WrW8Rfi2789kOpVkQxAIExpdBrQ
Bohh4de+/6lAA1kd6iv4yED/GEuRPe6vvBKCRurRPWkD9Oo8GLHIq2ZdoXReXEZSThZZEPVKewWr
NMYmngF5WVvG13xLtIxukhrhdWAg0EtincSqfWxnufghoG91amYb95TzNPzpfraZ+5AijnphjjXw
GsTCtBDOiIhGJ22AI1x6xOEjyZ/8xu2rGfH51ULjiPX6ndS1NUk54uMIv2sLZeO+LVJ3NoP/wzIY
F/11jpcXCc9EBlxnzQUepc5+1Ggao2NSVasbii4c0irJqTgCfEZ02oYKvveM9ZB17x7Y6hS4GwmM
IEu4AXkyfG9yFyn1XNx/WVtKw8TN+Dme5ICIsRm8OdAH7lDKhI+Ekbujusg7Haf5AjoY87KqGolr
MHJX/xPe8tZV8AuSnjCu9m7B4OgI1zrodIVZE87aZ5YDhiCI/hwMbKA7ZRRWFZibGJE0tL1/K+01
A+xO4OCLPJk33loME0RkIur17qmjxbdh7+RFQ/2YNhCAKBVqYvGJ4IXCMy1pMiGVMiJsXz8gv8Zn
khVm4QlbJQNhMYguVyNYe6lrd2ZplWmXzLI1xYqUnhmw4rnalILE1pEDaZF0tawNUvNDZtw2XBVa
AVw5NnNGeXHVrhiMY2OxzCx/EcZ+53YLE46NyC71wNltCy8sWvNifwkcO0DQzENO/GaTgK91L8LC
dB4kSbDa6NOXfN6o28gb7JoChLnZ9PoMXP7DW8P0ub50Z9uBmG7ITvXt8nutdwjfWixnGp9uapmS
N4IPFqzZrtyGLPNeWvyWhO4Newdtwrtv9QggTbCk6TTWgIOYs13OnKmxZfx7SO5yjTwFzwRyVfvc
E9rQN5GuFJ/g3tnMSiiipM88WqHkp3Jgkb+02Lagr7vsIvvfwv/XZ1kjYd0jAEel8jtHQZXInIMH
Psa+gNUjmFDmAlUltvyT90wILKEThXFLEiOLE1+9pvS+Ho6NVFYBHbpKtZHG9lyTE7aPmlhFr4Pf
Rtn6AIxCISiQf0dFjrpB5Is2qkffaSPPGuAy+iNbLPyoDo5SBotf6micSdNxYZAVshBIUeSEKWRj
1eIr0p8+d2e9O6wyJOhz3kTObWefP2t1VG6Uh8jMa765mQxDuWwcvRKWpptSYYqU5Rvn2khUjwq+
A7V3JRr9SoFH/xXYlW0fMYqmDRsRzdwUI3UEnYjoHqDDcMu/hXsDiRQxFzrzzonwlt8d/Xc1MXi/
vWHvE3j7GPdS7iiswpSJqbMZ/DDUbtECONRXUqIlwBVRcvvdFs4JOla4JHhqy9tXoHKztp04zuA8
YChjWO8UMXWsKzq2j3dqR8IQcVOvxVEIDdiWTcj9QwpSyCmTIqd3dxS1GlOiGHgVmb7jN9+n94qu
a5BbZSoR5X/nHBq6nLgNl1b9fIt3etQgtmDWmmN8gKespECjU1FKYpvWegtR+xTH5VncBJCj7DC2
qhqj9pqK/Dm5aUXnfeLIL3Rr+fzYu8FFG1NF+iylfkffU1EVAB9fYkiBvXSGqoutcTsoQ1VPSCer
RDmARNKRw/ZtJo+01KztaNoII1ChmkXueR05K+meTz0H3CNqTSf5nvtL1keUb4v7hvQwsYwJQcAw
nP5wdTFEwWlUrGyYkO9LVGhiLekx+yv65xmkmJiwS/pyEBh/6Y2kG/LHV+nucja3KWs3LM6A+jCV
uUIg2/cJYnREVkq0Zw8d0tFIe0qxVPmnypQQlu1UVzwEp0512r8UBNoLYf3FLt3jd97F0EFgEPCk
PP7JmuUH0neoQomRtkPS8mpDFw4S7Ui3B3GoVYXSUUL9Ywsub1MR6cf8qz46LFNZVDNbV2XcydjC
FT9RxrOp7Ls5YG9mpfLOY4N6y06EZATTFzUhCadweESf02sHij9glgRB733nZAhZgOcyE4VBzyUm
YWuQnVejZaaon1QUZmbwuAhVa/uZPmKjlHTL0IPPiQSnz2mbvPq5iXemNrMjSFMRi0+ELZ4YT4PP
LLHxP1Fni1DvZT3TRZJhOB91Ks1l3kr8FYS77KfTTwN15t4z2vj1YJ+jHpGxSM+0Wl4DUsAZBusH
zfBBUqfXxJt4wbPnOXb5YfIpnv9C7rWZiLI0ip+N05GPSeI1jNax+5XEDMJpr6mv5kOOUSwjXrrg
4xR88Q0wUsRVjRFj7cjcic090L5Vr8OWmcn2srAnAmspelaKVJUIXwLta8wqev/5Hm9z6rnIvd34
r+GsYBLVJnlhwwHOEUWwhYvAYKxoGMkri10r37R9voYxp2G9+/hQop2gQSpG60VC6QIx0BGIoQMV
mPTnonc+rdmeXdymrm4fLRNNgP1k59MM/GEPvl9gO8y7XosJiuRXq9K75KR38dQ9N252VGIrvSk1
gt0yLf/VoYfamSOEZNp2eCb/Ph7jO7tgJ26q9AA/fRrw9LRKsXkBoB4lz86t5fcL1LA5+G35Am6M
b0i+DMzfk1709ie22rSKGH6ABV8ayhpUrSjMo6rELXV6Wlh4SIlZs5i6itv3IYwgnYDQsV1uBaFD
RHApFX9FZo2KfgJJZDkqDNmP44nJzsfED9n0jcCIfyydosOxMmOF5RcvGNNP/wHPIxhRbCKw0YVE
QANUTfPwynmr4ySVDDVXyDwjLWCiibrpw9Ty7vxMQNFjgJVtjh7rBOm61vvNJ0Mr++XMU/9UFsBs
dqEWZHISJJRQIMLKIYLWnQgaE/fwoJ4IM5S6OJ9vL474k+mVJ/hGK79SV0to8bgBOyDsYJJCvtaQ
AtmCFtiA2DjK/eVaUsTkUuxKJblx/6EKFy0wK7rYxOcCunu1MbVBQ5S80osrk/zSxN5j8mjiyZuo
53kLTPsRiVSJOOv0lDPztJFBtanXvpk8QDtf60FWrtCIMi/bXUjcseYp5YR3BPNi9SOnSiTYtrDh
Fdp8s9NVVOBZsp/kx3MCNwFhWT8/ARCE3OE9o1poNoE8Ye/+IRdOnwA7vkmSSfJf9fTpLeiIRUk7
ZmLdreV5FQMP5vTMTmHaLtRP5Sq24Rz1Z4l3s2lPafB4M6JkscJ+683hpoRV+9OLmgSt9R6BVliZ
ftCCEJmixCd2tzX0A7CL4XCw6h1WH3s8MW7yrn2PbAOnjz5/dimWC3msvYju+bHPjVkErSo6u3u1
YF7iIUuofp9FmCJmlYmGsPgtVE6+DlsqGlWFqUjsNSFBv37H8NDyQHOyCYzTwVbzAxWvW0IMhcl+
wrQluTFBoKARG/4tamhagWYRxnpbzZqSGgSDsRvvo+xrRoxjxdx+XsYZ3h3GBBhge8u4h/XExFos
ZoutTaXb+dDcd+oJ5waQlss1tdGQ5dSqRDgJex+430vXNqbKB61xU7BT5Nag866jYJtWPgx6wl34
HPK8uVbU/kVomq8vdaIC47jhANKavJDOrKtxXaMbZUoxeuYqdvM1juCd2kzENazKPn2nczMq8dEN
EeFseCeZb45glHbQMprXXx+b5IH63HRtM+oruhRpnBda+6n0pofyjDHHQNRnYqzvSkBCktTkgx8i
HDT8U5fZqqdxClp+xobdxaGCBKEu8JFh2NNQZ6G5EdwH1lqcElT2j4z/QrP+gbxemgc9yZmd/DDs
Kk7Ey6ol8h4pQjjVA984nltyV7wsukJ1AENYuyDiibIPHcqp0ijYpio0kG0WLHWArew/WVNtpVQD
YkhWxVs6eDEDwpG8wCAf5kDcOhQOaoqfExDe1SyrBY8Tbi/dchYT2GtxEa3eYaeas1BugssPu2IN
e/Bk0flLnR9xs0mI1d4ommL0CjtfYMyp9KYh+WyB5o/WQ2WwnE51S1SFyvWy6SQeqFjTUBofI5cd
h2i0jN71iofX3uFPyp6hwMsNPOBREFB4/eej9Bk4yUghksx6RB2RILyd+akfB1ufZMkFkNsB73KK
7cTTfg3IKXFDYSJZpjHgWa+A6Kfq0NYXoeVB9gPPkOBqclqorNSr9ZlUFDVPH97CnBx5rcb/Zr2B
4aUOOEsETOun1AKe8nrX4A2GVsSHcLpL192AyBRzajDvO3hn8SiUIclgkCwNzKrBax9BOai4KsN6
pyQFWpni24aRvv9QkB+JB0DlZuY7Fn2wjw2PT9MBD0S4c4Ue90yQxMhEcdTIHVDyxwPvYeBtELEe
wHP+VRxmvB1HcpDz2x5kud1t5NisIVNthwsWbpM+kdT5V9JMqtqhL7fk2OqjnQTxhnANx7viNGZG
qPq2RuENPI3MCPZ9lGaeUE9QME+lKxD8zX3GtP1BjqyLCDxdyCqBlv+7offQcya+YdjRhxuGwjj4
k0piyDh1o2DE24Qrk2q/JZ8gz1s7wKrSsm/QYv7BelA+YK8c5M4r3+qsVi8EWm0zyICdJyaHYm1O
Dh9ANCTugxZQ/giIelydsO1Nz3tkNbUm6v2u8x3fNOlePiYPAYId0i0epZQF1S/UpwJfbdfTP6j1
3UTv/TRb6YFb2k/oYa/VcEp7t2YdAUPYbMusJjhF4SxbBWIM4TdiE4N0Tm8w+Q0HPbVkfI2178HX
XY2spBZynGdHIAn0IIfzwyHjk+znV7hZ3fSjMH4TgWIFrrDPRW0vUfTEgqoTvZCOGEuqVY/P2Q+E
zspIuaN7Fx41IwyEvZINvKo43kScrF4h0980+MwyLFn7WJWfrwwil1eBJkTQ1nA5JV2bhMZoJTuJ
MjetaAGPr99nmcDvZvJHSedq1LM3EoSRCnrKas5GXIrZD71nCc15n0Xz/qoZuFqNgsNmP9+aLRn+
eR3fRnA1lw7nokgU67xxHxWDSV1PyhyCenrOg06K2X06qQL4lmaPOkIHTGf0lVU4eGGzG45J/Id3
oMk/4ZC01jSQ4toBLxmMGcsWSow2i5zEqsHfU8IB68uCQMRha1fB263//rraG1G+eLQbnDGB0LOv
FdEXjnECn1u/9qyaudCDPoabgomkkkSD3XhvQLESal/ba7hyYz4Am9oKC9nWp/7NkosFon80BnTw
sC2hvmp/DpbFH+3PId/2NdH3cNKDfk9Dg/uB7cZHcoJzCV0f34fFjinNmn7x8QudPuT+vTt85Q4I
gPs+D1QgMB6cEXT932Lp3g853f66zwp6vjeMjOrhQ6zCHnsTo7uZoy/yGePOmLFvx+Vo6JvabAnJ
pocdsG76/V/kCpW/SY+v3Kmz+2Zr28pj2x5ciot4v6hPsWw9t17Z0Ko3CIL0fhoVM2+adp7ADHma
d5M77P8qQ8w4Wov3Qy8fzu0RC0VzFwJM4vjWdz3SEYq3EfYzxtPivFBHb9Uqu4fQP+9g3A4Xo4VO
66aGuxQsFGaUeZ1gwNloyRbTHz66UTtVKvV4Xds42+H6Z4CqER7s01slGFKOlJC7xkXb9mhQ7/+E
YXIhV9hiS64Pi5xTsprKnM5D+c9J2ZrfHTEkBZvgUX5yWlTcHZ4QlG6xTFtnCZ+Z5aJBwH+KQq0f
YD8t2kWLy5U/2L5tSNKXs9TkIMxxl4AYxiIVyhuTxCztvSDMPNsHtJ/VA9vgPEsOdx1VOe6y5wdm
zzTV+e/WzmTzHOP7pkxNqX0u3uJPKR08wnSxXOgVhV2U/w8yK/7lzPybPkHOawHwJ/C3RQudcs0G
FRyGDoR9RCfnKQDqEYOrUMbWGNWGPigVbw2b9wPe67bgVdFuLnIgXwLCp0ic605joXfj5eugI4XL
/K7CyXm1VLgHu174vWQ2sA4XNw1kaB5C7rc8+zGnWWOGYeWHn0k9dsWdwNmOq5ODy1UTaDVuzpaG
p8MKTrpQV0nRaMg2GXf3QQ6gBqUjn66Hkx2XjVbjmVxfijoft74Xp31vBr2Z0ZdI86c4GwYZCTKd
hUX3TUdsev7UVoofYBa2/viFaM2BjYEIqoYn4PY2KpSNWEQIrosoQu1HWlN9qAbuI3jKQuEedy+f
on59yIaAqy9rPKGnXTwShjv6WMwYzH0M4kYlaJUDemrvG09ZtZGK8yjCsWE+zWxfgHXtYgpv2H8Z
dB6vOudRzJyWt2LDwkXHbs9qn3R2IfetK9Y/HHYCFcXXhhMtTuau3JpX8KjgHouYIOAoXyGMdpvH
VQ1bM/ab2V23vxkekdKmuktQQ0N0sNVT3H0nRKehZuHasPEMyBKi7ezu3/X6fnXmqv43uHhIrkW3
Z+hGu7f5azxS4FWU7WJt4kNtMqQOsReO9I0uB+5wa16EkIUCzD3Jj2Rcr0MKlyIe8H85XarfzRMv
CJ2kWjHRDToip1O68lYHJO7mPCqj+7I5v+hK+WgoOtAAIALWMMP0OEGgsGrzDYLWdWl7FQxdXI2D
83yWuSVfk7g0YiCMk4/afD5be6A2CL+ztEsiD3z0cOi2mgYDwv1+F72UfaQ8SDgsqEJAF+gLvtzM
YbgW+IUftlRugqJc+ZDWd3jbczkL8e9KcHhD1FBoj6DLkjk04jdLPUEm5Ks/xvi4ElqVjCpFuC0h
6yIYpDLZqBOzHErZJO9v8iSEy+41ob3mQJBYlxiN1rji3+OgyJtbkkNFgfB0RT5glL2fdQltPzfZ
C9oZzc8k2MUM6yYFx48W1F2k/HEXPrNfxz1YmD0ctPsWayjd83nXkhyuyBk2UGOTXlDGG5Bmd4Wp
1wr5g3z0Ikhwto30Y/kojvq6X3WHCI1ChvD6H965Y8FO3CUruGW5J/YYDfv27GZ/lsl6JdA0MEF/
ZJVZ38J/V6L94VgzvNrrMVfVZQzvN2c+9rlpEnDMMi9mswaBJqfRQ8bW4ECDZL1gFdxpzWomRQnT
7OQ+bops2Q2AoF95wR7PuHwDA/gDIM8GWF3luJY2sn6euyq3svJrzTOl13V025Bw8pF/1VtbqFup
fLIFZPrbar7xWVbW+zZH68KNaziYfERZWZC+Z2uYUO14rng/IGDv7sn60BizfpWM/7OaBIdIbhpK
wOkGzy2fZW44nmtNMFIQE+V4+qODpKoIPWYF4V7CIMYNRotPcuqIiyOkVcpztzxSHcNRhZCv2NQ6
WoNuH9Af+agr3iLjeJi7gTSX55o2QllfQVInvv2NFNB0pyJWBANWnPyCP1d0Hu9u/WA5o8Hqx4bq
9Wb755/L0droXQVM3NgWAiwnWjdkYbDj40jLEWdcJWk+zlVnum7YrHV2UbZQ+decR2zF5RMStAeZ
JEcsEdislawJflGuN1Vk+yx7+//I+QYEsN0MN7K7ZTtZCAiQ2u83Z0ODm033rNscYLp2T2nJMT2C
Blby+xh2pWlov42yo29tSjEzGVsnO9DuzvIxnQaKAYjivV94TudeP8O8de3EUJ80aAn8W0d2BvmR
6F7yJeaYpMA7h1oezHYyhZyxklM9A5OUKWEqyCwDmlCN/z5nv1nXkJe3vtb2AQV9yLZTwVBMP2XN
oQL9f65hwgE7DGS4/etv0SP8wvLcBo1Op0KpHXR9C+dGKEyXqk6A6YK7IoYaEslE7tMwjYsTR9L7
NYfWy5S5SG4NJaAaOJvv2Q3vHHoNkRwEDZ8pbJla8XpEa1wtndJvnaqidL+g72yWkLug9UOeZPMF
jBufihYlLydrYtufOaHnW0uKTgDnxqUs0xCDoOEsbmHdQrbOIGR/4hW3HC9nNKw2nV1Buzl7wGGP
alxTqxzAw01PL9SkIBNjmI3qqr05Th4rFVosNhk9gOE5kowAbBjcPpr6Z7C0HetQpFrhcg6Mpiyz
kAnZwZtY0CpDOGe+dTgTq6Rm3fQSjWizsIbHnvxrOT1dKBbDcsZGWtOBMvYgg29W8+4TUwsufIHP
CUaswn08iOLq1BifvktNmjJCxfgTqPpIyyBXpKcnjeI5PdqIrZtX5CDQ9wJdYShppN9QaGOXESZc
9yrczlOvP62zVqIMeahXUvsDkaK6mjDb0C8fc53hIcos2s37bO8z0K8GjhJNN6JfNwejDD3rJ9e4
KNCtlfWgfrbp+xl8fBnCMqO+DgEOZ9YqFm6nmqoc6XLyoTw+6YeqaEh+kg7zgxevPyxdzWE6P+oT
kB3aiJ9MhJoOxlHw+mBdGSgw15PcKldSsRoWeosyxbGgiDSSc3YOR/G+4jFEgQXU8C0Af2Ae/+Wa
W6ulci9TL2vGp9QMwpAlrsfLDV1kMcYM34GwuNDgaF0BRevFVH861Z3LApp5uvgdJvYnhiTr124i
3Po2WHluzcS7WXnRw70Rces1UFTDAisUzMsX6EgER3iAbJs5XmpUdsZoFIz8+u1KCotYWVaTV+PC
8yTdcNpwMX75tPn8vMylQt/P9b0uFr1Hc9iXI9epT2wzUxrTJPLMLjM2eojUg9kg5yJB5AXB/A/9
oKyP32gnSSYMP7+jUmYtOleI9ckDtn1+mEFPeU16CefqAuT/KThdeT+hBwNKGlSI3Y8YdjhGpw8n
cXrRTzO/cBtmEkTgZ/UyJKKAzQwtsy6gmzqg4dN/QwC+JyHE8cBQEKcqBq7IFqdcDqXB8lzv6nfG
LZ0aGj9Qeon59MjOnTCXLi0GSss0PllgUdPnfDPs4aGq85Oy8wkT7sdMmIwOKKH/M0KgiDuZ2WwO
gyTyMxzxkQyBEJWopoiFuIB/Zx5To1bi5zmWG8cGOON+bVJx11JJQNzHzesucUUjnXnBiZQ1EAWE
TYhmoxLLX/ItofmgG33FLbOmN/F5TLcvQJ60anhbEbN8qDBO9TUkbxv1gkgT7hLSj7oYr4Ki3aCJ
SxC51THqmii8lYMGPVj1MHxC/xKLtLY/rTcnd7SZT/rNf7wB2vY+zGV98McQHB6pu9s2vXYCEZU/
ZpTu0xtmrULOzpvzp2tNGGfnwGU1BPimbSSr4TmVgrmJer144lWudb0GmkosCpR03GbfgPOavbWO
RHu6d9TAjEmjWlQKOr3NA8S3PrDrlwhlpobwnHeOdc3uYeP6bk0cUHk8epnvawNOAMo182IOfBgM
mPXrHUCP9NG99Q2IO6vjpdw9M2VSJp5BruV6UWK/b6dGdVbzuONGGeS1dy+1goqHJnkOVz/2VOL+
aaR8yEJjAbpLaFtQLc8IHqWhdu7cIHHs4LARs9bjmOaR55Y1m2ZstcCGqf5c68/Mb6MmMVMybgjP
k2waaJend2NJa3qxeOjVy5rkDkLWevISokOcchkN3XPJ4TkPk4Ou0QJMLEQky51zyG1FLpDofUfF
xpj/6NxqWDQTFmEZgsm/RfSOQAj4rG7c3DrRNH7pUushqhk3y3YR4lnk6pCq7OmeHLMrIgmvpYCB
ivpOO3zAdsBZkpDXzpY8VEZTWy8QsmlBerYDY3/z2ICQYnxJiU5F4F0qvJxespPp/mE4yyP6wgQ9
vNF0FyHknWuy6plRFg/Km6kQFNWfOmPm3Ni6f9wvFAL7CPk87mPXQgjGXpisFMBNOLnMFD7Xu4IN
cif3mI67W9OMbHJC7qfPA6D/RiqGiUbmQ+KYs5RARykJNB7toK3RpD7bNjas4ULAy468GYvDxhJd
gP5ug9q8FdmlGUNgl8hTvnwYPbVZgMEd2LfcPdqSaedINwG4IPdhHvjp2Ej3jb6NyOyaHq9ZrD9v
b/D2J75GbVvacSlBb9rtdmlxoHNYQKMBpErbtT5RHNHld9u01XCDo8cs4wrdMq0bahPDjc2dSiCn
S8PzP9Q4brca3tPA/HlheTyL6CfyO0uubU10ZydFjMc6ZzIp4LusJhAbaXnxVA/0lZVuYHxiJy+s
vogmxzHlgWa008IoJgalZH95iBlTiYylDYvWQ/PworIArsrubHdreJtvW275O3AFtnKG7Xgl3c0f
Gcs0nzd/SYT/2+LGpfvPn5vGOJh7+VYIl65fEPafOXisrdAM1L3LkFqH1Tzd+6yOpWNorcOC4zNN
qjRJKMJGN8czk8ECoqrEwmgpLZMWGCouJgcyMAB4jXxZkvaGW/7i41xAygDUjYPDYxF24Vud7nPy
Yj3fiJ36ZUdedHcpYVSU1B6B0wAD8S0eLgBafCr3jpecu82uBvm5NtY09WTvGpFmPLGroDTYASyR
Few+7On/5y8gGkb61rl2vgLHWXSME+SDMMgBbx7f/3TqBdVYjiMIy+rX0We3rt6tw4xzHFhMnbel
6aRiVRsdAElOEk5kmdjpUue8etOJOfJCXmPWrpOgwEprXNsDPcfcIZKb9nlwQoDUt159KdVkPT44
bngJBax+CGQqEdFlio31IBuV43bokgKfn4ZtgbOIBrpOzD/opQd5xg8OnQKZcZdSl28KIGFWsg4X
nSZ/+aaLsXn3J3eZcWoxz4sDJUxFarwt7ozyS7rOcy8EH2GiWuv00b+CsITy8IVmkEpXauZHvJ+b
Tr54NhRjoafAw0y6BV0Pm5KBZEjACVj0dzTsbOgE60jjufu0e0G7YqeRRxH271eqFFfvYbe/JQbw
h3jN69f2n/YEYvxR+lm/vuZGbtw2/EYoGQIFiAJcOuhFlGzw+8+406XvnDB+EQDKFoitJLdeyLLD
2e8Y3h9q85qin5JSFDwWebRD9tFh/r/RQosPIhnDEnU6+MmKl6o3jZH5zZ5a37jiWG2ZcPpaHAtA
FMd79vNMmeY0bi7Q0llxeLF8s/mMCMTToLQ+5VgNwmNraJgEc5ORdhC5AMJEwfO5fzEQxAlOIS7T
Lfn88f/BpRwyhLRbDHY3j78NTsnB/TrnIkmpRlmSirBcDSSIpPLID2STL5iOXYV5Id7GMUw4cw5i
g55BD5MR+yzM7CYj6dWd5Z3It501M9kMBZHE3k4CxY946gfkW79zbYeEnW8yj+m7eLOls2J5IZK+
f1kPiaRBSkE74wNcdpbUtQDTnY3y3Zm40U1xevetgUi0ef1fPAwaVcxILpFu3fYXL9445al32J43
rKuQMsKbGRfzTDuKM5Pi0HKF7bCu9fxS0gKd78Ov81K6itRu9JkyXh+D+0RUUN00YdXB0VMFCNNS
BZ8IzldxpBd6QOlecwY/INflCusfnozzkQ2hd4AKhAmYrtWrEEssFa5nmNCiUMcFQn2kCOFSNFLT
7HES30WX+wfcOr2nFrenfssETsoVGYoNmDAv8Bmrhji3iLhbRQEi3ZlfUQTxU0nvyjAyZV9W9ntX
CEyZPNEFB7ONA4ZUNY7L2oUGy51Po2ZmtUpqDTX33uJ0NeuxhmCdUN53/CB8eNNLJeynBovvCiw7
vBBif3J343v5oz2OF9CSspreWfi1knKF3UJAgWkZYqKEHasDhlO+7hI/1MQ2h4eQRVOGATHD3rNS
VNOWGppGjpDLutp7HHQVECCsMFPeqOJgS7u9JrU9Vwbz4+2bRtmCctJOStgAQAgc1X71t0nldOyP
DK6g63PkHXwsyLdyc5+JA8johvhqVxTezLD5DdVcyI0Y+EeTaQGYw2a/qfDkP5Kr7PbdDSOaK2qE
G5eQBYFL450TZVZN/CXuRgwTsycbvXAdYVzkP0KifvFcZrx7e59CXRlJi9mx8J/FHPDHEllXf9jH
QVuRxYawd/y3k2KEH/nRyWms/oVeeTeDsMz7U5h0fV+rzsWtDLEmBoV4Puv2mk0eRb94LflGqQx6
QsRNPTha63UzNtdDVhnTcaji5sPvauf1AyL3z+jCVedfC/vbq1yJu5AIEV/azYo5GzNy5k31m5At
NIPxmw8p1vteAiedB6LsEuKTfDBk4OpSWZn7E7ZnRJxrHYb05bWL6dl0QCE0sgjPlVGjuit1QM6P
b9Lvqt/er3P5mEeypvBcsW7fZhcAdFc6HiV00MPSG7A8FLNQc/kG47eovIJAldbUviGHO6x328EV
moVSuUb6P7Aw5M8PGXMQKn8FjlDIFG1NtqRKoigQ0/ZlHs7o/MJ6QEphuTR5GVYukRbdouZ/duy5
ikn0tDrG1wO1uBofFn+EkMZsA91fNr8RVb/vfLneQgy3llktwtoQvT30V3BwAOaT6D0RIu5bZn4v
1KF+Gs1xRqXqUEO3CyPkO3EVzWdtgXIeulxCTRMzdCDwcYN9q/sG+upNxm/HFMbGLjXdG0kc1FJU
0JrXbGbmyL/UnunL7/mn0HqfNoU5I8R+vj5sYtY1cQ/kN3LDRG0mZMdl3CZiFAMVJDNcbxxqQXjX
dVoRh+U4pG8TB0RR8mlf9JcuvwY5az4tMXHXZnXMiLSRJIInRZP3nDLIqEXhke/smzsmq/e5+QcZ
7ohfA9v1ZaBjlWOnv864+/K20V7CA6SHritKK3qxW5PS9cuolk2Fl/UMLPlHgWHSRyOgAgA6+MjU
Z0p3k2HtgaDQFlUBxdwVV/55r6c8uZl5R9IFPkcGOvCBGvVdALjrBk/m1AGgf/YwTcTyjQtTToqj
/SILLu9ywA3IRCY0FbaF4ZZii4dMhGTGhZTg/43v0q3S8BvbtkUMavRBWosiNJL/oyFmEuzpN7QN
sKb826z0lw9ZwcCju7fyNjdr8fXppDe11XC8vqOlTtIA+kGih64ZxSsYsIDMxGqZY+GmWDb2jAPt
Nt1i8JCruH1ijNsLKToJJpQ7/Bv8JhuGtKaDyLXK4lxDicHCl4oP4bSemsy3D3DbIpwk7ySyn6Fb
kIoMR1BoqOkAODZ1kTqM+5vfUpvPgArVI9rhNpEBKf0yxNHev/qqnyHSAYBzZTqAxTk2P2KP1tix
dJUZmTPLtNJOoG7oogZ96YWBZhmVVQfZ5XfuAG2BYrOU7B9KPpitz9IBWCBd9PVi8y9Y8fkYe2Rf
x5vQkxxuDWXlZnSO/THDHb1LApiMw9Uz+h27cGWVj1iCubFnP1QARBiem9XBDw8oR79KlgspCNnh
5kgHzjM9TEYc4p7dnF/elIduopj60K9zSXLlH/kvYR2pa8+MJ7Dm2MfHDSiryMcGU3pDluVCutzv
MnEkmH8ig7SJQaqgd31lkpP8u3aUcyUa7V744r5FtUXJB4wLu/MhHDUHBtza4wX5q2o4PMk2Hzbx
fY4TF9GTQeR0S31PfdLzus0r9Sv5l8HixOALmpecVHSEfkpW9lbo9NxeuRE9w8KgjMnrlakN5q2K
vb98v7Uy5CG/SXiAIc4gjxzLVygjByZS6PKk9a8YAr6xnNtHR183naZ9mhR8LYVhXOF4Wvd/2+JV
JPuzYMxbsb5gf2IWb7WzTXx05lr9CubD6h/FDeOWqzLTEhAIFQadtMZW304LhqqAcofVO51Um66D
7vCJdUahxBAIgzzP6VEwWFYNLLqKz/1adyDDcJZ9tOCmlMrI+hYHBNwk9K2PD8EZnHAODOfFWRls
Ik7AvksUgD5uIr4ohKeuNChRNEya5AbYD9r+ChCawfDFGUfMT6gki5RiJcviVr+iRKnnbiPoxqg2
z8gVi8ZI8YfqQsilaVNC2ZU8/G8Bagt2ubjHuj3TFfNqRk/2JJZzJPfOAWve+Btc1JfzUaU1KMAu
MDmyGeeZYt7e1Y6T2cJ8cfh50FEd2oqvxzaspo8b2Ld7a9Lny832h3ggjTusELIs2SF8WggPUTu/
sAX5+xkCf7d8Y3AKNKgNxInj/NM399Wbn9FNb5MgBfVUDBWhZkY4XsnDVuhr1daCKTyT34c5E0XQ
qm8+GpY7UMI1im7d6RY0kmDqyJw68Fzh3x6e88CvDw8dupkHXd6zoKgEQA6oHLM4VDBHRXgovzDt
/aK7PI2zTlMxOxzur8nyM1ayYKb54+E3ZWGFczoFAkZWweqp6R+FafK4TeLg5hGmrjDcMaxZ9/5K
5Or8DplBGMTuc4Ay2O14FUCOT5BtsjcPHeEvfMdARJz5BpvzSc/QDFFPQy4+gTFhpK8DQnrHUVsP
dlyCDBqIAhbhCSwbwE9u45NXjn1gjIzEKT9UXJMV3uZgHU+pKr4122JUVQsIYWL4t6NlzOwRe7ii
5bubvikEAkyIp28qaqcxxtse/khW7V6lTZLaxTOGlstfq4GpC+KC2dMtnOByDmtUc71EGQHlLfAi
ZQOP4U/MD2GA/zTHYAFXXSxtBD2JAP6wHm5Oo4HOmMLpXMSNpdyk/u1i4fEtrRiLfsp65w8BVRwM
vjRandvDGKfKuEbM+QSXvL/NhM6tj4IR9NASbM6QQkaK0/kLqn74teg2vHYUQearKFAd5hefHEd3
STxoQFFqoRAwWnL4yuVyFjxSl2brUEh55mxbC6aYKda9gRB0yd2IOfniLJO/gK2UyUOlCHZtBChu
KKNsN2unuALUw7kNPtcvsFBXNpMvSJK8UiMuZ/WqpkPKSuvMHSHA/X/7T9EXqDiKE7lv4DWa9c2c
xQr+Yy0J2GXmf2ml1/HfteEA8AQWl7x/dXDC/44TXUsDU7jfdeIKgl90v4FYRugQWcgHR282IrzE
hYH4W67NGngh5TeB9QNtBxttIGwvrh8txR2UeehwIUrLfkAKZI5eOycwpfHIkmUDeLAapzkV7ikr
JpK1+HIJH39mlTlu/5pE/q+QocWg+EAXUqkVtr08Qr9QRePV/klH4/B+aitrAzhauvxOJbHsk66x
m0Yvbwf1M6xsfmU7eYiF1jCvdy1EYFrwsbpnyyHnoen5YebSEyw/YHy8ao6E3H8mFKsX4WI3ckGi
CMvIW9Och228tJAH31H3KAuWffjVzYj3UZbWn0BFZDmFv1Mw2Hy9xrhza/o06zY2Z7GGu/Gzl+MW
z/b2f4quiCEMTzIuzoaKXN7S8pGhWJFas9FQxx26bApF1g8CBi2/Z08hk3N7d6WILkf0QqlTRGZF
Nvsv6peh7MjlnWfEqxMGCR0dPx6zCxTdI9xwaWWg+y39LwAuq3yf0BY5zUxPHcdndPVbmOJj72bq
muuY02FW7TOsCFQBJx8rXRcgM0ZPmTjlqMFhb7rqizzmFIFZkbxrYJZal241LbmWh1xhHS8CnZZT
XGVWJM9gY4rvsX1zAttfaC1If1pOupqdSkNvvWs/5zFG9jAOhVztcqTrfbxyF0nd91Xb/eSeX7bn
XcXIB2Kzs0589N9AtG+kHpNP3a4csoDyC63N3EdH21IJeAdJFHGOVT/kTk94EZ3xfhGkqUQuvHWT
EkeYaPRQ62yiRE8MN6L6zWO4KltemTgDxgxOQb2Wv/JPkiRCQ5bzakg59NP8bSXL3qumB20GgxCd
G/G6LbJh5sZFYBFDlutxPjzmg4ZEzARyV0UKcniv5NWPc7od57aI7Ydkw+FzWIWiOBDdP6h4Vtk6
3vQ/j551HBwvQG1Cl3B+uI53nyUjIR9v/F+2bf+kCRDN3UkntnsQCAQEJZ79P7MxpYcA8OExofQO
UDR725Sk/WmOjmMVSL986C3+KsGqwoK0XSjVzNlXUI/mFSYy7jdiaoemcJTT+0oquOgimiwfuQgo
SOq3wJqGY4z3ahF9+6qb0Phrr7DvvMnThPHYALSQVgWxGV37QlJnK+otpFrDHZ132LDO912jJ2VU
T0HgL7xnSZk9BpsGWVyXxJsorwdSW12E7sUUt5FOUwSiRsEpVSgf74gIqZwiRxZgquhtP5ymb7QW
pVVTmaW8lKG0oRNuFoB5e6G/DV4B6sP6sUYgdY5oJb21sGK8iar1mw/JHZYhjgjoTbQfzk4bW3zV
HWaX0Qmc2i1KjXgwoZKZXrGskJE453Xe0k4qdiH+0/mzeRpMZEdFpH2gwqnHk6tvh3opO/l3XA+a
EeF6JzMzVbjv1eO2HQrjPjaax/xZYNcIFQeJV70PGmIF83SCTHwgB6EuDCxYVp8w7Q+FVz3aXAqB
u0HulnMkmGFgyu/mh20mE1UGWbzOBl058+bBor+/JVm7AaEhPIp6Ode97g7A5OanjX6rPIdwJN3g
2+1FoVvRPpPeY8x/KSs5kEBORU/m8gbCUT4wS9i5gZgfpBHrs8wc6qfnJ+MQqO/I63jJZf5SSsgk
XAD2D8gXKtf8ZOqgRPXxOBgCfcIEic4G6uHGEgDCSgMpUOroI1WnllGANDjctwoOsF1xkFew+pAC
6S39k38TuwUKyqUstcTZEioHjdiYcszugCRj2x748A3uJTxBSaGvmd44eJ0C1Rbb/+fQGnXsuz7S
l0sUq51UZ5SlAB6IMTq3wbW4fCVWEj/Nhb8bZ2JI+6Lgml6uD9JAFLxwyoI/BCCV72Uss1JhRPHv
HOSTngLA3qH2URBB+7e/OcRibxDjFBD7xWyBRoy1GnU7gkTO3nV138zItg0fvuUyHNlaoeg6Qs5n
+qZhEaGzRWU16NCHWxUKqkn2dB/6akton3GC03r1KQ5Os2ubgWAHsp3ilYQWpulXcgW7AzSUJhoA
Ftwgx6yNAvac4ldTX5UG4XnmW3LlfuRiYFwTphfbssceQD9cahBnEuZfzP62aGs2OKcc3KYvwd7e
3FW4cN7RXKCAWcXJnn2CC6fxskElvBzOHN6meng8sB60oAUCiHFYv8WCEoPsOdDp+TiMR7YpE7OA
co5ZrhDDE1JtC3G+J19N4USSZ5NXJi/kt/W5mjXkbf8Af7CABAhgjUkH8795kBHBKher6O1NNLtg
GBqTL7sN+PhN9b8brg2PS+8eTDI0jhFYx9nurpeGam5UKm1QYkI2Fy05Rw4rQnT4ZOWTNnG50CEc
FITax+vv0zZxb9ufaR5AKSmxmHJWZ6TM4duLupxcLXgagqNr7yTSirn1Qa8ogRZh/JpqxVNtMFUw
doy34aLJJdBIzBjx0XOXVR2HTWysinjBqHzsgPWroeZxeRF66IKTXdycMBergnkkloAVe6b72ZtS
/m7ekYerLssd41zoZMTzhh+uj+w1xjbIIspJKu2K/+NQAmviREFgjB6w52+VJAImsp2baiSysvun
f270Pjly6ZJ7Gj01wvazZqdGZkCBvUDCsimS3dtXS+VKIABK/6LXd6aCsaTIHsnF+o+sbJMi6j5I
XTO+aSnf8xhaR6kTJPVW1cajAGXQodXSrUC65bEYPKVdzR/KekK/itkAuHB1FciqcwIquhdnwj9Q
m1/uv5m6+FUnNF5Gjt7XsAhbCCtPz1pTT3o2IhSyRxrOa3hns7od+JtEUcCiSYLwUFQ00xMFOQIz
As3ozRQz16gn87UBk/UE4+Ww2ZGh/hx6R1u0cGpvTGZtiSrnyzyiFP/PeePhGefarb6KVHzPh4Rh
TubgQ7clWybHMPoG1AS43Ghm+5hkc5I+ahuF/t+dRQdNA3tgnc48HwXxnKxlexMlQtRqwwunqylB
lTShuATVKdYax7Om3zeI948imJxgF6IrWHRul7jsebMpiUIUtDCP/5d1Ij+tXWeaj56ZpqxoH4bC
+PXpGG7OpOvx4Hd1zbwPVYfFUF6hd/D/ZDbBPYPDY5anteNN0jqq3CrZZJ6jK/MiaIn4MBLfNBmg
kNlUZbYM9aLHc5IfCiBKkBHO20phiYXiBcOtuvAAXUYGN2zhn2kzaESgQ/E/rDjnh321BEbwLA4P
0AbAj+RsPBOx9+2JQiAxdrbFTvzLxnCZzL5FCMiwXqYXrnvQ/Ex+kVe/rMj7zfSWDmYIYcxtNshg
vjkeFYCilOJInSAVYOEKo5KBcKg62qh4B4++pjXBKLtlm0KrEUulfU5/UsZHJC+QLAa7eYplY49v
PZz2BXiJhUyCeq4Q9UIzk8htq63NB+4/W0k50AXWjG1DtHqi5Mdi9+/cFavnx5LcZVxPvFP6Tys+
hhqGOK7f33ybXd4Q+8PcWUQbFUYKv2c7XL5DqUvL5YlrXZQu6bFGR2XB7RB4JQMJPpMaZ7WiTxmE
U/FCupVxSy3eWwgpm7G793UvsL9uh4Y8pUQVx/uifDhYqSPT7rIYuVp7upTSJ1umqz8JVpzs6ypZ
qjk8WkcGQTijdppuRc8GMY9UjjjPeFSfmGjfdODyoOr0s0Jqkxt3D6i7I04sl8dljf4ruXyALsqG
Tqe7pnM4OJp1pnHjl5k3zhS3XWsqZUhmii5K8FAGTvKqQoo8atesXCbodyjHvl7uovchSiiBeI13
E55QdjHGIo+78sxlwEwDpJRGb4ECJRiSf/i7lXtnxvmczy0EVEqfPkpM/W2dsRsksQ7XhmSbe3as
7H4+RbUtB17ByeEukynuNTvq+o5r69sBE0jk3j6xEbUJhuLhdtRtOSmoOFQmdK3gByrQsK2silhC
zoeSg0wq4bb9SNn+Lc/l7YFXLzwCfLW49bhuhh8msn7sHRKml9nGcxdGLCjr9lrifDZo/77LS56A
lyucOaRHSt1NQSBcL9du+xP7KzpXPWTgQ76l2qRX8/ZR5+kujf5aPcpuDxbfjEIHFTT7MqDF2pID
uNeDGeoUWROz8q2ZOXHuolTfzzDYAnVp+1Aln+SM1cLcQIxzbEgqnOElo9bsGQetq8i9kofpqwA7
drwzJbejSgE6OxWHnrxT7TBY3Bhaxbv+Vek1uV3o67EM1agPjRVXxYWCLQssC1twW+O4VZLDq4E2
a6rXe7z+7JP4YMN6nO2UpXsmsblZg2fxPEYGe3axACDTYzz9vFmwob3B5TPJWPTstrZDc4A6Hjt1
EgL85GZP0BBpxuDMn4g+twxL9xkYLJthTAQAX386q7EQ8jw+vwCi/t7tQV/xZ18UU+jYGvzGqv2e
82jE59jYcx2PwywzycZxDeR+69mByDfgvIuVRsx5CgJ2KOwhKcM2SB0j1URZImmu/LZdNAzJb8Cj
cQmCtl29IkZhy0+nbSrSSACKYM6PRKgynozqBDjp40bE4N9vyFm/IqiYMZbY9S3xtnWHFVF2fNFf
m54j9YV/H3CHKcCpQG8gl3QCtPoCrqj4K/5QYqhmr7kyLNt+gHYBPiCHQ4SOxKd409SEj++ifl8G
tj7uskf3A7zPlOZtekhH6ssIw+GCCCbvm5/Fmr02mDYDnwBo618jCG8IsnPtt6ZhGgiF7YQC3Z2V
gqgaxLKZXrn5bgotT7LJhwEpydZfRHesjUfzTQJtun3P76tda1AOhF0rKpyPAhDrrmD8sSkgIERt
gSGpqCR1jy2fzUmQr7YAnx95zzWG/a3l31oUEK8Ng5ycQrkgqkYiI0YQ63dML3AMqzlqSi3X2aeh
NuLNPOl1Jy+Pyqh42KGsWC5LmowS3AJGdA1FsNBGyWXWsrJk20xre2xEfsGPy06btpSqevLynL+u
sZ2ZvYSKLpfpPHOXw/J6hGFT352ooxtHadS/vvbUpV7dEpUbTJOJJUg6wgciwpifbyonop/FVt2P
OqOTVGOPP//EYRyRg5NvdU+0KEqFcIPXTuj//GmulTpzQKB1qHK/Rb8FBOAdTAxgzvIepn0gU/7P
dnjjZO+4c98rvPKP/paDcXmCxxQKYVemNXiy6MFlUktTIb4YVLhHao5f0WItjj+uT3dHGmxdoCBQ
1m9eZpwFmrkL4s1aOmUjkSRsSusFI+ON0pqL8hBv4HigEhGqNbDzjvgixH/9AykppE5aT8sGdBjk
X7uRrD/0PQixF92g55vkdIwFfk6sQXG6FBAAWbqcqQTmfk+x5RTjrhHIw2Ck0OaE7I4GEG0AYDIe
kHZYGJzCfMo3vTJji9hOROffzA1EUiXq1gfcbXzQubIlLO3Ibpdm2Ttq6u7xYwAajlq9tR/p0GI0
frVpzRT/n6+rurAnBbhMYVQqzW1tM3Dpi9T7OdL7IDY2k3PRCrduhsUkXNKmuFKENmQfzbPHvAGg
rzu3tWU7fOec2vghsLb+JcdqB0xp566msP8kWIbHAseLbVqOLKWyZxiNRshXk57lOC1BlW3U3q5u
tYkwMS/gvIQaMwh874t6FKNR5ndm+2ehwX6fQEbZwquzibhg8HTqIDXB2TrGTOMRFcPJO7dHghBy
raIgL9Ftzcwhd2uNvkO//rp+YyvSnfH4zX97s9jH/500g2AY9GH0sq3HJbubVI+2gybvQh0Df2OO
zUWyyaeQzzfJ13NegXvm48eQ4r5AA84OyWxZ5ynPqiZ2dkfIVWG2jUHhplTTdLn6yOYWQJNksgxv
MdBeQtTW2EcXcSVAksmB5uk3ZXjTLUIId11YJad3/TF9I4OndOmZAPOOm8EScHjWin35vSh6iNH1
2xl14d4/XTaEtngheCKbo81eyWHGeHCn2IE5Xgq0luoSBadPDt1GmKT3gX+g1RXy6wyuU/tXdhia
9hJC4bl8GkZu4YmbFyfcyRu1xOptOYf5/kwktYeP1ib3ksyhqyIt0R3zJkCO88AEVtrmEQ98yoYZ
wrJcYbqKvE+4Md0lOqu9Y7HcfVs83jQskzJGxYk41bF34pdkJNrOyICa4eCh+ZD1VZp58qtX9fVF
KUgVz7Wn1uYjblrkKsKRwuormVc4zRLxOiY+7rkQK+22Atuh4luaE06J6Sfhn4yF2ntKEveVv3D6
PEOoRyhTN71zw7LP72PWOTiJUokwUfIBSu6Hmzt+Swp/3PoO5cpwKZ5sHjpBvzGVDhYQmbjFchHq
mQvlBBwLzBRJAg6vCMFhw/F99Hl/DuCRqYPJEjV4sy6fdutX0FmXt6IlcVtFUVZkvT/WVf3g3tW/
Y94mB9dv0p+gzhd99X+27LlnkzFr34zhjCueC+que2tB5Stgd2/JRmapQ3rRquuVqudb8hmn6+U9
GoQTL0OD34if+Z8RYo7PDMkB+rMkh64zRNArEand+dEJ9Z3euCp6W9CB4+2GaHFKpgx2GX1M26K7
bXhyuor5qXgwKttOnqhX7h6qzAJSbVcSNBBxYV32enzFMkczNn5Ik9s7itlFT/9F+BhAAjQ/hiyC
RK+jtO5PIYWVMNtVa+B1ex3+Gx4VQkJjvWmorHTY3iIE+wtnr3U1bvJ7DghcNWMtw7T3xDzDaKVO
rbhCSDmJo0e8yWAVZBJx0cw3zGrvllrptIa3ZO/qfVP0zas1ar8gSimZ9nio78vjfbSuaoj9cPr4
1jtkBRYdjFO3mFVocmyccURG/Uh9WK4umeCU7CeXrY7S70QzOl4Nn3LSCtImcGr1miJJBQi3zJM6
kX17VnUah9UhjKKRIZdxCWSwkF9tVNCh3nrPhwNfDiS4jIBRYRWNqpeeIOP9aP7jL2UmBkt9U7es
/9mFoJnieX0LzSKfr/+wh0TnpkwriGuh9jTuY6ALnCJm/pN26Jgm2lnZCDfWGRamNagu7MdwYooo
z2R3iYtIj/PMycjt7y5ZaLClN+8aiCFNE0PmE/nuptDd/dcyTRy7x4p3vV/GIvPpjf92sjdYccoQ
1cm0XQ7NXb4e9BH+kyRFxKlEyi48EfP64BpxawSD2C+qoCikJ72JMW/SmTXBVrqTrXyhCAtgCD0n
n0TDm8fOgWuHsRee0oA4lRH1muE3UjhJ0BUeTfGXQjbNJz/6JZ1Vuy7vUIvy91TPAeBtTNf2elwP
n3rqJkjVafWKyNzoGocywqUD6PCPRjRv/WMQ/cNabv+aVN0asZrpKbt74qOS2BLYHRYdzFQbrw7H
h56jIr+puiRgNVtSJqZ+sZlht6B+xVGA+K+FOQoEP1dhfkGmUNKqnbz7bMWr6a6zh2dhPdaSqBXF
6QndMROri1hNn8ijLuJ6qRSzi3bfz8kcajZi6AfQA+zL2I9dKslmn912QakiICnsGf2UKFJOh0Fu
oomx/ZXijaogkDwc5soRX0KOStLw8xxIbkS4OeUiOrf4Lo9RFJQ8evlb0YVSBCMp7FbGaT6jBmyb
xmB/2N1Fz+FwEZC6Rt35o175nLjpHORbBaGAqKX+EdGhsJ2YUY1k5lz9XkfxKzvUw2XqzXtxp9U6
mk37o7OXkW7HNH7Uz8OkJqz/oBxcTLi/qP78si1Rt2XOCRiS+8f7+BuxsuiHAGzbhO/eI9/YTsOW
+8FTVstVYy+0xyDEVPQZ/tPydhvGPARo7jrOVqk/Aoi5+pC7kfn6ERSbkGSevhF9MHFXKe6mFl34
dWDMinD1zLMBsBeZqocemMl6FHvBLqFnrnk/0ROfK4uXNqLJ0QVq3wD2GZLIiDQvSEBOcDmQzZX1
9CJWwSsGZPHcnkAhNrd3dqkHKdNmSx8/07iRZ866WRUUnZYRk4h8/3T6+XCyJnIT9BZVEacSCABi
ZbzZ+uc35FFmZAEAQLR9CADBee87Kvx8e7UDZgBkHJnwPvAoFqYd9tQ6a5brHDl+Idf9CgcuXXoD
QQQe2iLH0VijHamj2dNRezOQfajw3r5cH8O9VWOBAcFfommdHMp7pZ4p+e4ryizF+bkutQl136+/
37qQHPb9bPmAfbppzEQx9JwRQ37PODpf2nd7ReurRk6E4lqP3WHiXDVqp4OEdBr4SRqYbcBp2h2a
buxkmDqi62XnSQK7c8M4mssxofqBsemaEaW2LflQH/i6PUkip0mjf/PK8T4PFiISOPb7P4DLzW+w
5rSB644RcRLLF6Peji09hsfycb+o+iICYtvxSDBR/Jpv7mZ4Gb4BdzvWDyKYCwgmYjJx9ffY0Aj0
Jkc0etOREPmmpUhUdPYGcq+mOWmcDWd0R4o4eBeOTLSb398UIRcEABFlgzKCSpQ4HHnzpUiQlrpT
BMZdq7qADghqgwq1sVrEssx2+8nBotjUf2NuAa23oZteZwknRa9osLHzrsQ0YPJLQZCr6Bf3HtGJ
W5NHMpRZHAUV6J7KGZfZRaSJ8yQJovKc9Pwlua/J5FU/d0mpcpDcRb6VwM4AkEkOKLbVq2EyO8Vq
AT6t1kVzV+ClidGD+agv1MQl8o2FIbGRSyjSkacA5HgPIRQwROmOINqNJ9s+g1P7ktAPI6yAX6n7
TBR00p6qdxPujikmRp42o21PVJhuDltCziHNrCjPP/EB+Hqw31EnEcdjMZeTb4NQYc2XLQH5Z8C/
D3jDhkIEW6RmgLHPk1E4EaLa2fu/0MYxCfB30CdY0vhxNmlt9z7q75Ze2ww5lRe2EAKCi9KjOOv0
BrFTfc35JwkUvlo+j1WrQKCmQe64q9s3AEsI0sibfCD8p2sQvmVi2LjFKpEwPWLO5rD6Z21/btm1
nJy2TXOjsiqiUNVzizG14v+hRUMJpe+v2/HiSgsPgKDPJLsQYYflWa/oOxuMotuTZzO6w3GOT8aH
s0Zjl4Oya0MGmrRfeP81s40lnaGTRhQ8xBziKY8RENa5vQXJHdJxvurQe6B3l3sbe3ojNaFnuCVc
+el9z3LsqlRaztnQoMrIenX17A3VkNcEqGfp5iONELqpSKnvy072L9a/RT76kAsRUyLOD4onFeqi
C9iOXYHEwKV0u5tcyWpWI2dGhTKmTqM0CH0cCQk4utXIOSVqlzfw7EILI4icXofTQBI+N5QJIxm2
Jpseur0NC66NUEwZRz5hwhEyvmgieyvf66+/CYibG/qS902cmTGwAbT0ZsR8eb4nk9qQNCxFPp34
uNVy1dguoTXlavGbK0qBKrN4kns5UIUsmQKFVQJ0kGrte4TLfHnqefq6kKptkn3vGzdpdb4ah7/J
e5O7DtUxtjWVtZhJuY8VICoQx00NgmThskTwazlGQ4Kq+ealnBpQE0kRFe8qWt1LtjCNnUzZcOGn
QbmGTkn6AZBUyGm2NkFDwWDuEVKjwOzfyMpswhDC5WO5nBAmmlnt47osqt4vbIJFkhX5SKZ3slSl
9MvIPJEln94LLqnvamtvCtvq6AbOwZOsmYOhOYQInVa2YIwGnBeh58buxJoYV1oVXoFORb3LZWzn
Kl2nvIYEImv3QzLuEpufsQsfn1eeXuHtmuq/dYfUIB1KU96M/H7lU8+90wPnLxtftDu+d+b3qhpT
fZaDFtx1ZnGWGiNfaK9e70Fnvq6JHU1GI31d3dwe/7wycDn2WJekc38/MmY6Q5f8TlM7mO7mvBSp
BwqbicI6K0iXEjFZgFtL9RWdF3HIVO9XMYBhIZbXB3eRjs6uSMAb/OUZp8fbGUnWYqXTgyEEXFOQ
znGZavbnPFfr/eFc6LdYdrfUVRh5X+qfICKd0f9anxAujGZrZwYTty1xNo71Ab7h3q77J6g/r0Hc
62icPVVGDM6FK2lD1BjmEQthgAySb5JxtV814OSKwJsVecSONXXQS4P5MleWf8dOGthUMxT6+4Oo
n9hj/KXv0QHuAsMavd70x5KaRL6yNtbtfEJW2iY7EyK6GU3Bq+6/NQpmo2V+1k/PfdLv/nHq0cbr
sJCW6icBtUpAQuyAo+jbJ1qgGhZ++lj1QH7w1jctJWpEaUkeoodVpWnaRW+ogyg64iBo5ndyOR6L
ckDgk2sxYoSy6t8cQxWzSJSnvPikcx8RlZp6jnfFrx7RcaHGXAhA0uLQ8WgieVOZZjv9M4GhiKnt
Hl8lCjYDqXww7DuNFzvkHPo5MI3HoetPllpOCvbrZqzQWUwge4xoRNZBuXERxbmp/ostSBfOXFkO
4B0gHT4YxNwqv4ITXVbbdO72cndu4WtAfLHYA3X3Iwalo434qFFabUidNq71SIW8GOc9eVkc0zDV
GvFTq/cezQCkIzXyPEsjuJdau5trEBXDRsvs81WfwbuY9+Hh1IzxUiwrXSp5gf/2vc4XWA0=
`protect end_protected

