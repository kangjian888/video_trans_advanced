

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CvmaYyJzAT4gGJRlCkE1yXt5Lv9gJbr2gC0wBzixkhI3TupXRLTg9s4Z9WVWp43QDkUuM3VRZjAj
RVnqESt3JA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hHyS2uxRkJ6sHR79RwG8dxYfMwySDoNzo0ZpVSoiAp/93R212I5J1LxM+7EujDw/cO/x9djlyxbz
erzC6/tIqQ2nS2hUZANmmER9YkiA1RlXlIqDOWo8pOFHNj1c4jf7Zdq7OJMDPvKF+fLgmk5Lu9Y0
15oIyfQw7L+gXpW1qEU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Cfhh7YIOGyVJiZpd5j8xa2ugbHZdDDpkNcw6vvVCCgnGCfzlen3wlGk0omzzJqyVapnfg0aPFCVf
eH/noQVGu1bQkowx0JKcNE5x1v5DKH//UNI+lq09SNF0WKlMcTAGlNSUzO8kgVv9uNbKUHDXodcD
5iGh6bHMhVPSu1QKpTfJlIMd2CMz0JfDQiVbfTaAGKvrQhaqVte7pYpnqiXM7povPwt/ntWHBH4s
XSF4J4eDVLMuQmQNy3vrqFdEUqmQFtLWgNRpG2fwo19Y2lRzT3ux5SiA0Iv55uR6x7AG21x8BZlD
JC102ufirdrREfWUzlClY8zmr+TUHpTF/SgPMw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UWceDgHVHZAg17Yudaw03bncVn75AJ6y0RYlYeqdZU3kMG9E1W6q5REaQAI7sMZSrC2g0zavsx4w
utskoq80P2avoebtdvBfjr/nBCQqUN3AvM3GSk85froboZgk4fCQ8UtEj2Qk7ob+ox/md7d9P9dw
2YULi+eG04dUc1g45wwF0ZoZdARk7Ml+fXMnm7zxmvqVieAEsVq6ETZN/P0pwvIpAakLTayKriGC
qcrb1S28bOuV+Na/FX9rxN6hM5aK7vSdFqja5GGs32r9UVRIkX6i7uqS9pWQDR0Qa31W3z6wrRrT
+2wzEwNMDKYuWVIM1FQo/Tp0NKa1Y+kyjahSGA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tLsJPLnIUk5FSxPTGLkNhAFldHrP7oFH8h39nfqyEmnC/AmGzR3fePfCEcee3I4TYySABpWhyXIf
m1jGiCuHfIpFkF2EJqjWmBev0bD33cbw1av2xtJRFa5gaQjxChO9URfjedFvCQWWwjlxejc9nD0N
O0V2XUDQxd573YmSBuByzshlxt3bujEd6Xeeb8N8NI8c2ZsfY4693LGdb3k6gtY9ZEoo4XuYVt6n
S2tNFVJTfQjyBEXbuCPqpwGf6bPdy2SKvTE/s4rSIVTO08J6bXDaEOBUGg13XVoJJqrayiJRVuQL
LhoiPzgOqS6ude1uUaMHE/SN9X/vt/6uOsOl2w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jgk19ieS+ZYiySHKvgAHMus0OAx0HPJ59p64LMaYK8CyW0wSM8LIn++sFz9tsOBdLj2gb8IKpSVr
SOX9XXXM2pQFSME7x8q0m+EPg9m1+ghIpW4bU/w4zVq4NBjYydZCI0Hpy+X3op0a3+eENVEw5SoK
4R/zOL7aV/2nZ//wkaw=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
L/BPRr/PHH5da1O06dKRr5ST8eskM6lzR1UPuTvZQ6RCsFEjTD1HgyqjW7/ypnIq7V5TYDC553+Y
rJnEENzDc6RSpzenrYxw7NrURpUedIWlCc/PEf5Zq9gu1ESkpND7t98rc+uiAz7zsn/pHD/K50NR
q9l/gcWkOCgArmADo1Lw9usrfZ8ECIPKY2kLxeTYbh4fsrCpPQsQUk4NxX3N1Q0h3RRUCdHSFc0O
lvGip/vd24OK8zXDMaQv4fPmgToFQMUvLrJXErEUeRlkpxkcX6g6Zu4RMWwwmkNIfZHpc5K8Q3RL
MMc5rARUSXbNbpf28H3iyAMZ0y+EgI0CrKwooA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967856)
`protect data_block
2qhuWxpP9pIZM+URWGll5ql7GGxc4WrY95Ns8laxEZKTklf0WRVQgV3Tn/iGIuD6wD30aHSITOLM
g7M4vSOcaoUo1qjleFCcZeRsIxxerAMcyRC+MwHLQcj7Ymo5iIY52euSUr1RaoitP5HTKk58R8ic
V1sow35FNkzpOeJiDH6kqCDHJKZPXMNTFU9Lxn0/4gK2ID1Hn/p6RJUYk0zRm/08IRoD+8lIsw/I
v5ZfTtVIfbgslwDPlibfn++f05mGTdrkF5/FnqS4xQlvBU2V5d5bRGqnG9DgY0MAITsjZDTSwYiB
70wnOgsmsoZyL8NU2QsNO+g/CZRKyNj8ZNQOUFRRZS+k/gbnM7pu4IDNwH4SIZn9isHJjrY8hVcf
XWBAI42UVE9qkSektXobSwrYwYqdip5WOFClJohFYCX1JsKv1K4R3n9pxNKfCHg13R6phhM1MEoZ
SY+hpk6J6jeVVNomKeBdKi4IXXcAeBuKoeGxnWzMj5FUIwGYQ2MoBdo6TU5ik+0s6p1+VkTHvHDV
ShyLO6Kx//0jSQGxkTrufsHYnhNsIfYKbQhnlwDMuDZhpEdrdiDquF9nA2vNYr/se3mi+bsaw62N
h9EdAqRO2fVWL47tS/oDhSeC8vXEmEqsVlTXtv1jKVsJ+BF4H8aAjlvVLbZ9bfsNzHjeqS0fY/2Q
8f31V2zUApLjlN039GvvTLeqSuUbvOHXkN3kIcCEfQL8ORL31r2P4wBsv1siSIsJL5Ep1H/I/2Bv
0KLJQ+X6VJgSuxDhlFmPivM/NRXM34aoxbcfUDlxImxYUoawDlQLXSj3atm7x7O93IfvHpcS3bya
3JjHLiAMTpogAq/0t+uiHcMvdsV+De2Ka3qXvUx5COQJtpOnsjMx6oBnbRGdir/Ntk/nfirqULww
mECTroJppgMtozXIFAanRPvCvoXJKyGkhR6AZwHjOhRITDxyp16++kj8kG0pyb4qnnu5bdjnupef
r/WRfqzMBQcq+mOwJOzpshWwRiMGxRzf2eHuU7A6UW+mI+rCYdP+WHfZr6fMtV12WuQWDPfCuWMN
PWK8U5AQ8r23Iy0mSrJ5RCTpGQ3c4lQoru6NB0IXWmI3zMCAq51Wh7aoAW8hIUi+pjHjqw2UPQGA
A816eH8DjLX4MGsLShSn+PkFABulPXeKfF9ilnHnvLFcJMcjMsPL7Ere+JmZyU8NNz87Qh+skW5G
JP0s7YhMudP3wIXFgxKOybkJPg4JpMTonbo9TP2Lc/gGTEYpunUtlGWTZqKMknL8pSGONtz5xnuA
KuIko1GY9g+3Msit9QTA6LHgHEAKqPm3aCI+UNTyQfZAZqZPBSk7nnb8x1/0XbX/Q8UrWeDgrTKv
HMlWfbsjjbN4dfakam7HMz1V5YIWzZBfAwLEmKd/3vKr+IPZ65do3wRCcv9syqt5mnetKsPeJHv4
TXP5bg6jPStgL/cgrX9GUU3QYycm8JM6LN6c/I7j9LVPqDbar4AuayZaJqEPCMJoRSzGfDEQhMAv
/KWIXT4qLpzVU+reJLzGUrTMTz1B+A0wZsjHzxoUNO1ApToZTAziP3Zc1NtYaylip5pkB2FF7oH+
AgmEL3l5r7FuSIoQrvqHKy6xD6I0IFQHD3gkk2yMvA0Dz3e2mjvY+hCJ5hb93LjUefQ5Qgp6FWn6
CZ71sSVEba6eX9nCuXIgJxM+5IJq56BzHzqBdaKRFuQaXPZkB+IL+QtkxLX6xWpCNY/72C2NY8Uo
WUgTUqH5AXtTgid6MiTujIqvT1agVsiezKPiO6ckfm7ih6uHMcjJJ2Wrsqa93aU7jBAqwBMjnKsU
7YajyxaZ6WY7kTRfSFj3xdReINSqHQjM3vzJKeA8q8nEPVfjmZf/U6OmpCwTw5FMmwXYaoyJmSOH
vbyV0Ai3edSjHkJoRcydT/sYX3WQq0EUEPktXoTXdha8CbAmoDbDl1T7g8/0Zv/8FageQQV0u/6j
kkYRP7cCCkY989wmd91/qwzSSxQFVguRA6TQuMAPVBw1hG/Oki63yPD911HcEq4PiF7qDkcNfKUQ
DOk3e852ld4bMTEh5P63p+V2jql1xAV7ifaez0JD1jOW7JPRv95bFe0RBVsUn8a1ypsIZH63Py4B
TFq7JcgCAJjPB5RIhtd3gbNymlLBEAvhRIJwOwqvRNEsCjMsxg7DFily3TPoeyI3bk5wZtCch8rT
R7vsuTQ3CyypfrubjSw1d2wSmEs1rfh6SacS2WKgPFQMHs0PInVlyrmsTBXt24IdFCDrzelGYgzY
lUMIAcmdndRStnVkjGSiNibR+ECC05GX+LUVetWnn9XQpIV/g8iYDfrDxSlCCaUv8/FTN8m11kD3
Lod0AStRH0Ew4nZ2HORM1BGMfhQOQ4wFmgu3yHUj8hJw1NV4e9TdXOw3BW1lZBprySrs0Z57yrI8
RN0gJnUWCsdgnkdsgqVpghtacNQXiO9uL7XiWI4Hh1lPsQFmrURVpSk512ia4ZkjwvTa99wbATHW
4EhVK3BRWwrr9ONjQyBF/zMv3mgeyvQ+oL95NCyBww9OvObJGPjYMmcYytetPUo6MM52dXOlmmyR
Du4tHEoGt7CQZ+XY18FcX1/NBZ7qejBjMjE27dGX38ve1361Bxd35pKJjm9KmvGBRsYmrF4HwE2L
kvpTMDIbRr0jl0TbsXiKHSdrR/g5cu7q9JD0dyDuY+1uhUB3jyqwQICWVoe7kj238UmsmOQUwYXl
NkjSu3IVT9A1CKLntfh4Q8fEzlR7e8K4xda6r7RmgIxL7Z/zoeLEVC6T6ng7PNjeSrAPO0R5IAhN
JyXO7SGo9LMpiBWkut9DCxpeXvNhLRaJTT23/3aHAxvt2rhyVY+ikeOCdmcQmGPmWTcQ1CT0GVLL
SK+QMp/W5GdONXXyby/CE48mtBSIIifpb6k+qUz5DqmO/CGTWjF/kYQOrblMEX52d99vz3dcq6b9
bx6w+ykdeLHI1zLgkUxR1n2BPZdGsZNj3iA0jZmS0ixjU3KugP1GaSh8vUQnT3hhCHPWRChyNSeH
0fkMF5cMsShf+AaShWp2HUShwtkWYSa2tbp7VXsjOYE+LylGfKyPKsyy+yPzIkpy8wdoaFRIUZ9r
c1HtXwxEc4AqvlVbaRJasYkX2zrJwJf9NnEYZuLBG1Q8mIzhXLJiN70fBQtK627XZRM1RRkwtRa/
k8OabMC+Astw30QzexyIYNi8icm2jXLdgu+Pf4texG9dG1xlOtKHbHbV1Hiw3Klixk0OivgI01yL
9owmeGDUXxIyks9xsf+nv36DJYo9/XTjK1xaOKV1FT4reAsoXaECPRZ3B6/Fs2b8yvAb26lMzJNM
bCyJCqE6msMaYFUnBhP+9K+k5uWeEZ5nElLKPTH2PL80lJTWuHF+WJM1W9zVkX6m8WecWHo/JE8o
II6RfDoLKYyk3Sz0BiCH61pNoE3c0B7gt6ap+7nx2FbCF4i2dFQrV/2eqRnVn/sfnhEuDBVSUV/U
wASu+8B4AYrESzO8TEcEkGDBM1N+ne5zFIyetE/ea4LYDU/MuwRTdJVXHM009c99Yv0rvg+WQFSA
fHq1+nG08Jqb0+ViyqM0GyEFNOnlTTnGVjw8CMjaJzZ0mnm6jrhkmFFRiieg0LLq3+kK7/mTT1+9
BNt2AYSCJvMmU5g/tqKELkffnedPdswDkKEsz7z0Jsybs7syThKPbYh2zl8SCK34nAdQ2XgLGznr
Rz2ALULCSipJUYq2rAV1iqw6WdSSUBXztZ1EJlQHJx9RjtnkOom0y6PBpXD5RLVJ0pzmkxRrb2Zz
i2pGnoGuIjXVDct5PPZluppkhw82CtVWQdhz7oWF0L03TrBE4mnGN6lVXvmNvB2scHDXft5/6QMQ
qAB2rtPN7UrELXXQa1+TsIUhxswIsr0uPIDD+zPV3CsXGV/ydcw6Kf/agvvkYBVzz6E0LMOKLXZk
0S+wJoauf+FgPYqZChbu3tm8IS0RphkJKG+m7Pwd+snFwcwLwSIIykOgRyO4Lg83UzR7Zl32R7nI
O6iHrbVhUAXF6mvGGLezuQIXL+wYHOlBTI471daZa9DWridHe0LL69HV8Mz7bhNtjcIClLrjds7m
E5pQZZFeCU/9O02uHRep9GsjooivsKCy3fntRZDfUO4mdSYgFCxLEc3bDEvy3Vfknl9nhMzloOWJ
bxyoqG4BIyGiDPFPHHQ5UHpaRjj1dctW7tJb3BdEz/2zQVLKDg5s+eHEmD5dCQDNGDH8l1ATmqf6
94dBHrlk3E6bnsPlV0KArjYfEqsdYoQ9/IIttd0Q/MzzXNV2yGIG6zxsofkbKdjnnwa06eS7HRyR
Ehtlpen3TCuWXaue/GN3RIM91MUpks7aFPK80wwQtIY2R+8hNTarSLvTD4RuSh2m0yw3PesSkUt8
tZzmGxCiNVT1FomyBGGbroK1pwmUV3mIfcCz0Fy6BKYWJX00yO+Z4MU1Zy+6ghz6zEUYjIh2NG8V
wiS1tlATQnZpyj6l72ingkbIRlTqesv+AEUidFADHaU+1Ll1hZTXRX1jWEKqERPlUDaT7o/UkLoG
m6h22RSSZ3vT8ES/bnqrksTyvVDGQ8/Keq9l09QRJWlhcmFIuqjb6Qk7J7XziGgvFWj5IDY+4sBk
FXLL5IDTT98Umu3jNFLYdsEAlouHWj03CkRWLVDxC/BW6ZNywHKqJn7A/I5SRzUUfXloJ1cpfwEP
iSsBST+nzRSwy2YlOAtlHp+3vX38XcxHTkk3mIX7hPpzI+Xbl/lbJjDVYqk665o9co1PmeVqR56R
ZVbC/7imgNAWpvt3og5gPCTOSQP3ryc/pJVgputWIYfZ1PhAUpbMsqggKtqLh9gHuci7QBk4Icnq
MthMQHmBvOzPQUie31AHW9F4fEwUf9zwfl4l0vd7HlTbD+mU9RpeKJYZ4JaZ7OL4OHhCEGlD4vuS
cGqTOShllcDjyaP7Wl5byWx6muK8pfnOPOO1Fam9YcAt1Kcr1iQsV/tJFSvE9sbi6LbycMMF3p8D
1W8qVZ9Bg77oSF+W7xZnYZdHI1/5/afUobpBeGxe7xKLtE9CHEy1fuXhhd+6WtUq3RogKOCWwwm9
VQsGyo03SxE2qMSQyz+xBKotTdXwjgxTIg7jfkCRHg+avJrZhGBr4EaC7qdbEcZSyQctbkDpR011
sHwMwbkhKlOjcgztBdzfOU5VlcQvS1tp+Do6pkpg25xwrJTWLG4C+pWwPZrGBmSnpv1JvMbPX1q4
0OKioZFEM8CQk01E1hhWwhhGkgFEgp3oM0T2z9cldmy89MKEiT+2mmGE0MlKa4VCuzduNcyquoK9
fO4GvS+ycITcEDeguQKpInkRNEMOHwDMnFqcjv0KimLMA7Q3P9W5g+xicebqYAQ5TSiUw5S7BApA
cbAJtDwdfvXgYuuiX3okF7j1PhHd9g7EEoJIvkZK3Bb6JaGQNZrZL+yWgmOyXnV3OOIHdy939K0c
jzEQTGvqdzhyFwXIP+1DEOmD7wArYbFdI7vUV/G+pxtgVebt2p0soJYvpc95buIFhe+DGX69V1Iw
Yam5y+zzBow3Ksi+tmun1MRzU3raqjxUV5YdC3738k5nR394FQNwJ4BE9yi+LhqXl7FjOkYS4UHL
lUWZx8ncU0zF7hcCmlzQw4SNWAY2doE1+V03yLqYkwla/yWukh3fZ34aQiYA0YRAcdnW7/teinv+
1oNoJnYcQGDzN7802LR3dBCFEsDJkPA4AggL5mI9DGsX46/blJjwXwAwcicjK1MPz40PUaZ3sHEO
r8Tch3rxgBJTBDpdynIDdrYskwY7FkLG7FykoLDrIvGr7lVPveplKMzHsqXwBokkbs3BIXBEYfyq
W1v3M9qvlzqq3m6Bk4S82H38iCiDTxcyg6WB7/vQwUwS+gQ+44qK19WqdktE4VPQPjyKeguZY2o+
TCYCGD3yQY69K8IqpZeFv+bSzvFKgWBvDCfBjSwh8LfahFZ5nOB2ggMqstWkY8S3dwlk9L7U74s3
9hppvY5+ghUYMeTCA8hW05okQN/4w1o4ZsO0NFlLYJW6EF79M7j8ljI64VM1jqr2GKNVnOBcXe2+
345oYM+KZO9bcdDmalapn8/KDi9ytvjM4mJefIvD9QBLDeoHsmmOY0FiU6HpkdVEjB1D3oCa59pg
opYN3XI+zcRDLsAMBb0PoYY8adjlGbazayzNYyADmZm0MbF3hA390HT2L2PtAPznVeFTxrYlTskE
Q2Ei/+42znYjnavWCM6dRx2j5eXGJBiJ7r1Mm7u6LEQ2SJnEj1QGWygXRScZPoL01VT8pAG+YUKh
8wPd2aLVEhQ9i7qtqdLe4KU6F9j8d2PeMi4NdiUZNhCuO5o7n25MlM9e0KG5jBrjBp5QPxz9Ji47
m0AGhUfu50YV3IPacodptxqfJ9e8sjVvHdLRkIQbSDQ+zzwE25hRlBQ7gNRp9RocQnR7+UyZwPLH
GoqK+B6qvj2kqdKvwdyplJTL1MC57lvZx5E3Esfdhoq4N9N4X61Dy/syLoWaBlsf/HDOnlf1xO3r
qVLDlrZCHfBzrOK/o6j0QA3MRj0HOCl3dyZT3YbFdtKyaXCy4Ku01koqvyY/71J/nVfGilMIh2Mm
u5LIKpbEqgfX2ZqxH6w65hX0zh1xVDfIuySOQqCmTOjdq2tLpL6kOC+rK8t+2TGJwxma0GCsOedj
av+g5goCstEMkyTT08os5CbjMEQZ5EwdMxwx7hsIBPpXK4IxExUS9I8CY8F+1fv+uzfFsS848Pgx
4xklqzOn4f66+ON1k45fRCQUM7UtsO5HbwIaXy9pQ6zpfnz5AFGFUYBHIIXdBfVGAC9vUjM6cIxf
xN4WRJI45josQk1Mv84Ah31k+TXiy4pQBIakHTzFHzb1oVRsvvv2NXkyY0UhgCOPxHl5HbWNz+XX
YqMONLkGwWd+eI6lN23YUkseLUqYD0G6Ct9K3cw7kcHZ3UkIBzT5InfRj9pgZHVqxSEMbLQ+uBnp
pb/xfKnBXdSRs4wLBvbMXbYec6j4ZnbjGqrZGAWmbeIGUNxoRObH9UBiDgkmwqaPDPr/u4/FcBTD
UTTeVQaciXPcvmJk73f9wkt+8wcLUlqiW9hf//MmhQgvQXwjYnw25w457WCcKzudeM21KfZyUFgR
fYNic0y7TWi0zR1EZmToTy7bkP1SpqFogmuEMt3pdn58utMaldJyg4f5Gsk2HHAt1zEQtGX4hsmQ
Jq3mRoOz8Ki4umCjugKkuc5GfnldrgcLm2vGNeCqGiGlIMCJFkTSnOoZhaf5bZhveQe3b6IVITsy
524uGaDDDtLpsdTUtxpj//Zd1RJTyU/cGBK9Fe5eUMFoPOd2nil1v8J57AacDzNs4hqqaQvkaxx3
CbS9KD4znjx0xSFMDv6eoCbJuk7GnjYRHqA0EtU1j3K9Xd3/vbtr7sXfhizmRjGjk1ESc+ho8oRx
Q86vXL/11kMo3PipzHVD4UMrKtkMdbx91wtdhVRMzWlGhwBHFa1+PgLRJIJVnlocCrUJePX+TLVY
QtuUhFV86oQM/Kf9rtNn/JWNxsrRGeGG18pRQ+vTPFldORUREsCuoSkBSBBI5X/RogO108zoLk4Z
HoULdqVIUoJLq4fTLVsoHQqb055bJkK04eE+oV+DExIs1cEmIrToGWXIB46gf0DmnEk1sQszzu2B
cFRvbUaMn0wGXfBp3Ub9QDkxg16+JWUr+oLWfvroR3kBpq6A/WRIgO5f1M6BP2fqkZuZVjOhGzyq
AuwH2fcw0KhmSpeRCdfvqf+XAMBsTzLPR7YN25qQpC+mTbSKrAca/dhA1+62MQ99Ygyci5EJMvqj
fguaOdsLXAm84yshgYnoia3YHbv/Fiwq1hKvl3/cWLnSOsUCpgZcBjyGCl7memd57TvqU7mn2oeA
L/gmlL2RsyAb4EZS6aPhBBTRibOzYkS918+g68GYoQfbrNRCPsv4Vjjs14ta6lOzMd6WpNUZsoPu
0atdzPJLNxcqCfgvzmQF4txHULvDnCEp2swS8AVKB2hQacAOZsLy35Io1S5CEXiKnZw4ecLSKW/8
f59PqswPHA9b//jEHRl3kF/Vh0qCeSl07kUs+btmJixTnRqIOcxFppmZsXi4ItVfJwbtaOYJDdcj
qOB6DUQfQ2Lz+5muokoOSAdS13bwxkR9aRFwHV/2zPUC8HH+unv2SVhYb42l7HVNbNa61KQ5HBuo
coG28H4YtE6vIAC/cd7LsKDbkaTA+5hi8X6kLdT0753ervc50N/QvaQ0XyxjR/KlVGuh1tv7cIaJ
yDL2lummRnT+gjSWzyz3Q+Tr+5dsvKd+tppZH85qyjF3T/D/AutRO8Pr9MVGal4pgYPbndNiXpnH
FK2dxHY9Wz75+TwYAW1DQkMgFe9klG0pNt4+6eupFVXZMebD/xOiNiqnFlt8MXO9FvJOpLP71p1E
7GkefGdqUxaSbyvuETjb+kQUjPX6AK+ClmI5XWhDSBoLgcK7uyUQX+vCdlV9TkieL9yV1Kx+MANV
m+PqPj/wo2RRpe5CB2grtgOgPg5hBnVwa758xUeTBNymZ1r1u03+s2y4qs2WDFkiIhl0imtZkBqs
gfKQP/FU3gb9YcB0lbbKJl7wwM186lVKeyoAY38FiRUpn9+hEOKXhDz6eBb1gQGVdUey6KZeUWBU
nDE4isex+fbVnO7UOMMdyGIQ16cdcRohHrHyVLi0IChtKS1HfGuWK/zJE97cXhx4oP76xnE3BOxK
YjIumFdCi6ynZ9K1qgGd3ZmhH3AeOypDpGzQYqACh3JNJPSNTTBgtRLdIu8f2MZQYrkpRgsUD66Y
ew0fLAkpFil0HgLNM3Xe1TiahDUYN+eIPRlglmtzCm3a3E1jLTFZNVJWwcQTwpOJmxyMZ3PWHRwJ
KGETcWqeEHOi4BiOq9c4xPOU5t1jK0Jq2KJafBVZdq1K1bjwiUPiaiJ3Bj0dwAxLbktAZ4cyNz9L
K2mrsskoBXYxJs2PXd2ym0xwS/OtUpiXRPdzq25JpVFl4uVF94GC6HhzpdBAtxb9ZGCtPRTQjeoc
7tc3GFP+f4KEUKPq6SEWKlqvUefRCSEfNBBbhR1oCL8HqnKkIaq5hZDpgOGsFk6OOsYMvcYGnPkq
jUC2elHMoBSpwBWgZVjYrp+hECs00q6KFDYdv4omy5+ECyGc9vMXMPSBD3635DFXL0cflWlamub6
5lsrSu84YF8xgFhwU1FxI5olau6ZufqBhq4nEAasYusWxlfzNgx5QStfk7puKJ9Ahmq52xxgy1zY
lNLZCopt5bi5oXs2G5i8xM9nujOWbIrDe0w/vbvjlY/yzzZMN3eZJHEm8TMVb0HSRx/Ejpr2wTDB
2BiPICx0X+UxPdl/Oaz3qgt/ruB9eXbfzaUU4WTF3+7HkXqEEIM2Vj2mg5EMvF/Q0BpIQJNbscBu
MbnmHP1aX58chmYPjiC8BxrV8q7+ywM76D9fMVe5XC6dvDRZkCLD6kXtZzZKsiklL1e9O8e7V2qF
V/cWZPNDLG9FZToSI7Pvdso7pEmn2onatFJ66vhViTXIWPc8gjnlX4hAS4U2i1vkHvmtgf8yI87f
6rQs0mI7z/1iTOoXnNylk90HxMRjFGGJN7x8APsyEEKHsX8HpHaTDKbxCCcuT69/1yGk1iTweUXt
EQTBZzviq3KBtHdhb7DhdjKiowsMfPlJx5zd3hcQRIMbVoL9gye45RO3i7Xts7nN9wNzA7FD1m5i
dXui/+sjdxzO0lqWml0GpXo++TuuWElEP748xFrvT8NEKLFT5aKudagA443nvPMcBe4KGo/5JqVY
f45TDPKK4hMQO6D6guhmcylCFeAhAnEOnv439lHYxSNlny44jQVt3qR3bWcSq1p7SrRSQGocz+7t
tEjRVDOAlu7sRgpqvgdLCBtytb3DKHx4LtNFEmv23t9mJrgu6jCCBx0n84HIEAPtU5x8MuPucAaA
ym+OP1eVzkTONp+C/73H8PpmTq5ZYs43cLqzkKIWIa/ZM13/ymtXMp6eF5Ylcpl/ex0yjkKCuQp6
B9yMCRLFhj7RyKJTq6/IEWABr8gxZxg1ABomRNzB9+FmhNc6VB4sopuYRsThh9aIiEj78Df5gX4k
xa3nImkEzzAGYSu3cIFaDbxRION8UVP21w4bTILYAye741bS75W4y9efSMtLXYymWUJv8+mi8mYH
2zBUUerxIAmqdVS7bYfe+fz/DDXB/zyV8hYlr6fWK4vW6trryBFPW/2BqBjrxdncdargK9F7Iw8M
kQWuGoXiJRryhfWk5snecIOXhFH+D/JtJL1q0es9FqZqQbtj8Ks9C7iXZAnUnx2453I7COI77RMR
ga7tU+1paM8mrg73FVI4WCIOUzNyL0FVkLnz1pUnPr2g1yIRI6+j0uLMtzH3bEMJBaA7G00Hk2F1
i6CLVk71lIs7GqyWtgRuExNfffsGiu41SFPZK2cjrKbboVw5/MUMiQU3R98wolGXWssr0sGTI4ED
Q646D1iQwoTt44YpFWCy3Ftztg3uq12GdFV64nHZ0ARVnPTdVMYcPs2lnPTxTbxFqc6j9lWvxam7
aUDCXS+liP+mB3EBt4PZkTaWQ6jUB8ZCLFdvecInRESDSN4zosq5hWa4eXlhyN1P3a25Kckcc8pl
Wy89l7Bpje8gFvZ3u3WRmJebQzo43hxFTfPKwwgaeGHjN+JHg9/LaYkdkOnhzxGXx8vEurZDAwoI
HIx8rNqVYjTk1n3RNIJPJTxA8glfjh2Qr/8rEo0ULnsfJ2cZFzvWgkaA4CyzNfLytxnhATfLRWTv
7jAjnxo/HakrDVaHprb8z5QQtnuW6njaJrMB5VYwv+FTpKZ15ZMeCHmcnWC31qDEacAvPVQCHW9Y
GXmVFzZK1i0J3HYK5++fsM+KCotdgKVdnBxm+0s385aNpMNVq1BCVnqs07jYJgeStnR9p0cQ0g1W
Hnt3Kjyy8vdpKgjhRB3rIN69yIoDM0AJebiQ8zAo2OweVgXq4Xf9MP/AZIU6qZtXcAHMAQWTCK0t
fXpEw7Q8cvgvELcTk3ekwJgB4+K896pKRfkNAq5lrygpwz46WwHNM5xZBdXbDUGResajJjRAbSyE
xi52u6CpEmqTSDVwHUkJuUmqhnPocFpky2grfkeJTVnhvo6llgSEdYR6KXzkGS7u4JLltYISfml6
lPH+CtXWwsrdfWIOdaZz30AUOUQJyiPyq1kVtGb9OMoNyrWW+TX+CI8llHSZ14DwtRjMFX5DvEqZ
+aH+7cJhkIbpghUGA7brp1eBVwtKkkg+z10bOEBPgCCeKKGSepKiAqwEmxxZ38YtXqy8r9ZQAYlv
LF8TRFUSdLYg7lQU47uyJuiLZ8DrV7Kzxl9HKV0UGPtSpa95VSlh8L4VS8eoI3B8PR6GId1U+ze4
tJAJql4gbr6mLB7xEiKrMowK9N/fnn6OHIW88K5TwhbTVl5AgBW3eKcfsJMj4+YTLP0I5WnZ/wbt
X+Brcav4vVDUlxupZDHzODJpLqgR7q3/co24RiNBH9jDjSKq0zI/VHIlc8lvziFYU+cgOAAoqRQF
gCiT0JGy+mpY35X58jaFbvjaQLUikGLtpVXhBEZAcaskQ3ZKK4Upt+HE4nPujhF7a54C+zgjG7qx
7U5r+5evp3JTQXVD/jNpgr7jR1A1jeZzPZuopZnmE9B00nWRSZtBtkZ8OMjpVrJIMeZDb+KG48KY
iDyQsxBrELzwCsxqswaZogPsHPx3AlhqzNTBegx3L69NGinav9i9DnTn40mhSIJzHqQh55OegktZ
1nOTRDUUuFQFp7Aa6mwdlBJdv0kcKaS96nmTIXpM8rv4LHe8ellIMqKsADzYJbQj6NBJxLbcmj19
MZbjNLmLAL/mP51/yZ5AgHn2egIPM7zTtxoe0ZgTZcGe2+Kn/TOhPfv7kxMEUqJZh5xNfFDUg49v
AKSObUvqqAqE9JqZFFzX5lnHD7sJE/4DJpTCsgNp07eRhQX7LaVFlRiSNu79lFAedv1hnV0cMUo9
XUa83x1q9HV6/z0WIYTMZMDDIy96taNnYTatDBg9l8y37CfVLTkCMukm3SWPcubx2Q2dgtC5r46w
aE9vkh1pZgWhDh+fBjJnqNGFmQ0wN66Mm+Y3oRxuXjDb8/xfiTtVxEW4FN04HfjfI6LzEug9VPqI
8lEzAGI3nEhLVqUSxbHvDDO2sJ2WTZW970qD7Hnq9S/HAvNbFye/H/9r5FYIanhUMXJrfGGjLt4b
9wLMuwqHIorG3NpQpcg8uxnb3r5ktE8Qg6FhVWBAPs3kZYhtLN+XAN3LP5BCDZsDCkPZ17TS3aql
ul0SFDjBXiUaPoepDkuJ+my6cqcI0uAasUWjr23Ewc7xh2hhgStAlOrw21Yg5caHL71QJORU0m6O
zRAJmZFgL9tMS6EiB/S6+umaS/gQWvzQi3RKYQOgGn98nt5xL0TLcu9LfuFPhhZCv+gtDCIxoWCo
a/oNUcRS3Q0JFxt4+jIKeD/ZUkLrdQdDXV8pEPE3pmVXZEP1DzWMdBu2Y743F1kOo9ZD8+CaSdfW
OHOZV9P2ckQsBujm/ZXD9JTBV5X0T2DP3/bB8I0HoQZvHv7QyV8VzT34wp621Vt62fIQ1AwzF/x0
bkPmaev6LpNbNEgukv/YMl/C2acp+1Vx6yo+bZqKZlgD5ut22J5ZrbMn3TB1+waIAImmVND1GKjB
mzhmNHlgYJNN0lAcYnMeNkOQ7OV1i3RJiHoMZGlHZNjg3N8B3gHeK034EIS50vdAWc0uVTaaL7S5
4OnFoPwEH4cRYTs4C2qaEn7lWLw39CU7Hmz6Rp2l4d1TaE4sV5Ab088rvCAdbPvcU6/EvCOgTDCR
6F1D2I24usqtKUl1F4t+Qq1wTnT3TGsd1GwPrTPMFnmIIhEY2H8WmgnbZRzVWidQBTAz9wCeH27i
D/GmJLXXWctt1tmqlwlY/yum7y44uYBpgBaR9oAghu2sZyO6Pf/9TQyYMDiKWY9HuYoiOeDc0VPM
EfJNAMzou/cThAyKWrIonXy2JX2NvOXEjZaJWYHXuscBOA3ypgG8eY4gacgW5YgPA+joGxRwg4Eq
fVa3bY1RxZaWoH82W6r/L4+4zYtMUopM7FYmGw+MLEhuiUWPc6bv4zYmxUjKCoF02N0nmuSzl563
pf7R9dZxTzVAaKzxMfgIkdS5vTL5iK7br6IGIqd32OU0ad1w3NH15YoPIDdM7TISs8YBCCJegHa8
07aEmg+QZkPm507QxQdjFG9EWuPqC0NVC7xdPlPSiVNvXJnGzQLXSbWQG53eJEDuW3eP5C81J8NF
m1/eKHpzmD7IUopUZdKevzCOCyCn5TyTHqdWAUuuVV8GYuIAREK7Y7eZMoYZL1zJ5dQBssFCIOSz
NoqWujB7PGvMTOQwyQAhk/G4fStYnaX3Q7/Y/IquKGo9ag46OyFH7p7zymeYIKFZ2YuWdXNf2Ex2
r6PO99SJnIhG0YYfexuhXQ5xnAMVkhhgfuwaC2uA0xDkk7eQ6nW9EzXa2M2boFmzLMc4D0XRbowF
VBRSoyzEdjhqDouXeZzcNJ6dxw7he7laAhn61Ntut15hHzkMSXQDroJmitdpoqhEM+G9LTgSIsGI
oG4y4DyU49UuemHzD5xigo2mtj2Jhmkku0pcSNqA/4FgxAkAz0yeOSP+kqtWYIdwyudhZsUy9o5X
npvM++jV7OnLwjVJ0QNpYUpzw2PztZcHeGnUwusckuq7g/pE3LoaZ7xaiHtp9nmOtv7CWENVdRwp
Y0yI53XuGDB6k6D3RZse7nQptxGqq0DFflK5cIcxUL6SEp0W10nND5ZVRyyGFSig+7GWtF8yztTo
PsE3GAPOXImqgRIm2g8OMnhRyveZ3t6EReWiKgXIk+3S54zbiU+u+3EOH/GZheiHJ+NjIaraM6ME
dhGljPLE7GmhKtxfIHoMe72jIlgdNexcgVE29nAcdONeMnlaiS8X0txXaLAxgHHZSOCiQDQSw7Pu
oigx56VgQiIXu8Iti+WIUZPLsonFXaH+b8OvfLd1ROdDl+QCZphxTy2x2f5reOZq4c6FurZXBbJ3
SRJ2xRE5QywqkDneHdGcZay658ThygVdl9aYzo377nptRZfWHYR7Q2KOjQR/UVEpJZ96sfQI06+A
/D+zx3Q3rVfrKiX/MR6TKc3ZeB9ENi8iRjR7JbTiVRepVvTdI5DsyZkJVPHnrmnUBzyjUKshbCEQ
hWgbYfq5R2UgSIi84wyDcZtvkgWYSNLtQ+Suw88kNj9YBFNiM+1cGMK3fIr1DcAwFCKKDU8lFkdR
80rwzRtuIPm0ZYb+reJwZfEzYVhzxfnxPZJWU4jJfWPPmbC4d6B+vM066NttT7ZZM8exBOsf3zX1
j+tygFTfXBlvNqs4RgSaePTuQkkTCBDsOP1c/fLvKtmOIJiZLiJz7Q8tK/FsBtmc20CBPiMihZrH
ad04Uj+j83kaPKTzGK7oitUp62jiQnQIX1dXTy+8bt28WHT1s8jMM956xbQ2hR/CUMFloV4cRyMo
HeEG3npPvA2R9B9Roh+UayNVEyR7I5zjsp9YNiVTqHCPzjOb9cYV7xRpnvzbhe9FFRSbD81CGPiL
UASPiU6E1wkpu7saiMZdVX3By6F8Zv+GE7JpKGgYERgdKztQvZYuUGyZzKIrqOmv/qmOYlokB7oC
QA3GegpmNdMV48/U7C9VLaLErCvlyTlTsbNiipWqJyn74+cjOPebSt9XAVK5OGlqp3Lv0ADfmYdy
StD7GTOnwad15AirtIKuqk/SqBwyunUv3m5pL3Gb4wP0AIplIlxB77k9GnUxuF2eLDxTa5jTPS+U
BfspoLEopV98GNGJ8Tvhnb8sz4lv/KH/ewDnC9BoQZ8ZA+rHlOp66q4R7gXvxyJTkLynVA/FkTbz
q0S9UjRrT6h++Nwyky7T2E9ZEA27KxnnRStqEB6Q3ALfneFWVjlCrIHviR2NMN0pYrCxXcs4iZAn
lEEVE0xQGXFWpmsMhh/paedJAnkkpNjgj543Zcqu0pfwWgRiFCxo3C0gjz+KPc1er2pNTJHwwl14
vesq961rSPgr3VuXJ44i2M6pmi8+XXsTBaV7vNaxlMDvGb8042OQVh9RVSLJamXDYc+47WVd/V90
c7pnO8bFEkqAYoB96QDzWcJVb0AcYS6GyW+cR11WOvyDm1jMEFKKYV8mfv9OnmJNEfcfdhX2j5C5
MnoCSK0DYJAXtdGXp4LcHKVQi6Ev5OMAKoJHm2DxYW52mGVzmKxRDQMAJLSBeMoe34D1q8zX6gvc
9z8pKhdGVGo+BkZ8sd9PRalZh4y3d90q9qnMF3fbuzKSiUaq1+n4mCxpXRI1IZUFHfKtEZtkZds+
rfOeF7EvE8/ijGCy9a74XuwUfxqe3MMGhLgoIQrUiPPcRQtrysgj+CLdFxEcHGQF4pRfgcWkrt3p
P3ZRcTUDUhmgSHD7DFf3qhKezlxshX9IGeCNChyb+ndEOW6rDKxFnqmTsuRQiNKA+N6jhUZspGsj
RHQpH9ZA2tqnMTnxaCim25fSnkkoyuvFR5uHCL4q8IBla9ohA1uQ+7lsxS4mKVr3g7eWSCcJLoJ4
oFr2xfd1VqxdMaJYCzFXyZd/qSirBIeBPyO87FDLNcqkgxrR0yC9BKOus1SHvTvWuBaVwFqwp7pY
nH6f/8qiwPYgvWP+qC+m1zgXVp61LNIHi/rC0l6vUnCLthsNH/7Bd3lKGjCaP18knceLtdzYra9I
HRkd1ct6d91vRaTBlBz2UTVSBeO38jWKApWPBrTeCRV4uEh3kRCJPliTHh5exo+05YTimErBjy+e
Z5rhd1lVintlBqr+v9sFLZvA1f1LNXVvrBbSpI+iplsuyGZknqnTLSowDV3KEgcMclKCYGkYy5cX
aOdztIepg+ZQZtlS0nBqVsmZu+UHGeetCqjASO1TAk73Jssp4I1kdvDiFlxfltE7v/p4XQj2xSU6
wRjixfUIlQKf94Ud6Y8H1cgmd4Vm2/VYD//LxOmddzigDhTARSmzrTtrVCY3K8YKGsZpASEAZ7fY
4Wys8OBj/Y1x4e9P1xPoMoooXrg6tnx43V5hqjzjyrerT1XGqvdWGguV59NelJjwPiK744GBJuv3
MXmf0/sXBVlpfqE6nR6lwTJ3cUAWWQvTYfcCbcfm5ctY3wahMEFqWYt4ozaJgmsxjUa7902P6kXx
nqMwi+sa6Lw6jTRhPa/3wiMYoubpTg8dBoVZAfivrLicfxfIVB0qtKQp5zQMPDQ2oypOOcTLeMl2
JJ3bLWVUfxZLQC6MlCtbfhrme9xqBu/cRsq+hl9ujwK3Zuppyv+35Phsy6OlxZEhQQGaIZ5uIx9N
z29ZJmcdKQ92YAiOtCVNfAPdEovwHaexVzdM0AiZD1VJNT7+kVpMyVzAuGJ/P6eOMw8eyPbxFhsp
RNDSe5GytOpYNzmCbh+aLqc0IHW3fwyVouhEsbLsR9H9VJBzrEW69l0c/Pi5fx1RITvlJndXexqG
wqdZRWTNUMukOXT8xV+ZHMivANKiblsgJqRCv0Mo4tIOtRQYSNCuiTyQG27P3er6KVug/jAsLKHZ
ErKkC9xIlCMOh9fgnM0HPA6AJgLFijMLYx1F7fGBtb+J2Et0ZB1ZorK1mFdJacwEoA6n729QZa2B
/UMpnh1/SXJ67+JnfZbnmWTIXucz4iau+i77e9AXPCLcgCzlIwgOMKlrdUSOIj0d2jPM+OeUCe+Z
0CfiKqenzs6yCFDX9mS6HxesRLNHzMh4KZVQuZNCICYTWim4BaiVQ85tuXUlw14zKUnhsMJePn8k
F5xVNimoD9CMCJWSDgYPRtI24aAVCpFzdFYnEptwowUF6bhwND+qX1v+m4IZwWQQNoCsrsuKfmIL
U/RDVNCjalcMywnE5kQe7pLNj//Sc1Dt0dcxjN4EN4s7uGn+vHB3Y0NCLeflAlTDwOMgtzKhYD3c
Hz9px4rY1my2PvBIMKRjBiZifsmMvyRNi6Ubocdxoem0hGv9AHKxDBfqmL/sMOdKQPiwFic1x7UR
VbJ+d1elhmFH6TgqG+gCVEH8JV/tde68tj6vb5mnkyv2qZvB32AuP7Ixo80yeFWNtIxLYMKYw73H
JAvm+CJ696BJ5BKxPKjTr37zInRYoGvaF3KY6vLWJN1fzfs60/7PkDQLBJ0g07FZkDHvpn4iB3WI
f+czIlygh1H5H/T3RfERcUzFuHBhs1aIvZwW/JyLlMEYzMiyaakI/mgBohvBq4l+mqOQbmpoaV8V
Atgw48nvtWL8EqP9LzERryyWsk5NyYT3yoaCeh/p6RILaxDifZUY6p54bblUM1MKusDd7MHqz34X
N52QH3MNUTvWAuh/FQyW8LNJ8Fw1BjphQKEnPdYuoTZ8/91kcwC1kCvBvjL/Cjy1GdV9Ugu/Zw6B
ochkDzFJhViwqTTV/w955IckgIiKRQYNFQoQ5rVQ1zF3BBuvKROVeHyALE0jYIKqucQRR/t/0Owd
0MwQykyyuWgpFWoe8YcXDvyQvEyk1oDFNjPCArCIhUfczgH88ztE5RMrYLsCZVT/u8f9ZtjUzkG6
Z6OUqYiMQgZ39zEUekijfc2N0FDB+wzCajVLZrtlDSmggcX8sIwQBMqVPqM8b8qLAWNP4lJaDTys
I/GUghZPLU7Fb+UOXBmhSfdJMU5Q5Jth64TVTnMbpFmOQTaKGamM5Ny0mkixZS4YU0owymTIvTl+
lVCIy32aAEx0ifFjObUwRGK2ua5irfIrW6YjYxHJEV9lpRHeiJELGUYdWhBEWnLyyZ7mZ7wsc//k
oDpXv5Voc2dypr7IxMz0JV9ZmZfaU2PlPxe+RwuYF6nvGm1dxY8dz8adzqOn0yz5aW1P1p9VcUrT
bXSdjKIR8xY5/Jvefefc5DYiOmM3mEMK8Y9SOTMdcPgsnurd54fF+vtdjjmLqOE7MMbvqXeKxzzH
aX155EamAdavAgGX6BHQqL+4q4p2NifHyi1+Pj1+n3mF1FXWfKejrlzFuPbgWEdGE1/CRiVFO2/5
LBbcFXTcoiWNWGusQazrd1hknHQZb4kJ6qxven7r8ZA3otU+XR1UGXtDpZXhbZ//n2NsbYzMFDmd
zkzT9H6ZHBVhj//CaNEg/W5raXvz12CD0FFtwoEjrCCPSDQ72m1pdyMoXpAPeJRnWoO3Udjib0oI
hoGF3eLypp/Y4ey0JJyQFZJ+1rFymAhlF/cIDCNAPCX1Xk97XdhxPE77q323HlleDtIADk4om0CT
gSKzaP+3g3cVw3lPs4pG8oFPfnvZytW+KUQEA2FwFZC3glvy2kmmgPjkcAnvZqj6m/BCpKEBkXNb
yQm/opaXdj/8VQ+vva5kK+1cpzCB7YHZ5HgcYCOXd8qS8RB5rrNZzwpDtlbxp72+7uckaAZ9fgzN
fv8htO2vo8zRRQpbSlsJZWN22nBbTGkhEmcpaCdc3zmUPHrA1tYlbGBz4dCZsdb5oJd/4uSTpl31
r2cf26bffxBhl7AikmOOB5nXP4YEcPlybx4O2hUG4Aso30hsRsB+eDyfWBMtdYY1tV5Q62DiBsRg
AAXZoBkuDgzq7vlxpfIeYlOEVcRSiPhiAwP8ufHH/KuWkDGrELGUw9U4GAC+qilLptBlLH3ojoDh
OTh5f1WC0cU7urYHsRnaukFHJWz2ABcycmC82+5zc6nsbLVbPNKmdorAQZPTmxJGuewHizi7o+Qn
bfCqqNLF/XEQe5bW5ku99genJfkajzUDrLjjU2Bl1BOiZUNpqfBfl8UMSBVRUwGgOSIBcftUoXHM
Qzj1yspy1lTYj9N5s0VLWvjz22gxbOkt9dwDUU3oZ7pvdMyJnmaAu/Pie1Dc2AYP6uVNXZbYWuPr
pyxv19LkJWDZy5Bcf47WkgzHv/ixKpXwnOiTkE4UjiMBuM/xKXKPzCz2N9TlNmA1d1rRnqnqKZ3y
YQzIUQAbyb132HcGYz8C0HJeKYJPuJK+AF/llnDbrVhRM6p3mhZ2pJ/J+CNDBTFKH+UytEsdyDLF
c2xK8EO+HvMXnSsvp5tHdLgXzMGrjUQBgovJqzQvcQt9tHF2JxZpHkoaE+s4X2cTgpE7acWQrYn4
Sy61IVxVcUTEBrKJpb+D774YojGGbjleUKTzs4WjZcFTU9H6pr+r9wBBJRwUtz/MgWeCdIUpg38f
SAHO2QeKCkVSG9zlD2qGu4K7j8jV5QC4LmDzdxGFjVHCfCXOgjajDT+O/kYcJVIecWqe9pp03iKX
MVKMkuf+3K2RV77ektz3EXGmrIRmPkWLgtHT3MEGxr2twqMOqmyTJjfwJobIb6HvdOtnpU8Qz3DV
arfY86mif/QXsRAX3wyAmVNL0W5QBxDhe8xqaklXMNQ7yw8kFWQlysPPxvWOL738b8lWfbxRn1/v
EkAuf5TnsJEagckfCCBeD1bYHzayvqi4vmGzguUlExjSu3x7/qCIS+swHG2SL3VuODnd1cZGMRkO
ofGQjX1Omd2pOt9mViBD0+1xOL6Jx5isgm5KlQ7GuCBiaoXQhuGddD2hLY/fXT9eWhqmLReOdZL1
iNsbww4STx5iV+3Ih92OyJLubedpE1J9Wxn5qF36tOrtw8M2maxwY7Vui3Zs2+TFY0nEq8Cf29UN
W99f+C4YstkovaqZ+c6h2f6zRe3wo0dlYUBaK/4XG8DEEadEPr/avRzWeNbTF4zU85cekakawcV+
lezdylacbaVDrBA+yUliZfL3gtp6jk4xRKOvlP7CS2CNEHbUL77dScDyHIfwphwrAQiwRS/0Palx
1GdnLt/A92BlAe69t58kHvUwqFW1lRBZaPu/rzqHbm8ZxroPBTSW8itueqbRx/xjeJnJO+6kYy01
MBwZk68huJyuvUqpGEHsx03UOg7GVEqIRfD5vbw50YA6z1XHN/2FoIJtFOl/37+g0ASVVYvl97Fr
YZc+z8yMHPbUy7SvvBTgVD1c5TMtQspPnVMVac0Ga2i6MjmLzvQLcX9Pk6uWQt7083G1qApwOaNv
sCi4FJN9zYyLv4CyjzZwoSWzyrNw3Zih8lMw81km7FuZsSbmAX5pB605Nh7bJc1EbKIfcYGAVa7R
qrwecrxGXU0lWx+RnQVxg7aUa9YQN5v9p6T9G1u8lxEaQT1ilCnHrLaCwauQVrduOtsIyf9EQoTt
mj330t8jh19Yb5WVSWKPGkSY7LpffRsO4RJ/U34bbSV6Hr4mNdaVKU4T+HvoqXLeTuZtzz9iCn9c
ZXiv4JqkepBhVxBfez73hGiSvdFUd5Q+8l3EmKQCDXIXXxlALAD+plKdWQnSHMaJz2VKwOYmUxkm
NeZ5qOrSP7Qd8OmlFhpLX56KGVsYdRZjf7sNW0iF7Z9czDlRYyrN0lfKPG+DGWlmhdoXHadwynFZ
RFhMX73w+t/0qnrz1fq+rgNYg2K3gkqeVBCUxULCw6M8uYdcBoHHg7e32GEO5Z5XHuJ2DxgBqTs0
Whk7FeN4W4lWUkfeKF/YSCXbxY3nlbYGKQX6XCXfudPZW6Ui6I3rxlf2sas/C+WauAJ8+/Bc4gmI
E+R+7wuLs67ZHeitqdpB8TvxELpxt3hCk6juxbNhAJTem8zDM1Uuz3qxM0YdpZxKjNlXG27GnFln
RaImcPyYnTkRKeaunWvJ/h2TUkTjggLcQ3Iqj8A0tJ99r2QOxH3+IXp/jtdBZnTaXfbkxVG4xsdx
tirPC7cXiuVzbytkz8Jzi7H3I1k9a0hWdtTbkbWI4bzWWy19PNzQNjpuvcbsVk8TjbKQOszSarMD
qMYwn4NglLK6Q0dMVYyy6g30nnleVlq+nDiaSX7ig/I1+SSNN6A47DaCI53K836jtULcRww5+a5b
0ICTtzuJx0B7e18KxqJQTbj+Kp1Zj57hUJHNah2aVLgcTXZiYn70X+76CYV1fZEx/eVV42/cP6h4
lJpH7jsLSgOFzYxKXcfLq7d8x606pPwTo71DnBylLOuNyMMDv9k3rQiaw7EzuGLd57oibdmxh54m
tzU330DKv6kOpmIHz0QAcVZ2VmqfYDpHKmZJwswTIv/+3ZKrpcQiDemjMAKmVvhz8kBd5cxJeFhA
x8HDYMwn9QDh0NpFEyY3sJPJIuzk6b0NHeiuqhKtiS6H0pk3css5QjzYLSlqr82Wv1hDvXRVPvJa
6C7BPl8WmaKQLo0y56HM1iZZPHDZBJxf9GiQ3X4j9XKuTtyxv/oF++dRDvXUoyclPKyfuCBM87JC
7Lj7f9U5AiAa6mG9L3dJfm7PYsE/uLHDB2BHEqEsT6YZHp208u4sYFw6pg6RaxpVpB5fdT78MRrg
iY64l2jhKXdprXNZFf9+hTdqWwcsfyLivyVnYRirPNzFLMlup9Vhyn2zZECjpDv/LjWapGaKjT4l
D2hRHViyf5P50fcnTy7rJWd16/kw0Xn8upiLo+jfG5MZjkQdzEXPBdWxdbYA7YL+fBwVGnzmqI26
eARwpYXIfaKQGas/iHn7LDwJlUahxlzT2FNrx1YTtwR6RqKSs+/cY9tap/D1njCEQRRCqxuAuzQs
ZH0gjpBNGveDDfKRhJazDicnokL5nu9X134eWeQ/It4pk7MFzgloeHf0MgoySmrisTBTr7XwHHw5
ZBPwDRbJUUQfbzzGD6/kHrxfkGSJDUzcRlQWsk7Hj8dOenFYNGjtRaXJPzJjrWkBFJtX9m3cLJYS
dsotRimLKQl+7qdbrd0u/qCJJgct9fD23CboKt3jceQc8D8nrmyKTqmTfLBsQesF+JInstz2Uyqk
o2j/uDF5a/al9E6vV7wgUqYkZDHEAOtFbK9I7N9E02Xa+L+nf+Ru1OZEDTb8GTqQzbA4QJqcsI/c
x/K383oeHtZnLTjtQpMGHjc/Ks/K8Iy1Rj1Ge19wgHw//dMRFdCbxb5xr3OoHWxLa2l7SNVKg24q
Ttjzobe6WCq4ahuzApc9JS3EAD0sV1fmCO8yUSz+pmvSGcqiT87m904lUr1TwWvuIfr2IlgIzCr3
mhN8zCWOQsflHUOBn2bCy7EfP/NUYrElfJaqGdeqV6ffQI7B2zWC62djTlq8QQ6yvv/K3OBE0WYc
O2Jbv0y27vN3vT1kIXdK1UEmGtL1v+9nEXH+V0e3WtFsG2yWFMT+MezFNOSKZgfRofcyRRPtcBkt
Tvw80TQ6rC73mN5hgWnlVl70J+PwzX+o/yvPRLHjDzhxlUmXke8+puGp8P56cKIOnVBg76GLpsSk
Ibl+EhuDQcu1LPPs9E1WaBvv5idoxl8I06jJAos1/wB7Ut0R4eo975S0JeABUWyr+Aisk3X4kI2D
6xmSDDVtR0G7AdvS2sd3CJqaRkiQQ6M1V2rbSvPL+c+2VZDQkZD/e2GMS/OCIfEg/BSgAI+GmIzO
b1nCGzbCBY78XqTJVmFlTaCeefFDwa1vgKsS472XYGbk5YGpdyjn5XO87C3bNQ3lNtFZbfSkqyZE
tyIVbcH/CVEQHykV3J4YkmjaSlNaD+AA/vVLqHswJCTyl4SW4ZIPNHI+e0l1hvFKeJua9/49sEB/
vJuMkS2wEEV2kGLjp3qNAsOnGeyQRoxAQNDGFhMB4qug2lZIWR7mdgW5EYmwGP/UZbk9lRAoRutm
962Qk9UQ0T46Nmky/ECedkFtwOAh8MaWxqCYSkA3zEDPq73S6QcKMU05bGJxoJcAqd+cbvRHzv9G
vt085h1pYLf1IsoWRGGNm6RsbN3PxgwYiSWzDdSIOVTI+Zmk1lOLCqxBICYsSgWb5Wy5DUnh0top
cM1Q0KHizbF7Ho/5hYw8JTglQIj9k/H7gjZjt+9bLK0nHPfLydxSA7Zq8XSFsYsjGVJVJ8hkMZhI
xjOicg2+Gu1dhyz6vhNyXtCrByqZaAPFEO1nfmPX8LcSNqcCdnbzyykjEj6TsvK80hTWJCCfYd6O
r+UHgNYnuzDtcXtaFV4Hf05w82IoNgYxPKEgTRmr//6bgz6oaZMEuPqtkzkil6cKFROte1907Z60
vGt/Lv3tuDqfPf37PWmxR0gv0RALMSQxWI/lxVYKiEgS1dlmdem0qkhKAQdAMu6+pwn3BJBkQliP
W2PukdERyA7J9HZ+erHYBcGn2gb/ERbovmvon5ztaDMpn2klUHSf7U4W1P9gfGahWMe0fGn8XtjX
tIXwsoqpydFsKAFxraTuLgBYx4ynJ9vdXEFOyz/OMFXHHcTo4spdR54gtTMD9I702TEcZEbzfBEy
fEGEEn9SGXe/2yky9rDQNvYO+rN5/VOP5/5iaO20OUBcgaGSMVlG+lH8lW7fdaoaZQi9N4DbzMPP
ywnst/VOxd4lvacXj27lqeeIDoJPDSBsadAPkUhPhOZ1LnJXqfVhX5y2GGRsf4tfDixQRjZOMaMD
JNw9sAzpBvYlEJC1LUji/blOKs+P2jgYvBs5SepP21aYO0lcUfcZKmEanyFpsUOxXnw1j7HVTkym
arASWXI2DZR5GlbYsr+GKeWOSWm0Xj28nteFunqUYxOEWVJACO3QYDXhIYTftkZJDPafVATPigxw
RVYjENXa3PM7ypaUubnDICyUV0JX2+Uu55/ghR5R57s5DKkOezO8/tyMa72m97+Xpl11WVblEUhE
WbdackMQRbuvkFuEW/+DY50TgJZdRIKFflYkuW0TGDM9V3hf07kv3xiUGTkY4SGtFwxPu3tW7Vm2
Qg7o1GsJ7aTnWoFB8ZpOMkMChZ8FGekznzwZ6+IJk0UTxtl8aClPG2YU1SefDk7xHyb0xAoCsWeP
yNId3FqbD1mKXyo/qL3Cdmls+7mXkKjmO2yLsCqhK6W4trkOeKqh/P4O/RvtLaUMIaG7cj3+PQn0
XrLbO9iYtEmjSBkDecZZ3FbWt5piB3cOpQye1eTqgu9NyA/GoeynaX59xLyKRDUCYeScLXoJKtiN
ZrdpSqGIcNBMpUdot1IMZnEJBA+Fx+MTvjhbam5OQkc6lfmC8w54P7uIsoxvsR2BJyWQYDqmBKj+
+xuN8rOxJbNRBCShw/xr+Y1UdHE3aparv49Xd3dP7PeGGHpJO4HJZl9SpyRhF/8nkputAZ0fcLdc
hIpwkVjOPny91xPvoTdcSSLb7m1YGLl2ZkfbYzpXF1Iz84RIshDZdFXZbqpNjLXG5S/IHrHabix6
xOs7nVfsa8iRAzVrHp6tv7azjmlZ3Q7A3XNKtjpkykNeA2pcE3u1JcE82vTAEqtvKs+5zEnjS6af
viJZ3yOQA44jgXNkQO/P78KPkwOPrDGio8AY7IzpKUYQBc1LthjcuIE44tkDDQHzCITnGT77ErTt
j6Jp+7AVR2T48W0WGeHlmvyEW96Hpn9tdHktt6dDNYOL1auqaMWtPH6Z1E6/Zd8mtWSCQPzANkMH
rMpqUiDAkNeVMYBQOERXgIBFvYgHPESkSX02PaBF53X2xNuX6AeqcQqh79x9Owk5+4YPdn880YeL
MgH1RenpMg2Bw5S2zmiH8wnomQ69NQtXSOIjhn78MFZZrd2hm5D8n5R7hcYiK9WJ5Tfxvs035Knt
Kc9qeUCN7kbtFM0LJutPUA0QauCW1g7Q5+8IkZQVOeEEjlQsKhoDe2D4cVWedNiPi0139gaw8t1C
Yy9AdXq87/lddvDo+fbfsgoHPqxTwC/5fex4hp9CIpDEP0P8M2+lzbqxFD9dpWYVRWhpA+q8gEyq
Mv3itf0zI2EiFwgZiSIz9VY0wzGp2a5hhGVyz4byMWDxDIesn93K7rjNrN0cbd4eztd5jDZ38EeZ
yNDmjiEwvsJQT/84uQ/wwqbDKb4Z9jAkSzG63HSll+Cv92g27sF6iy8KKgvuaYXlEx2MCQGhZvDs
TRNm+PCajT8EhvEHXHiZo1bLloNNoiCN3/Mem4oJe/qe9hiYODAvx7dN3r0S7tyJF09Mn+TQgYR9
23Rz+85f8qesYdE4fA+p9VEEGGtoAFnGaoYErfJqXXonmEfhCdD3Isp+rEpcbMLvjJd/s77gehF2
/mtvAXhTDy4SmCK4RittFMfDOdj8fezoxBQlOhuqkqQqctThJIx9rQVFn/nLfduUVHlor6VL22Ap
qMOfGH8s63cDutWXzximUurkupf+bxYGw2dmzx+/7vMewdR/pbx3y1G70JCNakMwhuVa5Z2K7uwl
TbTROfnCZWNCwf5OqSX4DhavK8SLyrYUeMbwYEQXqPvaS5QJFy3xggqLcMA5bMK4+yzIPbag6olC
XKzs/jLiCKsmMcwPgmfdlIdZvBDuiwozAw8eVYhKBnYKle6pbYW7PzvGo4gDnlhvODtTcyXNP3Ds
D4tioo3DEsRhmQ7npxkfqWgPIqaB1yjH3jYJ7J9pLOdBsIMJ26I/uTw8TdExiC75WdETFiKbd2Yl
VNuqEgICnq0Xd7lH/ec8yrlZ5G/HWA+Mtr4LQQZ8J4ZhXaLMCT6+esf3BoJHoEu5fAqv8MD0md5K
NoPJ/TS3z67zuelfE/ltzbyyLYN3Nk3/3nzd+Rf7ORg6UuUPF9UDPOxpJdY8Ovr72o4F03wtZig8
EA01+jdGAAu35oMFM2OrCdeX6IJRvR9a5iqQwMC2H28RCNc30lIzGgxRGWHQBaxOnvIenCwhQxlJ
QzUr2NhJHsGC4KHraIgJjGAWc4A6JfjeBwdGcCFAz2ad54bqGUvxTzdU7E3Ut9e+K1K+90dP+rir
CuRdLLY8SJfPIIAW+EHD90W3dS28TyRW71uUUwIxGoPuDtXgFQAITdBCTXMVfr0PYHY6FrJv4pLJ
VfSM1kJwYn0d0k6IMZgbwY45zG3kk9E1P1L9oSAAD68RgqxVcuGYsOHFyb48uxjcus+TiBElWvNN
X/toOakZCCUSULIWVzYmRY0pj/K3Yhrjq17HQPiJHMPMiK/BQ/MKgjeVm34GqrgoGlF3m4X5EDe5
Cofc/TD36l/eZL76yVeJpP3jBtkuN6aDm71kztGEwf4CMKRU/AU7MaVCl9qPb88/zaRVEgT+8BeF
EPZtGBmvn10OEStNOnhnGhX3lOf/oqdhkVFLHSd2p8KfhKSnA0Xb4W3qjLoVgoy+9UoJLebWg2v1
DhN2mXMay1M+MZHhbOs8RFsjWpLdDXLSvAFg6af0Xk3y7FJrgxUqAYnfCoJl3j1Sflkf7phlhPSB
Sg+TmwnPY+FwF9dksZ7yd+EpEkwtctir/hbY3hXMXzCCk0pBNRy8y1yk1AHuaJZmjVv+61WqFWFF
vFRvrYOQBCYdEElX8K0Gcb3e5pPXTCf+m4kZlk14BgR5njjsxN0OjHnY8NahavOVa47St4YFFBwy
c+UAEKUtO3FBAQJX0OQwdOF3s5HH61Y2Z4n53PJRPbRjpWEpqeYN1cYme3XCweaQGzIfEg+K/McV
4ov9S6rOmTS7gZimJDyOr+xpeiKJlQXRb6vmX3fgQx/2VcSbPYkyxhYpFtlni16BowGed3x+30bf
ad7e8PaWj19oNW6tvooEiAYsbwbTZAj5IMQWQWqNNtiGbqbt24U5XEugmbrkM/SjDXJaOAzk04Fi
NWBYNFupEt4mf8jj8OzzOGY/B4JCmpPqAVTTiCOE/MNY4ojiNwdGx/dvz4Y20PA0lgMxo5U3cbs5
xtI8gZPWsxtV4DR+ehqCPcegqScRIpv5o/WX/GKpVhMjTmOZo79yryzqeVcAJ5utv+KdZCxf7LHP
8IsmmDqVDIq4QgDQxW0IsD6cxeYZlPJR8F1o/849/IAqzVHS0ng/YhsfllAGxFqgMQLxhSwI/1PG
0seYJKu3Zwd3KpbjPcfUZyJ/hSFH5Q5jzkfUq35SsCD3+dug7q6rr7C/CsmJ7OiXq6uYAC0lGiwr
MYPha8C9LucdfjfdlIKxVrdsHCsytOhdVuVtruM+A0p/9/X7aq8UfQp/dWuVEoM8Zf5cgsq2SCO0
WIbgNg2/j/NTgVaJU0KB00r05tcwoeBEgqmyH1ioKad1A5DUV+peefqr/f14Yh6tN3uczGmjzRcY
iCaX09IQPmhuXKhM3q5TX3fwxL6RbVig2+eSeP0G2EF0xUtfJAOJ4hUGqKuHVkQwUyllZiXLTU3D
w6FD/6hQ61KtjI/zSFPcZFon0+AznS+w6wue7ToxcCK2BCIOFD//CCMpoh2SknDV16PElaXZKe+X
VP6k0d1cEkkmT44BgTOpmJnuGWAC85eyg4gNvrC+v2hz9h+MjIg5TLdmybwMpTIGsQ054p9VvFv6
f38J9OBFKZzZmi9CYUXMjbWiERTeZSeFFy8P3bsja7CrjxTDDVWTj0FRIuHY9lyYyGSJLgSaurF+
fy0xw3cyM9k1G8xVqHFRP2oiZpFR1jLqDxyB9J6FkGL1f2CPHmjM3MKNoRWXD9QwjEx5t3/9/3Sd
42jwPDpDMGzhAslLQz/P+Qsjki2OuhfenwVherGKGlQ1Ig0vjKBoNmFszyHkbVPlr9ep57+V9VII
bx/ai0whjPkKHpD5p1XqotCJNlTXysK/AstfEXIkwnQadNj5X8WLpxY6P2BDLU26ttcD59D1iHJE
NAlqmwlPlJYtZZgU/KMCtaQ95hi1BQgFOJRfYw+pDmsjw8m8dW5zYNko6oubMUm7t3hWxTM4q0wp
hfGjCxjpT1KtL4LQPMrgImSRSRGfk+xmM/Vz7aAaocovTQWhtm5eUAtixN4xZdi2dhM7/TUUA8g6
Xmr1bWoCqyAmPHrrGeDtbLIt6q/A1z+fIj1KPkCOueFbU76arQxaDvuGawz/Q3lwIl+LgFtdfRDK
uvPE7dVcgVrBBrelXc2A0PHh5AwuHpYDZq9Ukulqrzkiff5TfR1EMjoVRsCR4283HnBUJBNsA91T
TlSJ4/Pojq4xnilpQa9eGzxzrClEX2QcuWXOeqOmyvnhFHroqbgNbGN42Fja9A6KOMnDuWE5QiMb
Hi5uCa0rd2GO/75QQfyTFT59DvZv7qP55sedoMFXhNysGvefFoKStdqa8/RubJ5DAh3eMLrqt7R2
8LViAnolqI3TXt5jFteMIVzQV8hAxq2wGMNuhebzPFz762upJaiaibeeRJPkMxx+2prvmmMinf58
kLLNPnFovlbZdW5wylq6Eb4j2V6zmn+Cdn2I3HGcil4NCfsgJIwIjhxUhLrIiytxjFesh0KZhGij
lU/fjIOfOG7yabibCMWaSCRrVAImfqbvCo2lgoZy981HZqp+vPRY1GVMPBayzg9Lwsvi6jXP2tlE
GPbp+jWr4urIFj28KosiKlhBLMir1g0/m86V7OZFYDU7vqWKqHxYneX3YiFn3sLk/xR1BpEZ2Yq5
nC6TGyyaQgio9NNgmcDFPO84aF4G+YteY0bh4XSzv05izD6YZEVBKpKyyCO27jdu7Xp3RMHNclS6
WahjeIiXLmBjAR75tCRoboeuqg4yfc+wNg2RoRUd0L1nU1cDYUsJXFDHFz1mFlTnicve73qRxLlU
7b1eJZEEasNEawdY/3fgA0XUAUhecz6sZs2dQ1vWogJSIuVAOqP+yyhg4wK06J5YadjXy/3sbGRn
szPgc/QZIEs2COEZTyE0G4ieImX1M9DdP48JNd7pC29Gzkr0Qu1WO1G/JjTA9fMeS4nZsvuxFJxD
i79VnlSZeNvw51njuIqHMkD0eK26Ek3gwdeDqFJIMlwVew6F8M8tonBhfrFPXHahg0juioEXsxqy
nmwz5XF3ygwOm0PTyK7pbpwl2AYl2gzKtbC00KL///o/ygBHqmcVU/KihZG73hFf+bZOxYnkRCe3
8c7hz2aSbw8UsagUCRemzuV2bnLfdfKinPs1Am1uu9EQRzgSw9bp3e4bjGuGO7djkWrhWSwR1mD0
EX/teLH3oMb6/ildb6znpQDWiI8qqt+heArYPZrvORV/qm+xZZm0kcIdNV6mg+JK8IgiQPyMeRJx
RXaVNzEGVdbtT9VUKTIFNCvAFPUl6r+hOVfWNMtlprRvnXha3hMLY7RDhZ92nJOMPHRS+4mNAx6Y
r9UEpXgY9/3vHaxMNf0V36ewMnruOrLVkGa2JjgNM/TY1RLld3nheWMs3ce1XNgE8QxmogMdftzN
yMQC63hWweXt2EQvMS0v14B7AYoZraMJICrKCTFx81yR9y0vD/m16q1Q8cVLd1F6wjF44HBerD+E
OIrlMGw4u1aMDzAfaTdZvr7esVlTRKFXkMMWZrZXZbybmfheL4hml6GfQGTEiOkz4SQH9qANXJK7
DSMlD/RwkPCA2AdYxpGobuKBLuhrWyfBTfx2XQ5EOsUiS6QKM0IG1U9Lso6zTmnj25CU8AGSranW
CSJSlycYdDDXD+axaQL3Bd3aQ83fiKwkPTYof3M7XzsylcCU6rlISjGkxfcbQTpbQQw3xgWRLX4L
P69UmyPxFypj3ukIf/HLEb5Ifk/FvJK7EO2IP91QHkSdvBTRmI1pZLVVDmI2+tJqWCTcY2eMUMO7
OESp1Lsqp2/XZUz80USlbEkCP494fhId2AiZeba2k2+kYmEuDoQUrrUA7TqLnSFHOs9g8hrd7Gtf
/VwdVYG5ncEEqdJOzWBkZaun8qNZ2RO6T6ANRHIEkEnLECfmrnNqtOI1BYkyexOS4xI9L7hnahgi
S28wASQj8PzZigzxAjyCEfK/Ru8tS2jeQUeqgORAbTGoaD71QRaiwODs/ELNQ1/mjKutgpvKLLNH
TycnFepncNCQvmVt5Gfw/gwQFEwCUGhQOP6AOTCrR7WRlnwMJkOhcBK5vPv5olYbLypLH1VrlgaM
utBnsY7HbNBzbIvxnWqCZ5BuNqe3nU61U/aydnyF45gEWwcAyTtb5OkyXV4Q5VtXdoX6tOpTPEs1
z6kSSP5i6pbd4NbZUEvcYCTgM+1alhwMlexK+uUCTDN9sPxhKixdPXCj27n2u0U4DCYKA60cKZwF
m7LkJ7fuVFkU2RQUpOp+KaPG8SzTyFZNBSAuWW3ln6P3BqkF9WoPck48S+RmdFQIAxxKBLauXTKj
xcK213LdKvIO8b84Uz0RnxPKdQFbR9FCrtsqp9oyTYReyd6n6uGOM3TuvXlZspAwFWgQqVC63jhs
WYLB8/5x79rUCjXgR4e4DrHUP8fVyLYbvPGjhRDyiriJFGtl8tUJJhRKHDC6h2YFTO5aklu3yGy+
c5J9A1f+QpGtS0VB4x+gw1qFfmZvENUsMNzOryr0oRv0M0YTVaxSPzpLbaiFrDR5BG2brEKtL5Y2
l+0pTpvcakS5xyX5WQSMfX9s4zuquWXCRAAr3/xfL0EA3kHd8lfletgK/Qg4/TGEXsJlEBDM8p7v
UhBBTxAhqaagLBJxHXQ3gBcmUlXn6IsMdQkPYJJrbnI0UITDHJoqt66+gBUhqimA14s+9KvNSUqL
Dut/HIKG7gQCh1RpK4m4I+0aWAcNo+k+MbhgpdtDMju/p/IoK/1mUm0B9D1lK4kHcClJtxsnaybS
Bi3kIo8sz60qNjGbS/j4Ub6QAxA8uQ7XH1XsLTppAYLA0+gTe1GT3C5FbbZ2JMPPlcKfgpdDTw2a
fpJ2cVo9uoaV0aPsaXwKwOmBZeANNjBHM3wZBf2aKhepNUYDnxkoqFudcQW5q0EX7VXy8u5tGaY/
nhDrceVc+Mw0R9mIYyJuoip1MVM6wJmRE6f03rWn8Echhzq6m9jUul8qm0RLq9jiimqnoPRvi/cY
EtuunwM/0qMbTdCcMiMblqbRdd/JZ4GvdPDv5L16HyKiYw6YilTG5G8Q5YCQXfcfGGbblbbeyaZP
mNSBl+HjjGkkjUl8yYx39FQ5g41KcacVhC655COM9VrnCDNwYHAKtJnTy4IWQ2UQjIqikGXY3q8C
V3P5WrQQY3HDns9Iax24jNaZH001hme2Tns7zkSKYZn0TfNkh+g7DWn5/on1s6AWuFv7/IVM6Lnz
cUCskhjh+MyLFI5jUtTY+vl0badrH67XO7KY3uOJYx+hC8npkHQJ1wxGjdeyy1TubAGQwQ9cDd5X
bCKAQNrIaSf/HnSjaaX0obQ9E4Pw8pO2l/vlaoS7htoc1K/4Bt/nngD8DqkvlC+dxLLTW/fQ3f88
NiJTT8DSuOBALmKiYu6tfF9Sxc7JNjLy/eHb6VutNe/b4u8StV3jIzh0Q6xt3VOR/iBvKu5AJnLn
QLNFH1gXEIeTvnw15DOqtzV1QjREoAeNtVvmcv1Abv7NwrPl+Mn3b5WFi5QDfjuK9+giwLKNRY4X
2sk0rs+6jzjqjmoVsYj+PVQIQB5B3F0w8/IA4jje9eLGF91RVFu234jONJR148zhdXUkMrMc9Z42
pEVFsH3pJ0uhLsI0+ifaTGwfXxLqiR2nQyK7UUJ1KxbhwlPO+7jVYgUq+RdPZLdszyMVqW3kCZlv
qBLCgQp/IDkWDNlXj0vegJ8PnzjzkzycQkrBw/vrWQPaijFTi7TR4QlhGdMJtw+Cn0OErW+YNTie
xoEB6u78+bG41/2L0gsgwcTsylAMHze7XvMNwitRT5uQpmhK/XfJzr9mb2iEOqzxEyrJYnPojv2a
o87z8Wc6lgCI62nSc74ihfEb+SfvqfWr1pCgfYFzzwpVYGYN2buJ2vC2nV0pxH1RgF+Puppk0bQn
2uH+lZeQ4O242uM65T/yCVJaXJCBjbQxe8NWm8SpHKjV8ogVtNmoy6O8D4pX8LIJn53zJ47QlQuO
qE8xYMu25wLy0z2RPsyQ0Cil5gHUbq5MRsDVBIXHhynjTeepGqCaPU7Azn5Ark1BSCsKFpSw20OG
YtOu9O81aa8KDCiUwOW4ncIGSCMruNJPHT+f2n+UKTdyTkS9V4B8qkSYOxuPuuqw1WjQZApTLlqm
YiubEnL3XUbck92SB7BIBYMTw7rmSQSX/ogvJjYuWKRPNyfl7UWMv9PBXkQzDRuedA2gKm1VTl3O
zmEDagD/6c6SCFg8PUtukYxdWxQhuJXeKben/IVkN2eSKdshpd6tpbiMFtubWHerJZvez9EkgRa2
qZUpJ29YHZ1N8AjHqmZ6Q2yEWx7ci6Oxy3FQfZh/ZQNsEw/zxNPO0v9068MEcq+M4wHyJxJmUbAk
9Zh51NmIX+616+tzLjE6IBnaMKSF/pqzhCppcylRnrse8Ma4q0srpcy4X3vFvHLWYyjXnr7jnzja
/Jnp80Eo7Qj6SDEd8Zpq+KCaOzYkTAgt+LmU+xFbLsCD9RIiUQX6cGgEDIiChKvIuOrhNa95iTQA
PFbaolbCy++Opy8Nm9Vx9XetHikizquig0RHplxHmPFqF4o5L9FTBxyR0rbbKhSr2xC0OvGEq4qM
U8/2TNknT0C0tTkj+9AcioTosptznHR0PQdO7YT1hp5UuqxEf/hHAHT+d5pgKspBEa6BJDl0Tybv
hxy4SAXGFwAG/aXjRPqEquPJC2B8L2OCzjGXQBT4RF0RuIOGPnv5OHsH0NSVZHhEPRSE6xezbqAt
vE8B4bRHToJAVIvWb+1KjEAtbDSHj6fPbLQ+nxjwtxm8f7cK5qyXgKyL1Vwz4ouG5cJo4+1Yc4T4
pzRIaCV8NbXif/bzwSyylsZdBWHtTk8rgSxX8I0TNnsB7OjGtRZOKzfpWaT6NzfrE/KJrjuqNekB
0FvXkIkmdCe8yUCOAQAfaKPcwp4nOEOn/xqDYBw5CIBoZQa1odjFSRbBmG7TMMfbFQk3mvDMZ3Rg
NVSLtifktndoj5uW42QNEF+vHXYShOD53j82ReVCcrSiFVbYSwHTzykobVYMw997CJ20nP0WomBQ
CuQpcfWxesXwd42SIprTc0DvyZ/ywG9l8kuMR4S5np5ZuLSW1R7V/999lGXIHedlFEAcGewnDshy
/OssmKU1w6ouXJxYWDzftGVKWLd4szsR0khe7nUgbTk6dTX2FRlpkVwDsz22H228P61dtzgmCNVC
SlTXa7OEeaNKmmQEIUyyWAtmqJPWdLNE2fNF1CjcZk7HheFlFkT2zMwyaER6IoTX1ZKP5MTiMUMm
yQN4H9ilonZTW1REdzcGLPldKfmdP/e2HcQ6mwHnzntoO+MLNsm7y8httupJOm0M5W8pXeUVWdqj
qCp9SfaRS/tEVo2Z7En6uoIm7OkEgtKFDt1e+Wm6VFXBE8pxuCAroLMmA104kJaVDL1TbTTzM+Rt
bVt/l1T/NIpulMcpMUcdMbNf7/3JVBOQ53cgBH4/LM61y9vKtsKyBtkWQbWm42DOX322wl7qbm8n
amGmJYIXANAmeEnt8tFSPIw0Jh+qLyF+7scg0sUt+DCvvtgfHuNa0p9fmshgLb1ag0wEvmXNUwwJ
pfQFxm4lpiuce/rJ22ASomr5jxjMh+biiuBZ4IKaeznhRRgfqhN51wlhA9tfsUzuUTyaE0T4VEbq
5Vn5GAOs6RpKUuL19f/Wtk+YgRJRjz7quflGAP5u49VRSRF54T1t4X4vVvHIXSclbEueCZSvP0wy
vWx9eEVs2xUisoEBYawdDINeHnQJNywYMtY5OCv4+W6ItLDTX2Bn25ztg7V9vz/h2Ay3GidzFpgn
2MKrZe6gNXQlB6Gs5xtRF9iF37fo2RLJUKU+xB5B9EJGyCs+gqYpgr0t6X1V1YylFoNiumI02N7n
HWvhy5bVddROSpdRT7u/zq6hrcl11OzpbP7I01AjJNH+zR8aZw4NwPL2//ehTC4BHU5kp9A1L3SX
+x4sicLU/9RW46ONPqo7GDxa8+B1Tz3JGjwamX9k19ncsj9GTFpLXe7XKjiNnQhCt8D4kPadcHr8
orqTVR66l9WGTkBhF/2h3lyEhkkb+LC38OgKnPDlZA+Xw38tpkBFIxQSDIJ6LNTbXYIiFFSM7SXH
znLhBLn6gOvH4ORKqh7yaUUXWJrAdsD7sxrA8u9XeZhVJclw2N+DH1/NjYGX1UToHxmOHyzXvqIj
ontr0MtmcoV6rZYcIwJS+MEo6kc+e+tF2WlhBwg148slek/bsvVGdemnR7IaZvLMoPGwycj0trjC
TnYootTQt3P+gOsXLDJ+BdVjikNaZn1nujm9ceJzoFNkxZf1g9tLVFWXSp7SRF6TOFLrf3D+Lpzd
WD4Dfn9i1rw2c3x2QeS/bWMQ8uxUBtZiZF98mW+uv9LnYVBLkWGxwMS0KfO0MJK4iiYWeCrcfTYE
Dghy162iZaF8C+rTLUD/36qiuR2bIViRKgDdu4W9KHlMD3a6v2DFQBegN2Mq6/1XSWGIeHaV2EmW
RP4UOGVc/l5fhSCtfZd7U5Uaggv0CVBKZnv3lBKojAAjxqRm5z3Qz9ei5vVDuEDc92p9RUL4r2jA
lxBP8uD5VrgqBqTH4tvhHYY3IdHEs4puMWuXgQPJubP7d2NeLfdqdJlUAA55m23kdaWhRrWTWmlf
TwNgMUOhnAErVsrVyWueJr5ypbmoiHOXay+/8HBAQhmfMNtfDLYANXclsPH/eFyWNwQpuRBet8Pk
SSMKf6GkJOAEvvcAEW+gEmZgcGowUn7reFiLPnlv/ENgUEnk2gKMWCioarst8RHwaKnYVqobRC8w
Psp1TCafT5X5EiXS3H3+eqTbVrcZgwUOfMO6hRhKMWNua5H3P93897Hrj0wl4juIr8jB4vQeQNx0
7s4kDd5hFjQ6G/5s+zVi37J7tIxYV/im/PEusRU+naiU/2tBiq7QBFDvnECh+MVoXXmx6TOqEmZY
jxo29w5KneALj/UlKbpWN9I1kpObsr7PQI4LUn+KSComIFVnkWHXzWfCFp17kTTU5rD+MnEubpbE
O9Ca5rByzytKOBQVP0/dyB5oGxPy+3kg2o6jV05Qe6FaLYu6G1jRF67kXK0D/jEWUBfI5icbx1RH
EPqqcglf1WTg/lqsGy3k19GvoX0055o8ixPKTW6d957bs2ZvHkTUplnsEucrjB7GipwWzhytx5iO
8qJE+jSTGt/SIEgu2qNpOn6FLKpIOIv2Qr7KxKO+8z4oF7r0rO6XQdGLGvK+Q6tOx9W/UL2av+Tk
L+o7h3Gdz6WyGIHGtI5oS2IKKZEhkWADQjDlESArswPjFUenmXUWQjRNmjZiNZETXfGWUqmVEk4H
DfWffThgP5BU0771BDn75eIDddCXj7IokdckQNKebCP/GchZndnj50t6N8hSVpd5DL7oaGSKgrtq
LwB7QuDQkvIPjYchn1eRBBNHUagpVfv0Im5n/0Wi0gMkipjiQ6x1eFRw6tH9jW9L4IPRh7sggwzR
EGWEslzEqJ44SQXJNjgJwjHzDjdiJ/QQpT5GzwJOsRizZBmvWbtdRKsF3mnPan3PZi1g2ov5Ty8/
tcUVkTsopVyU3I/E4BU0m2Ba/BWcrNErZ25CXGQF5Vu/P1M4tQQc7uXJCh8URVP/7Wp5QhuuruS5
nr/ihqtdM86Ms0kJud/lM/S6IoFH3XAk8uJsCLhyjyr0qMIwUc3xTPRDTFbtVoOhCc6KYzBrXc1z
jk2Luo/RuSlH3PEDxCzDItpx394YfOpiteXGK7IzB0vngLvnlgMnXb3mLcgIpxkmGtx+0wFyskYX
Eh+0G+4CdVVGVyDivL/ElHpKn8dXJunMilaHXxxmFFMxUkMCOr3qJko1+F2qnm/bdyZeZEiJry40
R9SkpVZYD0QknIxFVhNanYpW1ywgQWIC0o7XLvUvsIBzqXV7ZaIe2ZsYjPhzTf2DmmgKdr5k/5OT
YOowxcKOtZA3nVZDMr7TdWMW85SRPZNiE2vATXjrDKzr2F/VSVnzpNWD2jTXlJpBBCCuI+b2GRxD
KrqruIEDp8epbQ9JvNSJzV2IDlYlMRnkixMxxbHbKJnygE2QVOSb25QHXUue23Aw61YPqARyurbS
gDc56dMI27q51EIn7J0BMuj0+A8E8D9P2N+V6Vt6C2hOTdnd+IZApYRtxwvXg/++pl4M924OPuPZ
w6SU2P2yvfN0FuZijEpb5hQS/41hXe/NFgAv7nRRrpt/vT2VL3GVF272AaHUyo4SVVQ8aEXjhO3x
Q3RCSZwXzmMDmAwmyxIdS/onI3NaDuK8vhFPWpGrJUgH1AqiugkQpN3DJLFuvttzXx4lqO7Yq3c7
R3QE8kCY9ih+HtU0HR46vRrZhbSpn5HOnIfCMO1pYJAOiX++f3CpdcxKnFzHyq3o8xud/VBsAG6p
I56mOovbJ/mR4v9YnuckTC7FMFD3qnLRPTZfD9/aFpBdmyG93cy8UoiRwlNTSEa/0iAZ2KlouuuA
1M/MfyTImu9lmCOoErthkmrq5IGdsE1lSSNMQ/ADfE2nBdeYfux3xD1X6JOyrIJQdSDH8NotqOJI
pTTT6N/2Mc11H0qmQdHPFTafm3FPI800HeOKWEGdxyxjdN4ynFzL/U6UP6shSFKwUIbP0aLT4AFQ
5sr9EGMa45S1EejI2kyzwgLlY3JQwd8MpYmPqKRl+swmf49bGjpNW5oS4m5TkZkefQO8LNeAIAl9
KgsR61ZN0mBFYAU4IJ7NuKhappl69+Z6+hT7R+yzV82nj5zlyhy8p1QEIQU/GjK93Wa6qGfSXIk4
GV8kGU0eJJNJD1Fa2mgfUWj96JzbjBV+N2YJrfMtKT1MrTw2H0k2XkfxEKtHSu34ZLpgfiJChBoW
Yw3Dm0NpP8SATwuQlBtubCInARXITLxG4efPYX0DfizzZpzaqUkTn0Pa06L9fahq6IQry9m/iSA0
NOXZRxaXhlXffwjDSE8ccOYFetsxuYF7oZnWDZHL9ydTCYWWipat2r1lWiGzU8DUr0KHRBfUbMtl
+XciSswG0ctIgG8MwDJJD+2IOEh1Puz20HemG+njjctaYfwmIVHvHfHHG11eSvC64eNLDB/x7yue
c5lTWIyhVzKAQJ+zKad9+tipm849QWtBTGFotD6nu2PLjuBFh7kdmLEKYwvQh4A+WAWREIGI/HoQ
gaM6dMHUVgD7vm7hAcF1JTFdCVn4NRPo2mCjYZETI6ByBLzFKmj0tBxi902Fd4wI0XbzwOrXQZ1W
TijTJzkO6HoU/qt7SokvqtQiM5XqdaHVS7Y7WCqZ2TurgfY1TZjuRh3aAoXXfoQvN2vahteWEtVA
mSF6HUlKG6NzO+/ILD8k/h7O+vOniCIZ4BKSSUpd2r9B0iS8HNQ6IAtXPARNKlcOUGieb6PUgyAQ
CsF/IP2KpZ1ymr3L/pQwcrbsE/rh/BNZ06hkCXxqUAOynWK0Qn9KVYX4Ge7UNn9rgDhJiVEFUAG2
7rjTdUnnN7tX0tCT+WxNAg341vMaLzIAaCKc4G+EXvSWXze8Lq0tKoX4M3xtO6rtrv6U1dlzB943
28HQlWqFPmmgGAaqKMJPLh5y7Ovof65EDT76tiALzg9+IJozEi1rk426/yJ14YRnE+YW8iZPv0DB
VtsijTrnY8Vzz148WqEfzNc/g6OHaF2gtpWwBrXxElFKilfC2VkgXh8wkt9QnV9oT9Y7jnh+vGLv
QZi+hC3JZk6gfgB/n5zmnv8klh8ptXZxniB8trfqQUUG/aUrL3GitjBgPx9EPUeBk566jnWz+voU
NQFbjitMfxOt5wHxaKqCSxS8RkNTJ33BVhyFStfN5vSHJ9E3gO7nNmP2z1BZHefPyQ1Lmz8hzgg/
hlE4eEj6Es/zMi+yL8y1VDMe1PvawjBsf4vcP1hsSJ6+k45qCOThfzUYal3pVGauvjTSl3GOXQG4
N9Ni5VWNCh70YIkcN6uAz6NUfIVMTIaMNDtvU9SSJRcs4iUkoCxLPu7L8eLN5VEUsfEKYhmUE3Hy
0tL7FG+Vi3E6kS2xXdVx7/2hkqhYYRjgLJko24C80NFckpQRPlhZZ+oaBC0t4Le7Xda7K7pMOA1K
QY+E47f9CZzpY0Xln4T2RlujZdPGA75E6NGDUG3SEzfl13BHaaVo2cvTlKLYDAvN1fN4P3d+eJfG
QTRNlVxFW3cLhlUao1fSc/Eu6qgS8tmZ8dI3xgNxUtvXoPYk/MMCNi9Np36+wJFKkPlLsFi7ZmZH
ALgaIb52M4P/6IFCW1PwzQEoWBXjYPsnMgakLBNGvwQc3ZgJJUZB9hBcn9TlFiJHbz8TfZ4gAaka
kK9rVu5yqz828AMlO/eHbybkbuVuzv/5krXC6QQiF7ZRMKrSkEY4QSWO1l72Bmpc37JnlSL8L5/J
NYzyrO3i+TuZTfMN/mobohToynnibGF0bQgdXDvq2TNrwklO3DKemiDeL8kLwFf71OAIMv/lHdAf
v+wuA8nzEPbGL+h+/roAaCBmgJsBSu/bujKp9vKbK0mheWzGJxzUKhSzL6iPKCYodHuVwr3v65tF
z7tOZJO1dinkvkWVj+PQBwM84jQKdGEHkthPQlgnaIHBe6VGIdYdbcp2jMxY6PKHnQI+8GNlZGuQ
Gw4Jtub7fK+fuJLj+zaZf1IbEmLsWeNC1aI5ISKihGUbE8V4atU5jpRgX2AGz4hs7GyVLw+0p8CA
YDbD8kMhsijQ/e0pptdzros3WS7Ix3uqSrHZ49fMkLkQc29ol8tQFyH7UwLMkeR/2pJRawlURQ5X
DJNM7lo8JycZVT42yXGFi/Daa9HgL1GKKW7M4IkAf+t7sy5BvEUY0SmKsD83svZto7aghK5sl3I0
qXdk1OrJhCJKOgnFn/YCntzlFJ8KHYLlojEPwfG7Tm26q66ljld2VDKeUse0xPhEQF/oBFObJM85
lKQIsqbCxENgHoJjTMYQKSbYSLoCW06e66WL0ZhV0aNjUgLZLuc2+kYnu38wS2prMwE2p8FyXKvH
LtUcIWcL48T9KAjFnkuHQp+qeno7bsjJ8OWOc9JHWUd2L9+/f4fE3fwrHbJ+b0b2sXbgwt+l9S5O
QiBFuwqVDBvslTdzbvEyXL3efnIP94b9d+h6VPMyPhI2eMVGzgzXUnIkcmRzeTDckLEcNICkFnCv
TEE0PBsjzACY6Ut8i260yFi6y/ptEDHE835iMvfaBgw9FN5k8gBNP3VD4751N7mUPruvN4Mn/L6i
/LC8XhA/0pr0MIsOm5B5MmvlnVsWk++wO8OYMXSQBmXKofcTfvjSZzfENiAgU776GQgVyQzRx09B
KPfBp1BuhC2M5h1NmjSTt8JgFimfU8qZ4Q+WznOYXQhqFNy0zZJLuyBagHQWk4KWzlSx+ru91lZQ
3OeQ2C99wBcNuKN9C723P3W0x9SBos+bHLM8NLSv0lZarTeou+LB8k1pS4EtfPXoY0HzFom//VZd
P04B/B3KENqZ3j4PztqXUVmuHskGmGR0Y0yqP99Bgn50hoaL4BdSpotVJ7CLCoQhGkeaa9O/lKKJ
On6OBt/OM7jSJWSEqXQ1cUBq5C+inaUUG16CpAu/vUDOHfDN31+bsOAXXuq1FKLtCvjE2KNLkjNO
UjonnCyqrYXHQBVAM1VPkCxhMRERcyfBM5prQXnoefyuSP7Cbhrlm6vV+UvdULS6KedDF5H6ccCi
jcONH6PwFbXiv8WcNlMU4cJt2KaDnNjWs/b9+mVCJoSZVojECybja2Jd3AjPl4GY7AotXcwd+/aq
3lZBRL/4MzWcvLx4Zx4aDePY5q9PCXx6mtZpj2RlcwqNffzOQ39Hl/VysEkM3Jp3DnmcFoL3u3wq
1mnQu5gGIvtoAAF1walXhiu9qinzjLNrJJtK4c0N8psBI89bTafJo5n5CmlMMgBhLOh4rFR4bto8
s0Eq6ARERyX9XW6WvFBdNtXO9VlbL6sDj4lHL+c5LE1ScU3OLegaAF+9YGQy5tpOXx6DMMLvUd6V
m+P4ScX89zwvGvSO0L56B8dSS0D+Ww8Z45AV5lEw72mYWjuGvDF95Cr6ZOg9t+1mRyCHEoxSVa0v
QS7FIj5zuvLossVAKDZ34d8bf0hIUp0pCSNiH1Y0yQm50veoiOgyQ9n5SaOeqUAh2UxziZz7sNvT
PGr2rgllzglPoekLCXRrep4FpYe331tiDyB8FWlYBsh1D5fkCHR2UY1VuqH4Lc/qsYmVAD4Dip9P
SqE0HxtotjWtH/aeyxGGS/vOm0OGNCRY3T0mgeqaBNNBYV9LICnKeIypZmlHUjesJQN71favMTYM
zMSBl3R+LFhNkEqZIEuIPC6sIWcLtk+iEz+Nkn05UkWZb71CrzWPO9N7irbawUrsHJGe4Zl6HpoH
QcUu939Bj3Zr+hB1o9Q+SnMHeZVJk7tAtkW0KOFNoFHs/BmUTHPaveTOT7lnecDUhFL1OLdkXf7F
kJdT/+MI8paQwxGsLQ0o8UI0fkIwKA7d3djkqKkqqPy5Mc12k2C2QIAqGjBJd/XFbmDLSbkD3RSQ
OLmqtZxn6SGHDRuFZK45CeGPgXhAGlJDj5YGVUmM9w56+xxN5zNVNqlFMY9JNX3rwRc+DjiBvX2n
3E4fRpKpheBdqidyC+SE2NyVvKLZe9e5l5BZgem9FLm2Zx482mY8/fTZdbvTH1GPguliz3Dn0Y8k
kCrUQBd7gZ88oIF/9s9X6uRyc0uDooh4Nm2uIvUeSllsZ7lyzUZGAaYgS4o7sR8Oaz0JA1LFOpra
bSmGsQA9HWY+BtSkJhj1qTgmCpJfdtR3QgPKBsBndS/50iFtGRh3bKcvyBdQEa794dtSPW+7XNdB
gmAZQfIoqKkJjU5ugZRX/R9UVJOtgF4gpobFNL059n5zF3S4JhU0omUFD8+A/Ds+AcM049XD2ylx
Sj+zqxjn+9+3u893BIBBbxq0lmgymmRFHHh3sDYfudMkVtm9Nj1kbRtS5svMBcBDA4qR21uoz/VB
z/opa5B2gQxLazNwSVxqSDymhb2QIqQAsXkeSewEX2aUi1m+se0XHJnjT0nSQ0n4J2tDikSy3XMg
zBOfRKzjMtb84qXFZuq/GAdi+uNVooVD0C5vabhYjxXk/gbEpnpVFbXMdojrDVVkb/508yuBlxFi
ia7p5wIjVBLP7THOZ+XJL7biN6SYCA/5gD3rSzCEXcJcwxUBSg1heVshXJ+byB08KowRWyxmtrIA
pFwjARPYZhHBH1o5dEIKUSQuZfcOGenlICq4CVHXJi3Yy2cLXO+8wK3/C5S7+GcuSzg0A/U6QUSd
UuKnEAezl3K6mmk0X1fgS7AvvQDYRYCyVmZT+kCVSvgUrRQntWSBzFGQ+Z+eWE3EAQGYamzgXv2z
0+5arqgh8spGnpWBJk789ZyWM/+CrQAWGpLMKkYj+YmCXkUZ7kjrjSmMZEkNwY5ia5DnsKtfb3ay
ytQKHeEpKQiqPEf2A9UfSXqxUqW5w4TLXv9RJ1oB41DUEyEMBiRZLPL53GpUFdlLXvhrNJyj4jLo
Ag9u+UWZElJsdQvMIwFcIPIyaPKIQFJKtFj43qOcEowsm/Aq1D2gciHRzi1wMRc/n7zm/IdG8lD1
mYHT0xioifTP7inxYW+8VSDRXPaQ8Ll7l9O1pJ0W5IdegnLXet8DuwdXuVMdO3CqNChtbJjqRkM0
d1LWP3YxXSIeeogOOTWPgeXEkGLNsNM3JFzm7Odi5rKD3wkbquvMJR/C1joc///I/W1ORqoF0/h3
W6Rs+Q8Do9J3e5QUJuV6ShZBztKh3xMzWNgEYrTW7qDpTC6tafrXyZVVNTTiIe2ZKofzcAZUEddz
LAICnK26mYpRHl53afPjGPPv1qxsGymarmKf5tBAvk5QBSNl6olmdh2+jDWvZWIRDfoflhpQXD/N
JLKSRPfL0els42GWRU4EEE8gYMvTB/KLCqng2doA17hNwEZVHWOKk1HKAE5JGpHiMdiaXZFxQTcx
doNAjn3XDlVivUfrQux7vMRVJsUrYYoHJ4CrqpP9S5NUzSLUB7OPqjsiXVuGDFOs+0CXpI6D9RRF
X1Hhv6/P/tEWMgMAlxBhKXwxfmlajzKylekENlfnwxe7tKD1zV8I/7sBXWmcCMW5t2TfMKc9CdLY
nZJD7twF4eRMC44xIpOqZMWkSvA+6wQi073zcCOoH/FWgcleE9wx3JLPp3IbogkUjwixRKCieb84
aOWbxl1PRpKQxolwIO+dnFTVHJpW5o0KStYHWsG0GH7M2EY7Q8AsuMmrbysHYr6nEVAKCzkbcRUP
gEswsmGT/dDYorFdceelGAF1ZxmBgDnRPB3m3ZMupSsY3ujDXF1IHcW0OHkyED1Ac9C6CXD2Hzht
60rcyEQ60VSLwvFj5G8aqK+OlQybyFXs9dxnNna8WPiRRM+cw+jvU1AFwFaJL2N6680jJ6hl+E4w
DdkS0dXfKB9e8eGPbsjX68bUY8PMsfEmO7C+qiEto3cf962nB26FKX2ux4gVLr4NdA0J29EfFBEN
2d1RevAG0BP+t3xjm9eoYk3h62XYDjbgSEmxSClYmv4Gif+r3U4hSWzS6qcOK5bNozH6xxa+1KE/
LjvYwVAn9DznbXvwgf0DfFCLdWs+N6cIYfoJmui4MOTy3XkHNiwO/1+ZfIuQJ9MNKjxF5L4ETGUb
VUI05qZ3o/J2Jrr9y6ivs7KP1cgVRgmoLqVC0ijY3uR0EpxJVMJhktVKedRyajWTBMJ+IRmlx8xj
vl3rJwI8l8Yzeem0TXPQCPbyvtMdyx0M3W2HZxInsV1i+VVAFdZXfam2OVr0pGGbYENg17X0U/6T
wzsrsevbOJw/XthFVI3iPPpiN80DqBwmH1LE/1KPwNzRlO5mfubB0LPbaUDyMaceXgrC3iukzKI3
8OWDK2gt0Z/Sh9p7zW8OEdm+7U7nXnQqiNSp98OrFTUl033fwEyMGEcmQh00i+nbfvuSRtlZXGs7
tFr9CN/JC/dXbSfRkXUx1lbaEpIx44PejbytKETUwen/miNHsUZ+BUTS4E5vOp0gcCv7k/aJRNRw
KGOua1da2wC5XCXnqfGtwS51iTqnl0PItYIBa8O+q28fuoZByiRHKXdfwrdK3suepNZRBtSCr7PN
H5E7V98un/kTG/wQ2MzuJpHgmw/uUPGfBihiWPFzIWOkahgi76lP85zv5VhvtPzA88E0r5QIIDD+
TKz7Q3oY8oe680s4bSjqDvD69eM63lwF3X7sy8uU7f7BRoo0izxSqp8L2NvYl1FAjt/z4dCfGWoc
uXhxYfB+M3TrJu98rESvxljxIZzp+UXZGbnEkHX3jb/XIe6/ZOOcDM/9GuhlwmDfPFuW4lFfS1r0
o3nq0XtkX+iNoTX24DBoZf/zUeBz8Xbn31ie7HDIaSX6elLJA+VhMKhmbrfBUio6uN1CoE7CqpEh
q8gQc1YI3J4tJq417Ztq6vdINgeNEW2uhwUMMyhdcBZuRlK+5esiJUdn3WX/9r1K26YMQ/3nD5BO
D2vzjOifzCRjvAMsJ6KeWzz86mWUeyZjwSu9AWBy+mwzV/kNxSGsXZfvhQd+PosKOtDPSgyZaJkc
en/Ixf+sgUqfQrCgHoixEVJt8lXmcutgSUD51BROCmS8fnDwEzDYs0qoDC9HhKGx6wk4u6Lfqj/b
nt7B0Vx1G6sMpKFVrWsGQeu5m7Yl84dMx/4E1rCTIwdrG8LCkzrjhuw6jnpu08ZzEoZN08FPopBy
S7RLjfExGgswsurQWi1+MpFFp4PukOOx7YdIJCSg97AC4qkv3WCj3ykP2ZGoQ+Ic30t+TnaqKFAJ
CaZBWEZQfMavDSVx6vEIE7i6uQud6itjcS6EEwPRXhMDomHSlD4CUMqgaBQr5EjDJcfJB8nxka8R
2s6ndRSqm8Nx/pxC36Xi6Bq5RYQMzO1kaERusdbhP5MhHp2R3lh25BlEz/d88ij4svuoBY3ocwCa
jentLWabGPRpWp27iEm0T4JVZdggwqKs9m2YAl38ib8SE5VpJR5SKalFyQo0MqmdSJ4yEWmRHMbx
tgTbLX+QaTv1jh6uu2vGyuANmUMOqtOltfgKSA5AZssgjzcMYXaNKMZWYF7F2oYaA94q2btEr8W4
lJdNOFLUtXouw9wkVdhm9uK9Xgm0vql/H19ddv3yRhYpY8rVYwTU2tYuOt7KWt8NkPIfg40FPcFc
csUtAKHb5WR2yWp+ymvWIWHmpDV7DGbrUrYcQ79y0/TWEfRSNZrHnNKLZoVWs9UZFAm4BvydFuoJ
iYgv3SX45mWsm5jpp75KuBj52OuBaouDsNIROyiRHGD3jNdD7RhtBmSyur/JRVfMhGY/mSPTMgjM
7FwYKulI4HbfknGIFgRKzrHh1VFqQygKt6sPiMcYnry48cqIwmjTy2UYMEFvNYYvTfgPEgQ50Ccm
XD+el0qFPPRGVCqPIvWiIQ20lJLe0gYcADjQNRi6tte5ifnnQTYW93rq/lANidBq+NrluhEWMBog
5SNZcBwhxl7yQJIuMvyqps32RUyU1iy8rgu45oWOVfBaf2wZZ4j5QXf30Gt/sR65962zer6eCMMd
gEmvV+HFHKvNsVZUjLtOT8y/lgihBlnCgshY7kbI7+utH0jsNymDlyrQBb69hnuf0Ywjp6Co6nJa
ZOlBlOPcfxpxmGBWFEL66dMwDUHVFYf4nLjQCOVmz2KNQZYWIcNUpSE85S+47JT4pjeHvGLBNfPT
SjbYK/A0P9GQgrLNNvRkZXnjSqpBsqgHZLooeA0B/vXRTL4ybp+cU/nIpJ4QVpidjcdzozQ4YXsb
48uRjaZou8zMHODu1tJvpfQtPoNPn1ThCvOZxCfJY41iqUSVpgGsJmFtbfEzQx3HlCOXcguRbUhA
56ASKNm98B/NlGcKoLWeCbf1niQthZRkBunURnkk9HZkVrUECSb49mANXHuvxLqjfMK06aQe4p/o
MQMyrzpI3Q5SH9LDHvlKQE3qo1df0I5jpyP+DNORmw/gmAkYgyEje005GT7F4xAyuZ8UIsiv+W3I
nSz29jNSCHgzMqbnd9jD5/Z4Sv1p8/EgkrjdRCJ7Bv+U9yrn2/8Dxy/f1nXijouh10/QjUkt6YIQ
EZIIyQj1wvJokWH9jBFx7KNXhryZwCBzMYejttH5KjC6d0duvVIvOeyojSugL18atlQewJ+jcIuV
9pDLuMtr+D167CQgCi4+2AII0DPdRxRrJQQZfvvCwLxqhy4zQZ7Zd02PG64vHjRs4GGrJFl0FmTn
MM3NQhMV5fMAUec57jzmjmUIUhdJU+PA/4/oSnUXlL7IeXEOkiYTVoA72jUV86eJ5YHEWTOgfKOO
Zh9jP/5clDfzo1aESejo53kpTCteh+arVVjLOBmjvCg8HQOJFgNCpEvCEoS7hgpHcdpr4x+hjodA
wZgblFw5o3+PtZZmyx6SrRJneFdcE3SizcKwEvJGnjIK/9K/eSm/njSASYNnoKoUNnO1o2o4lP15
YVB6+mj+ojAyylYlR25/aQgktbH9BWtBqiArSfe+Dpllp1EHBPBICXoIzr34RnMndASd5+V7XubS
p5o1+rOdi5oH+OkZLmOMln366t911LHR8evINgct5ZLLbjmFIlCXoFEh61gp+i5GX6fwUhBUQRZT
iNJdZ1/xL+ImISQ3ssFMmyYZxHi4KKmuFYII2McB8+WSMFvU0vqoL4xFcE5s5PjcfGWeA6lCOPfp
iPfcDI6SBnmh0kfhBevLfKEa6OUiHEq2twhX5KNHVOUVHDYKVcpoChBMSkHbHzm+fl5UMKw6XxZm
J+Jci6wtQde18VA5d751V1WOz+vUc+PfnqJbMlqakdYJIJ598HEPWrlaVIUvJJ/8p9nzzbYQgS2L
a4fIb/s7ecdDgTjCE9GX3NshE5hhgfK432hvwUMXUsH0kFFvbOsSL+/IJAZCXkL50VQ41llhTtGB
/hxqoUWQNqDIiaS3Qi+xIo/JdsKssfSANEPReGiotmWBSSLGLtzAp84gJP8hlI0nKfC2JETg9zPQ
YbXKbKH4v8bjX1y7ISsOPP0No47X0pV37zKgjeQWfqLv3IlaoxfS3LPVu7J2VVeKNdMmcZXsfvJA
dXrMmyJpiZaWYlHjEl5hWO8SE15E7zrbOk9+KM1MeU6exE44eUvhqTeYtRSioyZULDEng5XQndey
2f0Ld0mLZGw6JJok9RhuSsgQrQ/CyoRt9MYRvtuRnasUkc+LSYNlMmnRJSFCmEK7Lialu2J7+nqn
uCCgNL9gOfGs77iHb+r2WD/2p0ggUAeWbElTkoISzEXD/pUO8PVe7DuIefVu8LueYrxlELQ5OVC3
o9AlWpcxqnbhigCz+Wh4BsUfzruO76DtvdoSOAL99BPYYz9pNB77me9CTKVYKqYkTi2uACj5USnS
RELyYP5J4Dz87e9frHnoSezBc2OLZWZsaRbc4kjYq1MJwUUxHUX9NslgEGmQX/lzV01JPfH8BTrd
PQFBiQMv9DuHEB/3jcnWYFm+mI+/lx1pGmgnmZEaN/zqjXOWjZCbUVjKRqyoWcVkZiIkcvXrIljZ
/MCkPXDpOk0EYPVFhltRmQlo5W/DUyJdV7pXAb2GmdstQiT7WUdS7OF5YeEdEkdKxQQXKNX4NHnh
U5rHO949iVkK6osYVAkCTrxDmE6MQBd1+PiMDwvL+VJi/s1dvILfHV/NPqiNG4RFv4gICM/g262K
kcABfvzJIIkQ4lyqrSzdJXZhl6WAdaKyXbpkB6gCw6+Pqbp3pCWH74hTIo8u6aXvYkC8yiOxTFOj
MPXpECgFRd9pGl5jmEDixNTQ9dMGbm+t945Kotw6rdGxJngaeI5V0FV3eVl0JdynU0ZFNFP4TVYI
WKRGTzDBs3CXYSfi1ueGjF/DDRaUJuFqPkqW6ENp91BRc1bBq7qFpzXQK/gdBuFcVjWPZW2Fiu7l
JLhYA3zyj3uLMzku4xFgwqnYcN8NGt0Cwrcc3iZuv6T7ukrA9fKKeWyblahXqXJjf+vpfdsmgBOI
DfNLLTsrqOJwIFVUEZH/CFby8D//WirCrgWOH+/9ov7c9RYR5HXVJ7H2rrJtSSvoo/vDxqB2JkST
JZPWf5LG0NBLZ5p61CnHsxPXKjhbWGFqbEfyrFFlgUoJlB7L1dqvPyROcD4QvZfYwg/WEhH8Yo7a
7zp5geZbR/cdJmDz7GeTU4KlbhuCeLqQvNSjcUyoZ6V9yAxd/iyufXbpFSdRSDZNKc1mb0afu+yW
iSyUjFshmjpB4aI+H0T+Dm+6Y/3eERa/QidrNwi2GWcJhAqNq+G4lNEFR+IdXvtonxQKYegSzvaY
CT0VJ6DuO2CRGWGERF+y4ZKf1SR3onoHZAUVJ775D4qsl/CcQ86fi2JJf5ZXGUG4s8e7lpfI+qj3
kwqxtV3Pw6HP4SDJ7qIA4DPE9SEZXSbjQpJ9mmOjPolcoeCA39am1JPRQ3Cf/WAcJeZwzZcQmnAJ
p0GP6DOEFzkr8DC9evhY8cqZ8DBK8PC/gCoxb6S+pZjU2pqqSXLwefOoYGM2tBw27IFfjdu4C8pG
H2ukNz0IKmy9M4+KfLcYv6KoCp0wB0B/7yShvSYw73kwviEQqSX9rzBsV1l2wETvF52v3mWakfYL
QV6PSe+PDwe8+7YWKAyOmgUIZ4MYQZyxvPXJRzZKK4aZQ+shtwN9Gk31LRsOCMw8u+JtZ/N3kKmd
G6GzHd46B8ylLhp6z+s9JWMT5PgCidL+q86wot92YVW0sCe+/YxLcuwtS+idiOBXX7NHFg4FM00z
55pxya89S7i4oLRMDhWuFj+mZbcV+wlZJk3NPPcWgSSx+6UVptQw1UMV5UTT5a8X+nXp7UYTgVUS
wLrPZEbMmeomoKHM+Lrh3Rewu+QxGbjw3TuxqTRcZyMqNdQVn3gmCn9lRCRxkJnFnj35AQUaozuY
aHCvH45nw5FuHivaHnM0fytn04nxsVHONavI9yICw3oy0DyO7XpMOZWgqouH3pqIzFz4LNRmSv+/
HcsG3f2RKSxZvVDdb6GReSu4QyqINQO+PMo/0hbFbNtALlQ9hMC/hWbtI9CFRbKEUZJrVECCilNz
oaHj1CAAfEVoqWcvu38dtjOGLThahVo3diSp4NeipQpwEhJ8uOoV3FKaffXy7mi7U6bwYZSGPZcl
sbxXdLv3IzCi9P8NWVHbif/LRP4Z76U1ZPg6RqbsYWftw6/5+CNsACxDa2o2NchK2elCirJqNVS0
OManKxi2SfTSjp991y27K+vw8xmuJ2ALqZrJSYcNt6g8CM0bAxi5o5GSy/0MKq9OH93ehwbNtayR
UICRciQoGYfwMuUKP0XVwleU/Lp4s/FqBlLayCI9EacmsxiVSHWLD7Womf6vHYN3zRqLR9xBZyIB
t30p0yqB8fADrJ8fkiPT3z2kQSpmAaD2QjYrlZxJ7W1XQCcWIfdlvY8XXXF2qfEiqadKQBru6Hw/
RfIji2dbGxhsnCWe8aGQDDL8ZDEZClcoo68MPPlEEgpb3cUIQDgkRWyUimh5xR6VgJtBkgYp6+nm
LgKsbalFumkitkQFWbi/hd05JmwXK5JDIUzxcquhRut5Z625A0vHyEcUCz2X4flUE+xy5NXfQ+Dk
VGNAB1gCO3yQ6oDUfPirr4JieZQ+weXZsQqf10JNQXgoaZd3UA4G7rIiDosHcrSmStKUoqsg+Ox/
4lDUZuuL7eOcWHDsyqSDwh5zlYwN1RtzRSrYQJMuL8EsaZKHks8FKKrKq2oeKZcIrWN47dYQr8dR
2yC1Bp979nCdMAzQw03PJDiYNGimGsNDgo6tLnaTY1oIY9M8ZIq060htNSp76KqhJU2vX1A/pNXF
h2KO30Tohy/BGldNIbGr0NiiMofQ152H2xO1zAVGKz/XX6vh6CCTqMClfn/7rugnYXUEHAxjhaoT
D2hFuJB0eUUvjTKuyayD/l89j8nESbmlJyYh6sYp+cUna0xPbGFgacbYydzBexxnO/6MUT8XORQl
B7GhfoNmpgyKP8XcqsBMbSzwR9Vwg68Q9EiLWF+ozkZ9thvkvzNqtWPlg5j5fyC9diY45f54joDW
aN6Uf+/EIiepSOubZEYt2DXMRSP5k55s8UT1zTRz4n75SKBXAuNOerTO0BlhE7aCGO+ixivDUPCt
JFV5gS8ho/bZCxhKYQpO/EgNSgmwznIq8dfyJjEXf98YNVNw7Putq7TaJ0mhKlZijgTg5mR0y92l
VN3IwtG/A2/IvpFmvKFWG5XEAygj7v5W1piQR0/7q3d/0sxlxxnAdNUORyjnGfJiOzhT5qf5CJQ8
fnuoPk4d6WbDDUG9L/7AMT/sS6+1gGYwOMBoDCQnaqEN4jK64SlGkrfHuO9oZTeC63GCPniAWJjx
7WWpjowbit7brUe8vlw8MCnKv+RByLr3CJjSnLdLUOeb3QsmCgRl0mx4y/q976om6OFYeFqkKAS3
tVFTZpxT4fyT+KxetEEX8ZyE3dva7NavIKOUQy04cBCW6rgRFrQ5Cj6QWCTg1hbbi5Pj66XMN23T
fIix12kSMKxrpISD2SKMjKK1zq8QuFykymUigsdPz5HWK6M4yBRoMCxOgtj3r0K2EYFgl7I6hnfW
g1EPRbGGaL3khMnj9x3NkBeA/oMAaHC6D4eH8CJixHWYlxK9vCjOj4OenbjzVAH3u4AHcOljysqs
lEJDrkoszVi3gB9S6gr8TIr5t4JX/vsg8xKvSZCUyDTziDqoBqeTCyNWLZ1r49/XEEi7lKlyg1Hv
a3EBdZpR0Dvd4kqDAM9X91f3nPgG2yAyQJZH7ydWhzvOySXCdevt7x8LNPJcGL/IerXtvhyJKmB1
z1LsGlH8odNAiWTZmWBJwdovMzKn/L76coOMqpXKhTDgMBa/H7SqsUlpo40QoHcN+1Bj+CT9asES
sZl8PCZBO6Z9Bwd0nWtL4JEkDLGriOI7PCGh522I86yL6VKJqQ+pTdk9Is5nJLbwexJp7flTk6Vn
dL+QI+lPuA3UvotuUYYEhNs2c8JMpdlc7bnuO7QY0LYJQwQ9IgWrMxXAHUCXfzD8odZG4jovYwry
q+YwgkXh+QiRdc+Xid14MZCE/YuZ0RkSJWto8sOck7jVFLyG4yVAC2lrjTr+7KP3R97pjG3C5vCC
ylt0R5TxvLuoe7b5A2JiBcLhUDwcUEUDL8hOZup6zJjOM1t2nADZVrUc/YhR2xAr0AF4mqyPrlzd
cM+JfKi9Iq96oKokrHlQHACXIMZwlDkpzgcd7a+2MzCZ5yyroG9gdmZlVHK2lM8SwNOuP3wtPuuB
Akxy1GgWbS3ejjoPEJBqc2yezOUrB8FV5uFsLdHVIPxXQms1no/zEg7dNA1Xptu4HvokuWNLADtM
sfCYxcSjPH4fk5lCSeJGmT7PqE+f1ySmE1ZXE06ibvLKwRJkoCdUNzzEnIbGMMElB4/eW5FhI+Wn
rBALmNZBGx9lBPeYarKzuybbvKTzMjyRDOnt0GQZUlP6yYFZOP5iqVE/cv/DCqjG9+Jrq9NwgWWr
joItW98/5klZ8KBUeyvB4Qu4Xv2Pt+l3UQINrNp0UpJufCGeLLkT872SjMbT545Zh5SxwHr2upOx
pVSlIsDK9cdT9cYRgg2sTw9wO3+c5o3MHk4eGn2JJwNKi/0kxR0wZU6gVGjGmpefB+/sBJVR2Dyc
PUHQwzljq50OWZqjNvrEgfxkywgECv7ZyOCE4KM7IWEc/LYGZkZ+7n8zX3F4Fjk1DT9TKXTSokhO
1PJa2qFQGgW08jkQ6ubnyqQFKvbNk19xI//X6GjS91SXgWUUeSfxsDTkuAGWf3sKQqhFnodLVEUU
6rbxTnHOODOLk+YBnWBMwxp0obybupm19oTbruzt5lBtlqZp3rMIS9a7AJpHiKRnb46cYpJbIXQR
+SRWn1eVy4JRlgJZqg1QuNwFSjIpAULndfiuuf/xWkO+GgnooWpGdd6V/3M4H4hP8daJvE9+VyCt
R4Q414Q0396TEk1ZlynQCGpcz5OPvgpw0UKTObJAsUcOvP8PcVlceoB9qoJ0A+B89+qumEHrMFrr
smFivP0adl7a5Mm5GFuW8yOfoEu479l3EM/rjzVloQqKtFA1XwXiHlsiULTWZdGD6/mHE7v4rO7B
q/4p0NQoxkiWae6d3UVg/Hd8q9t4XsxMXxWUJgJF47WDWq8qePhqpW7TwDrKf+GmjeXAcb9iWp/T
gY84YdqyTENEBoN9qFEzRE2OQvAFMZp4TtaJp8WebgCR/aIDQWrAXt7cc1euIzMZugUk/B5Q4yvt
geSVRdO7ErHkb6VFu9Cdkpp5m1R7I8j+FtvuAHNfdBlBzdtHWYEJYzd1PADLvPn3TXReHjJUysP0
0mpun6bNuvucBcWWsiwQp1GlcBBtSycZXnquFmUoIHRqL/eyxTE7/Rokf5TfKRfj5r59EVkvHKRI
onTmGYQWJQZfpzots20hCK0cvX/8TBdOsBUJsJKeVIFLG3OZCVdsQcuXs5mzAXmtGmlBcHpIqE++
pmQ7a6K+b/8RhXjWLQlwx96jjulj8gzEWhj42DP6wp6IwbWt2SqFAK0NuBvnsBVESuIJgf93NQlQ
wAp9lI/3kvaBe60/8FCg1Fl9+cXClDljbcxUp6/vMvT611NgaKrjVafn9LqkBYpV6+e7ZAs9C0G9
9DDfN2lwZPuAZuBlcy4suNVLjQRHUEkHGwIuhCoWEHhtpDqlCEl3MA8+oCgu0m6k1WeVgh5CKiJr
0Tfp7/iUYu4oV7WIb/MWRjYIS1WQi1AW5mPBRgdn+Kk8JExpPHWYd/8QuE55PU6JqWn7kF5jz5o6
+dGF1XWoPwsRLSmv2SiignEAof9eMtXSJMMA4EGEUUFOLxBX30nqeretC7naGpS8Ph2u+DUQqgHG
etx6sPEVCXfkJi1wKK6UQpvhjLsHqIb0n/QkBxK0T2wbUwkP0jWb1/8gPYmz0wH5mbF2dN+Uxdm+
KVbU0zO2baV7vAzFq9wTLqgY5RnrpS6MOCkb/0mscYRrNIfzF07I+6w86R+gebIU1vjgHVtAdnaB
fWVfRuFT6OTgIgAb6UZ2fRbW9WlMAixVG2FVi7ZaXoqoMRCfRbmL5ZSgBHTwWC/5RUd81QN8XJhz
yafbeRNUBj1PNMJa0BVpTpLnJwJsRHPEMbBRGFLj2Yui9Yd7McjEgwfP+ZTIETWo8uhikPoAlvpY
S58fc/Na1RoRe442oDsP+zS1ryyQIYd6mQBpnHnxAmLBk+1SrN/ZUUCenHdPSyvsGUPfQWfeYe0Y
NXoS/XJdqjO4DRahCiTGVcsBjRQxAd0ZLy0b4OfYvTCkPIqUV2AK03N+FUATx7OBhOWmgL4M+f/K
PMHuQZ5eVcL435k8vtpyBLw76i7Gg6FqSiL0WwXH64ECNJpyVF5fpWD7SsxScIudQN8z8vzQZ889
6ICfpkLbbgfhWMrxqEgyBlknkYXFxM/x5GKAJfunXjGDyJo42c7nm9wNjl0nKH8qwrp0hxf0MHUg
mYorK84NGMEEv2fIaAEn6PPzQxFTrYYDMBUfZNNscrnKCrH7qJZPawv1k5++bOMS6Uet60HwZWtE
Dgbd6fd/XGqTnLo55s5jC9UYpVIbWsdcv9vOocpXbH8Vrlaj/gcENZoVGFkeIEORQdXxDfGomymW
bDhINm6r4PkV085mKBdbYhpjpIrsyOq8kWIr5dTB7pOAErybm94rGr6kweBCg4E2Jrqi+db/+U6J
hegjHU/vyXdnbwEBh1IjrQ65Vk2dt+3OgORx8gLECVnkplAMIvd2SYorHQZ71TRQmHQAxDJJeMco
Ox3rC9ssqXvSXOV5bi8m7L5zoCDRRQ6Pw2EhZJK5uYjraVeL9o2UEOYSJ43kN1gg81vSttRETD5+
n1oadBtq36NXnx9AbUmWexoZyBpZrCfQgol/gpgTjRQOZMHw0YpzsPNrNc3kcKJzqQSKZ+cxakHH
/71/tH4Jn7IkG/QMyQoUB7oAbXjSqLG9W6KxMDl0C6guQyOhngzAdiJ9kmmHaxzcNR5XtfvJambv
UIrFCOgiy+wQi4jKiAFmKX9sNmagIvdG56BDkor0BnJI7lVycTqJ1IBdG4Fu9JJdACQZ9wp0AExP
hGu9rhZAzAo+Nm+YN4ef7Dck0UjZmpDMKy+fYoYruMr+ZHlLToKDT8iIAA7UKHXZ0XE+fPgSYTUn
YXbfi+aN1eNMcHSxzUx5H1cfgSoN8ar48V1tc3/C3UQFkoSWnjHDwTUpYy86Dw0T++/peDTmIwSG
vcUdwyNkNU3YrRQ4O6LyCbanQO1l9rKtJPuSb/9Bl+Tu0lUOOeUPiyWum/uI8vxH5qmdAIq/KpCN
2Xsr8r7vF1fYqXe29oG+h0V+0vtYWza6W4t4kAZ3s0uqCux2gjD0kUtPrb5y6BRrpmTZReOgipp7
BtEMf1hOPGvlZYHrsV2PI1kGKox+VwL9DTMoBYBEJ4TfaT8Dkt2cTTR86ViNSzogUnQyk2hN4sxq
kZaWz2Ium95q+BOlyvuX7CcgxsHWTrVAPro+ZePp4py+cPfz354yH1qpPtJY8+xl11/G8x0dJrep
dwGvyrIexA+eGwySSvj4cjom450ejdyYLigNi9g5JyCcKvk2/tevrpvRNENjX66HiK7GeSLJT9np
VgvBkvZvqWTAb0jiFTMTuK4SjMFW92wV0Ww68VRLVE3G4aKNkwvTbeWPsorrlzWcZk4RXa3pnjnD
LlUpiNw7cB7eR4bkD1kD+GhSSFzPHcrHvm+KnYnDcPaKkOrjyjpuSS0pUEzYl9YjAgB5oN3DyQfy
bURX8ZrYDFc9ritTDkrNl1EGeilZgBE8vEUEbU6AHqEAYj7cC6UuHwlEKNZBsZcgAliuS0FMYi6R
CTyFc1CAvs50F7uIESueWka3yBOLvxE/hK6oN4mDBumbdAL3sVI+FAvNWOjfaSaoMY10Xqwoj03M
UFN3MXez56M0y+t1MX+/D6X5AHUQ5uyE9P7xCPd/XY3qHGd7iHX0AcHddGLxtL3vxTCZkIEZlYMC
PTZybW1j8KAsiYsnYpWfjKbrqjQdbXqujwNKLJV/N00ffroLBBop1pzWdiVGj6VvM+LAhwA2o9PK
RCOogKAe8HEe6XIlRtV1+kK0VR1WZJNw0pnU0NXoEP1opyb6O8xlJmQskKMw5R+f3XfcqcZImjtk
v++kSUX0lPQaCrAkL+ALKgf7AhAxTDowPXIvtT3+CWxxY/IEu6divYksBMCtguNEzeoSwxHlP9cf
3N2er3Q/eIyPf4/gxAWJpjY8FDVemMzoLwFk9UoeTLvq9PTgFQDRhzAiEZtJwxBBjJb9+WLuDITW
F3kPMngYuWZFKLM1DNSJsaTfVEuA90MeYMn5fApY3Ob+4UeS1kUG99bbotdEhlvQRvBCNMfsHyfH
83fEuKqA8hD5VGZB30hLNv1d00v9lC/FT3N361VxtY1ZlPZiWieqD9LaDCpoqCoF5gMz4qTu8/za
JhXd4d/vgogj8gTAaTHipg8CkzxWUn0iKdJUm9j+LaYZ3KldrpWyFiyt+j7nBJ+3K68+yJqeZZAJ
GlZLl93QFP0DksiijPG0FrvhpiMxR7mqe+PSxmp9+PeTJmjFFvMJGFUQrse8oe8H+vnGoQpQEY/Q
pouoTWevzcLgk70W1IgcRUqzXtsFzBV2PS1pdcmjWcjMwHksi5LEcAb80HcLlS2Y1l70d8Yh51mR
V1DTZOFcPSYvsmAEapRpEU/uzA2Xs+eM/sv3CRSih5HYrQyppCBILNfE5Ywysg37oaNl/9SrrbR8
jXxmunQ7SYUG8ECppHR87r8/BVEOtlBoGwzBXuewJuqMBix0El73iAwwFyFZ8FZVZ0bTvdakjvFJ
3D/aa3YdyVHWHIwShOK2r/BwEMGlD7s5Eg7Hcu8n/NzY4P8ILx+7+tXtC6k03YiNtokk5U41ZQlZ
g5wO2xJuoUyf04XrH7230fAAjYcVT/RZ+CP10KTAfGKeruP59eykoAnaIwA5UXmd4SHuvf09IxT/
LvE2OfqCnnotwbiQ/bfArOWLlIF1UjGPLwI5tVwh9VqC0LRzppdgqdseQWim96fxd0Vg0Ugi2z6N
dByFOIH2NAUVnDmAR7zkHVkGYfysftM+rwJ2GhgZ3atQNTdMcs4x+c37V31ulWJY9JI/PajHFsrN
GCgrzVCceygCUjwd5ZRbYzRLzezDU2oeuLc+QNFyczSfLPd59TQNyXQjbq4a2ndGEbs0WZLf9dHH
F+RnB3nC1iVO8OIVD48WrpklVOSGbajiUbaqfjUsg7W92/WgWvYGElgv4hOsikPm/PucR2hRrmed
z/iZcdQnyZNdFplwsS/OUZ0MetT3czSeZM4e0+PGzlp7I8eamZ5Cm+hMToSEDg1tEDAJraIuCLP6
khgOLqTlaZS+HwXZnq4SWjxHzeZ5aCyERdAlylECwBDEp/8pRy88fHzIii0rIrW0uc77QfhfC2U9
qE0sTlNtBiOeHgGyJ7IV7UQKTyo1Z4dkiqgNoFfUaD0DiW3GEdyhxrKO48VxYxNm2TAc6pMp4v6E
ZNUkvmnGKWpmoolD8hTmHpjQbTHWallOtrsdqCdJBim+M887FcEk305Xm23KKKw84gO+mn7gK4VO
293YHQY8mUFMXzJd2orZyOGaMKOvP6Cu3nB5hiDADZ6FgITDZovp5gV/Y2AfRoPTtUOR55Ufmk4H
WkmNqIFw4PJ1eyponStSxIUVXPwVyyDRaVgpxmCuY0u2Qya6CcDqLPLpOIPxrmgvRNosvGzUsFnE
xw1MiPPyIwbaSWgOsT0OX4kLG8kp3GlxwbfOh3NuFwuxHYuJB87j9/uPkHTCH9Q5mxW8yWDKHyUI
Hy7f5CRGBwLCyEf+Ki9zOjl76KTtngjcxuVOklxzKNbu71GenbMHyR5lmH1am4KvxYcaj3v6d9CS
7jzfdV7Upm6QffkFp2CiewGp6vsRITxdsPgbc1B4jpS1EH8SpbCms8wip5ilMW/ozR3UMgO0WtrQ
/pQCm/A1ALFDLlKB9rEa3ZIXkkFdtyFmMC4np7kXMh7BZVY69WCn84qPzLt5vg8kU4/6tfOcAKi5
N6X7zQF7b3+1ALZGxvGh+JeDe0hGGUVKVAQoiC1CraS/wBav0CSLiTNHS0rGJJlR+4UgHd4E7Rkd
ComV4Y9sa0ndt++Q58SGz9ZG9BiXPJoDSQMsOio+X4Q7xICnRH/mHeZ2dIFjagCO0Tj4pONUexvh
ERdQyBXtY4B58q/i1xhyo08QQv+T90yWeZvkKfUHwAuIxgI4s7Siaf2G1z+odaUg01gAv9HPGg1l
NrUxVUAnqarE2Prbw69mCgQSQuH7idzbwD4OUyFqtqjNfblE6Gz8SVGaSD6KGlKFTNldxk02qLqS
Og/rxcgwYCvAxZ0PiC6Q1gk61iUqp75jXtCKtwb92WE0f3W31lg4idHWUl69zGX44WwcMOXcYCUG
xsS3QhVWUkBmHpRnV1hYUeiTAvaQNfpVACpeF51L1UrkQfvxCu0FVkTu7fJvQRv2MyeVNopcUyNR
Eee/DfGibY7fNQhgmMwi7oL/Cnm1upbXbW03kbbdMpHVu5FeppycAXQ3Doy8CRzlJfho+jr050DX
u+Zc8COcG2h3I5gU8NbmuH9BIIrRmWvozRoBhJPjU0OMtlUkEhnhtz49D5+0ck3wbY5E+ZHSp1Q+
gwqnRMIQYYFo5qKgj5cBZ8BahBi2oKKLk49dScGmQq/4aT3LpswXLneUTobSVAkJTF6BpFxoEOOf
pvD+XCpsYfyVyVGyU+zmP6X7Ri5NK6nvYEC74nOCtApwCdPLxYSjYfLHXSyYtsxOo5AplUPGlfnC
KT1i13OwIPnLsR5EP7QAKkXySvsJfrx/6AoAUbdncGBcg+Nz5eEbb9sCIvOMrtF14QQMgpC/x/IP
SdsyW3bQTLguc6Vi6spGDdP3xmQdUYRHeJ3891Yj67q/YgBfRC/k+XH3QWqz2RS6k8OiMa3ThPJM
5bOSCe0wDHpmkFxztIb6xy0HEmkSKx3fWIXaXPEtNqt27qa/mpxuKGarNLLDVjiG5M4pYDZuuzk/
d27W2PMTS7rF5jmOsf6ONLYV4Ll9caxOtMrU1haPYpsd7BlMhqvahbau5eOKy0Ia9/QOHKQ8WfOR
FPjako7cBU9p5fwXDN+J/ERz9ZgJKi6gJw8FVJuzzsmqxgEWzUiq/iElajZjNHfRQcosOw4mcLN4
NNHM+EZirN0Su4AoHUf5TrVn9K3OfPcV0Fw3PBa69gsTiE7EIrxyCs6J0VJgfOsnxGa60CYaFd7C
kYUtNDsNqt8zmuyTuuYV5HAVBaXsaR+xlUqzPyIaK7NRm8TZwSStpNR+bNiY2vOe4IzW6Ae701Jz
Z2sM5jQRDZ5qIN2LVNi1wWVsp8gQ0XsE3VLo7HdxtscSd1yHI7qMrQhIwUEw5U2CfbAzQGTcPNBe
z+A4IymzS4neR4aPSHNp4qUQDkXv6yPKs6gFH2DroZW0cxe3yU6xewf59BbYuKQ9OEgsXj/dCdpb
fe2f2LKZUydk11lBcUD/DO/Zci3TezGIW5NBNALFrEvLqgAZvz4gZwyhnV0bL16Ewl+SNiYDlnx8
ulnIWHPppih/CGxp0ilPycRw/Pdr5Wf+g5e+5Mt5Hlm5HN+Yz6qZs/rT7U8t4z1RhfXoRX/2XL/I
O03vXua4HACZu3EahnaD0jMXSnMsfykPRzRK/OdlWUSHhJ4jB5xKGZuVWdnX56ZAMvvVPASotLgN
PwhDXr5L05rbjJK+oFycT+HEjdXuU+mUm1Mq7SMJ2iwuM/1rrC2wQcblMaTXSJ2Zo8YRznZKO+Tp
bo1iEaw2IiTqyAL5C1++HIorspSgGdQUXMr4M108lXIW54T+d9HJ7Ct/CAWbzRYII//+OJpRjiEy
7z+u12PNZp0wb1OEwZmiOJx+55bLkzVAZ0ChfbhHm7AcMD/ZKI3oHsiDzqOLHm3btGuqoxI3xwOG
+eFZ4NJryj7QH+iVgfwoLitp6mLOLIolCVAhzqkoukf5wGBn5jxg3Wes75j4/JdAzriB0p3g8f7Q
kirKYOt4lcHfdfllfOEAzvNGa2F/6GxrtHmxPEtluHsIGS+ZogLl9g0BWbsSriBGgN0FLZpOQhs1
wbarjwfB2QoCknS5cBnfut/Iu1Oump5vpmAljw09toJCR1TDusRL85AQf4U96ElooDwgH/EspdKF
7MPmyOevA9PL5okuwt6yL1ZqOsBLcC3Zq0gWvmp4MumcvvRFQlHwZQSoOQ8rdTtXYxW3MKmjg2Ne
Q8QpvOhwhh/I+iTzP887U1Yl+G+DwQbSaOIhOkwRNDLmfqmzzuqviXdGnY+AUliQPPZoYm14tUfK
x/0pW4RkmZhR1emQq1n8rFNK0XpUw0nB0mIItfaFgdIXFkc9Th+1CTU01CIp6KAmRAV7ulhUlT79
W16KvKbtQJmHct4NHDYrRZg/1nYNmRkP6/RanfsHp2ZTAvVaAhjaye5hVH9/eyhQh7qb889XEHpv
KNGRKGZWIOrNGPBdMq1okpwD4OlqpXjdp4jvcjtBlLToU9W1J0QMojMVgKdPqcbwJ+xM0oGkp8bX
g8X2WAi0RcH3szaDmMYX1f98b9xH9yKhIsndR0z6l9RpWgLWvZAb1sbr1RhJVjabE5OSklUizDy6
RTJd/Y87LDatxxRnSgNHn7w9tMcuglQa6aLeFfyT6scbOpGmwI5b6qm24Tn57mUDowWPFE8WklfU
wd0HpPNurgZ3ApayS4lyD8LqUfJrAKdbfht8GFP29YZbllmIhEQsH58wrPLPekImOqAO12oOKuDr
sl7hnOU3jWtJQkeM8h6ttDtfOLqz1sxhRGGHA92OPUWOyFSyPsUquKk/MB++vskTSvCTyF9Z5Ims
qjnuo7kAlToKPp3m1o1b/aIirm5Xaw2ph1hODtXOK01ySLlzS7cGQt2CfnqjhmOpepU+3sM4jD8k
Ctd1HExImUxGFMjzhGcyKEcaKpV2Wbx0xq1WyLQlabdHlCZEtfYoyHqqmDDrX0yqgaaNa+E+SudZ
vgshekX3F5nIXM69mIop4N9nkHGyvMmd24V23dFEEDkHDETzdJ49d55M6WvfS0SkK3qZvzHChoma
8/uvQie43EEgfWDbno/GddPjw7pRl1W9mD35zo5s1yGWuxOJTiMGYZdBitbK87kQ78zwWNlk1IAi
L4/Zgi2/uunRKXJMLstduMljuUQERaaSGt34bU2nBfLHMzp1CJHgR9mrwCRn3s5X0x9LR8+rnhwp
7nLcLEBVqtjhduSdVbel4Yy1OUbqK8qeUAIcyjXP6aGFJJCmrNulssaBmLwG2zWsJmWKGk7HAMyz
J5oNu0RE3lEcLpyiCVGc1+Hy5Y/xem86WIgDD+Z2czFOHfXU3bXogXqlJ8cCqVZRSsZr8/Eujf26
R07/0WsB9AXPhmaMYJiFYow4+F/mO8+HFCa/BUekXCbD7PzSHv0ejvG2xL5qMNPHeU85qklIbpiw
AReTvEZk+dXnAwNazG9HybF38tL9opq6ZPhd5UTZaUKXN5J+JGYhd71DKkaZvdCrDxR6nRUto02D
J3+xQ9twut8zXrKTa5xvPuY1rwN8Q0IiMVwkF+GdcSQQ0pmaayVr7sqrSbthR7sVkPXVwkFg2rZq
Tbwx99C/fCGWFaircL47cC0JAcN3j+aDvgQip+WYZFGcehgWXFbsYR/k+MxJVBxfR8lQF0I+ZZi/
rTjkheCzxy1FZOAc79BmDSy574Oq0Zt8Cz94x+ryrL6UEPQJ5LVr5oDJj0zYMIezrFptGPvYtTAF
evt1pqPE1spu4VtEVGNjKKjR+Kf03NBh35CP67iCDBsul6qvS+WrcRC+G3OnkS+L09HZUUQHhPng
WM4WpYaTa9lcxNmdHj/G9GQgl+RNE+IKQSIsUJt+zLBUpH/SfLRGzRDtvBP/2LfFEIxs8azsdthO
V5pCBkuTcwFq/OzgBbSNPmsRP2mtTnc/3n9hZY0VJo+YuB2+TNM92kD+j6oymNmJnCwMNMPUihHo
h72CpIbGbCKDZWCj9d8oUAymvzjfETVt88KYj5CEZdmk8/ihNQI9l+QqtgiiBVMgetaP+03WkdSv
ZThMLDt6ZSdDY4fchySjGOg/R6dOjzmWJ2x8JIYEOGjrjd5AM25QrCG6VzNNnnksFNyGgHmTNktg
kYLGyZOeL+8qcH62j0+6ivnLQRSgJ1MS44Xuo6Y24QhvNBDK1GIERw77uaPnWgkv+iuTel+vn+Lv
iaXrbjPRNxlIqxhBb0jNozLXjf9VGuwtvTk/LvUAcqUsqZ8vXLyFpqNfBygj99xo4fhUxctLo6bp
V9bTzIGH7UboL3JMkIO5gawtZ8T3ELVu3W7/savgG4GJ32UJtJy/QrSKCn7t/gQ4CdBMI2fSGGKd
qACCVUNwMmFInVOo00yippViYO0axnyvQWxG6jkYE3n5+ycDcOm6NQBr935wiwQkwUYDMBGZWbg8
Ch7H4wWfKajVzX0NlOZgGEcqDlX8XMKU3U20RNTfrQRBJyf9nr9PquSjk+mSzjWguBw9qzWgwRMZ
SxjafRO1EUBhNjVjfVxXEaNoOaFiDlAzRlyInWrhJ1f0XaEosjCmzrZ/hAM0y8hbr58rgDRl50f4
hS5FdY222a+45Lwzql4JNNk0aY2XZWYcDdG5lEtLlD+n0z4U2+fN77j2scHSUqWrVhU61Tjq2H7/
Jo8/0sMeXOdn+a1ZWANbTlj5ittn0AsannNmoDMWWR75S3jg5nJRhzNV7SSkgICfs8oszSUSp+/X
Mq4X39h7r4j7rfzycI14BawHMdgTB47kYccFxkl+0qpRRtAYwoCRcVgiQUYeu3b+AyN3HOrhDKV5
eWDGk8pWKRrtNd4EsC49WE0BnePXN10dFsWBl0bmxYsxa8Y0APJZSXcusXwRYmi0n/8unRmr9Wji
4Mk5IF02lBb5qB0EiABcjAnG6CjlnwTJSmvzutoPQPVLeNqdbxoOfSQlb6+gkarc8OxLFpRbjay9
6XFPXG0UdmDNLBf2btlp2GMyPxlg56rywIM24h6/mjkMNG4jf0aszjJfsc4PpPjlYztjAs59IJ36
aLPi8l6u/xKLDyiRPTZs0IiXMdhNsKnz6Ovu7xka7WVnLA+gOCShlADxqeoIv5t17a6SMAktk2hJ
fjqGsD/AcNxb534Fzs+m7BEK67dXLi8/AIoCDLLNj1Lv+7c4QEF3WQ+3P4oBxHRgTgHApTICrjp6
2DO7Wqg0zzN2ngQvmwnRzmBhfpzuyWxv5oSpnq+dWQVHc2sqUFsQgcG+lGLI+F1+wu9hs6jeqQWf
aOCbdV4y/laJKqGMgpaKIoYsaRuJnxeor4gfHdWV6Upm5xkf8+fkKMR/xsm8F3vG9B5bKGaMIEZU
F8R9hAPGzVJfR8H8tvaNz9UM6+luhxA5RYOYmxZ2z2AXgX5UOFtUas5g+3tkm15AFu1nC3ob39w5
Uln1uN6Q88DjDVyC6UgOzkC8OvoIj00ZVL/k/8+LIjUZ732awM1IdL5wx5SPk3D7Gxom6vx7bWrv
5AOymgA80BkMdMtK6X0SvdIKNLHF0MTzZTdgCDseLsNKC5q+dBYk3CFLfooRXg/ROH/8OOl4rTvC
fLKW2wU/WO++Pst/liKeBO/QI/yq8iH27tIZJm1ddDJFnW5KCNjO76nztiB9Qar1xO81ulcBNOTO
XG0l3wD5/ajNAm8fYtxWmiIMleipBXnzxaBJ74YRa/g+3oiBp5auovUNSUCDlnAuGM7x/aTtbAqn
Z4W1hLRlC1UnHWaR7YMfn5JKKvWPbI8J1jDIH9HqonhbK3ZuJzrquiHJXqj7JuSu+tosrnzx58hl
3xetyiHHig8KfCEpfSPmbFZQDX9N47CZd9wEPCV76ToSs5KAxI+GlB4yc9jftka3E+R1Pv/J7Xmt
0jgcKW39qv7qGb7KRo2CilOcx6Gj0rTwTmxe1YPncijh2GIYcK+txiSmZmXMimMx3pdp7pbkRZdg
KAKvbXWEqmDWOP/BGLr+S9b2NO9DqInEkeY00bgluY4WUbFLAzIL753525Arszxp73ar/HbpkmJg
GZ9VZLnDWOg7mGFvR4AsYFzxWMCtvQ0BG6q8H64zMAQYYTZnXkET90SojtLZHpTfPzSKjz1S3RkE
Uc0Lwzcr3C0fgsVcU+e+4+Qo4C2GWVN6wTgzo9+ZnedFbO5B2Shz+9ZS4W1SRqK6u8UzL4g4pjN/
VqDlGNjf2kxwg2z6U8Ju5uOIP1GuU1KgS7Kiq0VTihl8/7ALxUEPXzabzyy78dy7GJfZL/bRVjTb
Mze6d2ehCZgRpo/zhrJnweWUaCxBrf0ih7IYmRHAeg2bi324Uib3D3jo16txrZ1JhIfxj7v5zOXP
eOL5zPsqefLYS4qPktlPLx2NcSs66RVGqaXM6bOZz3rFRg0ioJp8Vj76K7MWF7fMACWRn0h00CXk
eOTUUyLNVF3rUMpJkiilZ51ekpDTEYgZ2CjowU5S6O2pfEQaEMlAsyVqxbSZ//hwpDd5Gm/Dzntb
idHeC0owaQbvmSY/ZK7AcpddlOwxIXZXktiVTVrZ0pkHoPE+F/C01xIL8+1ajtqhP/OyoGHhGyrl
w62/+ameJdXMeUpmoLo75JhElss/7ufTpZKNMH83Cfr6Z+4bpEIT0IGCEBQIQrGZv1hwKsbAreCG
yw9p41x4Oe+QGiyeQa+xD9CWOYdXgW8DgOU/awwi7ri7Z2VOjWjYeC98x0gH+NodEutVEb0+qdBl
uRupkGIaxLg5DejlCZdMJI3HxREIsZoylByHpmWJSPtErzH6wCGBIzrMBl5KjsWyX0UkSQa8gVtx
YWZswJVmAf7upBFKLo+dxcXQvyH2iQkCIpVfTN2wBhXLVUNJdZRYsBk1OCHLZzookFYd4q28qSKp
XGow9HTMBmCUVFjcD0ypgX1F0lYxTaUW2CXChEiMx32xabpsEeZzRRH6aqB23N1LGExZkjGWCi/Y
jgZ9NU3KW7erELvI2Vb6xLkVO3xsS4N6SFi5ayZccu4S5dduz5uSHqCUrZdqHqM0IjWG0i+BM7dI
+RcPCUOOQ13t4ZonKT4VkD8IKSoxK9nk0Mje7EbsEKCGpi0GjBrxfm6YGfJJ+xAt9OM/9ttRiMLd
socMZs3M+e/TU0Hvh7WN0tXWuYFd9+HxA6m/nBjTYRJFJrWRfgPUUJubR7FlgP3xOMaRTDk+VrKm
pJHUWBwhEwH42hT2VdasZXev6zWh304rXiHpfat2wg2021S72uzqrvqitnxHPVXIJDzV6EgjRvnG
9LFLUk3WWkjlHL1PNost7C2sCQWOMrrzrWHjC/P2u8DLSjh6L2DELtdEn6kxikHD2O40Y9vvzTqM
RkHtj4ZodCHiDbwBt1m++Cucb2jSNAoR4d4bU2+Ohm1GLouj7Tn7+6R6vuOpf6Qlhgq8wTr31Sez
7h13do/3pi+hAkz4mfraay4XHkLqCBoFYWq0kCd8ax4R2Fh8Z7veZu22kMwqZNNiaZ0f4CQCrg/W
wamWbirQwQZG8c1GKlt3obAZc633xDLo5oIyn/QOIJT1PAEEFXLVN33oYRuAZhaDp8DmHwMscRu0
6vxDqXFhm7y1le/ffxW4jXmnwj9spnkXJBbUMEd1Er2e4/h8M4FtI0w3Bc7/0EdiVSzqt/Llsd2C
OdsEVU/rX4AbMzfFFjx4LGoMwd701NoDba29rAmxE7mwuwrpC+Ecx5pTh05uYtKTX29mo3kGftqi
un+LXe++BWsDuHixEX1w7Nshn3woh5xYtfgeF6zthfZ9M1tlBTleg5+TMOx/q11lAduZRxw4/Aun
kk/IBhWugS004OjijEwsg0iVvIAYVd3ifjs0Yz/E7lxTCnD8OQfTLI71J3RqgP5BLsKDS/Ejk/zf
DPIpUazTcGaUpfhUg59vAikGkv0uENhCAE+3wGX1rmwwAUi3zI3X4p+IYpnLqz+YL7N/1VnEezOg
Ds9ZBhqw7IRPW5Oep7VRRaJmNn+/h9jUKRryGWTplcNvwmvwGl5tNzUayfZa/Y5v580rEzyJu9HB
INB5bLhivYVUVgqIpUuT76GhXAaSpJweodnVqsX4W6U71IFFzDfY0QdjbxiVcSEXfOigZRB9GTYh
59CxwmLJ/7UsAx22LpNYzOK+vXWROb33B8d4MaTgBaQT8kWmpgednIaIzcPl9zHmOPBgMv0cjaaW
m5W8l/4RUbTAeM6/sbcJCkfLWjL0sOhI1fybTZjMIut6qGJsUuuIptf9lscUBAZvNYPBERQqyMyf
8cJDE85IbyGm44zExpakeKz5F4Z1G16AAVBVrDCU0A857uG52qqKWnS3dWvjeXbxD5WN+11lrazo
RKsJBc9pY5WqdzxS4rS21Y32mdOexbYaRaIk3jRHqBPDZ/W7eQY94O3fZVKVgIyfdaiAaQs8c6It
bccYDmsvfq8/EsKbSmxNWDMTk4m6Kvw7NrrTanNMOTkQibmwAKaB1r/qJxjHPaR3WXBaOeCI0wey
FI/dSoz+e+ZGLxePjorSsnWE8m5KsnAp6FHVqEQaTPjQbkuZMuEf1liVQu0Ch+O5vukqNuRjFlUK
ghT0eisYF+ypgbeAnT+uMuYmpQUiBlUjDtc/BhXzSXf0usGcAuwtSaZLL7cUMCxEyhnjQxj/ssQv
Jnp4x2HqcRwnVUGE5GF6L9q6Ie9Hdr8s6zU9KPOh6gHBkIVG5B9PfPdhh7UbtrwAT61QVqSyXflp
sWRyP6L3M6cI0GUsA+myhJTEI159Niy1A4PAyDQfrwA7GJOKYRSd0QntvbUAaPhw+eTuQJWRtRg3
BDUIFZLfweklpuTe7uBdOWatZWHYZLttSHdMTOuP6IGWwkbDQ4qMTjXlf3Gn4iNs11P5y2+AGCls
jvDFMJqg5h6VCxMtf9p6B69Wv3iyaiifTErU68OAN9FRHU/stxwQJRJJPO8anKbRkGp6b3kTx8k/
H7h2oKE55XB8Blsx5wILNyta75oeOVZ3Uc6w+EC2kyeWTiW5ZBXBq4lrggRYs2Q9rsrsucnZN+/u
p7gAzu6MlpE+4JNga7s6XpWaolA+sEecj3j5ydnwir3GNfS5f2751VrRWPO+2xY/D1iEV+y5bjCw
SkyMoNtGDoz4KhL7/wQEPLQn5W8bIphu8I0FTeA7j1LVaZdgAnMJo21S5hSaeu9gCVTrnFSo1+sd
j7C2uX7qccBJoafsLLGgasIUmsvrimvHqY5DoHHXjIaIs2w7xK0AnrVd2XtD7gQHvQ68jT/me1ho
O06tYMY1GbHeEKAV8CpaGHDE//UNPYJ1O6qKwIksUDb6BI7ISTTnTWKwkWw2oU5/YtWV0xH3Hrb4
V9t/3SP2RHjPohmDYcMy3kptzJtoLHe9MHEXs/vfJ+AyvjdhIrAef8f3FJakNjZKFI/g+lBcI7Ko
pLD2zT+ZFVVWe1EolGXqLATZD3mtz1e1MJOhZ/3CN9DinB9LeNgbgdBKOSxmZEgJlN3mUJ0a/Wk6
YrSs71Nqn3YKVMM1cL1/sov1b4lq3NM+UPvYAwBDzyCoCbZUqB8vq8IQX85k3Tpm10MfLY4DCzbF
+DKHi8cxLVjAbEAe75IaBno32Z3OQsu0qTEUjIE53LrSj8ERNRljXgN/7zFm1tHrIKqTudhXuSTV
zpw98+dkztzEK7OhggKB0DgokRL6vUJSnPHkncR9gtDuKJi9N5Sx6ZGhd7vNxhyOw+v5Ul8MaPYN
nFYGSdiyMD85DLvTgyeQOsACIstGS7RjyRlWrjb7NdJ28Y0Gx/mKNXTiE7nZ47puPqZ5Zxxy/WzN
jxC6hwdSLp5ThliN8HDMM6Oac3sYkqLwIN62V0roaZ+M6umaHlnCqhb8eaXQjjj0ZLIXS/Xt/X75
2150ayYQ8pLim1/IWPH4ZKiDdopSBPKgYoLJd+WuFjIP+i7kcnbapHIeMz8dn+HibYi6O1guHWVM
TwILAmARthHYTyFroR569sRoNY7m/xG/gRsAaNm/4vcog8o8ahLsbnPbo057Zkl61l53wPdX5zWb
N4QAX4OotuJA4HeLi8/V1/poINivroYp72w66MiYlLELFzqTbgm4G3UZ8mekNVTJyrwe8gr7/CPN
AuKMiG6hCVUUS/RYHVqZgzMh0TfeNx5hnC2fdsDnNzHj2iSM0vvjOAkb5hCqaAoq6JpLpainNJwk
W4mqu8s2H55rjoYrdfs9G6WtUbd/DDt6wF006YK0BL2vXIwjQgf/vtBgVxBxKHxuHMPiNJY9guQt
FSXgkU2M24Pzl5ohdyoFRf2HB98fhZc2w9hXsDIkBDRl6WmU7z2jrFfGYnQ8AmSud1hG7+DL7AoY
6p7ILXfkQXG1s9SiDkKfFrerjmH6wWMVhldbNhAPEjx6LZQn3Ae3AtfiZB7pZXrN3gwC2KESX8nm
aEeXsyl7X6KfHIeRxY27zus9skQsWM/cVeEy+jVj+xrIYzyrZs9JEB+m8hi4wfUyszEdJx8Tmp2B
mtCErQVuoA39WCDF6HtfAsXdY2UvTuSfgOLWMR9yL9fib/+pFlWBk86HlM19qiGKNVi6RM1QQgND
v94+Os79xQRXB6MqFaVwlykHU4OmD3kFd1q7W56GWbRnx3YA8XQvVixeENRR9ckfpe6zlHQaOjcX
Cixhpw3wDtIQ5kH6CNxXy3NLRrrlZfons5y6plGRisfkokAyp5N02grFkKDa5J8hYW3J0udHsGjh
FVsXdujn8Eo8N6uz6J3TeNdJ1CNc3fkb2D3l4ug9IXjsQRlLrqm4u2rXa6wBR0YDGbo/CgDLPNms
padXYo+f8ziVzS/Bm3jlYtqwHNUjkKphVWoVn7KZLX7pWnirpEWdhUkp/oWQHtCtZGCMKS1OVImS
1neqry/w2uxb8qhenCkrme9ykgxVZq/dQKRwrUwrCfATjbz/J8p8B/xddIO/IMg+hVEn5yrya38h
UIJmpnKeFhi8Ky2uf4yh4SDG8nMzz6WyCyOtLGHsTcbJBOEV6z2zjq+5J9LRCthPm43upG9YMNOR
nIfD+jmki9AGO9W/zoG4GIwp4ykfWXTK0bE3iIRuojiq55qHmrxWdOkwtx02czeVWHia3gAo3Wl5
zM5dZ9zfPsX8oDODIzTSfjWUgUGKDgAMZluCKvBRRKPTVQ6pKdt8xsK8PL0NUcn2dW2fUl1tk8oE
vCWqu9h4oeHfV91ZB6s/zOqs9Hip3jEtxKSCSriAu9kSbimPswgk53MOmfDTMnUSMicUMiKrnEml
BhQJY247R1O5LWo15ygnO90DsyxSTATN4B9Nw8+UP0ICZVQ4QYSuE0E1TFw2VeG8uSwKEJxAACrn
reE+uO0Aqr06Q2nj30RLpXIphORyOkwq9Maoj+K4RcxNnyRc+LKClZUNzEO2t6GpQ8qXQv0FB7My
UgwAEInXDDZr8pNFt3s6s0n8qzG6NgN8vQsY2Lrtef12bceW6my+e20VRmVOtqmnx22Roqc0ULK6
2OTPqooyQXBEuiLznQPq3B/xwIj0YlxLiMh554lKEcm5im12/xrYsl9aKhodUsalucpj3SQvt7ZR
GIt2lhoqS97xGfLwUf3hjo6zVdjQZA3Qio/Dmtx5AQOcDDIuqre/SX/oOmxKUQw6rFMoRw4zXXgo
cL3Voao5xMCFwzTs153zL5oJQDv4ENgpDDynUgzQ93xBcnFsTPazyuy3KWTKN6KqNhPIp0k9m/x2
wRmyzKGgb7z2SDz6rLRPF693p/UPoiLkORgbSvMZS4UCy+iN3m2nrPVaElSwcmhdEBBqYIYshdCT
WKrrkJHkcaCbt61MFpcge6JpOUriqcQX+9pfvOiUa1LMax8/cbA9pSbeOzWw5OHFQ0sXDfP2nP23
X4QFCbie3/0/eXGsgxRUzg16o//M7jH2aQqNSoqWgKlZ/WVV9jp4yw9Hxn5ek+DsY1tynK8qU2KA
mLtC3/kjQbsAnN4FKT+sMtXgI+hFHopAFTu6H88V52wVI2xM+a4Z1/xNowpp5h1zDT7yyTLZU050
t5gF79OkelVAHI6VVaRj0IFuNJ6VkZrP89Zl1hTFjXT/PeR6XAqfREX8EHw0Y/4qBhwFLdwTOQX1
s0MglgqgQ7KJKC5TaphmY+nnFDoaQQ/w9SciXsu+9W/CNHaSJk/iFaBk4FOHE0g2qdxJ5+a4EypQ
DfznetLOYYMYd0hN0JiF3aYE7IpwTa0HLSaHHmi8W8nRrcejw8cCHgrh/LPwQSIiY7f1EYVj+cIO
z/Q7u6q/1Udwf3NVLsgPWd5QzOhqH0jTRLLfGuGPgUpJ7e3kOsTJoF2z+z+p6XkBpzi5cIfhKJF5
dtfgKAsB6V9xGfi8CNparQ1OqndpwNFIWzwH3wE7K9Tc8pDuzoLc05TDK0jNC8QAqeC//AHC9yOl
32u/xdFC1bUYluRIDVl/M3o5RddnH+5AoWmvy2Y650QkQA4Rc4Quwe1OiRU0rqpAi2dSYe35uN7Z
JyIq7YV/2LRNPXx9wlZvKdP3lgrdUfhS8o5bzX8ExEKRYq0y+hZoQeau+cRU4yeFFtl1OTAy/NQd
t0Q0JeoFdA53NwRcry29kIJMFWIZ47Pkq3EvOds1yc9jBs/tLwNgZ/E7IDMLk9l6rxUf0ZDwKumx
24k6PHYfx4j3KA4ZEYDLwgLDcFFIDucHcFu0YotCqyR6KLmfHibz3kQLZ8qqzoHmFwfK6Qc+fvdF
a+/WgHCP9rvjmosVlRKI66fQiu7D7cei0r73c0ouhhKp87sr9dqBDfK99u5J2aeZ2SPYaWdHXCc9
yK2SZowOOM6+j1gGUHUttcNlFVyMJWjpb26qCPexOBWN8yV5MR0tDIAejL7DexsYwek/2E8WRAl8
B7+2TE9JyT23RftB8u38YveeDs0OmUjaFNNf6aceKrGxRZdpyt65LImR/qFIfOUM00VTE6NMy+Es
DBXUyx48JeA69c35tHfMJVeJcXx42+llGCLp6jjPKhP3MYSptEch2OlWn6PTkcWSp+x1y3vZ5dQx
l+IWIopwEok0TMj3k+csNK94yI2KocdODAfcYpH6OEDqFQ/fns/8c7m1aG6fHvzPHso0/H4Vv7Xl
IhlSvXjDeaLnJOYoR5N7XLexd/T4Zs7wE9Sj2ev9CD1rAK3w0D8gj1f2Nb8y+PxZjoXIVXUqdFel
XRYvvCh64A/8iCV/cq3+xIctp24GAxFLBazC4etSt1X/YEdRYC0jknbbfkgu1WDs8DF/DT5VMJQo
UU3Q5BKCQ0ckWfyFY5/cvdxc9JInNZdqhbK+/1v3ZuTsgVYWaHNJSqSLEaNhvhV71FZJfCcboUbA
DKpyEzs6cog0ZJGF6T4OoT8D8IuAKcnFWrpwstcG1DWNskixa/QzCpDVMp3Jw3KZ5bczp20h4op2
l3oXC93y5uDk37eQF1jRhTVpJCX0h57RNXgnRRTNbLeZKTEE9R4CErJAAAMHAuAcwaV57JDcIO7Q
OnKWHUnF4P5219AL7kmoi+tPJpdjePWTG1syeMLbmL6ICevDestkbsHPLykPNiGAui2ABnezT50/
RBkpbQB2v1yGxpjvyontIySr/X7HW18Xs7WxfSo+Ou+auufH0Uf+CeZ8MTnx6Uy88nXJUOcwo5kJ
7HnhnqkyQ0ptejVLNdj9w0i4San6PAjKux+hH3NB1MMJBYir+YxtnSHxv8eX2ZEzjZ2tdS+PRwBI
3mrzPpS0grH0Gw3eaWr7R+tYkRNgNCRQJiC1urYQ93I9wXo2b7RdnIn2cDpScE6PAe8/2vO3oDmw
3lAYdb0otHn7NY6giy+5/zBxeu1cCFJD/rAdcrGyXpTfJB5TCQ2fho1p7IHi5V8VUt1ueqTBXVdU
ObMABIrNmmf4EsPYRkuz8VRCsyPIEWFSn3KCAff70mMXuQX6IVwMpAYZ0m/0Y6fj0hW98pG3NoZb
XJPETnVxLX3Xbr8TYvY15rnWf93YIrASIipHPTOv3CtZWkeHSaBU2n8L2sgK1NuNLOnp57L2DIJJ
ySZz9u9Po0AnBhOidQLvz2XJAx4qGkbAUqceRQ1jdCFSUrIOwDCfkefjjTJo6UgdmoYsHpxVqseA
tWIylAg7MTqKD862wKYdfw6cCBKlfEyK/2Rw0LqMUJJV0FN888kwY9w9/+20qMCFqSkenGNLjLs0
NrgqLVxtds6EAO5Y1XFOCnXw4+YvSXkx14NcHzbJfr3L43l4KcI2hQn8rW8QSXjaiguXqaSCXPAl
bFpykSGceXpyHWyVibS8Pl/tL7fjdmx/+9fXr2XBPikjTz8RL3XOrB+BidjOpVbVlhABU0NuJ+Iw
rQYEOrfRn2V/k2b+qsfwgjSV0zyN3Uo6Xlo5lVdK1RCyE6vQeIzx0+rvXmWa8jZb7FVAesb0Lysb
D6iv3q3pLV6Oc1U467qLJeX/YMUxFwxvpemQUmH6Uc6IPQeDzIrGbubrz6PSI98vu+5xJ9zLVmC2
tDl2Rjj1G39tOKItxw5Nb8KP3TfCCb2ouz2rWNKdLSgtvlByYP04OfFfKEhLLx+6cunyZeanzOJA
IQWU6PVu67apVKmrRyYrOSJ2Ip9eD/FFU7gURUBbABoHiE1ZZB5HrA2zOqReA0EEoG7tBHkAoXx2
b7YYhedKbkqFJMkTe4/ovZAQPbBsYbkjpiiGokd3FFE4/Se9wUGZNtoA7jjnwtv2EUeY22gs04ah
3UMYjW+KslDR0Zz9GY0EjD4d0SF5jDXIgkrfIHDV/LN2xtIOrg9HBplztlcPg9JVezoZ7UnDN5Hg
GzQ5AQPN9E6KbTA1FSKBFDX/2nRs4TDlc3VuhTPuz2Y53tyHjmNZ3C8uIujUyS4oZ9hTGuJ3M1VK
8kc4ane6bo/N//oLUvsX384ZtaXl5HzH0zgBK5JD/cWKj3YV/XBA9Cu7XVO5XPjDmSr9WDFdQPYf
gaGdm6frWiAhNu/iX9W3KmlpyZ1Knv1jKBXLN8SQfV2V1a56xYdgEq2aQToKjNlmpGqNOIlSQMb2
Q2clo1wn0ZZ4/e8f/87yCLXcGs0RsOWP8eqJNDctsaSaomp/1cZewAbNTaAhrcM2nnTX96gQHlrf
bT4dK80yf+3TsQdMfM7+PySbqFq4EqeIi6WZSd0J3FNRVzTdjm2r1W3NIPoJYkx+RtT0iUsQ5rKm
hcK00Kqfw+giKGZuyPT8anZHRTyTOFGz/Ah+th0exevSJVORJVypKl31KB1fMX5MsL0G4v4cWogy
oUjDmJvKpVKZAhcUZJhIclk25gJp9xowhTBRo3bf0GLoBTqhQk50/mvF8KYnZs2Bzso3rjWxOXWp
93V5MckRQ4OOjk7iEtNoPjdwVBEitxIJH3tTwsgoLka0Bb+E6ko1Z+275AWBj46NHxCX8dRi2LIZ
aiEeru+88Uyn3qAfPohDx4c/3iQas2+6qVEiCn+/WZkrwsxrbLxnfWzMFVnu6APVw1FZcLvZDkUK
FzDZxsY7Z9zBW8fs3A/EDzo9NU6JHt4vriY5F45oS2pbAJeFltbAUSkcAFCmfktck4aOp7hnqbUK
VNwYMGuleliP/59w6Md8g3gakRUrF68HcFqxT6RN9uy9he65oCyQAwIlEGtQyha53NFeV6s9CPgZ
E+wyi7sCgDMMocWmmfRPW9YtWxTknvoYFT72FK/RTo1JjsXoll2DYojHTKq0g4DTQ+tFagYKNF3m
e1Lsd3wYXUr5h/T/OxVqzzgIds4M0A2LEBL4AvDLfsWRg34PDaKRzBXQywkYZPtDtv/pdAvDu5wu
kPH+yxbjH+nsP4MXqTWQNhY+AgPEEggacgwwslG/HzgX7KYU075FgSmq6ziwkOQGY/kTRBVI/B8X
HFxTYfNVcOr4ypz7xSBtxehxKnDp20R3qY7yklMDEbqD4M/nOZgi2c3aYcMzRp8AKSsgDIZ1moXn
AO2iJMFxM7nQ9nyf15to6WBEFUJ6Cm/0mpvSbcV2D+Io1AhQrgBG1KqllGTRWvx/T8D2Qm7GxIgF
Izpw/g5UByQkWJzk8nCoELobuAxwFNXjNhmZJ+cxASvvRbIYzc76BQqoZH07uTU0KmsTL4ZNkHd5
3DyWt4bl4rJLKPTjLim8r6SS5DsLW3J7ibFRNibAEpxBZWlyxCfBTCu4GcK6TpBfLRzUxPV+XVSx
XI1fY2aj6mj5UqyffASbd+Y8jgWNjTCXtupziSTxFty+edAhcR8leJ0diOZmUxDAG4OeAcXZyS33
XXUqfEW1o2t+uzJtia1fw1fFCz0mw3nlKi5PL3f9rskEkTteGaP1W2cgGR7DlR4sGmDcTCCY1p+w
/6oKW1Z38Dc50PE/GoD6st0U5vkrRQ7chgbNyfuVKFxXB2q04qbxb8pu9ILLEUK3tyDzwJyU5qpe
Q2n42j9Y2pQOvKwxPQJb0FehIz9rf4mUedVddjrqyBMNnxNomqPoLipZmYbnDEotnUYC5LoRnVTR
TxYELbm/SWgTS+gJ+lYDM8gm4rDpOTAWyvhSv29JVMikNIeABwBAtex/M6ADOvkeHjRz4VggUedo
nMgjF3wVvQBTWGtAbm+i56qAkacfZWnriFCJjl+4Zn1UlAX0fVZCV9CkoG5nUOdxUXuE6e08Vfp1
VgKAxTkLjPGv1RcHbQaFRHsOUevfZmNUQdshEVQFW+QnyqgR/64NE3zGu2fwAgfhVBj1SVPnZrLC
YTjLH8N4/5J0sNcBpzLZ5XvlXd2IauN57N++WqPgHVyVNuazSAK5RiXdnlj38fI2Jj/389L0649f
OmkaSBRJwyBcbepUqK30ffJQb0uKw94AIcVFzAcfGt46h+jTsSu04+4A3xcUwr1O0toHjLuvHMka
QeT/CTnZL09OAMkgheUTFC2Xg+zNeqNjwwE0JmBMDGfCmIsk3g28/hPiKgz/IjVq30knfpnbMVE6
UU3UBvYbev71zO1G1BQawou915p6c4ixTAw6TDsERGTryPzs69VTfrYPWVdeNQANf11UnIf83OBy
kDYFUZt+TLB9SjINlWVpnedAsHtYkZrEMKC+BWNo+yqpoFmOCRRlDz4o0yJUtBUPdeTXcRcH4qkZ
d9JyqH5YB4xuyQqbliNNvUGBwC0D45Ki11eZsDXNb8PFWfs7qSSYWZyly14K4A6qWEcDU4Ni7YjX
Hy7rwul+47prII3nu4sWPv7mEAVDtZbRrF70Xu0wOMfpf+BEfvOBwlOWYO2jnDMQwzq+KHgmnBSu
R3fR61MnQwjJ+geFc045qwyXQUWpast5WrQdeKp+ciYhQRbgz/vJlTBnd/73jYKGtFq0VZplpK3l
fvxnP/JjGml28Uh2h55ErygTMhzHFs+MvhrQ04/GZ/T3OI4UZ2TuRUa5FRKR47262PI0oUOunBTK
rfgJTt2r9CCpD1c/sXxA2ilWK6NWLJYcshRThnoLqTQKzuO/hN5F2N06KLyJz5kZDm4cfdnMlg6r
8HehERQQFenqBhuizOMNBlhchDDQoLJrTL9CdoBtVl7P5Ll+pZEhFizLQ/3ilSQ1PY5HIWWR5VPn
Z3zbKieCbBku46Y4XAxuGEHSxFzQptZ5K+yDnMAmk74Dm6MwRMITK5ph9g0WfZ4JOiexFrg192QV
Sq4GUJgF83cMCPABgoIIALZ0XNdrlBN2YwF7g127KmzoeGXsOTNwNOmdgVP/L0xrjgaevQ/b2cY/
7lMPJlS2q76p6lWAuaXVk6PQjMAcvw/0UPixSp90LkqTHfFEO0kCZSpiGJwI648J1AhJ5KetDHWe
fJlPuGGEdESoZt3bijWWbgvztY0KFSXbf6PFvuBhbYBisdhbXrerXNmEDyR59BZpNsi+4myiVypE
Ofz/bQlBkPMQNOr+U9gGh7wAkrmVW6+gMuUQ6kxxi51Uy6lHJA9y3ESrrABnvqMEHWOJvNYuMeJg
mEdP5oZERmujxKYz5Hicr+LJrGDrC2Y30Jm/bjyTu2Wi+u+3+HWPctSxdUYnH0kUz7UkhR6kgnJE
sG/cyUsmvbZbxLfNdFGMorFUSAocGyLMWlSR7r2rav9HTLhoE0phC2u0ZciNvp/QYmm0nfqH8ATn
qW7vrAeSRiibTWjmTeVIvwFe4ZAIyYqQTjiBDXxDkW6Pndx8kwmnPswuObwidtMCYURsC6iMacXq
nFcTOxV+TC5RCjziiH49IMvwsbTaUR6w2jthNntV8kWwpVUp90yzUJHD1Ix4/pEXk+VK3w0bB5ZX
tqybYSpU98AsBUbDSRym6+GH474TzAZTBmn6i4viYZHv4+v+Bvgt2aM9lyQWnzAgtznTwmhSor3N
5YLZcTskCJPYYosVoR5MfCQKK2M9FmpIGO8rqMxq/6eB1B7F/XApMFGURE+FvCrQ9JV4H1E20RDX
M4KlUJKKxuQGtku8/QJvBaG+yPMs1cnh/3z3JvPBQBV1i/fb1YXjKqR/9J0t78S63JoQqrGxfwVW
V22Eno5bgOMay4lPnCpesGPThrsr/WYA+PpS0jP/8uRC0UN7pymWhFh1mWoZFZsIFNC0ZstYE2O8
k5hQXcseeUx73oRgvyHfuCvQNWcRLT7Y4lqfI8hOXtW7DnWi1/h5fNnOooBZYYFNCRHUmbDHrq8e
jKC0RAFu7PPQkxkf7qcA1HXb26Ep7j4gRznlnyormBs21OCYpGrohqP/DL77BdYa8CF6QnbyWVyd
nYn8E0QIQK0RfnwxRmDAl07oqD2nfmHkdei1T8L49GLe1UcbXGh9e+Nk1hpSzx4ZVoadnSMlqX94
GprLFpBwDYrwmxeyfRldi16FgeLtw6cGT0Li1JoikaqD07mHDaup6v68Jxt2cho3Na32Xzgo+22F
8ygY+OWj00w5d0hL1U2FZr8wShe2ZqRBlpPEmOyHBn+xbTwlDZ+NP+Vh5V1e21/C53MRwJYKb+uW
QpJSju/sU2soHJpKGlbyhnh266oai6Wjiltk0QO3avtAW9TUgUJBge2WBWBofsk0Sxu91VqcMojj
OUgXX2bgQID8RHWVydl14E/EGYQiIC2ZeS4oEtQe+3RU6nkvS9ZBpx5Qbinn1Uur0JuuJrDrUrKG
vVSR2/P/3g7ffD87TdwoEZ0F/LyD8J87heTaNdYRMH6yTNkqOkDey57DYXZtQlu185oCkGYJ8pTq
ceP4jKmnWSeJWEJlGUP7e0sOyZtspGA+wLj5iSSSayXEuZkFMUI6ThCA5A/s2Mc6YtguJGad7BoS
jgfx6MnPqvdnps5drzc2MbM1kXqul/ZO13MrcenX3dAiK335VnMLaeCiC5AZZte7WlqJURJquxOp
nQ3QW4Vx/v2AtGoC38bSYiXJXJyk3aMQJ8oOEI5HDk9wpqRA4Fy6Ok08XaXgW5Wy0FRFAhvb/0I6
UTEwjm4wJllgJeMNFIWZNzt/1ofjzwd6KXtiZQeEc5Rh6/ZZnQRN1tyOiuww1N3Ihfse6Zk+PQYK
jWg5ZMJJWAHzI9ASDa6S78goyUgtOQDGXkp5Br6FY9rIbsvIU+3kWQLAaILCfGWcgtTkbJpiUldC
XohENLSZ/Gf8qjsHcLQeSbcXdFBlolnqFpWMIodcHVoULEPMxPr5SEs0rNl0ZKTk1qCS29DLrNUT
h2aaukP++unlA7AgpUBIxafcfxckxeEKtS2pVBOlHOKq3NWoCbD50ZnIYl3rdZcOPDCnp8ormY+S
C/BRRZy6AFjb2bYAG7blPXlA6TziKS8wDpjzwezb+G5IagDpmO2C5hySht3EADnjki9+5MOtClET
2S587poYrYW1xAzc93m3UvhfE9IxMcbNKYxazo9yRY0yjn4ULZX9AyBya0EuNxIAu6RDQpK4/O7H
ypomsxbVB8CVHvdpxJdCz7t52oS7rc8wJd8nRLJVhe+y3YMhy8RwJ8y6GrVk6B1sp1zOE0z9P0Y0
j2NTSqwDLwNJdCv/3kbDKtMIY01WdE9z8R3/eA+smq+P/Gb+/R1xFgoWsNvsUfDuMEbpeeFLpYhP
EeXrZ/kOnSRhVCNofAsUWdttaGKDfq8CnbwMimdgxm4XDavmbar6i521akUD2gzgCJqI5Q4kEswT
XRrmCn6vIybagTWQIFQgmGzowek6yB2f6nLNB+0iLvP3Edzhu2nwggBBlEupJBWGgYJRLOTwYg63
Ppkk3CS17wYiO4hU8CZFKk6CqxcBanH5mXBd4pgO+Ozkp69Wt23Fzf+Z5k6O/jxoEDI5lzqy2fh0
HJLQaHZ//UUGoAitrjChKbgBKh6LbzEaA5WLCDAqZ+1YqJ1DD/0peTFZ8VVVlonEgL1Bh5dRyPyV
BeBJq5kO/fHhoZm859zBvIZpEhi3T05ox+KcMojARVB5jEqmkygfhun8G3K/XnjJ99XbwF35p4xq
OiitsD2IZSj1urqbdTPlfOvoVDbvMafbP8DSBGG6LllrnxpLq/1EvA9E5R020R2kHoR8KbMhI+ZF
S52rCDxzG6fC4gZ70ER/neGeZYfwMoGbB2r1DK5HB2aQiR0xpTx9G38cTa004tMBLUFnPFEEqlba
SmtSJZgNaD3ZNSBlzKERXaiu8Zm1DTCHdL9uDAMeRwtpOPeQshU9s2UvCBHwk6dOFOgXLl8T/mwa
6o9zZ1+4VlOCM2UOmAXOgPr4cCo0KikDbYINvQooc+o/m42Ol8yOgUlNSJhWgMWeKkummYCjFUOv
38eo8/Jhyj80KEcMKGBpidI98kSmmXJq9HYjg8n8xNh6+QFoclV2Uc9nibxs5Yktthm7ddzIcQ6d
D803YrH9ODUXLAimoIhibjO/FGtoT/G8IeoTmUFCU16t9Xf5YhbIAk21r5dgwMw8aYMdyOxYQUho
+GBgSmLOnImB3JhVNZqva0ZlysyXy1PSkf3x1I2yFooG64XudiAeAlob0F3sV/fV9IRbxCZbdGk2
OWm0H8x0LB4KVnhfo8RLAnEJBvU0LjTelvtj56k3EA7eu5zbNFR/YfO3Q/vrA+nxUjfawGEEvDq3
zVBGkH/9RDkHKvoSTXl6j8ouoWss6ophEBkx3gzoK9ROE0/D/lVZaJ1C+ddduul8yigTSXlpAJGU
EHLbm9WUS2JbgLfblFpsgLBo54JVwQ4RwZuLImQy279Zn+PQUkGTiu4wD7n1wGPhIUMkPPCZ9uJl
DkIPwfC2Go3fYxw10lgfyrXubITkFfgJtDlRpmVs0Le2fClWfEBd6laUjrZSjoseQ7q+oE973IGd
gvSiJQhICaDq26/DTJyPSwizjqCJ08zN8GyBRVm2EzxAwxbhfUh0BpLjhyFnGi6MysIaUDrUFrXu
BpdVrsefLTHfTWSD4BSeQ+HGPBw6fSe2IkOIO06B/VXlZvgZ1DZLr4SyCrA46SDE9gzp/sOeAXpf
sP9RhjOfX95ffaB8UN5QdoLGGzA8UNGuMeLcQ6UhgZdS5Bna2iYbpyr9JtD3fnHqB2oDIpbpRKzK
usOe80v6NClJ31aWRzIN09D/BlCFD5HVceH9V1NJrENox70zAWrsY1FIM2y6Lvsd0te2uRG7I3pl
lM5Si4qPLJqJ+UdMllkTQJNkWFg6P5Ixd6QqwCobeAE51Ewwn4y+Evic2kelVx1DhOuhPq/y0hOl
WkhA++WjO7BPX+g65oWGjVfwp7sj92jMs5OtIsIJz+IYSS2z6z9OzEI3pk5HlgijxF6959XxQ6gJ
9Mq9rPwDZtYrGX/R9jJ2GrjwDHXq4rFbEEJMvATZbI6rMN9gxnb7QuzF4IXBMqpK+vrECKDVwrFT
WXA4suTJ3CCVk3iSzRhtHGhIS6V//ZkaZL5wxzFuuZb0cGN0hG5SpEIAQAfHl1b012qv9Zh+FAjn
oxhmj70o1pMiNgSGy6Shu1+/eX0jdiZ0Br1Vf/vBUN7+OYLY/INf9MtZpuqywd9DJ4BDOYL6CFK8
1PaLtRm9SopuIZIfy/vLUxOA+52QWheNXrHCNkRwwzn8NTFqUHe0zbdiLcaWqXCbcIRp+XBQ27Pk
49/iBbQE4x7C+cq8ncCGtum21q84xvcJquVIfwMERl8ZBOG4wWlcsq+fziAbnple1N5NgG2AauHN
N0nqA+JJDLO1wsfxCg5yNeqd8CCQBU0rjZiCg/bvwVw/tYUt/kW+RNPUEkPVPkR3QiXziLpHMnUl
yCi+rjEKxITHkqCQm7IOKER0P4cUmonsqPGUMt83spceIrvm2vo6+MPaUtfiRU8k5pb0/Cu+eiL3
ArjYtka5HN8kEV7F8l5uwtL7jfXvTsI049925aMRUiyfH0o/CJ/T4wnuaKy5HpEMU6TROc8LngAW
YGPAKRprh7tlbUpG5e0azggegf9pu31gLnhOneF+7jad1TYA31Dk/GdmebqyyRsJhNldgW7aQp6g
ApGrRF3g+QcXYlASeW4xvqyT9+4p6tGI6yOQ1Bg47FDEquj9OL3jkFkL3Tx4Zn6/tV5FbI1Fqi0x
z+pToME74CMCswZ5WOgiBa1DmJz8TGs61lTCaeTYoUqW1NyxvhFb2EIG/BmOMmYlOYJXo4TEEFDk
4GpcbfREn3L/aYwG8O465nsmSNQ0j0fFz0UQ9VOmzlsXcx8YVnQe2ogp+/t9oV5fGRvSXq1+PO4d
DX3MKdybmVXVHGdg6Lguc7P/aQU6s6URT5M6ROlYCzCiZXidP+3I8J2+xM1blNt+LSftTsbtT+Z5
T7AWijjc4uG0Ev9oOZPdRFWiyawVQvAXhqz+6moZfp7O1W6x5lwwPJzxbTzOwH4LXfpd2RA5Jlgu
5tV+kU5vsDQ8i/aHV6k0WDuuzUs6rUfh1xCQWvda9uEIYGg6PRaFMF5ow0nCxOo22D9AUI7DS6ld
Ck8o5Jzmew0/IMnP90Y/p+hqLhZDMmZfOzkb6mq5HBFV17vU6OJljB/D8pgAi8qa64lp/zLBQ7Fl
MiqU3TldsTxV10/tcF4YvpVVttF2koVRgEkXeX+2qcRxI8tQfILR7eEDcq4EzF5Rl2kUvQF34qWB
dbUCSpRJ/UcuSttpG7H9qs8UZEgxhqWyR82G3PGqPHfVaSB/wiRVFZN8RC9DKckPGDJxJydNS7x5
lh23n4ZO92Ywyb1HWm+uI/dqBQz4d9eCdBUd50nwDLNlg5vDGW+1Uvz1j9Azk/nxtD42QLiayJ89
iSCfxzApoa72r+e5fQFPAPXjUm6uTcXKIj7c2cxj5mQHHIi+rc8uKBWcexmTlhZKgZcR0mDolo/L
WRNf551OBcWiSV8fSHmGp7KEH19L7XyHfw8OFjwGqnQGelRJyjdFleyfleeVkpWZfx2agcxlSQ2H
zYPPZCFNX2q3HruDU1NGGsYWy9hOQM+QM3LVGBDAKLj6Sq9VXmtD3ir1RfiQ+J8vVsYFA/PLJJcu
LYB4fmGgxAfG7Sywt9hOhOB6/l8fHadHVa8NsxZoivKVDhV5QCIax7KpH9KcBz+QhSRznpi/dsWc
ROKpAIxs2tnXuHCAz5cUnvdJy2PF/KluLhlclojOO8C0DsBsMwikXu2eFMWO04rrkvhGPxF74MXE
LdeK5u7LVF9GzTjFTtNiU8D+0YrG2H/TCkIeEVaQE+z1HIRty0k6c590SPUUR6zd/4+Uugowt14a
Dj+c7hXVtoXTGxtVrJaS//fETq+HdFe2/6OJzoHsW3OGfsvQ7RJMx3HRkek+6r+tOyZMAu/W8FYE
GIRXPUeFW3Unkno7D8rNzfupJ2xXYrewOgvzr8uPLcKyH2bSXcCFLIxP50X9wxu17jkB5qEHz4f1
26yT0wK5d0Io6dyofxHIxuQmkep70ZLD5s/wts4FAe+vPiGaiHZ1vIi0emVl1kh+8wUu2OfU3ZAQ
YUL3Y0YKI4MoT9Ar+SwYdVaWAOCSevIMM5+ODksRAZzeP8y7HxADk0H9Dt0FNRaSdP7ifMT7E7pt
iAQ4XvT35u2mRoKQaJCi1bAzYSZNZUOQR1IgsdznvqOTXNqF0z/WKCuq5u9TJVHXuEqx5F9b8Y3R
+wk/yoDVfst8Oy6pGIr7sL00QA7pMsW5TTAtIkK4FD6tla67/Of1nQg6Twyqnz/wBGshjuBsLwd7
mRQ4+8uxrT46TQj/yHQ809K0Ejud5Bg0kPF8kWvyBDXl6ve2wOwBt7E9dPmiJQmHVDTJhlucL+6j
vEX2ChLMyRYuJKdFuK6uaDVePbxDQQL8V/ec9UMjCMgNNlnrgOuaiNujLYd6o2wAOJUSOQbijNaN
DO6fe8GQmdxkstwxIykrT97a2y76mbNQFZ/b5zGKPPGwrgp5vBNl9wUEOwSy1vt5t5ElvoaK+Poz
PLW5bHzFnRGRFh7rb7+ZHL8/xkpib4kHT/HHLn70f1/mu8RBgz7/EIsHFVzGASYhbN1KYqAeKxh7
q90cA+qeEPTUowBtfi6SStZe9WKJIP5ZNlh8PiCD1zf00AxCS2a2bQcyRo0LShahcx0Qi6pWUz7A
AoZdWCHdKNE2+I6QLm35vBk1lnSVBILbSSi45S22wAsE6Oej22DRwi9ALSQbZm4DOptSczzEBBog
BqwfHSZDBofRc9KEN9pArVAXiwt8VOYtGkBiTK+byjSlfpR/bR9qPaAlpehe9EAEX1Iq4jbyaS84
1ytIRzfRGa73SLXY1KTwPpx2Jr/TeZpN9LD7NHUQW4RUJX+Qj0vfjqDVesntcF87H4OFOONRcTJN
+83Nu8SFff2Yf8CKjnX3xugADZ86IOxyi2QrNudh8JOzmoiUwHw2/MHWMClV+WKTWmHUDA5EtbDA
4FpClXF7bAw0VNu3EkjS4mBozxGkkSOev/mpZI9xN7anh0ajz64KBVJIWC8gQL0uzEE3ZO492Nz0
F8IsyMZaE86yEBBFFUhbXxBSMrJccnfBrkZ0csFQDJhpEtq9yHOnkQ7y0HQB+h7rkwo2hOhOH5TF
MY6p8xZTi5Nh0ubrSWEw6oFophbKOr84ywRxXUY81sMVRp/I9TRC4TtFDx5UDoOIX6oqvsuRw5Qc
jULQUTdpOkEsoIJLzuh4XuxB42C+LkaGo1xxYTBkny5nWlF4xFb5noiHz2F+/x1JpO5xZyLS6/9f
fUxpcfRXHI0rTk0kG2ty3erKH68Hl5U30WDl5TdmC5Sqa3sTS0lAT+itkcd2KemONDC/ADt8NG0i
hRPbz3SS7sCz0BfQCOuDOnZDAWQ2Fb68lwsLYBRCquDAOSX7f/dR70iOjXQxbl1ygCYI2uSFV3mL
skN3FzhQNi+CngE/Ym+L/zyKM2uONVP2VjD6ouvpUex6z2Ty0L4I1zTCJuP5DuGnGw1T6knBF2qR
xd9YWyXFBcxGas4utCyHQ6+QXrGmVjM996puFZjlTBFEEXDns0OBWgw3fUq7uXgCnu2EiXPEKWsh
z/YCqc7H2iTDMPOb86TKfaHHMTsTp60RGsj4Ns86auTUK+/PyyH9TbkFtWiH+uezzdzyIdfpteyI
mCqT/6DPdNP+7/z0PRlcmwVLyAwjEdgarfbmE2/tCeOGDE4fX37d1++TAP/1R7Yt80D6LRGakJwP
Rh/2HHB14SEEn16yBFnIiVHOX+0QoyyrpTrOHpbssMjJ/opS3ImYC6dFRf+p8z7v9IS4tDYPTjmd
s35DjjlJqqfWQ3PX9AFARVAUttaiM2DwT+fGBB4sAT5J++ccRWlZ9FcLHuHjLRPZ4WcE/F/OUi1l
cD1B/YXTJLP+oYbWB/Z85GjLihMpYbRlXDw4kGda6gIJ2YDzFhHFfG4B2WUnBWpMpBImqdgxRQIb
sw4yAth7aYAzbRXusX1uevf1ls34ScSDy3D1zwlvQ3TrhDa65241PR77Pql57YsUAg3+vPRN2T2i
vxTS3lw+4HjguX/jyDK9RMVGtK2AljX0yxaix/gkp04FChyBVg2k4Hi7upsItQWg2BlWofNUPwKE
yTx9ZVCExe1iNOfYpAm/o6uec/J3D8gE8WXQHE1yWsXuwcdEXLX0YzqT4WOv65kRsQBSFmPSwLZZ
DqR2nWgLxR5vkaK2tY3Hww4xdfFt5XvU7Q62XrElDjbmkdan913VNdpubrJMLe/6Z/s/ZIJKbG4M
RZqlbrYYXAWVZ7jwmbkwhdWdGKxbYVSnK02FMEPw8lrbp1JCWaPoaxSD+Wd8HDwQdZtqRHMbTmsE
GquiZbSv15shdZyDvU3U89yty66geewfug8uvUaPuDGWVRjZgt6pyhO6BQ9I7kCMDDyv9iOzJdLe
saF83sb77eaSBbhfUkndRxBo/68EiJGP7u9JLEGzNdFi8O7BKX84/lMbpb2/7Ag1nBQ3hQUDHdVb
A4dmc2rY5X4Mz86O3iTn6Z86cO/Y83YHG12n0g7EzH0VLbjvFsSpFv4yj/CjU2x1iUl8OHVD8QWD
3ZqqeNOcNfG9osJD41Yqm3MamfoyzFWwfL8LLCwxzmLaH7TLoYrrgmKiXpx5/T6TFhvbnQGAAGwy
xG7XfVbEZ7xvm17xzvwpv7/B0sIiuX2pm5iSkAgpHJapfqVUPg8EepZThS6uK6zmpJjqMM6F3/nH
yaVmmnDDY2qUz8MISFrtNh8c7DTemGffWvJEv29vsj0RGbt0ftlJNWWLw7Aom+JF9nXUIm+i4Huf
7aokaySyftr00LgqkJiLqu0JIP+75oGtqxikjKnxDRQE+jOsawwVebvJ0RWcm3SsVt74HoJwMDKJ
WrGep2ptNIDyhyKl0bXPwbnU/T9PKn3DHEW3DkmMtbz42J4FzviUpeREd3ki79qNFH3erguG+0et
cYEZXKfQSRiH778pjd6AKPnBvzVzVNLusMhY1ZL7pO7WWveTY4GmmL6OPblbZahLVGzm+93/otoZ
uoQKtnE3WjETd5s8MhL3UKBVnaOZHKvmTkLK0LN49y2WgsBJDCDwca1AYAuRiqeK1FP5iEj8jDN5
noYFg44ArmydgLbx5Y+g7MkMgR+r8sxu04bxZR4q8fwquRbxf/Yrgmlkek0wldg0LAH507QoyXN/
NUbRPw5YYeGIgc5gR/PBcXzWirI1gbwbUpCP5e8JjBw8craYRIK8EIvh2U0WGwSqzHC5hNtgzdhL
cALmziaVA9PgIyEIzhxZDJV+teObk7RHUcwI3pcREGqQi/HkhNfdHT1SrZhBimRjyzUyGelezt5B
p8hxvkEXm93dRABpKQumxqN9lDNDeDEVB826qx0vgUWnAOB3RCflC2u4tiaICUVx5DXZHavfqpB+
bOgHEK3WlxugDGK1REuLBh9+AEjWc6TVipKuYECRLgq5XALZEk6rAhMKHO0bcTbnIhO3NM2cy7zF
WteUaN3Vnyh0DDJx6jFnzjPjNXrQ/Cl2V4u3a1PQnxj3lC7XBaPgr2jTdbo3zYt+Z9dJVwpusAmP
gBQazm2IPV05De9rjVDCaGR3b0hy6mZ9MhqR1DXKInvl0Q3Gk+pT29+y+eiE1HvdwI2sK5TDZhDk
J4rNpyYYffQhhXo6Xa5BRy5NvnY4DEna1qPiSzfYJqeHrZD5mdN7IZoMTHONG4Yp6U4PfonL4/Fm
0FWH1ZfQISGecZ6v3WuhivMXw01TRX0B5XUbbwdMyhaJzGoCoI7WFWnp2FgxXtdXtsl/KPZFGu1t
txxPYzszcoNXEWcHt5bgcmPoTjJSsBVFla9a7C87+odPJM1Qdtdom9HIZfC/gEfU6FprbK0P5U0R
AZqpL8xbW+1eBSLTewlKxdc6McIATgq/UQ9wyipvn+qF/GCJ6PLaKPPAHKwU9a2waW3N5xQuSI6F
Keo3w16vX0t11Rf0D0J+e8lL/r0BsG+25flCk43DhXK0cJ/Q0RmXssHxAJrUFRddh2cahAsBOVXn
JhcP0YgC8Ez6ePjwOcQDrmCen9OomBQfbIjR1wdqV8DzOpPVSUDUg6DWRqu/pRpuhqX3eVH5CFit
M3+M1hUyQbIgHVdak63IL8TJUuxgxZwEk8AJxin+8E38QqaXIO7CczKsV2unYsvhYCqHYCy3pXv9
4zfadXdkrC6Ssmpkl33ryAgAaaLkoPXSQkj0NM9dv5Fl4c4ulyHBDtZ2LpadxsydDUEb4VxKq+hH
6JMfjd3hXvvp1ZiJiYakJdSyrD5avAcgf764w66wtMnVE2vygjcdP499cVwdF4Bn1XjMGEWZEku+
e5CWB6cPXHFza3Ml3HGuxKw/i7JBSFWwZwZ0BxgJKa3E6og3RhgjXqHtyrI+DE2rXu5AjSvxyvhG
9ojv1u5UHDoDgM6FuPA6jSqU8/dyIFdsW319DYgsxxq+Sm7uUUwpEjF977pA1qJ3Bm0H6VT01FpR
NrwsV2yj96XRRsloxntSs5EbKwaIL5TPWL7WhHB06s2UNgXVbWmmOtgNROcsXHEjbRLKRk5YuwPO
4aH9lkibBwQ3TNIJDANwZtinkVmdQg7xfB2M9ZS2m2WjebtJf/0pGTdsMhq2MxBuuO41K+G37kBp
Bm9GxHEWzFFnDTsSX16+L6MeC81IqpFWNh43RMYPdkZzBAdQZFTb/JXe7SPrInPlSoINXPzq5xKs
F691mVhrMSk+vL3zWmBFFkYxbffsQiKFXPiyUOeX0giPE+l3iL/rtOn15Si6VX/GLK7DQwRQ593/
3ybmmMwENYTMymbIPvzOC0d7UzgwC5+n8KxaUfRlljCTZ7VV/2bDWGaO2bvHcb05TLQXqewuN9N6
HXj+7+cQxcJ+oEYIU5qcLqwMGLOGnylpiCc1DqKEZvJjCnzfOTLB9xPqwZP/VVIL0QCPKK5/sA/e
/MLBOgxO3eHD/LNPaMKKMZaqKBW7TG+IsHSmUi4Y6GzuXj8k2UPloCWLYkIJAcRBQbkXzTJ/1bbt
ORYH9rUFmVSPs7dP/zqVT5kQ+SEy0dyFztMhhF6ZMGl3zpWoQA4sxwoiLXGAzRRFpguH4tl/X1XU
DjoarbLBmBa2hc3KWQi9ufJ3QLTqzFDD6+7IYXtXC+vbohkI5dfqjrac+b1vIDkL6Fb6PRDcJLb/
Jtt3xprAnV3J6BEi7A5R7LG5o6H/yYhbYlnAWPb4XtqSwUQh6m0h2AySf9UXGMHqaLPA7RKGd8aO
eCjdJ3L5GezcZ9AhTBU0V4wefL4tY8Kp0YyZM0xI5kmCzhyxfGctED7GodUKDGc+KxSexlkhRyDx
rWppUizQhTEWF5Ut+kuKaA7tUNPw2UNAu5CoQMMFDi+vGBkgpAxXTWhg8DOSNmVS7nZ0fOlOkfYH
L9LWuq2umf39QbRkYRUeF7Y9U9wNuZFbWqHoz0PVZ9mm4TzLNeyewVie1/IQoVuG5MSyYwoinwoi
qAjX5l2Bnldfh9qbU2wvCcED6Qq3gEqmijMHcNu2BCmeyl2QnGKBx9p1fPfHok0TDNDp19UkNx11
+xkKrBSVfGOiNMsYpTvwsSE6wfLX5dHrdyfL/oR4byKul+Mjek/2w+SSfso2ySA4U9U1Ac7obTgg
DdKIJOpn0cb+QHa+EhTEHDKOS4k/KDNN0vAv7e2yz5MorlUWaiJTG5nPXoULZ05ULzXp2GtEid4o
MkzBzYvm3KLmw7fTkmafCsD1yVHdHoGOFubJE0eOwQNSQLshXilNvwquIlWAX2ZjpGJpkhKkctod
xF0wF3GyUIKJBKGIu4Xhe5JwxGl45wKXuCXEU7m7I8+Xwlucn9+iJx0TR5meVO5+PESGlzo7Iqqd
3AxGET1KeQ4xdrTW1nmY9WcMBUU6eVKYJSrXDaTJUYtSRBcjx2XDLrwHRitZjYyjq/3S3SrbNV+9
eGurpyUY5AGaSOlOeiD45fXYBKKtbJF0+n0rLL5yBT/B7+B8AgYCAdGRmrM7EUFvsinPAvCbxWYi
QMFGPRKSzE1E8qOvHe97E+HRuh3aHxXNlFcVSuqlq+D08QPgFPGTVq9BkxplI6o89PJ2/3ZDLkIK
VPIMpbg0Veiknfulheto4yaF60uFXRqcC1znNQgGS5o6FsoRFLWm41OZer05X1LDp14fInGp3C1i
DalIBfIfPDURTe2jE284+yDXAm7KAsvXIYam/h1YAWXPb/OaZfyMow/SRwHFU38BVfpurpXtub6F
t5rafVGkiIyOpQlaIdq5WW27fgK5iawBaNU8djvx5UDOTIgmRjomCEtJLThjFLSHJHKpdGSu8R0/
EFmgwffQUfjDD/KLDa2yOoIZD5L4pWi/oqV0PVb5P0noHT0TbvK4sSqNcIN545Fd4Ib0tli7kyph
W/jqRhPb4PBk8XYW0vf+zyjfDKtr84NySl0DmpeMfGwWXdc7rmgzDgk/fBTEOjioDuTIyGUNgIfp
ssu/vyogG9s1nhdXJtlrcFcNWzPsOA1iUZI0c2uL8qX9E3i7130JlSXUHG4+0SyIOhKEPUU3Ykeq
Pfn9sNn4QcMvvrh+Vvayu/2k1Uk6hGdjn3tf47XtAA91rhVs+7fLrIypK72Eqgzck7u20z4keffk
GBp9OrUgGDCcwkGZ6+cGBPflhSShOq/OUCa1t/RNzQgfZRRn+FzqZ5jxn4e1YafxzO++BhEvKV1O
GylBD0d7CvRMlogkZ+8F31lsZpKKOk2xycr+3CBrCOx/pErKbLmNMNU9Gn54Qwvp0nPXcJYymByw
fxl7Fev8OYjsVPR4pEE1dwOEAEDlqVUTlurcKyng3pEXjtRybsXW+r7JUxRFHg1vdcA9ITFF3ttp
DvE4cmzUG3ZC/4RUbrehFlFg0H1u77KfH/GS6Wr9wP1WyswIKdbChs5dXvHM8M+ndf6ywGw8JOCu
smL+FdzPSs9+vfyhOCexDuReUB+HBmlTdjMeDhMnuf7YjdhsT78W+V3jNtJvoNhSlttu984eotUI
VRO4/ptVaQzI22egIG7my6tXj91yByQaKDHRyS7434AOrmCU/guedsoHXUoXeyBiI4BA5uCi8WBy
1WYCeloPFC3IPnpC+xMOgLklNk1LwCKYnicPsnR8E4XasRg9CDh5WnTkUJDMunhYibzCkXi0F3/c
S1N0KIVk7JZYv9dcJdKgs7aD8V95hcn7rkfsR5jl80KZCjSaxTVmrXhiyPL5b1WlBhLqKKHXANPt
EmTwa3xySmd+06mMqRwbpx/p8VYn/yempdEPRx7+UN3jX457908nQ+s64sQxI+mcRd7Zqe6vJm02
8iczOe+RqeeZ/P4VjZc3D/Gc4c3aHC1ajrZa5WtSjzYD7VGGHQydIr6cd56g19+jm3xwMyXXP1PL
Q1O01nChcrxBl1kxu1U9pInf0hFLU7jQ61A2SX8HpJa8KXYts8qblWDpyYbhRO8SY6aba0Zr6x14
gfkNbWnQW8g1YCkHXM6iFmoW8om5Sq31M3CqXfxP4UrO1jJhLKzYpzBqLHEcJuHzWqhbi3NIvLxK
edykHBHVeBKwh7qLkCNBoKSehaZ61K6nFcNfISnQY+gRdPXZ2+coFqvz22OaHMgR0x/HsBqpSV7j
ugn7DWmi4e617Z7RZPmglCRe+uMIUaCBWm9+RSrn5zlli/qg7UoG2/4qndeLiBIRl2ZH7VXLhqd+
IzIjovPdfiNbwqNbRW1E5kWzuqeO8oLJmaa9Ve4Q7jYzdr6F0bGxOM7EtVHgdaXq6m7VoFoseN7K
/3f/3NqWjc9MzbStm6nFRXcJrz0j6gnl6KaZavDEIDX5q3bpyiKIPpeIWF5cJX5dA4wDOnVNawIB
OCZSPemWSrRwaQttAxmXk2smBGgkh06TBbO8yZ3WvW7wzppU+/Qo9rbKz1O+Pw8kh96KhWbKN1r8
Vu1FnsCkpJV3woP6xIMHaMnf2MwnB7fGQMjlni2bioMEdV+9PMD/oD7bbeT8FKEpQ/jgZSDcXQSo
EjYd4t8gGUIyywaaGYR9EuRVQW9QstBmSTU8RATSSC/K+cJKALtIfGvL1ZpjA1UAV60rO7S/R489
hzOjr/a7+1Cgz1fkHCMWo1FR5RRjUEGihOsf/OqxBjXhD9Iqb9k67T+h3AAv6wYsn4/b0LKfG7yf
afqVMAX0/UxTQXCEl7HXxl5Z/0iUb0rxZT2Oh8GUSWVDA9vhAnp76Fefq/WRgiRBIr9X+f4Nb/Zq
aWKxmVmrGBgUCE4W9Gu8OPLAyatggdF8SxCQQm6pjpmR4l+klC4VP69wUaTg1nUWHBc2Gd/g0bBL
63Xv2I9sy47czLBzjdL8Vf+JlMcrHw9TiTqyWuVRNHTgxXwZotDfQJEGZ7NhA9zzip5yNir3kwiI
k+ILfIlsh5iI3tQmrF+z5HsO1eXWx/R/lFTEISsLBKTb+Jy+ntD14Y78KwIjlftid5Y1QE3WB/5X
p9oZnkvh6131p0ayEUwuAxKZ0MYEGv4vaEmJB/ECkuWYti8lwLxdWjIibR8gPxVuUHEZ2L0XTcgA
2b6TOF6puybrAayXIDFt4ZF3xYNmA+58WnS1qmaTkuryvdRGJ8d3BKLxGf0tdWnGupuCzVKHEj4P
GNNN45Yc5Vvc9UnKBZXM5SV7wd4x2/8X6p+MMxxsRz12NDa6hnyX2oUVOOSjzzhI+BvaeOgFXTT6
KXjVmgES8a2OCNXFMzYgYDZRFtQ6VPDyh0hhlzIPQAjJLUjOjl2G90uaafMvM6VrRhF35xT+cCX/
p5PG6xW7NKwX4FvW+t/UhTb5q2BAR+G9K+mP+0vjF9xd0D1kvOL7qayUDmP9kidQqecURjofbfWi
zgAeMPUFIzRUbtpt+xqG2kDV+r7iesyRWjoeGzFxNzLnxYhOlzPtlnrZ7vTZB2tNfzaAg7d4pyKB
hYcBAUFB3XzQyUQe29TUQzI9Zs/BxAfTJus3+xJeSdiUGwNR21gW6J8CHGK6/9OPdywSz9QYf9gZ
fzPE92X/8fko16/tUqR6uyh7pzGQYk71dJOprGcSZwcIgnfEZFy8poIXNLSQdl3AnZFYGS3YHjCB
lp22tdPvSYKFB5PuHsUsvgiKqoa9zgTOfW7MZTmbgtCweqNdX0BnbP96gkk5IUxUcZ9kHnw7wTIR
Kc/0+4hVA1phIDr7Xb2hl+JEDl3rhvxlcgzwcf5qCrWh6bNYWZrsLB49hI7Wdsu54Fee6glfi6y8
UH7Cvy26aohuHf9Pc9dyKsBXVMmzvQHzRIddsS87w+jgB9ChDAeLmooMIJlDO4y4KAA53zeLgXOB
StY7rn3LL2AwwIgTqCUrtocdSU/m8aqDwpz5eVyhfWwwc1NgLh0HB6XVrCoJsqnCnqzPc6kccJXB
XLKhrcx43R/Y+TgVTwT6wyRX0w+wGr7sjtPkf5TvJ+gldfJU+k40WNu4G11VFC77AZSigZP89enz
m1meEoioLNa3i3vYQzb/mPKm7opEmN9E2cMKS29gXTqsbhjSuwRdUc7sV4bkJfXPRXpdc9LrMHzF
E7xcICU2eICey1qZ+lbL5k3u9PbpRFN16pzRZE+DgiJ7l8W4jQwu6pjhcSxh1qxwvDf4ETQ2tvZJ
jPHqiCvFHH3A4Ivzoq/4cgYQxq76+ijJo1sOdwtfsZZE5alXAqft9+qvP71UCoO13bH7ej47lly6
yRlQzLHo1wAmP92jys90ckBNkudTV8aTKe6WTHqDHn9HpyNKsoXfTCBrjSHO3dvvbvB35yZnKUKX
NV9lepZPh3FMUU+kYRkDjG9lz19EjTjZyR2wGZ3YV7oSoFyH3mPyPR6saAApV23mXlWGJsDP4meT
PUER37w7e09S+RKjWJyHOb7Gck6NkVeyNfbh2W+xepz8d0KVS6FCD8P6Ec4p4FcryBpP6HwqYvrN
82v0lXDNyZZWWPkI18ScA09HfCLaG4wLyzwzhSMsXT9dq+DNFytLvVUguEGBdbg84S97LUAB63bO
UVrBTY2xxYnoAceCCXIhzr2sYUafCEKiEaFNeAKWahVcN9K/FN8RRh8PVAvpN3d2/ib9l0kYP7Mv
N4amLdyf7BzHtEUMR0szHuu9BSBw9kzOauBoP9KQEQllOUtKeETbCAph4viYYyU8JP6XFjTzAOtq
HxU7DMpEikz6BLyjB6g+wfBIdr8LmdO3WRNSTNqSl7fQqmA3eMGjjyJa+rQbgICt5F2BE+d2RRy8
/Mvw1YdxacyfaeYBSB7A33AWHyoGeNWj7Hf4oyMR4aV0z68ksSA/USl/JQneP/YtcvqrgnBUZ4j2
p7xNfefRVCaFp+erlCFDfOqdwIma1kWiphaLu3Ti78a6NgdY+xbXFZdAjx5lyM/VSZZKmE0A+qPY
0Mic2AKOHbEh2o00pwt550fg9J2+XKSGQHhI8MjkQoP7GhqyKVcuMbN3t1/J/J236AOSEiAOKOYv
IoNupXE6uCostlrXTcqy07TYAuyeQN+jNcPc8Pc7UkjHMz4/ikzg9D3qGSnQbpBosoEoyWaLANgB
D3Cp0eduoEaHWVViyrK29ky2Y6HBD+h2SkFjVm3+9E0RclMBDNjZtjJEGbBB8x4VgP7f7zZbscw0
eQHFrkADKE7v6/5iS6yzmcD4pp0OmVO3pp4EnQ1BQGmJZHU/t7gOI4AJgeR9qeOmXD7RqyXaYmsW
qbZ0uyJetu6rAqM2Rp2B7KtfrBPBW3EeQJPMM/NHFwKC6EXRL08hJt9tVQi7dQZrjoYjaq7rfyHO
zvJB4cKBEg+FWTzaqrRsLsjRUX3Ar4dq9V2QHV2sdcfXdNx2N83gc3J97NA+5sVmwYg2lIfnkOGB
3oIy8C9QXJ+U/kWx0apNx6S+tEFF2NiLz+rd0sdk7ShuBr90zqwt0NrNmCs2vLIEpoOHSDladPZv
rAmgJfpIvhHSizQbNIaGoefCcr8VibC/HrZjWxL349zqWjoBqyZ8hwpy2/x5dDFlv3VvqE1Nvu7Y
K743yAWEQkacrHdoV7hFSzoErO5SkSeaXN/zs3xcEMLy/XRi+x+8jqOyCfNMGvz+/ctGOuTc90oW
MVJ1evbvl/WG+/2cZaBxHmVlSjcp+AggaLAagKbdzfNPhI898QA+dNIXU0FjcX1JUWeT8CZsCmiu
sQG8GzzBVGjRVPrV5RqYXFIMfRKtBWE06Vn5tWd0bSp2IW4fWk+s6qGk97iwTYZfGm97jPuOYc+t
CF8A71P/Lf8iIc994/vdpcAQftvLH5JXh7ybAbTa/73SHUpWyo5fTkQBll7OrIfEw5I0SQesFfZL
cipr77MT4tcgL9RNE4X+Exbk2og8DjmX1LGuoCUhAEPYRWYM1BCGdDy2apjzQ7qBLecg3D5XxoKZ
qetRGY41CbUX8JvqahQQscPDDy1MXYjiHOCxqdAUC0hTbflm5vZTTzj8QnDpcOEElwgG/+ZNBWC+
cw0Pe4znhyQv+OfWPCOVkI439O89x49F0q6UfqF1LjRIJXQ/P+1vpuEkZfeMQd/mRR+8/ZuVJGaI
qHEA7z8m2SdgenzUB5O0BNUtJB4XK//wuOdSNEfx7t3PfSHTO6n5tV1trx5nv/9uGKR4PtRs/OVS
k3ksuhIShtFKkFX5e4kS41I8GgvqZBfZWZyV4NZkUtwHz1sFsrjQZOQcFwpFoJpYG/tltVTUdcLE
gpBmFGOrWloVEhtqRvmLLXRzULhhO8sKS3tlWYaFlmNZurqrH37ooy3ujnpZpyPTBj3YxtJvxy+P
QPxirC68n0mlES51JhJPDrBiVCb/ZEC1bLwJKAJpECBnnwwyjLuix44VIXYQxNG/b98SqdMUo+rp
ArTjUSSoKWQKw8uOViUDBkHh3rLoPClt4eZm05F4wTfjlBwUz03QrHPYKR4YpUgMx2kkfbug/lgi
jR60fKobHn29vd0xd3xo2z/j62ujDbvOKr4nybroqjgqkOPE93pIiTr3RjQDrmhfUYudeHjPkdZB
/IIjxdVp2gURFMSpFmi3ih0nCKmF+2I9awExCsvS4bRSGeqRo7kNRFb9RHCrMfSAXFpg2B7gyIl6
DDIQW+4c1Zu9bznExqFVhkRKobVnV83p76JISpTXN2OA/SSzAgUL+HFj/2fuKIIS22Dq0MquJU6F
kittjM5oXLf1bZVSWVXnf+6GCGSbuMRFKkPlxezu7aQ1viJsunq9x2ZsXqXAe9L7wUu9dpx8jkIa
TlVjgRWNp1QOGN6K6mB3UyW7KWGMpv1mZKoRfRd/VbE1WgMqbeL5giBqaNGU757Q7+nu53kK8exL
Kx4/Ovjj4iCoE8BaqChZzq/eQ0f0L79uTBqufW1t6We91oz2IpAHtPYYD9L0IpIoI5461gUMM3Wv
2h+u5P+lrdlif0QgI+biLpF0u/0AYLQaro7vPMpQEthfSpqs9FavJYAE8aPZSMzxTAjjmtuCjXzE
u+SJGX0efPSW5YoEIqCl8r8s8Jg2skT3aYdrc8KG36zKv/y+uT8j7GxFDdT+WeB4Dov5GuFc6kCq
tATk1U0PhR977gW4jNXmgZEIvAQDGcmc1I4gPpH/BJA4rLsS9IvpjSV7pGlL6UWPwZ5exPX10/dJ
HLY/Nv7F2m4hiZoRZsYXb5ISf1YTiv3BePG81FajTkX7Y4w6jUh+wDEQtbkmUiVcjG0lIcU2YZJA
l9TBVFo23R5nErYDvYSu3ReHiby+ktLltuZGgHE/v7gsEu4ivjAkudSfXx6xuQPG8uRXdovycglH
OXW1qtxUEoKrzwoFVSiCIPy/cnRBEOWbucUT1jUgWNe5oo0B1G6U1JtzdzrEQpTCzKFo051AXzer
y+EOrqw1HmUcm6WtSyKMeCu3k1pWsqY18mzrXkRt3UrvaEZzLJHkXxvy3wSTjrjRZTOwFFL0xqHv
pjE/OyIowCAHS2Ds9fybEampgcuUPcxj6Q8EZfuFallKIRgvDElq9fHaS6boGPUXV9gca9/FGn9X
jFeI65nXaXn6UMz21bhtl4m/9l/dinkbuU+MJQfYXNSWnV1tAQBdf3SbUTC+W9z1bUUXQPxR4Pqi
k9VwwiGEA+FiUE7ias/wncKbTGOmK8dWRa/tXcltEzB7hzub1BrT6EkXQs8IEOhZPSd3ybi+ugdG
AtLyX5VZzic/aq+T0Wfa4wwryBGkgOPM6P9LSDKbOcAwNwsrISeY51g/lHmfD3aVvFtoWsG/dtUn
9P3swf4VgDiQRwnEKnI2M+ZzrM5JX1fQldW/T4Moc/Z+09rdRQ1s4nbpxZTcsexXpU2tEKoP9O8r
6mMnCpX8X9Ux67UPHnBJSyBiiT5kJAF327op5YKdpfEVVTBqZciHJuSCw9Kx9bBSCwJngivvM8L8
lFdjgcMLHbfS/NFea+4lPBM40YpqBesHOqTp52LIG0xT3bCfNmUBjJsf4uE6v2Nq5uJIpo2aTQsS
rOuD/+Ie6cEuG42ssTL3ruQXYW+09UHdrzycgf3qQZCNZ7jg4cIL/WT+bfOc0ZrDOIqk0fFvXfRB
NCuF4XwYl0ZDxmOnGHnXMOVaVBLF1rtanfwTu8EfNrBm9odBTFSPPIYVguZeX4DnqXG9kORIuZ/k
WMEY6cf6VzUArdrY1O2wDWgepBwGirIxLZMHwlIZysCNVQ6kSMVcRt74XRhDNpCy/6VOZCplCQnQ
rPnnSA2CE14Utm3QqSyceVsDa/CwPk+p0qNmJ9tRwnpwnTvucacjDGVjdcd1ig96N0agbyZF6YBM
2fFuzNYN0gKdirvqYmsQu8CzgBE+hxPlpwNHtkITI6q0y6YsjxZ+g8RdVtFLoEd+OKcjm5yoRdUD
pWY9xdsYydffz56lkMwrekHDirWACSy7vaqNOC7y+P4Yl2lQTFyK6EoYZJZKmN+yyQmXFVKpvgf6
3zdZ0UNtuY7UADDFnMA8Do84Fo5zKU/QXIK4QyddQPDVQpCfawfmq1f84ohFcLpx3jTbzQiOlfLl
zxihp0vSsdw1YwGAcMtfa5X3wLIZJSmecfWzvaM829RgGkdvFQ0oU2cY80Czsco5mTY2RbGvG2Rr
0Nw1Bni1/P+XdYvZTe+dNwtSJptciSM56LcM1TcnEl3dKMC7uK6EkOLuHc+WXQRgDqYnBc2/tVio
h5eAMfLIU2RAGV85qAVBps5XLve4N1A7ULjZigHC5rDGCVOPwxQH4vYF8OIISIE7zP3LUd07MGHK
RRfByDeF2Ij3P82fkeDCmSWd3oNvmXvQswXMOXF6GlJdBi3tW6oqCinNTBC3EoeNidBDGGBarUhu
xdjvA9ewN3Hk2UAJBKtd5XDb50ArqnOAzPZRZzPckiVVJYcMdb1/J1lKq8F842AoRbU5SK0xvfFg
le7CZoEuTbljGcyEq9oCc9XAhVKytXSgfiOlziIyJBS7Ivtm71R6FrelVcjwQBUT4slt3g9HFE27
6+KlDsOgdRIi7j//jBdLONxbBgLF4icMwI7crFDl9niZzgHAgLjaNJFNOEKvllMWauZ3qlouujY/
e9hfNCk90RNAkYket2lw2VMXMn7Y5Rj5DhgcR2grP6QiQJtmXsBKmhWeq8SS4yyPHTCq28e8UAIg
aaMZ759ytuSO6P+YRp9V9tTgiEqGH1Lh5EmHthOpGYbmTuufOBd05nb+aAchHncgCys1XrShUQam
jYVb+4H0WFt95aczHSS49vpX9IaskIyyIAJ4eCmxztpTEyFlpSlkFk7xWqykpsw7k9EuMOaYS/aB
UPzQfJ5kqlTWa87VqDEPYnhPl0nYrlvtM5X7gL/FZ3xBoF/cdw9kWrhMfSJ7XWy4cLkWD3n78mkK
GlgPf2I2nqCLYixA116Gyg9EyO6jVG6ZXP/fWEJjK3QP7tgG22gaiCRFEyrx8cYfqOPMdzCd2AJ7
I35/Muyj+q5Gy6MbLKNB59wYEYCCaDIfMXoxeee76yKQE/LuSU1arARgEnoD0j25pghGmGJAmAhE
OJyBDyrVqXOB419YVehWJOcg0BzPlwiHHGRmzZdrq0Xk/I2DbA1MryJSQpNjaEJ+1rZiBSj4EwYr
g3o709xaAI+xCX08+yo8NfjN15EJwxQgpKtEOGTSzIBnnFJ0vdOOFHHgWQ7xKnff/0F2Ksqqro5/
0/yOZF0eua07+TzsmYLmvlDb6aq4RCyYYJ3VDkVeqeZoGxlW0qhwVPrDpq6kWQ40stxXUlfbvUHf
1RVfVURRffIQCVxxfCFeAJY41sLIUwhWpe3M4JaCrIpVm5Ek8gUp3haZPYPZNGNJAOX9vNU0ffRT
QxxsrjDVEXDOruwIc82x6Cq1YaSf31GWzSfd/dhsljuPVvdIfHP286j49b2wPhe+exCgBl/6OJ5K
Mv4C79etEYrrrAF47mOF3pRQAvuRGtYTU4KtQCBNSD6sBqmoBcGZT4pfmFQkgbNWl7p18mHrbMU/
xUZ/pRDg8uvHEXX7VA4fi7nuKpQe97hWT21qcn5ZCufHISCnqAHt4QM8SubtxsAwd8JNqNqoOudk
NBtaaAaYiivAqMHnpJeqkyr8LFIT6aVuVVYMmsTJcWui4NrePlOnigTQEZTPF004UJOGOowMmvRw
0Id4Rmnqsn/BLEezj8iguZrLHvepl9ELQrMkCg5MLwFAxX5ChYGa2f2BVAosm0iPQ3B3lqkIxSLV
NNB3UhdUC1xGQPdF/H/lC0+72c7yqyqH+us7OQgLAfb+RlQOdD+b+flAvl2Mm9W3kTFqsSHhdn5x
3lsXK4AyeSSvvdJ0H6/UxyusZLsG3H8LGQ0pekUgejXLtnvXRHJnPbE5hgWq4TIqSt5iV1QQFKwt
+Xtq3v76KPd9KLwagr0XSYp/MTMZ5Rhzen4E9t6ZcAuDOqnZtRN2OdC7aIXSwk6xQ7ZWJbeh1bf5
CGpJHsdUFtk/EEWMKfPYG55mycvW2qiOha5VsTAijXLAyuo+e9FTiP1sV71R4x2iZy7vFAE6Y6Ql
5pBSf488GblBZbgFi9cmjHVfjNIybhKjzjvvYs25vca23+QO+2cNY+JHWAj18fZatNeFnvkog+fG
szEKiLmCrX4ZAWS5ZToUyby04w6TXL+Jovshx8jA55lQTpdIEWL9qdsSUTw6CPfuPJhWiFN//l8F
BTZR7LCB+PQil0QRwt29BfrAZfTfwf00RFiZitvnythsHzHj8PXW5F/hFUBrNpsJsvt0tR7S42D1
h6eLFjdflpR8AThzdYPGNnauYCxiU1dXX+aGRT2OV0hvXRyq+s1N/I8jzt5KolPebeBo0s05CubB
cOnFMHB1nTvqdUihiPgzCdQtyQ3HmIwGRVVPIlpCbnnoqcbGiFOneEu876cecGRw85gylH0kcb6P
7ZKOTFnud2DOu2j50w0l3gN20ItJqAKr/pkhcVTTP2EYVn5KeQz9yTLcapB1uV+IILgWOz3qIQdR
w/rvHs2Zns5hxNAaVcFh7Db9SPLOYolmWpv+vINLFP4jL+Bn00CkdeoTpN3llBipYzg+3V0aWMe1
hVtC2swPZalYkNHgCXRlMX21c23gA98JewjvYC/qEig/2bxpKzDmkZw/y61+pOeM8dEPUQnZnNcb
z48BIQuybF1628MnK8WpIJ0GgisE51WUrNeYDGPyhS12fFGGtKxEf9AtRFb6Z8jlqbiQf2bhhSS+
Q5CPAs1PsPvOFtA/I5d1BfZDdbcGN/qd3SbNAf10SVwwQyEYSvd6r668MXejQ53z+CZvf16uWTHd
fDiGEtzbYScNxq5UTp8X53d9fUCGOPbcyLhe4lRadKfGnxhhP35HRiSUGvZZrmyQztwe+nRwP5OC
53zZZMcTVjMyA8CHLpOdiHiBLD99ArvBc4kTP4n0EwW3RAOGXT06z9HEljXVeoTPsVOyYPLpHMRQ
tnHAxfy6i+9Z/G7g05+wRZMDffrPJSW3ukudksrGg3EaFKv9uux+UFQR/H63sY7lpUtDvD9izDjc
MrVfqVK3d2XyUxeMrKokeMc0CUnpkKEC2cXeHceKXuJGeAe1PkDlPdVgqahtbiuKWgxHslCFNtxD
OlZprcRGTE46UFCeK0Q/utJUW2vP5PEObQQRxoOwa7pn6M2t+WL6l89cAraUq8bcQnuwCh5D9BNI
L9QIQ1Xc/X7HrlHJC2aA7uE/u7LKQ02QqBkHPfb+fqyDOyDgJGFmoriJS7R8cbgM6z1b10AR7uaP
oS9x37j37OARrnW0662w8MGy3RS3nhGZabg6pxc2U+0EVg0MpPln4Ve4H7/2gZYE6hIi8L6eGjDG
lCY4M88rlWwN2B7z0rD6ScOrHu7OS1ek0R3QdNWxxEL2fcpAt2z+7agntcYl4ipe1Ll7jsnx/rFk
JWG5YKieSGBdHh9qssPxJZSPq5SAdw8llUFO/fDtDjtOCoN8EEN7MVoP3GBkqF/pfZJrIEMd+o7V
SC5BFSqIDFqrfuvfW70nTJE16T2lvgbzJrOkIpkFzVMq4VdOS+dx/s1S1e38c12dPC4mbO19mI/e
eTIArQiXf1+i3+SZbDx6xKy94O+RlEbqBlFU2ypBZZwtkJE/1KVqM/RGzZ2HFbagqnWoaoVZWpVT
2U/80AT57uMlLIFeB+Veau5+lISCrWFm/N2eCAzeuNP3Fnms+UEAapEAnyH2sVwpQ9dYYGpi0d+w
8r8ONQAD9obdlz7PwAxOHiPo/ZS0ffRkr6yYBe9rlnnoFl8OmAq0dbFWbKuGlF2pUVmwW0CW5GkH
bQrX2tTpUq6NInuoKlpa+PHjDGA7pKpot57amCz7IF7xWzzJzMoJol5GQCXQ/P616ToteAMHmZUC
Vyb67srTVcoam4kEmfN2iQQwzQOPBK/KphBIcoi7mnRYryT4FWZ19g0nmpVQGLtc4fYd3RG2biyn
huQa8RWPAXka5DjuUNHb5KzBx9UADYBTD+hZzLog+04CgpmTXJC3oROYVKcVwwaXtm4NQs57+S1e
F0hlLW7VazA0yULc/uxxsY3p/e+fmFO171jtfqQXjfiR0umMD0vGlgXnh9arXyWeh7A5v+YOWZCt
iJj0ZB03Wos1VyApKmkjLrtn2zjsj8V/gKt0cKjrCnu7OrEsDF7lgsC3/Z7NppyeyBBXQPjf3l//
eUcicyJ2eOWSmFje/FaPWcEU9w8BkSdZJ3u2uMMR9A4s1kYST43INAIqgfGUGwfMjeHLu38ladxU
hQ6/0AmmTlCzvWMIhOApkS4dDuX4D8dGKR0O9tMI2RN7ju/iRY9aKDob62TvzbEbAKMoeFH25vjr
8oZYwyq/iBy13LfO/iCDGBf4qNMX7O+lh5xblbc8l6RmlVrkj75ipp46RnPzZWPCBMH8u6HN3lGw
MGdCr7NPx3G9215LvipqnLTz6i+S9WSGT66xA9nJbb+UB+E9EQ3lTTzlbg3yg9v9fupDUbUWoPBH
eGiG4ssA5z4mzKDROO+lsPyZFcEPks5Ic3NpEWnKD+jNFu7hg7RTAuSEezr9v7GzEZIWj7frfMKG
XQnqfZ4DaUYcb6ZVa85ucPSyEXbumDj0HOSW9vdKpwZ5dVyi+XB0uGyPov+n/Ioioaw/mvVtEU1P
tT1KsDA8EnY/aGgNgB0QbxtxOkC1fnneJn3WKuDdQYpcf9vXkpUg8UC6NO4lskQg6hrbnjn/lp9I
Ukm2Z1FUVixm2c8A9/gbgAKGK6EHr/aEdoDipq5SBwVfnLBTczGajtTiPFkZqfAcGwozE7UfTtOU
Vjf72fJpZJcZMHg07f/Qt1R/ln0PF3TCo6qtyrkL4ydyN6CyYWWpleWOYGIufMSiUEyeLsXQrvFF
ON2vpigZojpHX7xWgYA2qMojOkuByVKD2gGW7Ff5dl9ON8QPmEVkB6Ko7PBrEfERGpXn0Wx6UIlp
BxzT+p6iK/IqJz/YPZPyFe123b9JgTZbsJhE4FTi7ePCsMbV9EOh6JAQJVWicfvtnQUyR9Lqr2to
61ZqjxF8gAae9UX0+6kw/aUs1GxJ3tQEUzWlIfBBZP1jrg6/sUmOfrNX/caIh9bQAS2+rrho7vaV
Lm504B55c+VQEZM4cf+07sUAsohHf0PcPEy9IDivIZrXywuYYhdltcgCcj7nxtJZ/W8n6XEwJ1BP
MWTCaCFgeFr1NALkmr4a66UwhGb6MT5PNe+MpXRjoJnX33r1NP8fLpf8SDe/LEUlUT43ltZeoQNl
7S1Ju7UO8/PCfDKUHQBoGNAiMOBHZJLDDsL/uqn2PLxtNsE9p5xvacKPMa5azXQCSG7NuOgOz+DY
G1UJHWOshdRePdlHpboVZBza8OnYBRrP40GTc/kuGQ+7TIk7NITToXMGu06bw7zYSZkhcoCA8VpX
hyVUg3g5LlA5zhLnZH5N2cTr1YEX5ekXKsjfkg5YAYEiDTeyoS96Xx9aweDk9G6JvVGHbkjbNxKK
bkinh16CpVy9RGvUH+vnbiOdJF7cX9AgNLlcq6FqBDqdtha7NNgzvUWfSKHy4zDJinbM5sv7ym/+
aN0tX60rH8Mc052l7LJXYPsOGyBWDbApLCQh8X4ZZr+HjjxtmmLc3V8yZx7C2zfDmmjE+LX+9Ms6
/xdNy6X5J8FmXu7oBm7g79QSGM17k0+PbwU1zS4eEtcCBIrsnnOjS/YDxyqkoJgN+tph0VrpN6H/
de7M83usvzdstnOcMe5HY4E5wtBRpIX3ySL61zRv21njI4gyjfiY/qG7+pEbK9SI30sdjApqrhWB
+kagkmE0S+Tmslg4GxiMAX6VwTA4AZtep2OaoVe9Hx0ttXYoQNTMQudKhhHzbjrZX14Y3sqcg1ev
wSL9LMWz0cDW11gQWGHcu3fcQjeJlUR1/RsBglqPtvFD6/BZ0lMEcxZWCLvhH0PR6G1twxTEj3Zw
gMEBHUWLIFQNWJustZNBJ+qUXqxgaQlPLmEWUaxDYE9tNckQ5GGhK/X3pG3+CMdpvU8h9TsVUBav
yOo5eNOnUMXpAMw2FcEdFQX2s8gUKN7ZdMJW8Y6aKYAHDbpHoWEAm68MxG0U8yFSdHqF2xa6Jprw
M0F3XDkHC5AQrovRC/wCZsIHVPx8w+KnITIoHbYfg+10Wd1DUFjqH+OM4sz4tTqKH66x1GM/1QIQ
mI1rxnH3Q5cdXTlJwwBrvPqXgkz+ZUeRuLM53x8WAo0McJ6UHvVVSSJXfaTnSMef15L/nf9aTzZn
qtSohEL0lKZbWO79Z+AbrKmoUoP3VyE0+y87Gt8N8cD0ub2rFW4JbYEd0ogXnE7caUqww598Ekrk
X+ywY7QvDmzi++0DcWJ6l15qdZ35NUUN6KMLUydsHZwUTbiwDLBc5HLoU03NPhchz1SSv8y3W28Y
5q9M60q81w7vJeMPDUeO54tDiPxT49jhTw+zpko/nkW9D5FzTqKU510jBsSaBhxUCbd0PaqvcVq1
xjU6Qsf82L1pfEo8u/txBM0IwvU4yYjaLEx23aroqW6h8fngAVv+lcJLQPc5yl0NBxWmQAC461TA
3SNj/VAEFsKYpExAJokizopSn94NM24rPtOsVb4a7Y/dtz0hQyGUcBnOJXCge1pYnTZYV/zxCorQ
R3c5pQZrRlBHtHqePnxT4YuWQR3yS1ZkGVdkYHJK+Vv1mOCu5OsgvIPkKU7mhwwpvjRBVp2ZCVRL
TVzadmTra7v1PrmbGiUoAwc92Yo9PiYq/1drtvziicEo+HosnlgFO17s9IRVEvtiUz1N53ePbJwJ
5pqkojRnaByqrdKY/bVNWOwI+6fFxNPhb2QPeDzvxd2Ff2VJYY0/+a/dCUFYoxAY0gBdyQ+jFj/0
O1BfPD+wMBQuzFK8f/dPXEYuThsevvUz8FidD6GiuqF6h9owzG/OvhQ5wz0+j24WP0NQM+J2VRz0
mKSwqvhsl0ossWBHUMUdEi9O7WiL9E3S7MzR1ndxelpkDq83ZhqLeXQdBZjrM4PPHgKW0gUqti1C
qYI/EUbVjnRBQvQolrlMrKZSjF5aC7gQYFsgIpNBU8xHsmSqKzaY7JIjhLpxctp0RlgJwccX3kVt
+EiaU0oGONdHd3QXGK3ZGCSu0claX/T0Avl+FNZU/GidudsYbBs6vvdHHCdePjlUCdXqjtZfrJdC
kcQKrnVvkxrbt8rS76LxKG2vdsYjwdqfexdcdW/9WuFeB11hcVgpUOzaq0Xi/H9RV/zMnT1/21Yq
dFsQ+10F1JyT80WEk190I3WIGtF2rUb6okH9uz38P5J7xbv9PZLpXgX9ppCtwPzioZ4t+iA6KyWE
GMYFRvQhYUOluBEx92r4yifRPk0UfgiC1G4iNm/npJD/sbo38LtkMkDkHOLPvDTW/0G4I0x4sCvy
5XjRA4euaSWk06rkIX9Of3geK8575uMuEzBYRslGdB1xlKl4wh/ymfLZtHnZmk6yVD4MlKbLrfvN
Oyw/mxiaaPq5gsDypgD79/JAqjCuqqEs/5+1OuHu1UQuLkBN6QthHKV2OuZ6+DGTOHEOsaYMJFOs
kCzFBsjHEXxtT6bJy9lQA3Dbf7EGoj0J97LpZEEVp8oVog1on7K6c9iOKaWl8K05qkHuQDbQnfUq
9LDMD/zJHDxdNaPapfotpLgZkYIdKT+hnBd9wVQQ5b2yyYwg4YhcSERfkoj31CLLRCXy8bPyl+9g
KAn76hiqpljIVE1ojocMfk/rqNsnb8VwOZVD1Ajn9uRs2nrMiOtpjKih53q/alL/h1r4JUpIleIv
JcfZcwxofCuVGR1eMVa7inzUWDAHB8nGkcL4LqLLIhZ5NTvWptdxJpmcbMKIg8yIp8Dh5zLHlNf/
YueEIqkallYZ3FkXMisZECnnsVqCyp6hZZVK6pu48j6DufZTPh9EyIn9P0u1oSEAOHiWYMxULGzd
Ii2CBQnaUGuHAOvLzcU8V+aFLekaD3gqIoydgPjRpZ3pEPNvWQcTUZdDUu3vgWkxw6w/UDuAPrjp
areLRWTQurq7jAjaDXFxdOjLfMmO1u9h3e9Z9r9v0GNSldQMy8iKdJS5pM8QUMzUHOmFlbkTxXDN
ZQpm/dgG6vQa8j7iMjjxntErTfE7jTBI2VKk0mdOCGZKFabRD1SClG0tZmsmnG4ZGGLeVX16LEv5
YXU1HkNf+lNIhpypepkqlMgw5MwwMWGtHPnaO+X7S69vk+LD6pZfhx0VXGFdW+jeWN9EoDgkgIrY
847inO4wOdO6kTFxCskrV8NkEg2FndWU+uU+/vqvU+I/k3uxePNGna9emRwQ4TwfskqDM03Xg85H
L9q6iCkDbIuZ0ntbo7vZUwoeJ3dgwsbxukEP2HDHmyx3y+dZFGBPs3D1FGEpLQfD/IW5ZT3pbo+i
9UhN07Xu7X7oXx6efp18TaYg/XRrf2gnjwC1Yoj3O3ZI4yw9KbKPzbSm12FnLYZhMUyBXzAhGuT8
M5vSOU1rNsUjUIBXc3SRWolR2imUq1UEn6MnnQuCwdE5q/3FF6tlILW1pjMvCiPi8oFXXInCau/K
rWo5kvp5c0IbT2V8HuDRLepTPh9tfQ7kL6viPJrznbr7kgxCxgNB1yTeWT5tlPra/IuyaVEdGX79
eITD2z0y4C1WrZWMtDARilG9Az0Qcbu6UsyA54IBZUHzMkH/K7AOHIJc9wW+bffJyFvl3N4sanhH
5jb0reoYEuEoAYysqENFZudt4ELOiWIEI5/nb+c7iiQakFWScG5mbqlexKnqfoITKcXK0I4MMmVM
/2NlrAG7OD7hfg4Ino6uhOi+EV0lvjg9PeYFrmDL9FUnswDch3pDxUIAd3toaEI5C8ik3mxcs8s4
3GiIeX6tRDK7nQyK+J55GNjkDk/kOMTMbHMiQ5rx5Qy+yTmzUOBi/RJYqo/cdTuEFF/NW5gbXE0l
ouHLHAnqK4266ZGQtZ6qkAczdQi3ckCweAX2WPAnlnMxFvAXjnlca63dNC0Kq190RmFBRqRJonOc
bXkLE5TFG0pWZoKt+tHbRz5bKxqkF6BlcMtzWWr14sPMJG3JmlozxHCU8RSuOVBXnwEKy7Wg53Lg
LD7FzBxOAJJxKghpa8MQSIlWmtamA30CyD/xJp4VdanAKmXfzTMxhG7jERKXjog9z/2bdr0Tteb3
hzuT7LOfz6R0qjAx2lNYvFwtQTPFZEUgrgDK/RUsz2sbqi10r3rsVgeUOc3avjgo9KV7VebuOdHB
LJmZQqP7m/+BXH5MuHv/DFCEi+NCV4y1d7CiFvedz+9HmGcZZbfAA094s5F4P5bNW7VBXicihdjs
SOvYzn95WQS+dkJlgobRuAh3cV/MD13tByJJ7FpUQ5Pk5qhgyChs7UPZaWsOX4sv686nEz2gUhYc
xATLXGsKee36VUCglmcAHYIRGKcMpbcdQbDPSV/MBG7BkgEgPrkNVEi80Lrs5wRuQSNgLF+7lqCS
AxDrBiBt63YDq3qBCNWVu5iCXomWVs6ascSOJKkdiQw3B1xNk6O1OAqbPK04vyJ1I4i3Ko8uEnRp
ujk1ZHtZvO/WbSiHDAz1eFCf4bfxXUNcVKXhk1hYY8lGoB44vwSE+v4dTLVkWqqHzN1Sdi5xofbI
20YOlFI1SBP6x7uVuCSUNT3kNTcljTRsKvQnAZNRMckoxNt/4jLuIG/HI3WMS662tMjZ5I4zp027
i815pfjvad6XvgKagbQB2X5DAWR7/44Xl06KqWEKGV2vTdbs1hlLWIPWBjXJWCA+S9IiVtiIb3uX
FmPPfOX00zReZhkEJN2qAjpFhg8eCaOVudpwMQ/G57zE4F5TRM1f9JUeQYn4JMdr0gq33h1afuqO
kiUeMcHMbtqXbFNTqskKFQ1YJfcwuOKPTSCsG9aNZuVd63iPu+7VWFoTV6c6BKhbO+EN9tnkr5Yp
iPG/VWe8/vDXJhnekWuZ20vuBJe/+UhG5nrSbKIH7rParnvC+YT7ghQPRH7JGCQJDCv0WbdOSED0
fx3hN8IjYo91MBb87WZBktdzcjQFrR7LX2K07DF2ZQdqFTgnLRLy4Z9rO6exTNZJJ0PYeKsnOQB9
9CVQ4qpOG/CnheUiDjcEHGxpsmD7BCOcXRLgYMx24DkDOHj1JbrcX9XdxTZChpqqRAVgkUB5ayHt
2fasbjJiDhLLtWhZCy3CSSv4CoL+7/CaHF4TeIG0lSq/tIx/rd27GMOftQj+cnDaEyC+EZKO6bw8
ozFBaj9yojAmT+KKClbkrH0k71hVDfwClu2BYBINbEueAW0wK+t+xA7xDrtyuMOINuLK1TqdNUqr
5XXiXk/UITGQ1wpDW9KFQiBDjBfSh/o/BJieoZGnIHInLWjDvRkHzXu/0ieMrKtp/H0nKEzQPS5R
y9cE3SkpDOGiqjYKfIYAbS19wj58bpAfpIfT2Tqt1rr9eZIjrqG5FQDUCaladPlqJyqLwgkY+baE
Yl/t+1YOwOeVcUuWQhWRi+HMiGtXzVeaws1kzC9ro2vQ4SQfZHflbPwxePfG4iqOo4FcpbdYhj9z
BuPR8AfBvgs7oTtEM/uv90zfS40LlbNpbFzBQeOszvOlxozDxC9fKbFwnjZkiYSRMZN13OhRJyCB
tzU1cTUOnBy2ehqr61vIUFnyWVBJC3b5k7gcoPpN5ZoMCGlZHC6mOp84tHsqSY+59x+O9PEYINqX
RLpJKj4pOII7dR/aAvF112130pRmKLGQSzg9B0dZLS3RXej2MyVYFC09WBlPRtQ81iSRnuC/6m9u
kh5mDemIL9aEjVHKaxZdQP9UIrlhIXi3ojj2chnxIR3p8KeRLRjMPnJOeS5m2whIbn8FG0jtvpmE
Hg+czlhaFaqij58aUTMsNqggHKAltnsLeVao6rzYrsaF9Hpn7j3uTXlWgaNc9xK6V9XF9AuaBrwP
M5S7E6VRbNpU4oLPHENVyB8TwL2uulZ4QTZ9znCReNFH4oynQIcwq1c4XHMZfiECZW4MZNYOiZfC
R7dfdjWlQ1QrGsuKyxOL/78teAErHb24ztjn37PHCIfH7CWpQR8opZUxwCbYngMbZGO2Pe8S80wV
mipWLNGYK5uubBYSyP8rIIZo7B38NZNS/0rj6V9WghVq6gTz0N4OJaZu8sNyHnAMr6Fa4fwTKeAD
opOKqazrL684q16DKGZDqIbjXX8cJIkuW7SlG441kPJ3i6Z6qgCLe8mCrTm06wzFJzk8torIt5zN
chmAUv58pdtKeTx8hct9/Vcf2tIjjtXkU85EoFFlOrPviovdg2FoDAuDBWFshMfFcOmrn9KcBfFH
PcOoN0A3N/SnGG7MfxUpVcb3AD08fCc8v+JO0MNWGBhTcd+fU3p1EAwc6vLUSuaMBRczOTxZ8EXf
FWzy08MywzKykAVX2U2uc8z6Rl0BdeSY7iAUS6lYttoQTmB/mEiQiI+Ku51+a8vxAHCocaEzoxen
rAcubvikL7uwaMtNX4t5Ta/ML9Art+bSlrUEdVOkium1HdS+iuVfGDmchtCOaaRyFU4LvHiSEEq4
Q6S+8QeK7ddBbFcciuVGe+CgaNYeSr5aLuzrGv8VMP73scep27oMGlOXQInQTa8LHu2YzxterNck
ySe1hTiYBQxEpLmZFd5f8t1bm5TsZCDGDrSJt+m9+0K+W4/5YV2qlLU2oBHk1uWS9yggD3WLwp+9
fpA45eCJhlHUAXG9PoL6WyBqvlB+pGHavKivp7xuJkOe7Al9+aPcpPD2vNrjQ6KLHYW1ZDUwR/9+
CNPelQMebqk+oizVO2IEK/gWUTJQdfgN5RIbjWBOP7MK5wwhkdNlVVkcZVu8SNsTozbI6BfXrFu9
Z8HnhJyoGb337I7d/idi0MOIlS8lQG+LO2bjU0WnfRQh7k4KAmGKAhYTRhN93VgtALl2ur7oZ//N
iD2UvLEiNWo63lQ2taLHp6Q58qdxN5FQynAqUJ9BV/14jRNMYmuTF1XvtKfjDFddzKaPZbRCbbSs
XcjU7rxQnp0eQ2qXyQONaufBWcyZvDh4CHX/vFfhekP6JTJnPsYpy6bPmSFHl2tcuJ3HOtgcgEAX
p4R2ol+jzlUDJIeMW7gxtYHxHgtIjA6Gg2eKYLT43XaGBlpmyE5n/V02dLgS9pJLNv308Fht3sJp
iiFfPxwkgSfyN8S8xYwy8jyovDAwuno2itiSqjND5BkWZNQM03Z9IjmvqNKZJevpJnxFfHBXbLnn
FxAW7ZHJwVqUKPahmYQFkbBA6ii37gYfsd2mOHK+mKnYk6xR5pX7BgWpV33krBGDprSM04zQgI3P
6kUSi0m/bpB7VHGkpl3pcXoCh/djz6FRauo+5BhfThY7ke0Ox7C3hnO47XqUP1EsO9QZ2lHTX0zX
ltSLw8D+D+Mc3cGwViw/8VNKzgEpgmRkZPNgpSIx7CxoRaxcmyBIjP0wHHrApRPtWBq+m/H0ttfF
OMUXHZ/r2BuRjFxTNES90s4WfJAdlnuji8RElOu3N6zKJULi2T/KEmRakEQFoBhaQcYtElWkvbSE
lqQZLI2dJHTeXdyRNkERRoDwE/U4Y+eaWxFUFBnYrL4QGleYA35ia23r61N958VE9pdSARWWf4lg
Xlh6a4dcHY8/cvriFJKKJoC14xMZKd2wKi5tgV39KnDvBW0+FVFBzocxCntz4PkPkAhHOw/PYGUK
fuPxRrUy8/bvJbFXCv67yCRRuXmOGXBFOwoyRdBVjqk00dN9SyqQCELSNlTaUC703bafAn2HXDot
pTrQPO0P/C8WCsrY/wJgVNM4y7wB/m4u6/93Niec1r7wgOD7+bRI5iT1Z5sjFsa23dKPPpcOU0Ku
dTSDWORpXr9lpx7ddFN9Uq0j49XN7ON//d0tG2CQkQIIfsKGIBiXgJ6F6uP4ozx7cFO3KKKiFCX7
Vi+t374bTiRf1uVB2RHDP1aloFpfp8K4vJQkQ55HFdAgynI2fI+0S+13mK97rOIXeQVD1V5LsoCT
Z/WkPT3Grbiu5Zpe/R0RuXSeaAitnmMzVS9dhTCqXRTK249fSmu+X8mRa2Sn6VoaIwMqtZtoS3aw
6aVVkcvuQpdACqz2ot+oKt6IOrTWrs0PQCbXMdxB1oAZrbGKUJcQHIEV5mxHLK5go2rhNO/gBg4s
25Wy9xgGH2gmWwOMGVdNtSksLcAn/jABpOa3lAGYaw2in21sbPjqb3I69jiKVUUQn8lWKTW8zq0L
jZ/frdEVE64Y+2tOgNFRAbF3XBZoq8ACxP9vkam+dOw1taHZSuD1WRNJMbiBMdG+7/Sxl/Ub9YAS
yFj5PbXO9+PZ2m+vdLnH5vz4csvp8aJUUO5LoMt4oX1CLlfSOI5AFdbi7vdcsd6b+6YVePFAKcxO
ZomB9wGjjasaszPQY0GsSQRoG25mYMfl4vMiuRf1So60wx+xpPzNTPNSDBhSvqqeANmD8r3Lry3G
51JqL2XqdDqUNEHzy8M+2SUH2DRHrkBpnDove8V91VvmqRv5mAWZ/YXYWKEd5eTtLWENjSV9E/5m
Gfnoo8DFEPAvp9vdYMnCZ14jcZHZnPNdoDh2fp/l+v49LxQBMgo/WiUerYbusUoTTM2KOZgSzJ/o
ZwkVfR3zpP6+O5xk6MKyhz34iwo6KvsR5haGLal9TKAB+eUbtaB9NGeuNMp19W5Z7TMIh9dexKwl
yAzr8G1HQLB5QMP9mNXDcRRldWh19jtFe2NqzQjXEs8AIDE3c0GFBW6mMyAbUS61xuliqMQ7Xlhq
DAddonTEfSf17kAvEIyD53bT+biu4AmD/hsdJSCIxfZtEXvxeFP4y2ffpI6F8TCJUJOPo4HPVReQ
9vF2ojXGv4KseqNFfR5gnIZkzj8HQa5VPGogx87+xWNYKH8w/XAYxcLzr6HxjO8JbYC9/G748Trw
LDAV04KdqGZYISHzsUO07aVd3ngPVy6x3lo7q7x3U18Gd3mZPixdzl9/SI9nQsIoY4o/utHRSb5W
zG9ocuOn21wFNVteTdjlswlnA+eVw5R72e4VH/vyH01Y7Q0kC3+IUpPp39bnY+scGzo0LA6BSOqa
eCWk2hQgHII/RmeUa83NBcZyU+jrQL2fCvfR+8XSckVjj0Ju07fTyjhcyZa6ATEPSwcIh0HCgjLM
f69xW5XT9gP3We4c0oOde3Yj71n0vtO1B9mxx7WgWq5w7CkW2kgmgNbqYGB6j9M6t/xgXnCC5spI
pp5KkilahIWgsC9RYtZxO8ZGILpbaLpPWPzC52QOWqSrD9xlKxSqt1b2f+341k+xww+h/HsHmBA5
Vq2HI0BKzSfJdIaPDv5rZkFwhOm+UDcCqrmV4aU6mcgJWok9OWggODwbbMPaCR+BH1jxgwR/PBuN
WmUA1fZfU6Ya9150fSGxWvn5p75+oGKXBJeQzAJKRPyz9apODwm+b3MpITxvK4Dym5mXPYMz92WF
B2fsivUFf0iX4gyuP1zlbsThxyxu8Jf0UhBtw2VifVv9jCdcEq2WSAMmJf2GqchvmEaNrZf4MAUn
F4wSyyYCpyBiQB6sTX1bleTXJP/O3dbZOADkOtFbjuQERCfVX4RXLTO7V9IphD/jLep7LsJKTe42
jq3cCpHrON/DjZnR49DsM9VooY/TKRdfpaWl+ITz6jO8F3zzzXg0dHzj8IIpZIEMi7+a5aHEEleE
FEXql+x4stdoNs3/pf6996bniT+yrWEJFpiWGckUHql/x/QZHNTNS02687FdKyz9VikrBtz26MSk
C7ZgJh0o42yqWi5xm+BxfOvfwLKqDN/YdBemagu+IK98v07CF8nd74BZgLBon60O/SPI1ZtGuJVl
h/kU6RAd6gsZ83IpK7TCIqvrOsYj8H+/bkT2WWmwonSzQ8dgsTQZ+ycGi/RnU2sDELg636Xh/WYG
riVjQeEkS3UMy0jVevUfRr8fVSyzgK9eK2A9rr4pmGjPtJSbbxWXOmJv2+Mo2jqsG7fiEAORpqQc
rbAOupSrjdcSdN7PYITqD+UXzw2CKiqVeMAHiYX2wygW9U6z1Bt11bBYGNRobhA54H4NU1qS3NKM
EEkk0rvlJC7Rbs4ETJRCAooA3/0vyGEPO6ETt/X7K6snv1WJ//ShHIJF8a1kMdTrYvbA/Bomzzyz
mIOWHXRz6nTNPvf/Mvw3o4L8qeofLdlJ0/3mHJRfmOIX5J3DBoDChTcboiY7uWlmcfu971jqNvX0
RTCMfuNE3drhcdb8OuRfl8IHH/ECgbVfiTnVJ3BdY2V4fWzcy22V2j/n5etgX94iPsJjzTC2Lkzr
eZMnx7XhPNcwnd8snSQLKy3B4OmRzN9qaOVjVE3B44iK3B1c55FQWWJmJr+agmNhKMM+B5WXOBEI
nhfp2pZYVANL5LrPC74gKYPJG3H+NHmLOlbeKqTVoId7pDFj2cf0c6+/+ksAZX8Dswi48Ym3DB9N
yuGAcG6RD/jTdOLKTgURYOQZEY2XRA5PsVIDmWxza1H/S0amY32ane/BEwB+QpkJS/2RSql2UHEL
/djCkE2qCKDM2jiNwl7H5Ku48N27kegd8fLDhXlnQutFmxUFf2aGpcW41Yyl56e0Odf5PXxs3p6E
7bhasooXCLwS3PJHdn30kasy42WRMlMgAzB2vyqJPYFYTGL0DAvZzosSZsw0w7vKlaWA+2KbLl9a
4T5CPem4K/eW5lXHSpxKVG2Iz+PBXJZZjF91oGmMARn5OHoVhynInCO5b210qzlNmd+iGjclAxhP
RXYYVVLoydtcTIG+nDQy7EfgTRx5ElY7+3frF2YGsbjACHme8hvZ+qX50jUsjfPRSdw7JMpWjPwf
kRdOSUlJ85mZyOdQJ27CrjNc4Y7d4RxD4sILLngjUJweljE0h9tP3RkSIEQ37jVdbACc5+deR6PQ
CRNBysJ+dUZ8oZlmQybVaQr4CzDg0cx24d62adHJc0PEMzoLuGf9/oc+5tnM2HMxzA8QOcH/OFjW
A4Zp0kaIZXoHq8d93Rnj1slW6aepyWtbnmzXDq/DZybYvcqRKXs62MWSI7lDxrfosDhJY6JGiMGu
AsRj0X+EqyNpyLbYICmIM3qA9MpDkKJIiRDspqUIYkCz9xbVmNAtfnjpZAuOv5lwFNdjnTUtb6Zs
IZI3cBSW1k/XMWypf4wd16hUCowRN+8MGDNfAwIwFkmbeiVZgDA+KtDnLWMs4NGOrodBdIJlXnyI
Faiq/sEEYXOUYfoFNrwwvt+n4c/fcbLo8VUhS8wesIsVTTx/A6EHf51W3uGDFtyJ46t1++ZwfqN/
C7WPOsgge5TGdTw8lqc7ilbDEJpQyBoMjsZacNCFQlADO5fBmO0GrDZM/7Z2ySiT92xKywv1ZZgS
SyO/LLhJ2c5rlK4FwM3itrUTvjHOy3qRT2hvYYmpTK4BmdCY4CKXVBS1YooLA+aG8J2ngh9tLVtt
PthBX/WxG3LfbGADGJYzHrnMBBkqTLqS0+N9i//Kg3889fR4lcgtTLuBpkhIlrLlImuUJhZubuLd
mcBYQ5B/mm7nUzglc/Tnqh5kcuGsVsA92tZNMZ9xTiVGOhMgSWt4wpwBIbwEriZl9R13+d7usS8B
0Nw+U9n+9Cub560rLbiV+zbTiW0aOEwMt9ExpkA5zWJ9TlL+p00fujqz4THhOG4XwD8KA4C1SP8l
PLAg1bbG3/+wQT8T3PMMO90Yi6MTq7GaYftWdT/byME9/dGhYkajuHaP0bQ+gWoDfdUxTG1CDq7p
ilTn0KoAw8Q6W0kca8P3T9H0oOUowzKI/jdr04VP+tX9hCBL+9Ma46ACIPlK0vuCxxctHvUHBnZP
Yh460Bq5JmkI3vPrsertnlaTKTaogR4U8i8NjcHQaKF2f72b/9IYEi5t7IOi2hsQ9azNBtkYfSOQ
kfmBtELZyq9qkdIWNt8wzz9umQvxFbAQq1BVUsVNa6loswMwVF4kcoJRItkgn9Ok5JOk5UAotEv4
Py/KM/Mvf0iT5so5X1NA7VsegMB5TA7VXPmaRMS04tqEBYugBwb51C4w6EN8obSXInDpvCehCbC+
N44uJO26IRhXZT6L96/7hBMBGCunUQUr9lLconp7KnQs1xHS5EnNFurtnaiJQGYvDrLutAZ/dZGb
D5syuyDsuNZGbF7q2LV7KOxSnWo6ySRomJXl5EzHRB7WQD6niFwoMqgKoAvcKkHL1YNPlRKD7ppx
T4/mZEx6D3VorIV8Xlp2uKxEqmLHCzgLLoXd8huRuMTIPLIiuLRCC7eoH+d+BGjayTDgbtCv0Ee9
MI4+bUAIYk98dQmZ4lOvH9kdq3l/eQ1l65qBtrknbSndZdVNetvFYLI1I4cbF2iK/YQHrPdtzEmU
cOyHvltjF75QozKk7vtiZFrok4gj9cQu650lRfE7foY/bfrEQ9a5MA8dE3mqkyQRhVb+d5ZqYJQY
yiXpMFNvQiC373ReGE+iAzVjN5YtOHOQb/vddo/bVxyRmkWwypaRAZ7Av+inMlUEq4ZXYtJ61pCy
ZLGfazNRvVvalcP7P+MlY8zq2cVi3k1rWr7LYanDBuvqu81JUr/LLGz1oS7cx8grYVrHgZTUzVS3
bbePRXmjwM1G0QsYRKQQ5dOa9Q42CHv1A7v2skjfPNUuiD4R0U8k0qtz9duPae608YYHYQqbDeRf
o4SgtlQaHjLiWIwW5FWg6AvSRdgeT2q/RpDiE1+Zk8beptBFu0JQktn0jU4eCwmScmh9SCvmxJje
NCHt0+g9gopEnyMh05p2elTLIS66ZKM8SIJmIBHYgdCkLEfd5YY/BHG4R37fiqWOxKdt6ejwMNnl
5vbWQrSxNZ1bj53tDPsWCwjwJeoc3SpX4jCqMAEGQdwEs1SARbB68MwIyJt3osNVkw5/v3A3lpDV
BUD44S2p0WHNq98lzorQX/oPfe4IzO0rfpzqXgb8hujRneSJqkuJX38KFVRA6rjfv8umuocaJsY7
7iG0SAQhxakjfjQPhnW54OLgPIuF5x+bMQ2pAifPShdjnD1lGPv0D2Y6dIF/H2ka9Itf7LTHDxlX
v/vScU7FlLuOdiEP/6ypeqaFKXVkVhjVH4Rjxo7oBtfTqvRSjQ406AV7tGPwLAVypmYue9RtD5sv
hBr68+1IihuwU4lFj4iHBBG9EottIvrsovazbKWg+VpW1T2HYiiSnu/br5/P7Mn3GWtH7JQtD5mF
iasxCdiiKiG0h8FMNGmg0y5ef+L/k7FLNVxpoqrAJ6c9MWtzBDNLzr/x0k5W4G0r/h8uTOn6Shei
EVNWJ0AGy8ovzLY82GrGFgceL8IJwQnDb5rxkFSsUDX03sCwHxoo+W26Zxkv+t8KjOiwxNGK0R77
XDVqo/ko2tfEPsM2oRRCG1vH2LfHjM4uAXMF48/Wvym+Z9N1dg6w3WdHQq7JilF21Z4gyM/qGFhG
4nVgRlv1P5kkrM5iEYdor3uE7pLZnmdzHyl94yeF2ucdAMET564Huf6tgETqNqphCE+chJ3MtUSO
P0V5TbGTg1TkVWwaeeKn4DiBlOQRAEawtLn98/BMx5gJggY79IlG/pkmoiSw9IhaVoiACEzSAv3M
g96zXfnuL7Mo7ump6uif+wqz5Zc/+CqmsdTGYKZs7HXrSWpKezrH26yMktq+GOU9QOYwtimo7FAV
2P0h5RYJgwYSoV3M6ENQpJ2tIbDtc2qwFVKy1bbGUFVm8bi30zsvCHqaWuv6x4vh7fth+rB0XVui
iNw7r2fl7d/iMg6vTxmPHOhuEwDyvH9jspaXnq0tZcxkebNNKp42LXYHwXN1w/TqSJpeTCH0JTF3
eTbf+v0lTrwgphDVWQQD/Iwtk3ovO6QXIL5lZL0Asp3U+bTcL+zcZ81elrr21oxiheuwExALPj4E
JVb3cRHoDHJBS1NDx8qHtgRsm5s5lSgD5ZfiWI+nY6LKgjQ6sKC3nldGDyrHn2AlYgBsETnepQb0
GDI0v2spe3VWY+viy+yy6Or6AZ22gNYURDoZBRJgxXoM4hkQE0lu1f7Mkw3oBxVku0YTkKz69Jbh
49hZqats9AfNf+VpPIjH5/P+FQg3Z/xOghTtU/Z/MQLCc1nwXwcejsnSCmQvCEjp1ojaP1JetZNP
Yv+bYvSemLPzFNMWT/ugPXo1h0y2dOU6LzaYEhP7AFFlCBZH+18vY3C2HtdlCcx3nAKzRcDymvcf
DaD8B+Xslu5ADTtrpriW+DUmomTAIohlTuOpXRVuSB+a3aGgglIaiGu4N4CrjEHP4DezgSJHQE0t
06MWlRhPBJC8RQR975T1ERcy5AVvmeYj1H4CKYoxqCxnkuR7ybzT6ri4AGe5uh6qhYf4BfnA6Dbq
W/bCoCkzSWZojUrsm+UOSPkluvHRih2FKcmFmgmIHE2fqqyiY37YHdPg/+JlHKZIFm62trlARsj2
jfVNv//G9PVVDNbrNDtzTSWxCs/szjxNEDCLu2Xprihf028uBJZh16mH5sMlo55PQX7uQJSVZ1fZ
gCGpNiKko1A8qMZBWf5Af4W9qVJJ5ca8jJN3p7/Tl+rO8Ifk8NCkX7Gl53mc6X0n4GdbFM2rMnaY
4Esdik0j3ZCOgAgT6K2JohDNKK8lERqkvapKyCxT3qQaHVR1/nV6bxwiv45IBp53FIazkJ7xRtTJ
Hgh7A03xTLbxnX1caEZeCLMZ+PYWzvDiy/OtvX6aaIA4Ok+YsbyLzIEhNcsR1ILL2nUGTmJ50c77
lLrB0YrLHE0Pxk5tL06tVGqrPXF0H37wChFmFXkW+E+Kgu6W79DaWjW22anuSDtP4LRzfISv3F0E
pIeSYVkn3Wqf3SumkLnfRKuw3D3J5Dxn7S6I7BqNERja4TZbD6i0uRs9JXj0J8+oeVfMUwNkyU5p
zLMeBStsvGAAIVm1OUbkths4j/wT54G8oIr9nqAxSbuduBI7o0jDG6JMDdN5PExVD/zCvBWKrp2l
0kztolDCxs8PCppHmhBl0l0yn7eqhrzLB3sdfF6AWpw9l4IqhLUx8dqIGb2Yn9ThPd4AxcVtyvVl
pciZpEtorysc14WT3gjKCHVwbpsJJXCgqGKS0p6jmkO0Gufncvgi3LKGhxmdZTi8wkndINq8YYAT
eE5uHAhx7BUp0FysQhdGf/QQfULrXfFhIcH4f3ok/cIguDguDcJKK/znLC+zWU3xD2QNf3POPbJn
4q3UVuQeg3g1KzwyqjtafQJBOnp2AHv17Zpi+1u4oqh4AZzUYlx90GHrMbMaO408tMoQUmPsFq3j
Yo+aOfVE1qchgmRh4C7X8dwdSwJ8AJwbYpPgqmmbOJPRxkqEHqyhfL9N7VJLTcFDOcVWM3yKyIY6
iUdVz4hgPsYVKG8y0ATCKafDDj6aBfL38L6y1SS3KFrsAZNSZW+HttZVSrGdAoz5LN35Nzv9erKD
hR4bjtQQdu1zAUfm8L+cxbRQ7MCwKeUETItvOzi/Y7DMNP6RThPJlumVYGrAbqR4ebBPG0noZYiu
ifA83LIC1shHqe5JrRgjJGekEcwgCKNYgdcLtryoTkeuEHktR17lan8BZNabBni2/yImXtyr8sXO
4Luw4XrMr7+fr7WkGwAOKtaJkDiuaUpOMvXWKSS6UgIyMFOnZWzBOhcNs/rWa4G9ydu3mb/YYSof
Wn9qpFcOazRP7tS17fzJPkV+POdjAQlrxCtECC6jXsMF1YoIkzV1JNLJtV6MLA64Q2ny4AaCJ/v5
VemRS1XNyhVczi6OUXr//6Dhkmvl1SAB76T9aC4A1k5+QGBTaMOF2ObCQQXjRti7QK/agSEMoMDV
rpPK/8cXAMzyJS9wuABnzFVTKhBzA4glBRpuQ3Co/LnX6LAZepNxWceeIr4q5oUCfCf6GBbMwlQv
WqA0NQVXtpLmCJhGFMYy0ZIzosfpHmBQTqe8fpOafiRntiWoBVh+VetArSo1vB/VEFXxUaSNE1ee
4M6XuNGjMlHALH7t8W9+UL6serrYftKqwKiOE8OdRO3aKEjPssOmE0ajruuprJf295Qem8KwwRq0
Dfemd/CxcgnKJOf19cc00pJm3HufGZgrzgs3tB31L77gj+w6QqI2FKCjPEAi/qfawimbcO5Owccg
rtvnFgFS0twYPKpnN7+U0ZaGTT/MVyqLZv8iJA4l0x5QNFDQjLxTHUBKC5g+GhlRCasnTBFHt6n0
zo2ZzrdOPHyHpo9rK/wK5nKKcACIVt8WIaF55Gmc3EJy+xwaYQfp1FGouGrW86shJ/S/t/AKTfTm
kKmuZXdNohztgmpPrlB6nzXUtkKl8Z3VZW+3NJ3zbWdTZ1vLKDlWsUKa9tvmn9H1m76hg70t4Fog
goKuOy/iqZ/dPuCi248jcj02BYX4hRIZLgeUI8leAUK2Anu7IpH6UsMapLb23jvTyRV21waFbSpe
oImsqHFpKnjtVTqWgsx+WnGsfnmjDNqhwwo0HrkxfuGrJ2AZMfMw8zVKVEcDmB/813tsMkR9F4ES
hiow3nR120q7DsLS9RsoaeFUXIWYTGx7BcXabR7/Ec2CkGIMuzu/QYJUFgwH18WUo3TTjQuBuArD
alHTwCljU4Toy1cv51Tz6FhqxymMLHgr9eLNwrgaGbWu/wHpUgzMWv59dT93wVi+4TL9Geb0eCxz
uwoGStIffE4g1WieUXYYOX0N2mE3tCL8WCChBuzVjOeoj/yqtoUS+nbsv8M9W5ormhQYNED6z3nH
XgLR2Nvvk7vb4YTdUiOBEYGb01ME7grKFCMqOotX/2i+Ee7eqFqDsEUh8k23cRvJtGm0UeHLhMB9
IuNMOKyOwpMznbspevuEncNzBHf1/O9NLYobAUQHKDzdOVYKUqkikeyNtXt4ngQCSAx5QwZ20P43
m2UX5zJVm9HJingAq1vY0iu8AFM6qndmTzxhQA+romjVb5L12uGOekH8DuBp7skTIa7uCDI3ryVT
UQKKzkldX5jM5JO5IYesivffsd9in0CQC/Tgm6klAJe2wvDb5U56hIlmZhvckLtmJVe8B5vr+HDK
HSxncsYx7kKS5DS6cFRklGnwUUYOFU+MOjr/vVs+WuGAXLbXwiAoF3pSLyEXMOQ03Xei4h3HalmN
mYxJfh68JeqxUMlqgi+lEDS7CbCKMg0S52hvQ8EwkYmCmjgngpuvKowzswmFZdFsPdf/9lZ3yd6l
45hP8b/E1FqVwNfDn0z6qgESz+qquz702MmMI2JoKkUYcZpb3C20S9odUfE1ggfs/2W165QZ/REE
BV4TnaNYtd4VyX0kLlFOQcRlCbQUf7aM5HZr5Ob9/IEU+OzbvN9eRH9Jfg7zEHWtiBueEEMPf/yA
qBnHugfMwoqtheTG20Y5lxF6Jpng9otVb8Cjg7LhZ+0rOAxkUb4uGg/8q+c1igAVb6of59+92ugU
4HgU4gUzwfQ477rEOz7KmSGJcqEHgeRzvo6DlNPOCwyvHBk6P7DqV70HhVenI/LmASQQFMh6JgCm
L6TN2HWLogPJ1VURo/2Lku+FWTHeUpGiq5FRdhNecaVoVMk43wQaug6u3l9HZmvBYb+27wyntrky
3oObAKj2VsqRTR7mNGD49J0WHXVXOD7n7vx7E+DDMC4Nd3W2fVhHg9xulpOuqF+FKHEGjaRjlhHM
Kj8XGee9VJvg6byv2yagoJUsXp5vhTF6XoXfF6zlEtKOUrTH+7mvHJKoA3+eiQfohIK5qYpzfwjn
QjuVeXLLL2LYHqEbHWMPJ9MnHgVjnYKWZXSReXe9vPcBZD6c/M2rYC9DGNQorip3Qk5ouTeIVC9l
MHeb+zz/FTzShE9la7ZgnW5+mFWVdt3tRQUngStkYLIqMmHHQwYTUAtWSqYjYCtgmv9sNPCZh/Zn
9fzFzpYLzp8QHExgF4cOPgRHMNAUpDjbOUOGnzsN2besCsZPg1b8XPdLFh4V85M0qmMmQgSUNBbx
V99mUynRjd18QV3Fh0Z+7R3hB1pQGrSWgstunE+bvNmY2yPgWXp+bxjnn7PjejFkRcu4pTzo21NB
A5mHxJg2/GNDW7I11dz90vZPTpw5Hr1HTGIvWO8dMtPE+ytriuXhPxHt6Hs0HmpldDYJQFgmfPND
IEuv7R6PJCgq5dCOjfZEmTHWkokzbzEbdI2/QSQVP6tObbdzv0C5WlBz6rxe+I3aly2PI34NmEro
h+XwN5Ru8baQI0ePVQqQpHNe+h69Cug18suQzzUNzoWFirnqn/Yn8FZCF5SL4GMQvM7OxF8n6lnr
W1KziSv2TjZ55FUx36QFnF2a/odKaM31dHpW2KCHFVk0TnFYnlav+CEAkp6Kh3U01YrTbhk6+X2Z
7DPi7LBjx8a9GWv1/ULde6COoiiCkx6+KHUuC9/LNUqslU/EvvaPivbVpEriF7db+hE0Ov1/ORjB
jC156y8lebYxQftN9tgp66vUdoeEMFsZElXNoLVjiSiO8/YH2HoQTLW+AveVhP9wAa4Pi2KOLXej
udTyDtn+li+wn3GKQVdjm654NFqYruU4mKrmGRp4/QEW9YqJ0P2/36lYM54km7u9ueLzYT7nBXBI
HY6UZGIcdrlowhvyAN9QBadd65OJP+Ijn6nRU9KpE4DmTGaIy3vj/uMBmhOLJ76Df6Mtjqbs2peU
8m2yezghkoHfUNCc6LXxRGDklo3tkO5Bp3r3CUpd8GEiSz3tNtYf8V7ypNamZngjQR2lqNuTyxjc
gncUacyVNSGctT5zJHW4bYOwKJy/7C76xcTX/NGvFYcf3bcf5aXnZVbLm7xcaHe00rgx+ewcXsPT
+/gKT2HrfbdoanuJSUt0mqcP+Ke6qapMLOw9jCC7UtN2iFWV8dCy6zJ3Ig2OUHmy5AEfY5YSaFqC
sUWnwFkkrcx1Zr3JerghHB4BIjr9LopyQZ/sbDMNh5uEk3SrCyz8b8qiYfSSdJJ9zm+Gt7d0OJ8u
YzTnDRwrkkwHwoXV17vZvd11iSogjGEV42PI8OCcsgjIq4bXwxDRnSlM8xBkV0KF6GGGDZxQAkvA
VE1gG02YxaDwuggQVQuZJAyOnLLClKmsQO7Dd6750o7+85ybCCEh+pilhMHansTyvg0OT2bX/niO
btX2h8CKKSzt/F7IcBt+BvtY+hfxTMi1Pt1oI1J17rQz74alySEOtyAawj1NRilsmHCom+7nrFwd
TbjKyHcPYhI1xREfl4TNcvDTkUyCYhcDMtiNVROVd7/E8X1RAdtZ99QN6rJLob/xp21oJNqcXv7v
OVz9mNHGvINNpy4pffAkeNjPA9mxx3L5om2MV4AAUVdX9ylBpZqCTI+MHPVKfdHQ8qa/acFt3Qa8
Lp7DRajASn8ri2UOor49cu5f7IRscBapGf2du2vIIqOIggLnaEUsI9DS/TF6n3T5A5JEAucJlf+5
7KEaPaPXmxJs5mJfE1cKWG9W5+sqbOpp1Y3otGp8FU9mgnkBG1WFAIm7+5jCESnW7812sTI7B+sV
HA/yOameLJZw3iyj0wTtJET6lyIgO80Jj+Wco/LCMXnjjnH+T4Tie9ew9DPDeFF0PA2csnmS9LnE
E7B9lpWe6eki/pWuSYEiV5vh1xjVgOl0giQ0oocQHknuRNhM/KMD2QpQO+/kykjXR/pyg06Tsmbi
qin3YFUqp8SQYOSxm4H3n4TJKxTjio2AGtVtOnqs6q4dbf6/q7Dc3pxggCalsRGmCmpWqDkvJRbc
8VKVO0JlhHHvvK7I/xK/+ciEe4oloiqoc+ykU9gd65arK7GQR1CMW0Xm/6jiAKSjBIswNDLtYLXI
FdjohPCDMcwI2CIWeXolNlK3EN4ESn8rzzlr6exdg+90XFsySzcCGzQlE6Huf/+3vNHETNy1nSLS
/31e6C7lTKhmKeDZHRABx3Ooi4DBTfcA6GYYHmvgTQ0TS4LzC6uvwpVPlSOr0MtyhM8xDgkSGl5M
Rr6LMGvDh0Sxdm8++qO8sWjCewMkA2XzHU/Y8BgQBMOAkZFdUi3gt+aTC0sTixmKL3v0fLIBQbLO
Ds+6ZNpsMXjV9GN2+WZFljUhWSHrK0UlJgEsOxuPffXE87kSQCekFHiZNn/HMvxiKufsjALSkivt
CdrYmwILWRRcNGnd8cnzt7qfGUUGbbvF3A+Nkou8m6Iz9gsEsKUzMYhY8RbT5IupN7dg4sR3mXTV
l3169CHQkOSxEgP4rXoyD5pJ6PcoaNUoXKLTvR/wHcKt1R0DD4rF9YUBpCVzODtknNwWwlzY1WEp
OsGQY8B0qLYIA84DywIi1w74aUHsX8t1RjWxnC8ky5YmTY7vCBsJqbG4L8aSNASADa/mdIzb3lhI
iCcfr0G2paXyJtU1lL6a7Ft03e+tNwTIYsDFkrSuu8WzlH/f/PFLRoITJSKplMCQCeiKl8XH+/7j
6/ZNAbAz0g+WAHHeyf2i/glO3mTEFZ6aWeN5bbLBQnA/JEmdwoYFO4cVjHEr4BsEKpesBQhe/jf7
/uUfLh9Y0T2VD+hMaU/ay5jH+APOQuJo29pYJ3PZD0wPZKQXS3cSMZrUKhXcs7hMwzBoHOQ4Ovyo
vO1GzLbAkINt7QxfmrIcgAoeSzIxxb7lqArnyOAXdHS43YNlUSm7067A3sPeXqLtb72iMw+qBjDZ
ET/Nk7NT+DWBE9S5h9VL7jNLFQkazod03fh31vdwzJcvtvk1iPlyDfBj8axXqVNRM4PYmwBLVZyf
kkouuTBXfK2HaVysIh0d8iuq1fPteB0aTjb0G+YUKirLjq6+6gdcTrfazcrrOkJoC7Mtk/oxvKAm
gUlSIbiCS+s5uMvYVtmzyd7RlMStogJ0ycXBjlvuRidSyCnXjvnBza71QQWj7q/K3Mv9/l3nfBg/
ezXRhQ6PHBsA+fnWJyegz6LKrUVJVu1DI3k/LZYN8vaggJd4bLEuSR8dZx3yoelYakyv0phbVl7Q
vQhk+qqtmf5cPX/MJSD2qCf5EHA4c2dfQl0TNGA+/trbKBRMiMzEV4wbHHUkNv/v0dffVW16swZH
x9KjoWdjI++XdFdaTTGIQnhV8pJwRQnUpqNeN4V5uT7tnf7fP6qXRMeaCbnYyvVmREbvunZpXCd+
dysLlShmyF9Rkv4MlzZnTh9H08D6xOOPauCzCsPsR9PWFLdj7AScjl8M7sMqnPb60FEsKv6EOFPT
rij1MroKYSLNB/rEfe0Tf3Zyaw7P1DtWR/ODV3Qpq5fPKb4aow8y7vvoeUNoxUQayXqBLWzjv9Ps
cvrJKUFYAV+fpRIiLxVjBoObyFrXBWcIfrbnxUYOEF+Kn3Ty7jD9BELHlk/l4hLcgEvmsSmN8+Pk
CuXhiDRxzR23SB3fvrRGcOuN4bKbaVnuUnXKh9F8q/ra/n2RSfD8SHlhO+2rmSh5KbgnSqKsQ0TD
uCOChiUQy13vKG5/q6KbU8/MyvgYEx0kAQQhNOiULYLNYw1zpScajmJf1/2N+xeh1dJLT1IXdB4B
RaPWsjE/FsvoOPpM82h4VKd1nbcra/Wm9mMSv32gY0G7V5mnyjF3fWjGaZPewrd1faCagHZMujDY
CTy2lC2n6x43eYp+SGyXwIYbHGV60XFY56/BYTL8awHTvpUqk5NUmJTqgrjwL80/Odf6XLCkfHhl
XhYcMYScp2aoZO0o4SSdj50fJUtv+ACIFkRr4LqZfQiKPJMJVeaaipWwEYEkrcYKT8RJaO2BtwyJ
rUGE9Hkw3Y4EZT9eJQ05s67Gt/bWj36lrS81iCsEigcVAH+ahmix93NRvPFiQB/qtM0NvCbffPSk
X1IQzA9KeO79rBcjnTCg8zEArpJya3E/6anDnCLgwMgXbFhPFfAP44sVEU6r+zv3Y3cNNya0FZWo
7RZto0chO1PPxNMaExw/5mMWkTFEkSEKgmahsh6TguhOuYZpj/Hs74hhvNVbu7S1JOFTq7XUVMGe
F/M9JFmWlbN/nNnHaN2OQMBMjgGFqgHIodWdHTCODmyMISPfEKF1cZ6uHgrB+nKgT9t9QtQ0OCye
CdOqAmY2kxV3mYJNlM+AXdEtwXPw+NwhWRd+SorhRJZj/9JQjC1AeuGYLsgIWFxwYYgZRLOmgd3r
m1TVPqy+rgFBlKObuV2uK9tPflXzJ87/8p5bMlGZ1A8C2RWdG2v/N8//Ng0XMvuMT0U5Zw6bzOai
fUzZ/86+cwzjGUwXh3+q9WUvZdlYHVy+qTAolhVmsLbTqs/xPAcRfEZqclLUk44w+MD4waDsK5E6
H5Dfj+4Cwx/Mn/K6tp/d8QPbbZGfDwfq0EVLXsS+ukfAaEtbWr9ScsgeUL2u6Sr6gHvXSOzJ9emc
c7e44JMLf7VTJpnVoO8biqE18t3gL23ZXuWmxm2IOrhZi6IZO1OxkGg62rzuAk1Z+PyR96wdOGIL
kK3N9nS1OGvUt5MuXYmcEXjm2V0Y9K4uEAyMGvugRpC4nwSzJx1iU1z868kzMJ01bCQfVH9dGjwj
z8czp01WhUVKHDNh0O+fzOkq05ExJGV+V/jn8iXkGUJ2od81XTkBbTxQMo70zesCCkk9QrqUiXd2
ZIg6mW1NazS9WIU8JPsdAfDXR2xbyBeBzRhxvxPjvU1GxxADXCspK18tqry3Mqe5CZfridLf08B/
p5Qc8IpSI8vQvq+gWYApKUp7BagxU+iEWImGH6pqeZkBAMQFfG2rKNlOOUEfTVXmfznYN4qRoQun
GG+2cShj4fZEvl6wlZQ/2GhdQQUy064HgQDXQUNUVmepZg8pzWicON6f44LzbcBae437k1nve97d
WTuS3v+w8hucfa/93WB4dYAziFkGWMlIYamRPxalRhsDw33Kr8wZkzkRvT5vfWUapLL/WsFsxcKc
MdiI0HdrcvNopmGzQoB/ywp5qFLGyNLezr+yo/dxarTUtEoHUdwWOONIWfy/yZ2wu+VvrQIX5qV+
l56i1t3SvNGfl1yzB37benNwqw/rixFluDm+gQFjBuL6c44LXjr7zjcPmmmn2fkA/b6RkiXz0OCR
OSMzoUNaM/h77WiKOYVBq3MJQMCoRcIK0xLJP0QPRL7kobZBYsbny+tmRGTZeY1GLOGimIba9MKX
PuvR6ypwo8eNQGS9i9mb7LLGovNrrXWSmMRtqmm5D3ZNDWgSrPGh67/9fwW5QILdRpobvQ1QTb+M
WM3UstS+CFOemD57DmJIEs/ToH2qcaAAzxAzBqO6gDsv0LMJzQzUCdy10T4PV7Gcl8132lHnt9ez
+3a8kR0tvJRTpOAw6PK57tDx8qwY3JTO6+JRky4cvx/5RjFqqio+kmHwBy1VNH/VzaL2NkbY8eVi
6E+Vo748ZvvcsgTXNdMNoGIO9Rf8k3gRqXdROGU8hEUZJJb7B446SLp+BIO6Xk5K3Ar81GNdruME
o1gOCgQp43Mi9EvMzPH7c3iklNOsJctdhfHRfJqVL0pPkNjc8S6wHbH40hPJ0OY+lE0so1IGVsyr
iuN0gU4zL/XDKIozhUOjiXGttkpZh2RZaaJKoYPBcItiKgKVrLpduUXLWpEqASkK6XoynBoQx4y/
UfwyFhWJxtJrFhyg+f9w7A/kE8KFYZ1E3HLMUckcMmKZRA1OV1R/Wnb/mpV9yOlG8PXpMjpEp89h
5+vMRYHKaaQUfTscQUZx7zfpKRVf76u5LvHoNrKDoBeON+lU+8xdnKY7RusZmDtJwkCz7irqh0k7
ZnmdsDPrsGe2z26OkvIZIvfsyx4akEG3V//pg/ynOY8hsZgiEfIieWgT7OekRHOddLxyett6QzK+
p2MjaUCQJJICgU5vMQwPLF4QNUMKui5Rkns3eir1MgfPEBVPlZlhH2kyDUkRMtl2rZ68AOVxn3tb
CVf1TSP/1F2pAofF7SxzjjeXMDoRLB8p99oh5DRKKyd/s0yGaVVqZ4a6d00FLwOrdgc5F7jOjKEa
TWI3hUXgDIBipSuzdrIAxg6SeLaeeasr652UIXt6ta3hct2ZIK5ZucfszCCLkubvZSekSVksvEbx
1wd0kxFEKxTUfj8qIqKrVfxvS9boQ5tIeJYw47bzPpUqK4KUzFMji+qzMn7AqusJKjuGiP/wzAbP
9sDOVWXjN+FI6nJGao2mn0kKOZGboPGhLKVnjj9X1TPLfv4bdGkntbwvRC+/RVKkSwcky194A1l1
ZYdbj/oMCjGZkjnvOIJD6qw8QoNjqX683SuGiNhM/IKdUCOWhny+nr73ul18tf6fOWUZzhv3SB2z
orVZ85W/7BfW4WVWUBMy8Tfn5mOVbV+56/a9Ey4skGMJw+u3K2Ss0NPScEbb6Ltwtjr6DhnyUgdO
tZflOtQtIKc0hueunh5AwIA7ed46iopVBOIaxP602AEXvfISnMqwCKS6aS7gmNBvQ2HVzRQpOdiZ
IBl4ZnG+mjmz6zllJ6jbiNfN1VIZAv6PYyhWY38QFWDOryINRUKttosNfRucsnQzKCt/LzebuYOE
6TtbVoVZGHFLTqYJyVs3c05Pz8IqC+51Y0nfaiJLwnT8+3M7un2ZaqWFVs3vsFMalXKtVJqkQwCn
sYbRKFmSMo6P2/NyDNcZkvBEr/Vsd6IJ1y5Ioib1hV/Ym9W/Gkq/oLt50aYCCqE0tuqEPK4MLXTv
zyP4zg7jwIVu5cJ51dWBkcEJ1QqYkDo52/f1kCnTdp3wHA4fguHmiaIr7witILotBZ6m/ZOwzeKg
RZsAjwvRvNo6xcY6sCwoscy2CGrQDcwlpbQlucL56AN61+pq9ZtMsUStaoVI1QUmCUVm+xnxzcec
Y4PJkjjDDhQEwuu2awQml9M5OW1lNOpdvUO86XT45aJMVnLVCgSA4vP8MO0y4vH1ob2RtxEhf+Yh
BaQlkMHGQ88guxeapWxTSfZfYb53RL2SS6Of7seOX+NYklJceUq9IJhzi2QuLv7rMk/5/mqAbNZ/
t6eqfjm4ddVKzQNzoIrxQRmLSyKhJETJ1jAuuK8GhFxylF5XZzQS7/eQ2/hSsUOQFZBAlJ+nfHSz
CcXC60RCAdDMnZYsYK3sElewO63OqdWPIFzhqoPy/J7OAEMyvM5iUoKB5oR9MSG3wQBrAY0Z1Zl+
5SIQEPTyFM+C7VpDQJ4+hKOHoOdkGnFpbf203mQShmM1Mjh4bBAlY33onXG/fXw/LPnea8Q4IEkJ
CWKTHm7x4LA+BfUoz27GQs48MJBBmnnKXbemDpbu2GP5pMLb0uWG87ChsqcRWHFXGWu0Do8HPdDf
jNarLjJ3Ogc0fwaKlcANDEOX3RQOJfLkH5aASOWWTSnWKYNoJUOW9jCz6/HQE7M527iRiEsMXg2C
5ApMZAMlTnfg233wqWOvqPFupnwwhb8cOVlCIJYPLcLPPJQm8Ukbi4vj13NnbwEe9x7sDxXrnKzY
GGvvGPzk+p/mEcg1eKbFOtlmI2R+NXdxrmEfeKmeUhotP07dnbcHjCY+2+Y2P8KEfzxJhlpPfydO
1VV0WFpHyUYbbAzR3My8GAEJbW2O9RoUGAOlkR5w+3DNy9pmGF0Yzl9y12f3A0a6D/Wv3nOh7buW
dxQSEoHxOLVME0MgclaPmH007mCWSXeofZawDQTWFz+xGK0Gs8K+3bbvDnAy6LlUtSoIO8cPCECu
I7ZlIKC6truRcxqIANwygmhvwCtr22SuAZWYH5UQIWjDQIpaGjDP+nxulkZqg1Sqakla2vV5WKrL
JTtF9VehRfRa+jiZm9ijsDFx7jgkdm7CQ1N8//ifJgEUPjHJiECxXW6DoeT+yVKCurvDdtmC9e6e
76paptjdR0C6cAxq3zHNgo1ctO/BSsj8a6hP3ZMAeWCj2e0Q2rGI6SDBby3bDY+Xf3PrAsji5EBt
MwkHoiWC4G/PLzX8CVRkaKqhsiYhTp3vurhUMrQlpZ2+7KBgaOYl1DR2HI6MM/YqYWOTkvD+eFM9
0d7hSxUZ5EeYbSlX0QXjT2dV8PwywLu2cyeo8cTytfL+mUR8Uw+eOmx5YsYqz9Xy1P85Mim7D9I+
fujUIltaWgZ+YVaIPmufByKhw84H0RpsKRLq8ihlBqXmk1ytuT9MCxdC7upmiQdIXJDbnL7pqiUu
huYwAmFwBNN5zPfuzd8tRP01R6P7SEx5mAbgmOWCnMOgKhMGatfDue5uRJuKc3yt/ORzrB0xj+XP
+fMo1bFMrb+RFD+XpMXsV2UfJsIH2+aw8k+LTkxojfNGMXPGxxOjf1gQ9aAnsMQS8toea3cfbvse
0pcTJe1jCH3GUAh838xJcC92/F7hshklGORSxEamDU+Eeu9S3N1i3nCYQQk2e0Qdmlo+2Dgd1Oy2
VQLtSYhOjiEQv1H7PbWolCEGc4NjEQMMnjlEQ4Yh4HIjyyxUALxE4+cz2YtS9o/GMQ1O1S/0yLhO
jNQErCnD7LWzHv4DzjTdQZ32Y0pIJSgvpKCWs7fDCb8zJrB1ITTafU3ozNMLYEYDRhRDp2sVIXXN
tgCN0uAxhuu0EM8VH7Y1ykXNQjMhHgmyvWrCkGE9QZLsedOyeWK4sdDIVNXhIgEZZiArlTpWqcNf
JqEahhFKnyRAWfoEUa3AABiH15uSSLo0Rz726sW8KxQbAl2BKePoSV+6zOw5EhVdBZa+Kmqz7JS5
u5nbj5Bfu5uT6VapkL7rGGTgcjA7R38v6QiobHt9UlXPX+jxZyoCNamGdtCYErqrzo2002xQKafx
eH7vbMFSHS5NJezdVKSvR17M0INil814SAtJVkXMqE1ymmcH7UaeW4b0+/28Hy03+8BL63o/xxRY
9bpBrOKBfkfl8FpT2guyODE8uFSyakUEz0xIg5lsj2//vJ3PkBLe4MLzGThSdMFMYrizpbpJUP3G
Ifr5lXuRoN44kpKB297GVkJVHtLtN3je5o0QYBckfsuSaK4mJvziPToo2ItDyBzCjjDQAIxtv6Dv
yaaIGPlYVqbCp0A1oHJnVlj5tS05AOJnS4YA4Ok/P3YtKd+luXPVdx/fYECeo6rr5hjYNTz7TBTo
N4g1ZYBK8yDTUV95Ai5SHtEy2LDnvhKa1BQGwAZZCENG8SpMNAh22Xz+J+lt5yKF/nqTKKxbbwL1
PlMPrqnMUdVLpgJroDwdFVYvFrGdW0uhuLBEpog7CUo6fmLkfSbs8B2maEj5HD25OJIYksg8W5P6
rdi+o3XW9liCxS0iONc4wSkTPn4ZkK4j1Fa34c3qbotvdaFG1ex1o6hve/C0p/L0m1vKYNeqBsf1
cLfqRQ3FDfHUA9/Fgl0zxFyFyeKKzzpH8A3SttlEuilfSC9VHYdOoYfCDLfI5jdip/wM/i0T/E1G
m/WpA7cQ35m3XbPLiCBVT0wA7nIL+Z/vstG9GLVBbVh2xhxCEcer0ZerE973myrBNgldrcybfN8/
WAqs+czNaLWOoQR/F7WQ0pcVv8e2HcCIWuEKUeYi7Zc1+4tW39zYzsbZilJBpOdtjdzj/2Z/qlm3
B65wbCD3pxRZYuZPtYmvDsP3xE1PQlTfQE1wukNIKpBQl+VBqwTPVKbHBMj4+j+UbweJFeDKSaR7
hYCyuQbUTg889Q22V9r4tWNYGDODsa8XORC2pc4iVePV7WMeRTyzd6Oe15VUHxlDE4oe5bmI4ynj
wdJmuTrZTHqqYFR/euMtvZHY3a3q1F2gB7wJh4i6XiL7mFxuaCjz0Kcqx/Fm6jHF8kSbWXBOH+op
cx8edP78XPeFbn3f9MUpwLcxspLbLtJqYJTLM8VjzS1dPoFgr4nySj/i/temfMTloYIgjEwucxPn
BBkTi9p/U94Ei2ZwkGao2VAA/l9A9a01VWR3guGgWbHEN+JH170DESK9mxLeAL1szAjOmtXkYqkR
1c+EYBjjuhDxbCh2ShQlffBGE7Cs+o2vdrRINcGqYIUH3ztnHl770G8+rQNdL5bBYR2Y3IL3XaEu
gvyUmNz5/3zMi7ijsaKA7Jr4PTGYgorc8VWFodO7+gFQR+2xoo5Qaj84wZHy7CPrDExH0dPgy4Os
XTJiA/OX0X3NsTmn6rw+7Ml2ldtRFV+nc1fM8QYVDuymJDI38zoKadflexRzg+IzX4hJi4LNYuwL
wTwHxxBr5O5jBLqIsMWQknZGTrVQ4mS3A7NtGr1UXeB9pIL8MSq8ziYBXxNDCEXOzWtGvRpypJvm
TT5qoqtF18RlT8EOvofTs32GpkZMkW9DKVmB6/kzaPuQL1dNDaz+GF6bEVdry05Xrh6ZM8t6FAZb
Hn4e5IaDbINscziIZeLvIFVI61T6CEOhBggZDAKV1R6tswSMnhLZhriuYrECmlqgp1nSSSnoxeSF
/UANo9zISx392mX7eG9b22ewvljUohTPWLY/QSXusOFs9WWdXerjHvWyK/suCfR9fIri9ikSjepR
hjrk82XJ7+cu61pg/1mNZyiKUr3T6+kEEJ+AnlP27H5SnKIwE3gXoHEl7aq9jMuA+aLL0FteoPhc
OA7t7P1qUGojx/RNfMxd4RF+1mbf6hRRo3NHoPGOFYSoy1SVwkOiFksSOILU96/L4VdaZffpplPa
bgb1XYeaVR/5xorV7aDX4Kw48UFhCyYQzvkMqVlfnyLxyJyZa1Fx4GDysUq6OZrH6qqcxQNXml7J
EWcQOdk9iKYqZIi5QwnK7LVC3joq6OsDH5e2yqLZyx4rFEJEFsokYVaPaGPHTs23/B3cBNIEABqQ
Bav9WHbh9nfxatTuSI4C0YX45ymdJ83DIDby19SzoS2hzEQQU51sF9pJOMJYdRUjRtb5zmQYihXd
iaqcXexm3kcWLViMl2rOjx+d/HPnhKMjQ8+zChAjD31t9WTyY0HpmANUThW2J4aPCef7vbmZcEdD
6xpcsJg+K4Bl9vxk2ZoDVQlJp1n1WIbskVP4BOozCn0SQ0hpsXjtPKVgt0fAY4qCFKOgeLQUDYBE
4bP2Y75WkxMneR6Q8NIR6sxRLTs8C+eu3okqdleOSnngXkWU5rBGZllLWoXhJYWvpSnNaPdAVpDR
wtic1qC24s6Ffcy4QNWVMvMxkEX70MOc+I7mcR3GeUvXBZ0fW8a8iMUoV2yOsxRdpykN0gvKNq1v
ZDDoX4voGLIp/XpnXurK1fhecD0aiOM7wfKrrPqoQfHgstx7ZYR/wQ7MVCOmBc3uiqrQhzrzWM9N
290fPXO9gCBVpFJSsidoh8UbqyQG2YkGU5SHOVRsd4FnhNpikMcADUPPb4SUpbqBTABhPRJFjSvZ
KD3p7fBgl+cHZ11wIEN7oyy+VN1387iu0VUhYQLLF6mnMzYfhIxhDqa1iG6qXvu9kDzHvvQNS7fQ
KvodG6CtOUt039HmoSOOAUdVnMMGVEWvyKRgnFtLyABWzh/5OiE9iLgbUryjQN8c3YlervZiHeaU
dnTpOt+8P7j/y8vEl7r8UUpmFn8TsOHN8dE1bfZxTlZraXX+GqxiDo3sYE58YLJWSH0wxR7M1CLs
jd9ywGsLYhpcQ2DeG3pviashUbENPQa7nsTjN7xt8/MTvaYu94pCrzC52Xd9DazB4+uaPjWGB9Pi
06D042Lf/1sN3Wbu/lwqpc4yQZF7Nbqb311qTHXQxVyeMVVJLWBlX/mwY5gr5OMq51aDASXW5lfu
SLDBWIyZgdgt6npzhXzANwpd9YmIDPPsnbrrGCYU7aWewKTGC68nRt1TFSE2iIdFmS9wrMITxx3c
AN5ZQ7r3Hv/ati8UFraqqMo0nHanJo4aLEwYcQsvwN3QD0jIKSviKpSMjUVnyf0gEd9E3Rm3vjMa
in0ve2oY5cZFbNqyWsPACf1M3Tb8WAYxQfMpeHck1ZBWb9whSbEsB/EqO3eSOvgDHRi8Vdbrx7lY
Y2T/ZOudtJmzct2lpXryJP6QUX4qEhDn+Y4e7UlPg/R8QBMshfkWEZ3SWAA+Ju1OK8w7BBVR+YtT
wU7wmECOhsoZK4rqPWVwr2/lZids8Y8nj+1KN0KNtH0yqAHAcR/yv3XiCt/Oar9LRPN1SoOkY1A/
w2Io0+Kw3uxhnqFYZ6RCWssTRmr4T3ajFsmSdiQ8VeGbbuS85EuzV39IWZ53E0tt+dDi3bvvDdzB
r2Bkcnb027dHev5Vu9jfpRRUNRJ3HUESFRMqkGHB0KexdB9DwFxP53p7sCGZhQkNSG1WwbY+MNHa
TW0F5hywJAx5uaZdPlHXwq8BVflfssg1+TxMthMiy818YzwhYvIpmflAaL/HH10KKY4Yqy55O/3t
YEqTBlHjhsW21b/PobG7gk7H7QwFaOVY3GxZmnLVzBSDlkcYH9JMclsdXqW5bjNggXAvJ8/C9S+i
cGCFmY6CQd9LS5x5LAaXa9IlOQHmWkmQK20sNM4HKv+cn/XsCGK92c3kSkOY9F+eaLBDdtMIH9Bn
mXxYVK9MCukLwBTAvOftAS+Rihd/5fsDDe7iCY2rFUlXkXYLVEYZfWw3P0axcXm3sFKYm98oImji
JMMa0UCtOS3GvorCBzmK+uwJEQt42swKw0tmJk3gn3+4NvXbUzkVlox7tAfkKPg+yFocflVCCK5h
5yKERsAnZTpBZhnY7b7zcFkRcLjzYOjj58fitrHSDmO5pnoQFfY2QEdHWCbLmIrdHuLiq1JpRUy9
pjDcdUp1wF3vSP4M6n+XzR9IZSe58vZc6jdku4rcd4CNUZ68TVHA3ZIFgeK6fDkuIwO8TF1YzzRw
XSu2jW3esFAkIBkzes+Gp0oRt7quW+ThiAQXlRMrOQLe83qExP0z4ZuqPI+ILRKpHIvdnxQY6kUI
3VlVYxzsMVN0zwYHkAE6jHVNjgjnXlIP2mKSwh4uKDXNQyDXB8vF0AIDREfeS02U8evia9NhxPh5
nHJvnkuxFwL0eDXmHQNP7QdGABG6mHaAfR2xiksWIdcxcWZTqUuCVvIrrqFmE67EXkC8b7orFQFy
k0YUeCK7fkM1r6KZ+qe6U+215SfuWF64DZF1WQMp6QOfFb1GWJgLfrJ4iu1DSlqGxFPuxIfwfdFb
8i4ebz42wRRuZZAq81+WWWArBrbB4nLgBQgv3nvuBKjr4DQ+A00AJ6tuWXOp0X+mdlDGmVfclumn
3Gr5sLVQclfNHt8VhCP0krG7rY5ukz4cWL07zid4K9OzfZ6csXWIsTq1kNRHYSiFMw3lFGv/gg2v
OmRdJ9Z7cCLiK89svtSkyEUmgmGAdWO4oaOPpdvGFOfPe7At9GKG1YDMEdlppAocLRAFyF+pKz6L
nnAAE/I6p7XT1vGsWBJ4CChqrwON0zH47bkrU0M3PGchLY7XmevQvBGa/wZJNLttt2B3FabNqOyf
gcjljIDFTnYQcuN2zixIofJXttiImR0dvnVz9echqtndTcLkjEmAhYTYhMZmZe2gCk7eDJ83Zxp+
0i5rwhn/Zi05s0h4Yl6BD2E8G6L6bVL4oJWKqazlaqZFqZhFgaHolCihbcG4d+9w9GfDZgmPecug
TuxStWcAISW2cABy++1ZDS4RvCWtyuABgStkpSRCewhUaegUhlfzvDNH+akNd75of7Nh/OmumihV
Md8SbsTHNzJFTaD76ciQeLWnO9/OlzrLOLOuZUxgWkLzXhaK2qgMoq8UFEHwF2h8c920ux8lFHwa
R5477tOvF+G4E7Cn4Bw9fFwxiHNkIOhLmZ/xl/xzm3ntM7ioPTzxvXr6xZtPKFAoIAvwsuUwu56I
b5H276+blSaOcgbOsKURKmUX4MYB1tKy90i8OxvOvCN+EFjW7NJzg3utYEAkt+55nnn18dZKNm8C
sVJPY2XA5NLuXxK4Vr+rhGk5OmCrBXocenA38ckeNIA6QBpLeJWgMHFvdvPsKcF+maLjlCafjqZs
kNG3hQIGnCPE1TSmY/b+45oekapi2bxqJw8EThOGQxyPXSkoH/YI0V6SFXEAZnu76QhozrnJIYp7
MCfwCoBFkStcm2mOnUZiGOrXnbbpt3lpL+1LKQxMj4RHNyzacC7Ul29YyaflpB8PJCkX8+JRW0+G
tw2q7HbGideDKaJ/2Xsy+mShFqrqbR3d2BHPHNHy3ju8ZZTPl4SCaoL9ACTuRGrgzQBOmquUHgxy
slS3y6J+ywbwbdivw4YK5uwPIEkf0IXLbQ4OpfPcpMyPwXucf9vguBH4nZsYcNxB/i4JDxCMibiU
FV35z803juESQ5UCQxlKJDAkIGfghnPWyBTx45a4N1EfXj8ilnMY+c4JedORJM09JQXvVnETRBCO
hcN4K+a0bqYztrbcuZQ5lYOJVYIPkOqUzNHAOCvRSC3DYoHx1cZJsrou42iZQ97r/PMmjKhbTozc
qPLb329LIxsPdIF2yJVMWljUMqwuRagsqHaqS4Y5286SUh0qzWeyahmYlibgNVEgQYUWbdj/dUg7
Ym3kL1G76wvBjncROWoaYuF6RXn/r0xcI7e/3gbQSMLXD4th48Y4KjCwbaWSPvH7e+FZeqxDifVS
xji3xeg4hYg5/FMw7VvxVzeuaMoG9AfKqNcCs4JoBb38IKiC+aDeXFEtIRaF3MHKik2INDukk4HO
GsV2wK/raZ9Qsk47A4ZwmgNCkwT5Oqs4kq/dBRUZ/8+3F8+ndb4X2tMMRhljdT/VGazh7umCLY1E
+A71kozSeXgIMb2Kb5E81rr3gJifgMyGTKzidfE9CaMH+qxgFMcHyW5HxXAu+jlw85XyKKY9ZKaC
AuuMkaPnouQFa/+nKeFhMol3VZ7W8/Iay2Pe16CFRVX89XMUWFG1rc/XjozXvIvE1xV03S8p3res
QDypMOeDCD4YBeZsNX2s0YA+K04Od756Zn+mamprx8EOm8w1JTElOD1YFchRVVQ3lsa6qaGcqcWy
435KBfQ4mdKkvyOLCU3T+IPiUcsS4hviFluhtpjyRAyGfN0HBcag+/AmpRIyhsLGmnAGfWKpkA6+
a7YgVLieeSL6ZlzH1SG5Q0tU6U/Nc8jmoV42zHTJFn6gPDazdvUTMERlJIpvYX6Ppt/uLdQZOX3h
Z6vT7aQ/bCmwdpwJNBJeFnXu6HZwk9twntSaNmn4XL2WDgGW6JFnzBj/8q8C/pN68Onoq6tuW1P5
gcTNzGdyu+qXTj+VFc+skrRtkvpRG3rzH5nSVY29iIyU0XRLZ2l81xQfPNx58m81EKzvnrI/Qb8g
U2ryBRn9TPRV4yMT2sflg4S7qRT11rlRIKrWq1OeWoNmT/84NRQW++uUCCtC8XwqulOgdH2jB+Da
METlCUW64Rk8FHhA9dRXG8pE/waQPAJTos6wMQ89WDqAVx3/UP7lrh5T6r6jwIw5YtBGlijgE9Rt
gvGW9VqFpf3bB36461SZ/drcL/qRDZHeGd3Qt1/S33ctYb1dlvVmE1lhVS6H7HqXEkikvdV3pWpF
JSRXU+BS9AwcynWHKi8ei7LDaR9yuV6/efRJ94uGgclbn3gkFqbw/UDkPrvFtzVahOkUMJzCLlak
vmkjI4TBynNqH2f4v0rd5uzVGhycXDZRSsous6N8nUsOOU/62FR+CDIQYdOOSCMDhGvDuigJdXpS
N1e7DJ89mqEZAkN9JqLbU9gGNhrnFO2gRLgp9nnDdTsGvFFKfS9dFE0xB3UO0UCrMuj5pQJj0fbK
fpaRkDK7r0cyWMa0AabZi2LmsuvghvCXsSylvjB2cXUsvXe5Y3+4/MQ51Y2cvvIUCNaDeK2xjDhh
jiozaAdcanYJtRDLlspHyDkC6Vm2Vdcy39a3xGn1GPmVcnhsm7OH3Jqeymy6BOL6lV3YaUi95E/E
WLgnL/XTt/6999WkfZKDkdtLH9OzSYQjGlghFiVQtygeNrgdRKdwYG00MAJicPq54sMfKOhGvVo+
fVGc4XXNtuc8L+1JzR9O2lliOfcdF2HQKOjoBE13VIXv0xhhtJ2/4YMQPT6sE+iW2M8dDtSHEbzE
ya/4lf/yhCuqCTuQQwEGnSDQYLMM/BAj9A7xEdK2t12zkHPeX0xj3SNZslcnJSA1zsGxhhaBN1JQ
kDJhg8hj8WfieLvGgQqVi1yT7e7rkPtG3GdJ5iqJNygdU3esQ1GnZAC3kmYveB1yEXeu9QSCfBo9
agBlU6GgwET1PXkwolQ/szk93KRKD4hIqBEBfigLKT/MRayfYoWklqwbuj3vStsr0TzFb21xmhMN
ZM3+tEwvNFI8jEyqbS3fgjaUHkVaC1DcLfz9ylJLCAeztjvERBUzc8JQ4GhfsNizAwEZGJBtcL4g
ChXfQZFJwydrqfUSMuGwWf3are6/9InDJ+0vvPqtgKLF/BDPbrl13VFtR1DAET6Cn5GlpuYNyQwu
I3ArxoNv6kU1UTaOBakuggGJOWdiTbg1WBWuHFNUVzjhQYIiKIJRIMWAPNkez+EtISQzLWmxma03
RExOWaU5kx25Qeb8vb8uY7Hitv3kkH6NK907vqx9aRfR3gnb3dEgLBy8dFjtwKCmal3OtUgMc+QI
L4wLqDskVF4KqbkT0SbK7C2IqsyvikGPiWKU55vUtRWWAWsCbNgdKxEwqYX7F05yhGzjHS+DH7zy
XKDYSMvT52L+Zvy4LlM7FXvuo8Hsv79Gx6+OotC3DqCVS5eMqFL6sfjO4Xv40FINVqNuKpuvFv9b
kzO4P1m9+4tKiS81b4PcDA5YyuCPPtyO8SZJWoIUOtrrrW1C0tCfwbxj3mHW2JG2QsSuEKQXadCK
eM35GZI14ZXpzEht2Zw2rHvqy4/QKsEk+fGLlqpPX4KL7PDvsnm81geEAeHrIkl77qjlfSdgk34T
VsamOGniok4fBsddeM5rMa/pgumi5Cc38cQsInQlxiGdE3Rdz9eB8J+KJIdYiqNh1uQlMAYvqwIw
y67qaAeDgK4Mn4Xqp6e3uwsJDJQ/qXVwA8+G30pYiuiVOH54IrLW4RhEUuY0eFvn3FNuoygt7/xB
8JO8P7yXasGH2p9chZmLdYztjq6mADw0hi70xCr5ZtQiyaIKMC/HeD9M2mBIT6q65aQsW9i42PfM
Qg42YKsVYZ4iLwomvZ9OFzQHTyEsS7HR0AdUURv7JY/akAYoDv29R/JNA8R0AQWJ2ydJmf1cMlBr
fu14t4VQ9U7H4EupAWVhB5DKPR/W+1OwpyX8n1bEsYbZjGkDQiH4YxHf6P6t+lUn8YQAwyhWqhtb
8w4INlyPYQSIAQhjXGCz731+3ZeFTD+hFkX9mPIogN/P0QgNnxPc6h5n+KaFIBE1G038lNe51h//
biaAVPGBpDCu6w7wm7bBBBqCK4cZhCj60uh5ewkgPzO8pU7sbRXKggzPn2xYBc2eqsKRGkotkeX5
vXkVCv/RPFFa04S8AYvb+Mkr2N7VLb82ag226r5wKPDWdotMKBdXhLOxTOT0jXtgG9A5MQmuj/zX
Oy8IMGI8GslvQLyWWzgbO9gCKG+ePB5jCgT1AGFl6O0dJf/XwkfCg4z0PbGCvlzaHP8QXqA8w9tI
wS4SDiRl1itPq9YpX0eCGpJ9t3mwuS07s1QNrW+M6iWXRfAWgijqlU7t2A+j83o2myTYo9hiJTpm
rIE4jbQzDSLypAbbpEZBOGRWwQUy9H+ey3wlYcy1aWuqzzWJ03XxC8/e9z+ro96YaGcJbsg7dOc9
Cs/WaOtAgb8Jt+AsWHtC008V0RUjq785BpcshGT1zo2Hd0hqPH8oVyNFkd3zBWlA8a8K/lX7yIZS
+jQsA/GN/KVNPcZZTnbHjlz2LNxUTPr2sLu77A6Jt2VSu3quSHbNq4PG5+Due9z/gzAHBHlZrS8Y
g/xX9635HfAUgJLliJB5j6gf2bHsASMSKzoIdnflwdlbx8rjtE+PuLBiFsAZFd1O+VKRY+LdfBIW
hGghWta7Eo1JWlSDrT+fQ4bc1DHVMx0CnAbGRbcEoW/iVY/I4qmJBgZYmh6qjh2Km20zRG2CKwME
C48uHG/3sl3c8pTAY7kfeTyXu16d5YSvyYovzPy6y/NpQx0nF3PhBZMaR8KKpXbB1s2kdXegUqpj
OvGwByc8A3TlxyQezhn9K9P+L26eMPWY39aIg2xSzLHXepDVKgW9F4RXypTbeHNw2KEnEvwDh4e6
mVE/CnffIPNR6yLCkAF9vgymr+rsdYNKG6EeVQHLE5aMaBV30YqQpgfkO2q1jGELezU3OYuTrYgp
WDUcTdWboNTfNBnXYpYkhTMzK/BemhAyIPL3d2K/dihwCfSx8da5cJWiDeRMSvSpCqV9zkBLznRA
/wZvDsH1g+OvrlOT/5EZhbsWnPUDlhrdiP5jpgOUqRwfZYXl/vodpJPuzy/ay9GSMeoZp6ywwb+N
YCILqCl52vwi2fXa7Yr7cSPOkP5R1GGxKYgNLS/H5FFScXCaFDcHxAjvs2II+4NGc18YKp3azfp3
T66laF45fj7Nbp92l9+G8yVBJb+qgl9V4PsK/WObpESU6OUjrnUfXWiG2eCKr8zbMKmFU/r/0uGd
/cNKeZBH1XbIRtkdExmiVQ5FVQcLzWzUPNvP/p5bFLDrH62kKn5lIgpIOiOSBjAI7okeiwTA1Wwt
OyksuyIpYFZDxxv3YW7NOrcGolQAl1T8MMUd/pNlZSYOBE+bagaMGF4R+pxueiR3he++6ATXMWN4
DGbB1fHhAJLI+Yh9KO68f+kSIIgZizdkqNFBrXq2JZP14MVLhfuEPqevFW5XPYNnzEivdP92Gchl
PQNoZXqMLX6fowHXmYR7AHcTgNbOE2XdEkkIx9yLYCWhnuJ7VXLoHovEmhOLtjHfTZDrMdM3kKXh
bhiH8PcshMIC4OYUO/4zrGCV4FrflGkZIfjLx3h9TNONZpXh3F7I6SSiwRP1LyxdaLx4Q9/bxXiV
n/ZLRW6PHteESkcPlwYJPzormt9vlREfdDHQvJUvfq+gS0lDGEcahidg0RKiwU0+DCsJrGorbvLz
tI9kdiIyC/Ymyc5sj3nN0elefs97PyO9C9b4cWTZFnbJJuFSnQTbganjopcaPA5xMwyH1fPVyigi
9mfCTGbMKIODlsPxdYtSuBis80KXOj+9LjLHE3VcLKi+3JOrgscpRLNG+IgVCMXO008glkWKbIdf
kzq1CwxByzS1ij9YgHZ4Nqi7NwFW2ECa39PF1dT1cyxQ4cFuYOOt6+L5BQgx4UmgCqAYOGtXr+oW
JzaTPTuqaITGJAb5Slx49DKRieGBUqEjejb4XeAxxptKDgGlh9+zeZDM4o9DcBc9yi5Yw/CM2slH
2Yw6lDP54oaRQKhYqbxJxXkdCKaZe/Ck3xVqx8nme7nH6f0n/D2yNu8fI1lY4x+rvr1dKupHMn9x
61QYC+utbz9e37Ly4oHPFLceh/L2wMMTK4W2/2OntS73TZ6fIGOqjGPScDlT7JJZDjkTr3k0TQqC
1QEo4wT04AToTROwV+eC9LKtHS3VkQC+/7K0mkoc/ZGXJfvbVo460EwfvgL+ekIyZec+PQ39J55A
0KOTXOEDJUkdUin83wGsCrNX1IWsPPquOvtpWfqrYeggLoxfhQUZJ3/S6we/DGmEruK79VdLJLIK
qbVeEJ257JvjQiwyXbmHimSLf5guAaKuj266TJsyOttR6F0vXBEac7lg3RG3JGT8qDRIc1ZR5syR
bAgQUASoT2LyGcmVozNh6jwUYREkf3RsJN2Ba3GLR5nazPrGrZOxjmVESJuCIOWuCfOH874/oDsM
arHQtGFa5vcntDrxg9q7KL/adBsbbakM+moMtqHha5pS+4+4+igaJyfB3VqvBnEaFt6PbRkArRaA
q5QuMl0sXcAYAsLv9F82DLUetdZ58Y7X4urePelbfDVhmWvWk7/g1AvNLkwI2VNf1QdjrPJkRTht
+stYcVifez7FCU6WmHn3ttAdvmmBI5TP1AVsTP+IwJ1Js2bb5f8WpauH5cGa6wsY6z2tQnrchhkz
qMbxOFOLxf4bdfGPSIkx6VIFXE2YlQpS0Y/LTDxiPRg6xSNAOj1VGuEmek0TfEzPYqqQSL80mnq/
v9YKsKE+6FMk8ROc5B1ol3wezcscFXqC9V1S9zYZMVBggqYRBeuyAlq2ocSwLTY7gNkUlCBlUJeO
YsaKLja4xov5D6AGizxpDkzWIlmUO/uXYBwG4z9mtyN0J9vGLsFwlG1LGgxNW07nDvJI31vd+JE9
xF/Lloe+FyrZ1Y4Add8/cEvKpIq0Q1ryYeTHv+x5MQSCxTMRi5Y1Ow5crYKBZbzrckAWQVWM434l
tFac0t3m0rHdj4iqhT2y323NWAwqIGiLQ4gvg8lUtrN07qHQUV4I1fU1KL1SoraaTWTOVwcTbnZH
qlUyIsofr6nqyBgA2o+gHNI1W94EJEPo8RkyoodvLOn969DuX6C3LTtQFe2+D7C4il/mknj9Baib
0XdJE9FSt2rityfJbVgCS/8WkCQ03OOPvRrI8fVCoYynOxSJStMBfoYHRwxdxyRp9L6h2n74IRrp
RtdaGcQpuWbOxH8C6XKRaR/yu9HJyqONYRntVvgkXpRDleaw+ZwUhT018cXe4Urnc8PmWKSCwawM
nL9IbzDbmg/IDkGLG0v8oZZnFS87z2E5eHZ842rPYTE4uGoZFYSG6CySN2pBe2avmJIirkmo5+bK
4rDoB6TWeBG7rI3jRPPWvAbsSFdlfVP8ntpcVXWUMOdMmyGA17KFM6DNhxBsuFwegZ0pxr5lV7oL
LOAJwCIalGIjX7A7uFpgAISQGm9MKV4V2y4WZWmJFDnCbH9dJuybeywxwmlxNFwdmzeNWqtCCv4d
29SwI0rAZeCpjudbRZp5BXPYg9hPDKiDV7diWtd0Yhrut9cc4wlffuePSj8eexywL5Hy2a7W2vgZ
6zG9CrQXVQhEqRr4WGqgIncIeyLIzkBH1bf9jS4W6TRuNorBsD5yoNeSdklDTDNDNw6kBlY/MsVN
haugUd//ffkFiyJWBMVXK+HkdDxZoCX3NLcILMzcvrGTXFRkBIPxcbfdEhzvVouJTrkNq6jg3QbS
vWYNeMAnwYnKkyJgQNCiOzTGIBsKbLn2Vsz97tUf9VNapMXv7A9Y6bkXaf8nUjOobs6DtJxTxM+k
LJYHP3CylRLlyuX+EDCjKewECywz4ziniPmb/mjB/0kVSblMY/khk7xgf1mPsr4eZY1k4jN674v5
oTLfaOSf8t9HInmLdhLBfllv5asXw3Mw9PzgCBc166aRY4mQHrK9t7JKdIkuaAwoNViPvkeQ8Sql
zbFUKaa/0X6sIrtf/Clfj8D9vBp/ROECRbn0CEfI6WtQy2x5meDWRVvYtz8XxnTKbJ8fgnCAquDf
/bz+8wgSOT1NB1m9L9lzd7EwweQG29GZo6ikpQfSVqisFY+MyD4iVmboqgrbweGNON3y/twXZs5R
gYcJdyRIzwh5/EumIHV4VgEpiK7kPXKwbqLguLSzLiSCIyavIToMy2QVXPO0DdcuGGTHFvKDm6E7
yn/WXuQYrAFS4dA3mbrkmmB+7veITELHfSFV6sQaNWDZEaQQ8CNaHpZk6Wr5NNDrsceRKk2auqgy
R1iAXYg96mkMUkmkwuzC4zBDPbMZLg6MrbnEfbz/ky7sl5aL86NwFMJzV4Aidpsdvb8suBrxUWCU
qveUt6yheZDKLnpyFpFkSMd7bFmPUqXzfjPUuvqwmhlTiOmyTV+ful6Cr2bU6Tq3Yp5mZGBmZLug
WC9/6F8STXJrF7jnMKI9QPOi1hlKQ4vcVvmeDoU5ci01Yq5/FWCsMhrxEfDEy4D0lKKDoAnDSDi3
OvKyzKxhJit4/24uMNBdPt7EhgIULVn27Rgnphws0BlaXHpV1hZR0EILLIkDm8n8R8LDKCHPlCCS
afAqjkxTl7+AJAkYJpb3dEmp3tpr1R8SN2Xe47ylr5f96AwiZBFDVbRfMsvSfMudqNwZaP37Awcc
j9GceBuzmTiNYUjE58U1N6X4Gxn+vbo37Ma5CnFHJaP0HGTxyRJCP9GKEDZyu6qzxRyUxmTJ/pK/
22iZoK3PWGTJPoM7IJvozm4WTIyIPzD7hL2J/bv2u/bH9SMJHC+lp0eAFDbI3qUuO20ZnhbFefdo
i9i7/KP9c//AGygzszUnYM7B6QOxp8eTIMeuw/1KGaY/FnUf9Yw/EaBvHF1HDATyCKMjKjtZlMah
ts6hS823vHm8ehZ6EAJiXFGo1dnOxeX1ItcZzpTLLL6mjRMOISci5/vGrkIsGRrv9N8DPjR/D8oB
gqVB0wk/FQdJ/nvcUcsY6F0aFC38jJTxTJJfpS9j9ataH2F4i2RpHBydBOnxpKZjLo67Ofu0G6dk
f0q0H3LpQApEw3jTH6pcWpveaYIOuCEBH3pq53uiwhGuYW2FYDcjamPaW99To5Iqlh+LBjdyb6L5
lKS3DL5wSduEZpj9vs70KV+ofwm4+gJDkOKqdqQSx/cRAyeWmmw7qrnowMrlAXFioKHUFnNJjkF6
H9cjh1fVdKsh4uZYfYU5dqUjQhdSHbOAonb6JsODvzBFiy1bmEdGBKOPQuXHVCYYn+KuiKl7Gnro
aZaQzPw/4OltMArR19ue2yAAWaukaEerGaDntp8hm2WkVo6uF0psBYpH1bKN8iI8XvgRtRZsuwJJ
RfdVPxg9oxgC48pMAn0KAPjNpu2qRHsfSPmmyxLpUGKL2YHWSbJhsJFTDij5km6xbCbbuOVSqfbG
yGQaQPCSflwBj3nA5BE9SJOTqziFG3wP+2bKp9eZ2TyRq0/9AHa9vb69Rb+8ZghH+rVp+/s2E3pn
9hHq9Li3IQHkTUCmC0zDGgfJDcxy/3jHR3YrmqIokCibkdYWn4zhg+ocO/erN5D/Bh1uqp6fnfBX
VbLBcJ/JDkyylLgbMWXrRGKOFXD0eTIYtky45CiapzQc97eX7AEY4uzR490NkNLU8EtjZZZPV8LY
dFVf2Q4yAEmKRIGj+XD23Dpb0IlDwHNCy5JuuzXZY0SRJ9qGwOM2qdiXBx/HKY2wbV43U0pGNki/
tVfqdG9O91kQdFS6vJa9GUL+QVj0Ba77X46HhWuLzqKHv6GxdA46S7CvJ9WSx8yYOvv/c3LARCw+
E4miD4wQiAfgBWINICDlkFI/Ty8zY2yH2d+XdqJvPziHZWzChnggkHjw4qPjpS/hAZN2MXpvCzKG
TqYFQdlUbsjYr1/czc/AA06bKp2vq2aXP/eCn1qprv+tDiCGS4ecP44IR3JW8Bcs6jm+M/kjh2kx
1RQPRLTRMuAbWVUA8ZOCKnIDkAMcF4IPYKMSYsUHKqVhPAp5tdQgIDMNuVaNo9KCpHtm8MVso4zR
Lc+AqUenDp0VpsMxzBOOBkOA1SM7cYnryVIE6icws8QmuMJOXn2OFmbalbti6RBRx377TTy4uhgI
acHmoNPzHjycC0GZz3uy1ce7BCMXeKOc8tUOROZQ+48PU0meLRll6RwLR0tNWEKN9B1SchNhP7b5
+d/vvueHySUSNiFuUjahCRZCYpWDlCKCdu3pmblZsG0Ox4HLdvpxp0z9UtQjmqUbf2vROBMDB421
gNxfmFb4AFePeLNzrp4rn+/xkHDpboctCBnXlv3sa1ZC03Mnf7+mMCTrSJKbXsPxoXvaUMxFxqLj
elfBqSpqVUnFVqyltp2lATG9PlkP7g9WV5IW8ZtiaCZaPhepxMickazifYvkvicTsoGymGU9hmBh
5/QkcyIlDpL1LkyQJxcMzp4dXefbpgFLSpiO8JY21KpVieMSoZmTxgYxUIWlv/q7UakkpHamP9bk
54+sdm+7PyIS6Mc1gPuQ8ISaBap0g1/M+WbKux6PFv+zBV0LTnio1JJuQ8I5OD+RKTp8o2fCBSpJ
IPR9jCFF1Coo0GtqG4OkwPXj9PX/GgOsTH+rV1jdUfW6GrW/AKePmMfqZNQ6+ZUAeYBElAkNK7FN
Z4Wv0T1RHgJtjgzRYg6oz8pJBAfQYtslaAT4QrUVKSi20WWFoiC9N8CsV9+Mj6ZmwtpkvJB+oarO
35h9XDiaqU4SQ2FOrFIhyvx0usaY2ZTpcn9MEA8KSGDyK+Hnu1FC751ufY4W3QE6JycboN723EKu
4/hf3L/tTB2lf9gwYHeZTOy9i7rpH46SSd+wnu59WQ5MFrKr4GmYuzcMG8nmASR2801aGPYjy32S
K9SIQuGoaO4otgoQrD2dxveFWxIrPpTXrHRcVXIIgoGcfED/mR5QDsPknWQ2AcgVV6ayqMsBSSH+
nHTlmS5kIxdgCidDr7Rd/lEnnuNWG8hqaUWQI2Gv1yCAUphzFqQ1EYvofVUNTXLM2hukOJku7Lvu
QVNQz+uSy5Gl/FRcTiOtNAa550C7qUO9e70BO6GyiJ4OhMaXtX2B7ueclJPNppU7P2fY2S9kgpS3
JRcFhv2686Cywu0ezAbyX29HUyikucggpkbS53oBjQXyrEtWZMcE52C0ehzQXURTJO9C4Z1yUeei
hSxJio37otwCwT8+S5gZ/YA6UkVbuzV84mj8xCggE0Pj1A7ahdpyTHJubbJQ0c5VUD7q3S4sZwfR
ffEC8iI20AG/Ix/dDosZQmNxw1w0kulcFQAN0yBZXTODF3jSg8kkZeDqhfW88A3IJyGadnjXNeAJ
Ti2N1qkZDMBUpelLnTKYFk7CXbr/4eK+j1uVLNHoZshsjfGqHHD0dro03x4Dtb99pQGDfmWTuzOb
7jiNT9SIk6uh5ZayER3uY03LxBKMXP8JektOmXCZxZfZZ+ETlz4M5K61c6TG0NI74kDXmv1UHrEv
bzZZzeU1G2szlbmwsKvNVW89KHC5NkWLMQ4OMnBIyRch3CWWY5kGVeZGicNiPQwXlnyHKwnNwtlt
dl5Ux87e40fTbNcKiqEN917BRAvG8AkmkQ+QOpPR3K3cRGS9ScbOad4uPK90PJx+xXfTAUBTSNVg
hrX+GbPY/9dWsIZ/NJHkWrxJL5q2n6woA4gcsv1ujnSJ5VgP9/K1w6SrmOSdNyG+At9LHzkVO9dB
veFNYjVnVimjtrDLSeTtHnA61K5OtmTBngHsTQaqKj5hwafLzR4kzm3mYhpQX/y7GI2J3nd7Aidu
oSXl9sC4rxw0+yQS82XJRQBX/zF5Pwpi2ln6vl82UdNRG7TWnU51j1EdtIM4lFPQ0W5YuG2h9xQU
72wtmnWBkp6z4n9QNGbAtz5wk5D77tsQjDSXM9T3P+wy5TWRiRuq4oVnpEImGtUOqK21g7alY6G2
gVsPJWPA5JL05CIAPvwzs5J3T/s0o2pPtCI0xatvUBcAtOBVStp7cio+IY68ZD0jPVRofkWoHicO
qoOl151xouFwtoqu20u+xrgWoOA3VvytB1ZlMOS/RhbbhTaT62mKes6+0Y2OxghXMOz4dOoC2hzy
r66M39Ejidp9Uf19oNm3rGTrXF1mfT6QeDBHzk/Tl8CZeKz3sk/Cq6LpKCP8iAt+6x+ujgjDVPq7
UsXP8ivm+tSdwVEWVxzG5vluXyUW5Tuu64aUJG7AbPFxORESBdAhvEmHrLjej4S8uozCEMCsAkF0
80jBvEBIW2hShDUfV2BZY7VzWjqsAReVuYwGk/io6LOJu2h3I2fxhYjsQYuuPbvKZnVBSg+ckwbz
9FA4+f0hTUEoInkWWV8B/4HHgAuUr41aA9sVyib39o7+aCde/unZUsgQvVXnjq7MJkzyPUXSFEVe
XXQ2zPlJFYCfVb4GQtBydBeBNDkWENHy50JfKgrc0LoRKl6VYhGi2jgBIsKga0Fo+53SJBXWJku3
VMtUTwcYOUPw3mzUt0snHB1WR5jSl40PWcPJVxZvrNXYFHPjUBQABhJOk7r5LFxM5CWEulmYhQ2q
yTwmnXqC4YhihsQpvaZRAcipg8Tg5ziyaxwCo2sS3z4w6k2Lk970x9Co+IG79qeQUJlO41MD0t7Q
YagUaZjHKDz6wHJSgWyKxRMrRJhfCfdiTIKEaJHB0eG3fkY5q3G833S+MJFQ9S9gG+oFNkYIbg+z
8DwZRfmZin5fhnnWUN23b5Xyw8xGrmiSIbdsuBB5xxpJtVS2Z7BF7WO52zdud2dr17cbFp32NNY0
SBeWQnAcNshiBrUUPcIXx1LUybvI/TpNYeWOcG6vFZy3g6UwkHC6x/htA4Fz1KEdfFbQZsw/UlVk
xnNXXj0QeQIdWsm1wPQV6rk3dd4cNmOLZE4Esp9VMEDqAXcmkdMaBOW9Xa04pb5ptv+9vdIxs5H1
iGX60WY/ZJLX2AG+W0FutV42FmTeanbYrHiYXkpvcYbsr8JtJrvsQeIdXcFbtWrHfnLxD7wnxJib
lbaIkVs5cVjjCn75mL0PsQLGPvRxaKGcO28Sw1xB5xYwHUPfKY6TODCAjTcts9wvUq3Jj+7Y+Mdl
LDRE2TnTVQLRKIdaTbBJ8/O5vu75Ud6JEhVpY3PSWE6tNxagXPwF3RvNwz213I84I4rwr5QdF4J8
lQ3sBmP/ICZ+ujoog2e56OiG7xeFprII3iCcscqrm+zGtnX3rUZCTR9/TE756gIUaoZuoMXbHxFO
pi+M+yU5/sk1TR9BRAQT2SQOsNfUP3PzRVw7WM6pUNkmd4/Ch0RAW0fDUzL6VfuS9BnlJIBJJ7Ay
+/JTV4JZ/sIDOfl21K6DbD8VdjRdl9pVAfzsc9MX8og2RnBi19EEeCjQShssC2aZbp9YOJQ0chnT
7PGDy3Ij/JfiXJ3iTkO9+VmkNldy1KXo+2Y1BzWfXXChavkoTHr3IwkwIUeJhgbPXZL5JXPhwy1E
z//AVBal5r7NLWuQTLkGaQcj3Mhc1kXn8LCjvdIvfMS06Byh0JRq0gD5QqffI7fuNhnQwUumm6ib
DWak9iU3lNl17ElqAyglOjP9smkZZWT7KoDS8TCVicqXNFpWnCX7B6fEOhq7hE2DeiF/RKJizjX7
7Uf4z1OjOYPkusKaXlHHBfEH5QjH5xwYDPjLLMUqdglgLV0Xa7lyNircpHddaZauw3jjYhYmvGlz
Bx8qOw1uI3cNplrkZZqCxRzFojUVsze7OWS4P6NHAgE0c3AacHScfnGJkzoz4H5BxFymb3/4onSL
383+53DqclRh0CWUHAv/yi3XLMiHvmI/Hwh3EJww7ZuLPDPXbE9JQ6VxDqqDYuepJPFY5sgKV/ij
6mW1AWg761T5lSLkRyYNaEGqC0fKB7yIf2+2qPv5/4USPrGb3KoUvZTFaY4b1Lq+78ZkNatzIKmm
cLDu4GSc/L2ociR1FToN6sZ83hxLZXc3amvaMiVeWdE8QEbfAQa5SSM2AJiCFX4ABgANRenuYdei
kuxHqWlmMTmm3/bSfK+gf3/+rYZD/ymTcKzS5o7Zwgqy/paoFefOdrb/Yu51ft1uOLP9eddC3pVw
w5WPaL0ewHCyISt8N5da7S7NIaEHj7vACbEAWrCZTfvVgUYiY4eY3wcI93J3ug5+qlc9C4GeByXv
+aUn7gxTRq7xVL8vW5UXw4nrwpTnTq9EqiKQKJBht3vn/76U/FhN0kbHxrv0rIp1Zw0tnjM7VNlN
i57sphkMicZW1AZzUrhf7WDDvrAt/wy+8rqwu5Sh7fsip/P3MDQUvfUz/oBEHnSa9ZCUOpjluCQ0
frQ60JnnD6DW4Y0ql9liTIeUPb/jVI1UEeHFCyapBP1v9k0HCkv9xDg+9TnBrwoSNYACzXlieUff
KC5KRepEutY6FOF4egplDTyM1yv/PJePyj5DQ2qLfv3oC2dtQtUyqE87Y2EId77CsLIjc/2CN1Pd
cmY+7JILJ5d1mv8n5ytalve2vC9Ks2pfLmUOYcHrwB6otYBtNeUwy/H0QCJYFxOSCiW3Rrvc8hDR
UVG5OlU8OIdFgvzpvBkAYQo7ZPelk6o+zbsXCR6NkKSdILf1qBw0itqBDDslhGcgQ5PqXISN7EwY
2nQxHTJXHzw7gne26e8VEYB/jG+t3u0W14VfKpbSTN+PjnPMXH/VFKMtpC0bUBOAQXqItlf0GsY5
D9V5qesQ2n0tQgoeZXdjcoOUMQCXeYzVIa6/fUxtCaMDaLR4EFneC4/3vArWCYW3GnUfUcLhxGch
xeopxZwEGLBfv9v09Nsa7SlvrBQij8vQF3qDN+pDhjRZYAuTjdkznCKF1zeTr4xcFCm8rnt9hK0x
pT0IfJk04O77I5JMh0qhfPrTGv+GLZ0kyKtmawl/Ka1GiM8K9tK+PUiFAdOeWWdsh+lgRlUMVCVN
qSxhMZrEmUZfSpMfZHHNV2xePfr6jWYMTF9e25rpaCXXn089B6K+PRcAnMJbWkbHN/DRfJOiCj9Q
jn7jmCEB8wWM2dG552ucCw95m19OVk3NWTVkaNRJJk4OBWUY6t2JSmAnRwIqEBIlQS0gK9BWptk4
Q2HY/2h97OcaxUfAyX9195fGtTKUvwiiAVLfxIHcinLBov4A38wANvXCS4WVvuseM9M8Akri6n/t
bXrs4YDxgtmfb5ONz5fNu8VEFfXJ5zfkB2x7ZHzH4sLGFiFYujbBL1q5vx0w4bQNDgm+A5hD3fe+
IC2b/prMPtt3fjAZE9ZSqPXqKGUpuUB9nrzswDTY+mMcVWSOPqrESbVFm5jaRXda3gHt1P34VOIa
Ob0Wm0ZDxucGWTAr7pLzWaWYHrv6HfTME+KOB8qN5GFx5DFrCzMJdxs7s71Zt7Wb1awgLQ0QkGwm
J7fEJmUrEVHhbAArxJJgkY7H9cvc6oZkyh0e9rSN3Ylj4gxMINoT6IGq1ksFdKWN80oLeGIh5hDi
J7JaJ/NZPj1Diq8C6UbDaS5ziC5NUBrvjz1JnJPL48nnurmjG/I3YIP5U9ZHccyS2xkkd5XUGy0L
NboRIOP9RR9eeoQ4p2A5KBEBGmLrAL/f+X+Wb7LhDPYsY7Cs9Ariig3uP7Grt/YdpXOZa3LqDSht
gNzUrfMn73OaA1CPRYWmYwKYEhqIBaKgV6ZV23/4L7lI6SccgJGHMGX4ifQ+6qzgbvqYMo2cS4hC
tmpLBHYcy1VTfSmcU2Xsl0EJrUBljV7E/Ue5F2sja1toX5VLMEXSjV1zd5v+qQCHjhwCU2hhe3TU
abIQ+MuinnBmWI1vp3/ulGiGYQtkCTgHIzmmEGIb5elyBQ5NmekMYZ7E4lsGK9arJLdWi6eZKV9+
laZvWFp84YAiKAGnslZkUSSqHNPULzNBvMc9dvWxr+g0YE+7CjQ1y5ZmFyFB8PFBKE/HghV0e5Q9
wlODLrE/YOYs7y1Oss7UT7m9zwg8m1X1qIveIKpD574FT2hh0QcP5UPHuc3N8ZZR3mE2rTMfTwz0
xc7gwpyeFjnATZZp3IOB5cozDG+UutEKeYzFwGu6nAL87UI70aS2T+7HIx9gjGnX75IyvumJTEyV
oQ8tF4yhA7bVi7M1FVBzcWOdgsoky/UL7XFCtnF0X8Xc+jN5kxBeWYShjeOS1VIHtwY0VRzaIC3+
ujfVkkKcQpkAT2SQXn+lM9ixZTdQNJq9PdSHR034hbngDwBBPZ+WOGHwmuPOUa6xop3/flIceL0i
pDDSGSMUFNm6/168RUwX+gav+G8+IJOx0xHr95ApHETJHNE7PkA6fWnrGyn8v2V5GpTO9bCR2sWd
56qujAsel6GW1JKmb9/kiHYvo+veTUrGBnxk1D+63BPFdJ/13Q4LLx86Rfj63xUdh/BUYiDbeWiq
SytDbNd8DyeVADkxKrJS5QSjg3L1ILv4VvbusHNcaw4QOcgHPmFTkTx06UZ2uKzyZnx2t3xUHfQm
zScjk61wygB5DMyLb+jDKjvs19zPsjWC50Mxo4C05hQ9Z5Co1ecxx5anhSPtSNP7ngQEPk5z0Kli
qgb/HGeS3s6oOOM+PDMe1PAPuMoaJYyhNr8xzaFJRoI3L7uAvRL3AJPOoYXhn1rn33mcKBEMkP7A
XXsurv0TXTpkOs4nTJVDpdVeekz26wXGJwWgkuko6R0h0DG/f61n3FujHHAHG6wMKcrHvmlcUDJT
N6bkd05ra1J98ZaoSMr4j9Uc1jnbmVZnpmO6L4HKKGiCwwpBarO7cmoLbKZUlxGF1fQOgN2ePnoi
yL7smuVjR5QQhUzENgBG2ME0poo9Xkc4gLNdIhbF/3tCOfHa3OElA7c17gwcHbodKdVT5hrfWyKr
tSQugcw4Is76nkW6If0PpvQtRxl6nYKnLHcL68XItdNQM0t3qxVXK4FKMO13QhXB+S3uauKpWUI9
7pFiaDXAkakUV8s5G3f/X5/NeI8pB7w4k8bG7cJG3BTy1hrT3kbt2tnsfBEDquDGP4NNLj2XbibX
PjMux8xcwJSiqMKiLPUtqFq56WeJ96huGKl8lBoXUxHTzI4hECdFB1lCR85eBdTx4GtXe71ypq8p
OlnGgywSzc7f5HOTUK/v2fMDF3XXImeyNLt61LyndGxk9ZTxfQCscPNLDxO28LHIZ1nzvZzOWFhr
nLmWo0HZKc9XS46oHQ5lqMMl4GCF+OqSa7U+LIU8/2E77zvAY0yGt9MIL7007lkf/GRTvoBukzT/
KwcigAbmXc7iHEas9Rr0iLEI8c9zpJgy5iQ2NkwS/eMVQsVLb+kRi6/TrRk4iZGpmEiIoA4cnbSl
brxtK/vDI+G6I+yUaSISiEVwsBgPjSOqCgff6ZGvdIbNX6OIcEIODXYmSSSbYlgR0pNie3JYWCEl
UGi2odeBYPKYGnT/UOUJQwyK8oN38oVRUseyOUaERjkqF/pgmRpGBeHcCWzIyZRJ0wXQRDuIjj0M
rQ1tWc2a8QEaFxMox+SoW8i+f/hDxmNrckFdTaqZgnjAT51ImvmDstsV7obgLSh+V8IZCsHoxoZH
TObA8uCGfKw/F9rClzcyTeTMcV0+W2g7p/petpTWrQnQcHEpANuMeLRgbUG5tENyrazR5cEr1cxV
3x0JyC1wrui87CZa8uKL4nIHo7sWa43bWqfZP6pz7/s+BXowvWoCc0PuT5IdBA25TnaqHGP0JSU1
V3s+ISxxe/v6bIWe1akV3IX0X57zdCcJI3Y7jSsAMw9EIkEfBo2+H3Z8tkxMbvqsKFzjiYWxTYmE
zEFiGE8U30L9mdaT3A3zw8rvwGHyP5l7DUjxVsfCsqm2Ns+beIqrQHT87CN5AMl4PHW0QcbH0QCP
hFVwdUx6ArurvYyUOHH/HCyjRJhkysCz/SWFIcY3b2H87qUvkgZTDImjTtq0znlEe8PSckmUOwXG
j1D1kieZ2kgt48fROyFMdStJz7YSIiWq04my03tbWOzsEV7YgpxCpQB36ZvbiSTnHTU21GnDVnHz
5EdvGoK6VDe+qkY4iRb5axdC3tv84fo5k9xsE/KPQv8+GX01gCp301FfuL0NM7y/XDZ6nfvMw2uK
8XYs+4kX+stOs8Hg/oAspudpeN/XdlEyVXzBN4bziSda/zV3pgZODTg4SLgoi2E0SKAwGnXkfWYb
6O1GDZ/MqsCXLOeO/yTQ058lC05UXH7Mtwndj9Q/0okB7Jl/SHf39x6yT4fLZT2mPcKvpPSnmmpn
T++cRPdPttGjuCl9P5oXodyvtOROQJseeCLZvI2WdkRU0afADH+sry/4wNWHkg3bi1u0TMxfw0ec
XYOqZmIiicdqZUtFloD2QmAfocJmF+27/QQWIWGYvYCir8xV4Du44VXWpBovTEX7DCmulM7kCaSE
ChDBHCyy/T+AeJeG3cekPCHwCo3wQXrACHEy0S3mdIJm2pvE6bgAk2BgWtcifHbQ4Nn9Hi3GW7ES
viAQ+3qempJ4v6gR0w5h8urS7xbGJmeaQzRI2Tr15/efXwGs/ElnyZreQ5BKHbQIfcsrB7MEOIml
UW0pj8bQB86kDWHBdJw3QrtXyx1J6fvsEQhlyFsmiqlwMY8ZcdcFWjN/HeVheTwf2OvfeRWr4ivW
U0L34IyrVvrq/kWH6In/qaU/c4qSWxC7qDh0rv7pQ+hDKxgu99asvx0b+fBkrgXbLcdsFSc8Xstp
tPblUffaq4//mAi3kmy2kazw9VtHtiKV0jkk1/KFXzTpnPRQXGwiRED+3FlHChBCN2EDJXkLyB1D
QzcUqGOuCXwojaKqGHByXJihfgJHTUeAvw7bzpYvJ+hSzLyKD2NOCkVolRYRpI8gMPAQMO81Qjhw
W1+neZ7SSZmGgyJQYdi3lGYnuZ4H3KUqcbQRibT+S4JRW15azqBKKvrz39Bzcn1orpGODVmTjPBZ
IOGyRFyAKR/BvPpnCeHSSeUTor/xrDZRCO+A39vkHJMpoziFNNb2l9Gxv/PfTnIULr8i07ORXI4E
MWzSOYKdovkzZ+hUEjN8Ys+2Ds+aO3pqfEr4pjZRPN6goYTyPl5QOlUP8wUd71vtvQ+nSb105hWo
rzDiQukV8lNM6bRo4j4XtKzubFIB1CDzl44ADBk0AsabaBkEl4UMcJ9w8FgbT9QcyZOieqJQ3Xy0
nfrNIFNJOf1XByy0PHqVjmYjjcG6mEDNMVooN/IcJvAPHxJL7kcqSENNv3o8FzrXjQhgH1xQgqXe
AdkQhd8GsBCA6ElWu3F2mX8F4rrN3xk84TTiiOF0oKZjbpUdo/lPJx/EaaQVic62P02/FvLBkE6y
pBc4uLKJSYY/OtK9uRxyURTZhu470r2EUuYLU7JVc5/AyHlzahEP23ieHZSBx38uNXZklvOgASeS
zW2DVHg+83uK+Kuv7dTJM1Z9VqtnMyj+8Mu1+w+qTFYgZ0AQOZMiKfBDiGqgaoAbsZPBAqmDlTPK
rlRAwW13WU0Z4B8rs4qbRomNGSORDTA8jPE9MYmlQ12zVAmG5xy1otcLvzB0V4Rk2MPBMZLPcEE7
SrrT8mo3JXh8144M0H2+qptNajOCC84E/xTuKzRl5SoeOCy4Uk8+PpBMkTgpVuZy7rJGi8GC2/ym
i6k96IRDzKEyuYolqxulnKxid9KVo4vsuVJ+QEVl8WVsHBl9+Y/+qRtg0cj5o4UrXhMj8l388jwg
ppp0BhGVv2h2WJOc7Lsmi7QG27Kq7jQmpZ0stPFau9+ruq02ik82oukZsutpmE3o7MGeOA+dulDT
laQ3gpX+oubUBAqxP53X7iy+/jFkLGOwhxXWXFnqaZLSwcbwFbe42r+vSRSxs35buLvEuwwtC3dU
Ep4O8pEB458eagp1s5L/rkILzUVGDno994ioHycKQGPSW/JBxLCOHY5EhUQDixeScSMpa5H6nqVb
Qe7vnwYS3UK2BM8+j9oScJx+GoYRKLKHT/YZNnAwyvRa2UjgZc+8TNxornhIUzfqBAzFzVlJqVox
VqkLJIAFUfO5B0U2xgayvA8bqxnXptGO2IyhY7LhzmkIFkeppKKL5Fjo42mQQSu0mZ16joRQVcYP
VEe/wRYe9yA2etDsGp/JRpBJqnXAMiuIigL9e+pNuq2ojRzLF14hnyn13UV76aSGb5CqF8g9IIhg
sYYYt2FwgUeaCSWX7WOMXj6WZw+fqpj5oe4Tu4vMaHrW9Tlzz/i2Eb/gmNtbTFcGv5pSrsXXFtSc
cLxYXQOIypIgH7/mewMtx+kkZR/Vcb+g17sFJ295/KrhrIMtJYBz4EKell8POZVI/9Aa0MzLKX+6
c7PiFnRPQh0wKzLIFTno/nbzPvs1orszX+GGrrp2UzNlM4bJNU6QiN0O2eDJHBZK2uhjDKlrCPFP
hRjoy5ZKVeG73fNeDWbjljulmAetwyiWTBz2dNbLXSFccoSXYS95HzPdpbLC5R952qDHqGbY/9Bx
PyPsn2JAL0WxNmhN8d5la6eAHzh3XUAKN3NMjKeeBwFs4jwbpGmTG3llK0E6xUX2t6eOyV+W9jiY
tSmm+ezhO/PFe/qsLQnHkoccjkXcWTdxVqkcFCLaDEfqlo8wIg6aqoUkXI9luBwI5XpIWVeONx05
5vtLOrUu9oBYvXaEYFJ7z7lqEU7eWfj3xuwp7c/2ohhr3IYJ6UvRsSwRZ3zjOS8TgZsv6Gq5x0K5
0+eZaUluSeiDNzVQuFxYVbRyKNf7+xj3OSkgfWG+royykKVHb+feZ9wBh3EJGwiM9CJLCoy7q/CN
UdRYrARiJQ4SQAYOurFru2jOC3isBfXMQKGLqbA+XGjl7vzPimfB8REtVXeHzpSXDPKH3dZL3XnD
1U1JTgvxnX3Xget5Da910GqpiavRc0kktwXbKKCrXstn1ZKKtmig0HoPFKQI27JRQHWUoQNjS9aQ
V6fyMfk+O8LUzpTWD3jVeyd3NZPU3lB3Q2Olw1nXm37ERFrhLoSt20ISq1oOjwof9FosDUGleFRl
ZmB0mtIZOY7Fktl2Fdnpm/Mwu57TdtFrevbp1Z15zNK7DVVFE3/J1Egn0Z4RX5lOOR3GE9L4iTrm
jfuj655+VX4FQdQhzA5shIlWBUsdb5GR+aGNxRgtzXCJXaLw8XGNRLrcBJOe4cYqJe1LAeAqMnKh
TucMC/Jxo05zouR5US58uxttyzNlX0mN0Bsoc0jtQzbaHNUJxDsUjDkaX8G8OfRpHgb/uKt9kbHg
uIOqGJoPp+Id9TwYvQToS83GaNyxQZjGW/k1CeR3nenCQbt/M4Zf011PxcGV1Nz0KmiPzErAWvYv
3Muh8FlBPn9TIrdnHV5CF/CicIkSSMgSbwtO8kwPpXFoZ9hwEx1FLCIJ/2BW0oBeaKNivUfu2JO3
WRwxXK0krV4CT65UuizMkSxvHroI15geqlNGw83f92tGdlex4JpxZiifr3nK6Hpvn9PTNWkx4gTt
26Pk8aISAK6JUpmASjMTIiSOH/W72oPflaj2MPTqSQEmn7fvmzJj2npbI57uj00w+8bgZQpohkdv
AH0n9u7R49KTMdmA2mX4NB5NnBEJTHOodZbNwUJbrOdnfYthThjaeFdFs+1xac0mTMmD6sh17biL
JZmeumD58D24UeCsvsSKIcjjXlb+Ej+LJRbilZTPfU6EHZQaeu9hp5SMX4JiIyxKSfNUbzU/YNSb
bxxdXFiri5RRUDKhjg7BC33wfhfnn84oR7hOWtIzZtkY6j6Y1l4MBAIFecMBSMGVpBP0Q/9y4Zlz
v+XQW45W5Gj08OObCf8X+fvAqTTo+rNdvjnO9brD5cC3gLmyMIbUd5427WvDl75ugE/q+QmZxIYa
Q75tzvbD+03bdsf2yyWG8lCF9YYp9pmZnpDS/xf7Z1ZGN+qwB04lWcrqPlqfwEipFzWmz0XHv8qi
lLXWFB6nGd7abVbrsZ0FvK/KT/cmAsVkfK2gC1OyfR2FUT409IUOxsXgkzb+qZpsfvZ1p/xF6X7R
xhKBnrfWA9td2xMSyMcUhZv9nthHDiF7MnJuDOPCiMrBEY1sVCwpaYeMi+CWaQxWEZL1mdr1HfGO
SkZ2F7zm2xQ0yFX+89mCNLVwz0d+hj9Eh1hwyK4W0dXv5j4a9VDdf9ffTBDNb9GIxunWdqGZzG2W
mTWUXAl4Ud4Wsr02+w2WFgRlI6mDfua/yizbIm5cx7/LYp9zW44sKfciEU0eySQsUSJop/lsGVt+
921fg7IxEigUN+HevfDEYsBvGVvqP90H9NYygCGpJEy1WQUY8odEuijkz/WnEFbSJJrxJ/g1sNaI
nis5NzvU9g7KktP2d31pB61b+PN3/7+L8F3DlGd8stlQ1TK5VeIBQV+/2FvnCYL6ExOt8UpskHYP
gXiQ0kRxHF19iNdlrM+anY2XyA9qUdAVd1Acz9GXZ1BCbmiouOGQycQKyxvIhQmfw6caqgmbS3Wl
FSPzUapXoOzY8lhFY6Hc365SGsCK6R98ffcU5DQHpAWwUPgAZ6G9USicvq9W96rhFUN7rwVCQenl
DD9TSzdtvuF4DoAHWs/R68bX8wEtk/VV7AdfmWtgdvXTScBebDw4cM+f9uGfXOH6CIfsijLoQjXi
Q14HPNFPN9F/OToX5zE4ya6RR8b+yX4jACS/MIJJB+NzpxIfyEBrRw5QPPPaJs7dfT71C64hCuDl
BJ57BzMGaFH6j1qx50Of6cXS3lHoYek+o+QhqQgKIeFfh9fKUfGSnEgCHNoRESjTUNHmyrOrmGoF
buupgWW2Dc3szZKECLP/LbWqKJWJmroPxFSimVd2tq+biqFUDLHOoukFyg7s0T0SiM1D/nmFOBw2
Rk8QLBHiuFty+3VwB9KY+e344PsReAF/hbh+GMYtvIwH9gUMbw0IBpajMAbFD16lQWODnC6YFS7C
XKXawcXPXbh545qVdLk1d3bd4HoviD7rR8RwS08vE1o6VQEsP3sFOycK0qSFsDqM61y57hW3IkZl
HXlqg/fY4Oh6vhZc5DuPNNpk6ZqIZl6o9RVNx7A/mTSK63bTxJpU+IxVs7ZnQFynQx4vXBP68BTG
1bo7H+sMz8l3XTxX7kwPme5onrFCzSDfwi8BzXGS8XuRUh5qnIFomltOsEu3nD2F+H8x+ZrQE/yV
H6/sDMHM7+nYYSVkM66tBfokamUulSk6F4//kDaxgNtiOsWqFqah7eSF048HxsxfcQMVPCbRsi+k
cteSNrhG9FgZxKs+tVGdjD4+Ftm3Tg2/wZNGSZ8GulPO1IXyKhVI5J2H9dobt4/uAlFQxNRsxj15
gkK3hf5BG22gwuybh4pFuApilmEGn8i9sbJ7+P2OWtI3y2L2rJTu9shI5vKdmwstsPbUL+b/8T7g
bkC5b3JFFl+9qu0+LOfpRHH203lfPGg/BfKin2yKgz3YdsLBAnENA8Gw6c3L4AL9cSg5qAP8g+/R
5Mhv1bGDNzcxoOjdw8s4yH+biHERUBaY3cNS+tulAzN+AymES4HLu2rDIuukXPXm45KonAQianLV
30oUPdFjvdUWTL0iGjwu1Hf0CfiZSjZggN3somGGbiyV7epJbvsFAuCA1UHzQQ71O4pVm11aO/Sl
Q21CMIGoo53rmYj4Mn8cWITv9g0ml2hfHxuYpGYy8P+aoAWBqfBEla/ngh/lyUtlhePj74szdEgt
BXLJA3vurP+5rPuw2FjeMss/NTnAfrj8oQUjmGOpDyIoq26m61dbIun0ymDYGRCtsfyTAXoxkxWP
sR8tACv0Mnx7K3VvRym/bbYo993pa2egB2W9XfsLx8DHXtF/7vKQkrby5pzIcuoSJZXvOqT/1eig
VP2NRHZ+HuMCNnWpaXctOMVE/0kb2FI6QL0gaAegSrA0ZRO6AsG9BjaqKUwY0yvp5TYfc95Ds13E
Rz1RnEWk85vA6Gogb3zQDNLRU5teBrfjD+7eP4aETr27e7ZRtmM/QtLeE/JDoYpGqPS71E3+zPKd
sB7YyyydKdNngrqtczWlEbs6IznHNRjU1Cbm9cNBDYzS0gTVNuO5YiSQ0PCPTqpUl6usx8fCiJnO
PCmzfLut9vXiS//Bajk+rWye9nT8X2WJNg0FPBgdvj8B19nnYEa98QJEeAkYmU3+tSJvZkJH8LtH
5h+jzGGvvNJuDYn/AAlMWnP0m90aS31TAxIalsNpkwLB82tBWUJTdaQ7sIhSaTi6Y+xXIRlc5Owe
qiOn3DmkT7hzHb/dGzL6qJkvOtYKEYlAhp1/c1BTLBbvgorrBOes+8miotyOWm2my+xbyu/bbxIj
5f5P0ehdD3MXb2dGaYWnQAyN9enQUyzzyJo4BIeObApmQW6t5Zex+KUGro0dGShAQDUnjVL972Or
k0vEq5m4nsU/gQ4+CbKd2WNdk92+s/ZE+cAAD9mSDbJFvsCDHOfyprN/+xMmtRhcOYK1g1xWpB4Y
pRfbmWMtFdLSV6Fb30f5OJkfCvax5x3j2cfmDhfwZogawSJ3PJnO5vA3d0KVvjfAA96kmgHHcaI/
8wAr8UKrgIdNiCIwA4Ad73Yq/7eUiMSjsNwkKDYNiAoyiO+JoX4VPB/wYjYxkJUKGwV6Rwh3n+/l
Shzygga7tglrzVjk4Zme6g7++UYxkSuEA1SfWqM3qeMu0S72sL9GmFjDZmq5KomrpVYqdaLzjwf2
eHo8A/tVkAWPO8ldoKhxoodlg9gogILBwMpR1rKGVlsle5UdFOrbF82vF3Ah0AKioiTryX1W1P0X
hgsCjRSaGmGMuY2RouDA+LdS+uWRLfMF0elPWLyzFtEmcFu5SF+oZj+DSU87SSJi37b5rfESEjWF
zUSzihIwwyr6kPkqhnoxEOP4R8OMl2lzAwjJcTLNHNwfG93eoXhmrw5kFoouQfn50uIl6TPMXb2M
y6+rh7UBW7oAv1sblfrvD3OJC0zEvXvl6efIaz7mS7mIjPwzZIjGrwPtup1GN5D+j3XFmJ5RuLeQ
wrkeZfczFjG0k06ief9vjQ40d1O5MVqmLAHzfMSu9r/fxVet2m1Q+FvTh+qcm0xrhkdqg1KcVuBG
gitTJsPWI1Ymh4IvUxu0zM2H7NkInLsqZxcUiGc5KnDZ/cUcYUvV2ZdTXKommn2envp9uabUoGfU
O4MWrla2uHRxZnKfTYn6S0QUr3lAJnf34oGx62DpByt1KX7I72WMwpfaDzW2Mh9G94EbYKQ7tk0u
QdBB7yHQeTk2gfkF/QDewTpmi8b6ugeekAkNpyQTGoo/qx4RK4weJd/6YfP7Ac0O0tlS+1VxqH1s
DFCmcZHJku+fgkftu4g2nvXGHK0JliDPIkjcc/JTOeifssTI0TDhHNUFw5eIomEf/5/ZCx5kwQ0q
OKj6e/yvlrtmfJzF8O/wmFwG3tscpAgLVc7CWgC+x9Fj7NOhc7QeNF7qXh74dsMlxz7rXfnFITPQ
xgXwUuTMyZJBIviW7Pt1CUta5+2eEKL6+bl6lXfb8aEWKEoQ45jzq2VXeyLJKW48YQVm/5aRD0T/
yenSgSEl+2GEHDUUTRqwyZHiwI5/Dc94WCemzrDFGh/i2g3pnDXfMUXANgJeEochbaruXQEiGeO/
NCm6jChsyf3X4n29ThuBFbn+nfjjiNcIIGxjwfi3n2jjtA3+jgqk7y1GvlWtTbF0MmXusnWDCVhs
Ifn9iFazIbdTawb3lXoftJykkhyVbYggwT1fnGso1KLcyQ2gUvD6lVyHnk7SO6ZXhRlwlFJA/iyP
z1/3h81WY3kpaVQpCPI8edGAkYFPmWH+CjHk1RC6Rp4ZppG2Jm6LcCtBbBvNz429QHjzQgoStjvj
8dw4eTJYMBVwTpTShaXhHgcUQQ62Xq7l9OgLSx500tHLHgeF1EtMqeKMVXUJPjlG9YJs1Um4Mi0Q
KHUa5HFdE3MyTAy3IUD4CR4Fy7Z5DYf3E8/QGRRQpSSOJQP8NVdZUj22HYWZg+mScQX42OHIrNcl
BR9ZUmyDVSsnPjLTWNjP2ite+ujfXqrkdx0LUv6aKSSEQJW0UkNwNPHNo9QaLCrz5SNvMl25a5/t
7ji2feRr9e8CPPdtc1JkAWqVunY9VICYp/64nWRxfLJuPnJolEACGm3qWx4zdlAtkf02omKLJyht
0LQQakfUlnn56FQmjcK4hBzAeTNWtxMjUBY9OVjhiogWGQs+S0fHcH+xgjBkpPNLqqU0nL5yMqS7
mn5JJqiqF7BxdJ173VuTROERd9a7lZqwMQZlalvZj5Lbaldkq5dVP0kgCl4Cw80OvK75Qd/dqgeG
rjfL/OKR7Zk7elBr8bVrcCVE1Iqy9PxOjKawtbdQuEzdlWZbEFwQIUH6TJGB8thAXeNAUzocCANO
9XTJlcYTzfpp6NkFLmGCJ4p0sq6HF8A7HtS013P/bUM470dcA9k4yCCI2/SPBMZV114e1y+34kVC
yg2G7HtlHni9WBkyUmTt8pHVuVW90UTVQX3tJPA0oon4duR4q4Yf3bAgtPAykapLgaOxGFdmZhxu
EawotSTHTURrm95rw2Md76prFS8rRtqZVlzP+7p7cMMagnMxXruikXjmQ/7me9vs32OIsTRHJB7S
3Wuxbvumt0yh0kFLEcSc9As1wb34Ag4R64g8ihFXQK+PK5jUNAdMTI00bC+3s0sB7vBj+gix6gKg
GBkHVGFODilcfWWW//RHeH3F5oDajhrP/0MnGi0I9hiMKGzYiXo9MfVpdeqW42n8lsMSAe3dLGOf
J9XVJ3h6lPpwS8h2r6mFS84+/8sF1CS+xYLgnZ6h/foP33fhXtVpwYPNPVgZC3Iva1lcvyrNcE5r
SsWhxLGp2TJ+xebUMd5kE1hsFKV7EwC4sjZnBHlrGBpKWI13hLilHblyXNiKUufp8zQoRxPmiXEA
f62NZHNPYUn3gIwjwP/on98EN2Ahidq9yczmft1vfodV25Y1pwTlwZ1zWxq5yg4oGzs1Bx1pXMJT
dbUU61rZz0uGH764+HLsSpCrg11Ekv/Z0vZ27RfpI571GKe4MaUivyBhfOdWbLngIWtlIv4bFRhy
Kgvu/CQMVEunbtVhZ5UWf4B9EqYRj3bWLoVwsNjsLB7oUn+qqKmUI80ZOckLuSFOYi2p/Tz/V0xt
jSZiulHW5RBKU5VOn2KXx6CqXgYf1CIaVrbX3m5XEnCs+TLwFls0t/cnluIuw7z5ED80WLerQiPy
LkahPw7+dpZr3gP8KiZvyInBx2J/7qEpu1sdXIHj8Y3J6poCcu7R0rwjkKm9LooX8ShqfYkaQfFa
4RnQmlpr/31sDDPkuTTbPc3CJCOOD6hKBxGDP62h4ip/ESqiqVkn6LKy7NEO3+a4oIaBcps0x9Gt
2EvCj+lifTNSnVqD72BIVrmdENV8lTR/SEmHDMwMvLKTZ0flKFyapi92ZB8J68/KNI8SezCbH+Gd
RUC5AyEsQCUEE3o44WcaQUXDokKk/5h9PpZmKtaBUUJE8I15heRUwwS6qJbC2ae8KeiFnCjbRuch
1NoDhfRFsMGQeQtqxLhTUNNAPaQK3B9+QlWRGTkC6ddhc1CeMiP2RnPWt4+ZQwhAJSh6Vhu23EPA
KoclVDbXknuOGLctntJWJylGCb9XO+VDfeEyLmdkXD5KJkCG/8ojEujJl6oV5B0aYzbHefj5iCSv
kpi2PChQurbWcg//KZwO2lRtFFTAZbJL/nG33XHkHUh0LT8B/tEAqzS64KH4dAl5JlTt/3CfbSz5
iE0IeRT39U2P24QzlE64dCZViuHyFo1wJ+BMgJvG3wgbSKloz/IoqYGHcMYSi4kPEcrP4WCBvbmr
YmpSo7dob3oNEpG5fgqfti3B6gc4TnjjBFuPC3QejKNjWuVEGMIYH1wf76RfImy2KlUQb79HpvrQ
baLHLcaK5IRwLxSNlz+7OldlqxzqkK9DbhC0jLw2JT2R4iiaoL5PGAuAm/ysaJitA0xl+dH5yFkO
FHRiKoGpXfx8IGYr6q4FlrjB5qrExr/cbSTufuMccKCh3+MIAzTOfa5l1tW6obZ8OhfmsDQX2fQU
7qc89DD1ckPLg6tfVmSPsTC5KjQWukYbfGrBtP0yh7etdWOIKg/tvSIeemcJUsH3AvMb004QtFrq
/T/naL19+M4M0Ezb4nxk48N6ge0AYRKVVBvedIMhKI4zwMD71uU6fskyecy72IwwK0+nYoQaZk1x
ItuVI/wVATtxDB0ku5CrEAwHbl+tPpn9rMte6AUI1HhIjPbGTmN9llq8PwoIC1a9WA7T/BBvHKeB
Vxwo5S6DBQgx75V23Nt/2uCO9u5vTX+8Sm5GTwjmILoLFNeTjU0oHKlfhPbCEGUydmDdPjo0lFsi
nGoXA6m5HLZHfZ6Z17S9JqVYQHgMBeWbhNGCJ9PWNGe6vEzoPl0ITe8O8nH3Pzee2gbCmC3rRp8y
A/B5L5zpnCFsjs8MyHGQqzR4z6SpfF5Y0jKtkBElKlvPbOjvJq72mwjUFRRXclSV0BtJ2ZYzRDQH
xVHCAVYMDOD9aezi04o7gz+haY4utnE/CtrLhXcLgEizHj8/K2lhbQt+NrkicPmmAN8NXbWYsrwN
+xJ/c1Z1z8lI4g+N41YziW3waa8zF9c9Xhp0IS2lKdrMWivlBmlP/HjrWRsldAVDZwyqaCOOe96s
+tLldGMiEYBOSFrdZ8WQkZ2w+Xq5hBdSqhwVwRrYBD/uPuIWrqjD9TdmSlAAhZA3j4CmMlbWzm0n
NgDTJIeoWi8ouMXKZJxCpja4ZH59c3TEooL9zi4V6M2PEpaVIy5sT6KTvHqs5g8nEsf/+1U4mpHE
H7XhamKsyyVed6tJ5zCCdhPfTP+VGn/0KT1P2GGpwUAhkoh0aKfEJiV2voicXKvpd+yQIXcCPQlt
xyP/MyxUhkONJCcKFCEXjA/NPcRbU8DzOgmVTZZgZcJcLUlSiHF/93JnYE9IAtvkMqD/wpPAUG8Z
51A32a2h+QTILgI7j0iY/B0pNWZ5+OAXh0Up8n4oKVO07W36aW6Js3cFAuGXQt5aaiv3trregd1G
b7DbkoMQPE3LWdic9WZZ9uhHVVd0DsnVYVOacISxUVh7X9I30GDF4VMv9X2vpDEsH6nCR5mvCp3E
Mk7fwERpnTXorXBrEEk2qIeCHrNFETmf9DwVn+z5vZx8nwlOvEzzAV/4aLCotL9/k9pQ/vbIycr9
pRr/+g05vyaLRekO97R7geM3hCPQUvsA9UIuH1AZuB5vHo4zaV1Fiu8cZAfil7iACpBZi6Gn9eQl
uHwAgc8tI5rSnVGplQyZ7hEdNM2wVnssAt3J5PirfbAYC0HOzNcwGcbf9rPC2RDZfvT1mYSRNQJn
tI3mEZ0hd4HnVoLrQ5bpofzzbD3ZyoYlfiMKZWDlLmKa6Zy4MoZowK1kwCAWaXikxavDz57VY7il
cUQb/mMUdGZNanH4StnNT6Y1QSLjvx4F6H7DumK3ZIuVO6XwnD/ZmxEmPIeMu7QHy0iu2v96bBqf
0+MBRVt/EzY3YfRU8avSENLePK2ZhI9VfNmM1eGxJFPQOPLO20UJHDScSV+RCOLDaJxlJGGjSwxP
Ya2U1KmUuVMvHoSqYYKrDQkQv66cqHmGWiZ5mG0l+dNk8gwfj20WgHZFglV4/ta9kGGv61Rej3om
DPSxxffa9w4+GbdVGWmk+3IP/ywpm1gs+NrDw1gRNrAsc/ZKOYx7ykoNNoyuU7jZ55hEdpgEE4k/
PJ9DWNdmUVc6eA6SkXNN8uCHEASn/5n3nJW0d4Efv4SOi2PAryFjGWJ9HPXnyLMt8thmn3guTE4y
iM8n/1VgokjkmNolUfRX8lDZktiCI59Ma4HhrqdEzrGS8vYmo1X0H+0S5KwVK+YjmevGFzs8A51c
hJga51RR16G2RER2zYOXgjYUlevP2KuonqfoWCFiFx0Il/pjvS5/YioTVOTop1Tl6WhYyH+5Sl9/
Kk8KxvXP9RKRY7lD6Ti9gePWmR2JZOqBLX7Q4wmSvv3W5FN2pvDSw0IjmZ5iylY+IMXk5hn9OTxw
itZumYmoaOeZJcxKyvzNNj3pZfvmY1noqvKxXs7pdqQHbdGdMKIBzFJvzvnoHGT8FXI2wMl4JsSU
2u83ao8gnwAvLvfpjF19NN43wBGRAoIFM1VqjjU8nIWYgDQM9qndJ5Q3VAd0viSpFSYQwWR6OesP
QZDAz0qL/cOm24FhfMjjHX7Yip8CyPrXm4KnbeYl0lguBby727n3paqwFglqdlBgG0HOWQJ9gjud
TlVf8931uUB7zwlTg9c3bU8/aiOZRRmGHmTHBt/70c/BbeV4UKFqSJrMiUcMflslGvJ9ZhV+Gweu
LxNO28qS5ZJTcjAypDuIJgqgpqnMwlCiA397WLcb8zJvQPbuvOvTBKi7LqwGCUR3EtFMC66pmh1T
hBsMz2r7YW6jQsOn7n/Yw7hFq8bymAalEw/MlTQOoJ6T0USljBrYEHObq+/asT/EM9WzhX4uunE6
XDPAQHU2yP7XCo9BBqb6ixWg2GAaD8HW5sBF2rVQfrolwPMZq5dqYIiJesy8rMbcWZ9O/Kw3lsw+
rjKtowR21h1cLD169Q43DFey8Sl72jxRg1xXXteMF7w3US6Wkc75IUSd/sDX93os26MG8I9QyM65
VCgykJ8uKyK979lLPpypynA3XYsOqZkU3m+G4s3e7eEE/Cr3ia1fTTis90gXLYmjDyIwbNZldYBI
vLhWlM19s1fbof2gvRgimjVFwLu/6TgaMyIhNmJAQaMBQ48Xn5gd2SLrfqD7VQlJ9tIAfVng+VKP
7cq2VtOcLJGafr3zBeiJNeLn3DExQKy766j1ydSPYuGsuZHsQf04j93BAwN/NA1HtM1cXr+3N/cr
CSgxtXax8Nmm4LWc+g6JYF1+jkbhC0zgj5coSS262Mjj4m+ZeZ0mIaDTJhnddKBwknkVkA8BD82b
XsP4Hi2yNMu3ZhTA8SzR7oXFWMTkXFQ2dm3X4d38QGTABcI570cfhbE+8277FuZJ8BdDYHlrDhxq
hPenGUPWR3U2yYUGGg0FUyqnBR3wyo7zzhgEL4Dbc2smED4k00FliXiR52tPRLXzHzJYO8Ob9MHM
pg07lItlIr4yRWA3P7IzKhWvXyP1/JUIOo9IyMDypk3qx7RCi4adTKkPZ78hDaxwv57umtgYqWbY
U1VGRDgL5uVUN7gpVzkd4jPirCB1WbsVVMDeWP+BURQLQ97yJMWPVTsM2EwrB61BmnNZAmpNzfi6
3KZSipn5jK2CDmgL/5ZYk6oh4UW+oo/dbhkDiy3bOVIYaQAfrlsY4O3rpjhbYpWM7WSBl0Dhf+gU
rCp1ZK7NI2teVm2holAQRdYgA9StG2kt3VdzNOy1Be7m+x1HJQYmzTbwBSVl1LG516KnqOq+/YqE
ehr1WYizJNX5Ywh9TTNzEAN1uGWSgZb93Db5uueaueH7aQKfTMrjFnqZLh6+2QPUhgyE08x2oAiy
VDdpv5U5cpnAIDN0DQAOzfH8w7p9wcQ3ofEbBeJJ2cpYXCkjUI9T1rUnVDaZ82GvcChKZ2wCdNpE
827RrO4huvh1B4oWyQZ3nPysyAKEls59ydOi3i9McPh8mh05Ou0FhlM1JfWgj7bDoTjoiokFXmE0
RTbi+n6B1CqEaqJ5wjFVLIyTpyr0BhpQ/ygjQi4h2kD/GMaOFqLNc15pDQJYelp8ZU1G0orEtgMY
0SOroFM8rxbaXNwQ8yvN/ok0n1A0ZwEAiPS+Vu2zUfhEzhAOjpgCTVgHPSOndyiqDrN1givdxJoK
7+2qwoUhrUoyQ3r+ZGZzi1/oGgVIQ9dSm4am7oqsYF5N7zg07b/8nbNZWr56LhdAkFaINPq7l+AA
MNBTKYBxmCPvZfV+W6Td0vHK+Y1R5yUCQ1Y8hbI/Q+yR8bZu8BKQ3S/qqV4DxkgU2TnHHZcH8ydl
S6ZPYItMcfjg7HG6ltjcJVlNFHEdvU9iXKU56hJVdmmghPgkKYfmM/aYvLMmlxErDxUBCYWy0nQL
zuoUzG5t01VUulmjI6xVhtRe1Kxxjf5dIFnu7lt6Yao0rwvQEaWicAZQBYlaiVbg2UmbA78uW5NW
hOIcl4rkpFMBmZzeGuyzxbcHUboKEQG+KCY/FRL+jJc7rO/slJiPUXIycJZ02z63KbX8oH1g+z9Y
Q1EJZNBtvf2xr/HCcKqc2PMkvgTfAKXtjBEh5klrMiL/NLrqH9GTBjJv5+MLJNVJG85r0LY48xge
tuQ65iH59tU3hOvoCU9m2a7siU7RZm/Ub4p5InHx2rfupvtL8PRVAi8tAXNw2upzCBb+KduQh3GI
2ha0GMJPMF7asmfc3nIRl/khXGJWujFAlporCDvqWwS73W3zNZB8sxG2Asb0q8c3g+oFYX06pJkW
dzjCIFuGyrj4UGReSlPuPFqGSRG/zfWzEc72fIwIqBV2ioY+zBPq2w31Sgj8nLw9PYAWyJ4yKGf2
iEhFNo6mIf/0x91YTAAPQ/nyniJLvW8STP77Os4PfTVG4/J16982NaqExaIQNHS/d5hi8XIztIgg
AKtkjAqjrVk1XzJFzgz3uiF3PRuoNgyWGq1jq/smTjAam5vmM5EdL3vjw/SXVwoYWrrUWib0LvmB
PbIEnS0EacyjdOU4YCUs0IY7I3VGAAwihcJ5IZpC9wV+x20wZiJu8mLl+UFLdq91Z+q+9HKh6mpL
XM3qAgv7l7cXWUog5HkRxc1epVeqcfIZcbhhhyxFxfViPTyb4ziWrYKxO9AbxMwuyVaTWmGNm0QF
2YW8HR9zZqoxRAfcYCHWQbx0bDaOcaQmFsbvBXUK9OQhkDQB9/N0JQCfaxLJ6ho9OOii0/w6vS5Q
7j2zh56GPfeoFhcmsqnUquOVVIPww3IS2mel0QAVESmXZWraXC2+1/y8OcR+HSFYbMIW8YUSHEqD
b2AELsdKUxgmN1oe3hS2yGFzBe5N9+JVJl4UHuFKLSrD+vhCJBYBr61G+slJDlTJnkU8Pr8F0184
lrvE3OWgO13mlfrkqVhtvFCSXDYERzCVGd642uYW8ds6kHXJ3a1u2sZATrm3Of3El/HeIx1aywpU
pJLiCYJpBf3PURQrHbLSAyaHPmdYPasT/9zdlSkhWmBWK85fFpx5cHPeHsmAmCxghMLB8Ide8PC9
Gj+i+3Mc/flb8SgQXXOIAV+Zn3Imv/3O9vVHcZWBPkviMrJpUS8m+EIAz+2IvvW+3ZOyMC3Xiq6u
jlixBheQc0lGNe3eHieOxJW1ZZ+f7K/0ytUv1+2bnJRd71d6e55Rzl57eKfPfRRAja2kTb2CawL1
1ztQoapM3m39zFk3VeGfeRwsx58dHVcj9T0h8S9/60+QFk4a1bIXJ/TvPWMmCFcApyKPOAwqBeSO
lp0QD06rhnuTSeEIscHyhOYL2gQHr993zcKpAqdlfXRrWDAHVPr1RB3nx74+1tWJFTPrZ8O1dwF5
uszvgU19m55Zpz355vJg9BEKiA0OEecP3T88yBAtgcjQEof7kKZkX5gHYgwSrApICya/zvQaeLir
aQ8Wvb1Mj/PCYiKlS43DPuvT3c6SbFfKrTGonoqSaYogSxtciSRB9m8Dq4UbYIKdCWLXCZ9rcL+T
P4V9TruhK8ovdlgD5Aw/ANk5oZOuCH3kDzwPCICRaaMXPxCu40pq79V+ldy+EmYx1GW3ylI+34rT
gsrKXN3cvt3TBMEqBKIXYb1aDzBzhWJqcBcYBYgzanfOPOfss5d63INrS5ZEiW+W4MKbch0E2WVZ
Zg59kzFVyFbTKFPwEQCuLUeYjE9WxZH0p+diZkpLkg01vDiszAopNezjIFIU+80lx4mKDTWtqSWT
INx2nsKfw2YezpV2xn95gt2QpVgCJHWdcUsQU/4l8sC8LKTu0laS6CihJnAvmIx4zlk0qTI5O/Ax
1FfPxa8tVfU99KFY/LAccUmx7RtGQWZJXgP9/OZBlCPri6UVxlvnT6BYUiM48E01vZ0SZ+ouCtMR
gq8Dsif0IJG7lpNloAjBpRKgA1iURL+CcQEx5R++BnLyJaXD+M43Op2lfq9Hyn15g4ndMuu8JHX1
4r5Iea1L9qkvENmsBZ1oOdMGqpbHNqTRVDJRcDSiQUHyHnhpXbCuHiPiMyG3U13C04ZyWw0lTpjh
5M/B17nF+ZGtG8lqNIeBOa8iR/HP3ucInz+OnWd2/O32DqAYCbJ64jbFcNgAvFi3RgArzNu0MSsD
6sUW9LKaDIb4cSdlUN4H4sDo3Cf88dv8bfbmkcroyT3NZ4J4F0jigVY7KW4rKi6mpRQv4YCuYUAT
Ny7tLhrjVCUcSsjK9oYxQEmv+VAPcA+XqMZ42IZ0BWejdQHhru1Y8GaJL2kil8Pkf0gKVceJpLn9
HuYW4gWz/HrwoF30vkUMtmLwuzRKbUx9EjIueQck4+SYcAKn3WaM8mvrVoOF3RnmQ4IbeHFlx6Ow
hENoe0dvOus79mMLb7Bc33tzEid0i4BFwCIByukY3ObTXO2yQsEX2+CL6bEX+lXBveC+61ssUY4C
e7vBeY1npHvtFDxaMlgiXYew4fq9Cpv1ZvjmXGCVj5bLza7U82JFATJXPkFg5T/t+fCWNrAi/JgI
ATeIQFW+6riKaHz1FXjHseGuZpqGAQ4SqF40L94OaYVJHgCeSSzthDXkUsW/EiyHLnOFIO46APMw
mnIKEGmdiTM471LyXakt3V9T8tjMU/tAZcLWXAUfvWBXjYsYtWWCkMIVDKI7yyh3E6iABdP1RTjP
ReQiNgh6oGS+N9bf8VzyzUkyLUIeW6Igvekoq+a3MWciRumfs1hNBkvGdzgYtO0lGbeBxOMunmpZ
9kUuMGj66mPUgINu1xCZPGzKiScpBTBfY89MUle5eqT+fuq8iJC5umqOFaQs+mZgZh0qIAFdzD/P
bFSxg4mxFDFcaxikof82ceLxjZqWUFQROLS5NiMpR7hwU3W3jGT54yxrla/9uQbnxEhgvksaqgqy
X5VVzZRPZE2DWXjtJQbagMIDQ0NJL0UPdc2Jdu9jgt4YgzdqKQDXopLO6Oyo7k7nFEESW8HCxLYt
DWMtlg6koAWMLmmTWTGoWQJzpL65d0X0uWFU2mVwuOF15sZ9mi/dHxhAHAVFG9jfFEQiBTriay9H
Bw3m2cMRAJdpDQMN5cgRqNWuEBbtH61q02n3mQHk7SVZy95rjI5E9uDAJvZUOUhNgLALgY74asjC
+aCl8gXv6sdLXJ9wIg9lakzziqx30TzHG/MhgCnuSnV20SbPoOKZvmGXomjkpkvMEcCjveGAXCLc
99abVqtOuQ4VuGDqpRld4Ar4qLoF1YcMYmd4upFnxJQ3gsV3CwD6ciM7KC5jM+0dm2MA//ice7f/
RHAFW0lWx9uq/ma1E9vuxhbpqJ455F7Q6SpQZ+LYT4aLyv10Tdw0bpV9aH0n3SIOcX+jQwLdzwLY
ZlDzKlreQcZi1DAOkQq4eLuMsOfEgL6DdCz8eh0QwUntQjr5EM6+VGoYBEenCxsypf7mah4jh9FI
VT0ubKf7Bxa81oZeYOl22bscizvjEdvsh8Ys08xxjs//TDv3Ua+YHOFIfYB9lmJQPDF4dAi3G2Lc
YEmdFV1nMqipZf4tkhkOWGKMWAxA0OMNnlocwM/F99BfK4TLiK9UZNrY6+qId4+GH4B42mh4zmYI
ORdACBRIwvn2cXI8lwxGUegovVUVUIbP8fq51m3umZqxZwtWgSLR6pwTvGPSQmJS6gP6S582+sFr
h8H+Kh0w0dQT3S/vTpwC6bUrlluDQKUwC2lW1E+UHZtAOPA/sHBROSSKwLXOAbkmLuYisCmUnxqY
oNC87ToyyS34rGTW1FjT43vWx8naAO3hpaU0nGklzsgZYHmYEX4zubR6qU1r4UsYZgPYmNOl9gCO
CRHjGyGQHlwXXl8LnnkMqug0pruDCbMs7pq5BejmvNOkDf3+wKLLdpIbEMFGP9ZPlC2LnamwUyH1
CV7TWORl1c3nEDp+k7ZP9kD7PLOiJk+EzGASnQTEo3/6h0Biy7cV0Vaewszl/o881gBmUIGc9MgP
N49m3fglDdTONE7S3Z1AuSzwCryh7YdOOe9DGEVEbFCx/muk46pkewo/pD8ELFlmPSDu34kJvEyt
fKZKBJnJiul7Y3xubvGtiowcvLJXtlVi9gMfwlSv0dRlCaz7EhhWKLsdAmrxht70/dGp8UbPrAuu
jB3WAxaJWeHntrJ7MnBcLWzFGZStbTNncqE9omZNhCjGduv14iPtvACq1yrN9aSIRQpH0sEBWF0g
BmH9GWZy3ducPNarBl0ouSd4Aw7zcJfP9DRcutegWJuRxezXQl3PXq8oy1xImBJJ0bP44C9uPFJb
KWPG/CY6a08DcDttLePsWm7JAq7CNR1MrwL8TutDNT3oSE3+EbjgTbDdKsqikJWCwJp/TLyQc8wC
oknVUXbGKWuOaMfC/U38ctd8u3QXoFKHAa4G9jSgJ8/LyGZ7BHEqVJckbi0K0bBQpBm3J6gwecBY
Pq1fYEibfH3t5dnnmLg9amiNji711ONhn9tUKJ1dO7ge3CaG3+OY1TqLtNzEGEl4jzA2xRu0/2FT
9hOgRLzZfawyYauH3kM7yErO/g1ybi+z/Ge60jkRa9WiF9o5MKVoTEqCPwG4ojBVXjbK/LnrNYBL
neH22ikPZ3YD+hPkBfcse9zoheO8BvLUiH9t6aT2gYemvX3lv9vgGlEyeYHPFvEtIrUGxwrKPxNX
4OUnUH3EQkKpYVhAlWH73MxsXHENDAivknqR6EMkm4ZISd3MDubecK4soPNQSHqc2/CBjNjGT3ji
9N9qsiuZAHUi1aHB3Q0jBaGhNUofRRvGSSujMokvb3DKH7SxluMTVlgklWAZ3DnbAQSWQnwieV5Z
Zm2v6SOn9xrjwILMxCvjVsdVoKQ8FLPsA0TqAUB8cwavmPivqydfLxLRZsRCiADO9xVZPf5lEIDm
4csAZkpf7OqATC6I8CCaUtmbjq+BqALqz5T1t39EJZB/tUq/GXcx6ta8WIY6NR3nWcB/NGVyFBlO
sYQb6B5eM09mFNjouar/gPnHMaaNzQakrMUvi/NNaLyjITv8VroDNF5aMgwB4mN2BhMwwcGdqyA8
FwC6R11xTxa3VCJy8xLjpqpZytL7WlLfxrN810BjSjg0rbCe//1AQInKcjq+tfj5sh0wJDt8lACy
AdSgkG9dZ3RgvbpeLoqk0wEdzbCapY814Al8+9vSzXWSnFtcAvS2ENH500gSt7QblJwTDskYzp8A
UmqnCENIJebdJR2X4BP5M63f0QkQo/kOzzqSb3SPxs4TqVa+Zxx/3S+Vmp32/JK8U4FvOM7IUVNA
vNvGCGsGfDvYScxc5mWZObGKgAArChEemNNvw/z7p6Kh/5wdRQRcN79DrG2+J0+4sskBgzU2n/E3
pEuCctkdOrTCv3/Du3iuliT0VkzUiSByGqGmVxbUnp9VgMoAmCLS/jh3Vs3F/RiaVFhxItIGsx1g
qmAluORQ+vBPz0gKeMtPqLZCJYe1m1lXQ+q54iDzJ9mAn7P3Cuk397GoL/KHTpDuRNwAFL20A/wN
SdqL2nEFiLmiIjcIiU5w71utgfpfIzAMxghIdDZL44Wk1dOPhkR6+ltC9YXfHD6xXnffFPe2lPeI
JrhHiIiRCzyHWc/iBXE3D7fZJQbMTTGBcN7Lg9zKNdjSJJUUMvyMFoiycKE2GoEhkYKofLEPiv3v
zLL+y+QXm0ZmiG0YAUdQTklmhfNbAhDtgaskqjEUcyBEJICLWzU8EADMA95UEF4XRYrU21CcOHgX
oLtXMcnJf4qWJ0W9zuUWU6FpOsJZD72eIheVh7DHzRdDmOZae98ZaBa2VfH8lPqXbgcQ9nMjcYYg
u+9tLWQhvMOrF/a1KXHGwPc/P3TQD4rRotQheUQrsYQbgfOFbx1u6T4e7F9Y2xHrkzDknOavzzh/
ZV0axzU/cUleTVOJq5M2OSFTD4xrt4g/LCMDd1yjTtVqkYY57nJQuooZj7/Rl1wvW9mA7xS9RHJZ
lM7ocNyjLvL7dbirTuZgBxNH5X9bqsDrBwyczqQ4QMYuhlwesq/4OcMNuaNOHSDFk9K/067kitCi
Mqoc5On3n1lGnkHeiG0SzD60yS+zLEr25JiYV5/Af/0Gmnx+7TSwI0xB5/bWnOum+5103KguA/Oj
UY69kCDfuPM+lDd3XAPq6IcnDMDgHmZ1TObdoYuA0vqWVjC4y2VQkT6mJ8yXyWjlZDTsKDDVVPnv
8wyNZCmAo88Kr1ouQ5C1c8mx6ndZnoyk/ds/KYG2CNnsI3EAuhAn8CN6J9q7msymcj1vCMq3qFoc
zH+pmjoAYV8RNrqrticZ14ztQzTxHXU8BbCorp0NnQR5frmrunEDnC9p2DcSpgy/eUjyFoysDrAq
4SrGPPp/zkw2EqwfUGr8Qmy7DV6av9UTWoKhMspan87mmKYdTXdOR7RKvuHjVmiKwSb/bsjPe2GR
JNrLerFO/1J9C2Atj8OABdWEu8+6eNvLy6WOmUuiMZpsftvwFEWWB+zW4Q6kBJRI3wDYecgtq2rt
zP4RY/yh7OZStO/HTcPLNwJmClki3H+/Wcau27ZCKN+w+cghxhnOCxLK6EyBWWHXHxkgqnthej+o
E0be4jdRMkXjluqq2kKqYHw7J8tobKmH1b4p1xznFx6crMgBiXGavBCahBzM4B63QnTMKH26RZCB
TywKeIwL5KmFvu8+tbgBVS70sio3OVXpHXmsC/ZhNiecWYukgq79BvI7aSw53opDmRVqGqpe7lZB
v5CaQg55lzPkhyU9rl6BPedcTDcddh5PlKdI5LF+lBPHj6w2I5V8CO/RXP6VZvByUgfWocUzrQde
RbtFsIZrXhlQDCMy97pebpnU41LgK9jbDnKCPqbIL03IUwCQZiK8zJ2J04V6rgGiqS+/kbyFxxpB
vwaq85K/N899JVOMVUdFKFkvQm7OVth60SVSwnDwUs5I+nv3NAg5jxzpLym/YauRq5VLURlLnWhd
Gy6Y/IvXkAlM3b47nq4OGDLVjUYV2Rj/zZvD0VLP4FSNX4TFeanMgZ0uTH4g2tgWBS2u15m3e1Df
WTM/SlFedO5bIGzKuK5omvVzfrWqYFU5BN/E7se9DmBmgGT9Hgn6z1j0OxWkGsBqxq0uEYzm2n42
LF1A6WaICrwwWDfEt4hokDDLEPpPjxgc7wgg+P4yL/vW9gqWS5frWpZ3NO9nztjCJ29UIKc/VHJF
/8ZfXABm318VXPfxolvufJbN3xPkiMIJlh2q8jJI0/azw08VeNO9FdAQVa1KlTw8rOdEg7prRvty
HipoMbFGWxHxbBIUTrj2/HMlCI23kG78PNg5rYrI7JbTLTFFrbByizQq/XRs73gSJ84uJAGOHccK
mhTQtMitmtWD3NMT8HXX6nVr46kxkxUDMuYnQH/pmFpVNUwPDfgoLF5EuvWeOgFegqi1ZK/z0iuU
qpMOwXkpSN/ZW+VhkDh4zdmk269+iGCnlvrP7aPLizdd2eBVd6q8R93heMOyIxyVkLyOpCo/39sW
EoJAPN8X7kRb69VBGOAguBYrZCTQQwmvsk0mOadlvCmgaTKtzHnmoqveSZJsFhM6364jsLuUFtB+
pQLAMKgDG6jDMOlc7wpE+zbdsS6ryhaEnd2O+OPc+wpkHho2RuQc74nexLeZ2biB+Gdi7D9K56Hf
Jv7f8sdhJ2OBRtZ91SL0aTWf0/qWhlz8+FY2pGuLwYzXr2YzimMIYmxxBf4UcpPUUimRwaVzs3tn
O4YaAfqOVQ+de/w03yyK2GLpHQuRMbfk6Wj418vB/rwD44RuxjNoucW7m7Q49+DUUOTT8Y4D3Kai
jfehlhkrscQn41EBQPfE0t6r8e0tCrTj3yqVQV0Vn7AB1bonHAANGBkcbKqQcnl5GFjluI53Icry
193PzViuyD8028ToyRf/WDucmN9Y+ByFQmc1pX8SLCfuTq9uCfo25pW9COzOrrW1yANp+NGxBDyR
ybL3BVJWU/lLJxFvYEIm2Pli8WAB9MnzliLUIb8hYJBcXbgWc3k/Rt2a6KlCkGRTEmUpmAi2TJjl
d2ZtbsyE/DNetXZCTN9jb5Uc2aZ6C59o+pDtglCQSoHMqX+Hg2q1pSHnNARfXdwW5y7yH1l/0KV3
+Z0lsYGAT9M3Eb+AQibG3oA6SdSYOjD//DQ9jDOzmw/77qWficZTocMdQHUjtSJCFrb1q6/qKUSv
ulsYaePTxgY+Q4mp0CO9I4Hxmatvw0wlGL9PRPjY4GB+40r9DquUq4/Z2WerUzFYkSYjXDUS8BVu
5KSJeogvzDfx1CJcPAq6t+b3+YxD27Txstbv6AJxFyiMd2F38G7AKg4IcZCS6aTc9lg2/fVuYztj
gy1LqKkZ0f4od2hzT2MrHJqSF+yYCL8w7+08ERmmwOuQSjj4Uxst3aCZu7Nv0D2kkicpnPzdaaJv
+TI1uShIi5KhhJtZ5T1dooqELlKkpENxpgkdz5dFJWV6fxjG5XehNwNDReofPFlxHYHwmnvRcHPk
LwuFZ6n80wEfObveMPVmRZl/cu1Pr3gD8bR4ez283qDZ9QBgK6TlpsDKWcpAAkHV0QD/kOyViPIq
U4MRgHWoMRNQ2MlD6KXE91clv6dqiVLxoO4q+KMk6J4Fu4hAFNBK1at8Ikvljta4LIlIv584nSvp
swk8Q7NP9IXUgWo3SlmkpdXIua/ogKqdm/q47lx8DdlUfHGvoD4IKIYDawHM+BHiWHMYiRxnbdnl
eA4xId1qDEianUe3BvtcqB+WKu2AuWQBqqEEdBP/XdvIbaSe9320WtaU09vzNIWFhJy5taTQ2IkN
Drg9CbulTIwr/7NQNCf4XhtWSLggp1hbIJZPZFOUCm/uMlLFpYwtZp4E6u2cSiFVGDbC1l15uEd3
ea5typZz3UbjrJZHSenGbXEnF1LEedsp/XxsGhe3FRf/mj+bdZ9YbTi7XCcdA+eSvMS7bguNQHcL
nN8pOWguBogBLa+gk5NVMiXpSafqxGYi6RwvVxu/Wk/P922Gbcdl+9YEWefKrIS+F8yI9GtqZelu
rWs/pQRiMYBIwDSid/50v+ss47+ngn0ywT5QtyhD2dqQepLvhXk1YcRDViwOI/6NPj+1IlcrAi+b
YMfppQrlMwhjaE7BPXxmPvg4+JqijCqc6Tvtu0gh0lOG+PWqUuOepPaHj+b9gNNQKdhqv/094QKF
1xpzg95tP+jA1V5Ho+o6031mzTaERLFInaPFABzGn2GSa34r+O6TacarweNLIa7YD9Ux4KHOKf0P
3XKUTG0vNRSwijnjrwWN+LDDxBrf+6Kn1Kk117EBPK/KqwQ95ukD0f/UJG3Hudg3o5NJNoV59JDi
eQAddrQpG5Bn4IAxbWt5BlflfqrsbYEvHU4BcbMsaTzwGgLfPFVvtHWMz7mxBKKZSA5tavwhsiMb
a1utKvzhqg763ovJ8hXcQstHi1DXUtqBJbLr0tWsqZ6FdEMXbvINDKdWRshcfOVSebU+cIi7r4bi
BdPSom+LW2wnVmbeb+4dPNvuGRpRI93/UEHL+LN5aRv4V2+DLtyALQtZ91dxkGTD6lzWOhlxg5mD
EHqvB0N7ijvKMMqd1ThacEBuErFmBWA0IN9ORDWlXOBmafNHvopWp7H6ZhZQbHv2fOewE//Ge37D
0hVse5i93WDHE/WESkJfG72fAgG2gzLdPjUOshtI7EVRtjpPBWiYzj9FPcNZzlvUce69ICduT7DC
mLF/IHPHl6EEML9lNreDbyHB1FW6IZ7TRwfmZw2brQJGWri7+Y9/VIfC9LKNXg3TgXIgSuApG7OR
qtk/9pLHUkXjiUcNEwgNm3k8vS2JemQPybprfWIZDuuGEDLTHw+DB2RsWWfzWIdirLv0JhuQGt2M
FD7ziD7vBR9g/lMgphAlv4wpa+yKOvkBvFRXCt9a/CmFBlk4vMKcHg0JI+zPVEtaUW6IF+KEpdKR
RflpNVey7X4zCkepbyhSMVoIlPfOZn+Fx0reZgsd9KFMQE/siUP4FQ8Gr4jNrHW4N8jHK1g4Foae
emOtFJefZuvVt7a4pnRnM5S+fxOVtFj0xEgNdM4Y9LqSOIpFPu3pBX29npHvb4DWvKYKGHW8F95M
cpr8vnNYQZguc3uh4XMleQB/hScVs9PZP34kif1rkqVyLrVaCbVNUdOLwnlW44Bkz9h5eZ/i7Jzk
ZFTo0P+JaWJL1UE6O7j9P5rUWDf+pqEFvf7ihhIvgE9aAsCx27ucNsNmU71qDW79NUK+P+QyXQ7v
BzYCEYtc95ceYpy8MPoJEy/ipb3xrmXVfu2Argf5x//CblDEikBqgTd10CJjm9nH3LHBO7Ru541g
GEbBisfJj4mS/mB8TD36r+l1yN5c4PJtwRoKuFGOFeunStwHs8maPS76/QPSYMhtr/B7Q7WDLpw+
fTsA5uo4bBWB1YbFuX7zpCdPzrUnPIzSOn7JuQOpzGcBI88RxnND7nNbEeHpXa3q3Z6zL8XZtd1I
EiYPrm4sOhxqj0VTVdEr8OGg+BL4Vbu8FlUlNWrPJDVS+2RW2LsPBambaDfnG1EzEsk4VKbjmKkZ
NOX/W7nCLoh5rCCkOopHG13h2Ow5N2ZYJwWlxS3AOHY3QWkxlSVw+Y2yZYd2sfxhTYM7JE91/vhh
Afp/mWIepLraUqbmgIXMSKoAqcW1w7Ha6VDRTWxwU4cm2SdY+OQfq1TwgkLtY5XKEqG4xmhrPsow
KZtffq33paiDGH7Y4iSskay6NZbeyrqZiPgdqMd2Kuin/dEPmgvUaCsoZ1sSMj2poCAZNy4OlG7k
yaBrdR/c6gOt/mXPXHrrdhmIzZt5B0AkeeiNUlZr181GMQDrCI62A3CTimjnj/et53IMDbE3sHRe
B/UrbrpAhmjMs3maBUnYgFXBnukzwrLdgI0/BtCE5edWFxmPBEfqsVDEP4VCgZ0OhdkeUnCUnZPX
v4zsH69Uq2WZYU1tg5JoABj/FnK215Z1HUl/wsy6HcuquOxwmD96CT9d2ZGdww8y8b8FfXthafCB
NlC4AeSmoKN5kJl866nb0EJtrwNQ6a9JAJI+ESAupUKguIZePzbsS0dw4CQAWItE6lIhNQeENa18
2a759ynD6gZVEov3JUa3WXRoisA0p9HV55a4Omc91kIU+GNOeX5flnf8P6b4X1HfWwABxBi8WvAN
nwv9uUUjsiotKK+4UO4pfJhB66Hed6fLJrFJ1MVGqRcD8jTVgnZBE1cVw4iQl9+EfZ3rWMkvjzZQ
mEbkp9x2ppbo2cFs4bDXhO86LvpGYVTeRbmB/MHsDNQ0GNOnKfeKNKQcuPQO1NHXzP+t52eV28S6
ev19ED8f3W76zjtt3uUGEm6syDqTdlspp1ILxUSgboeUPgv0X3cxby19kY8pFapicHG/ASswRokU
H0jtEG9I5Og3tbJ490L+mahDt4w1wCIDikQjNmiTmMnZpRWdLBYcGpkyGpdurRDUSC0CG3OxQlch
cEt0DcTpDFbVRP/at1vHmOth1sE+KCjhgsGXhkwBNAaOJ50n/H8IxHg9zZKezYdePGUnhIBPMl/a
L+Hp/QlkyIj4aUtDC+l7EgWRxfzH/ErkjJwplOBmuiUnFpQsnhKRxiU7HTo+yjD7DMCQnjEEEGkA
S43SNgUh33/sW6h/X/chGs/4MQEp93RdJct+ZIpr86rm+i9pF6yCC7tHwGMr6PUwyAw4btVajyPZ
ndo+u1lVAVmX3ijnQIZg4Sz83o1EwhCmMSQw6fgzpd74zRLbZJFiSV10lh02U7v7BLVX/htoTm1J
yGXctyEDIT//f3bOpr8WIfXq6e0BDm9xHzP/NYYzdyUtXqVfNfD37ZKZqKjQBj9raoYCHn1x1cnx
q7BE0T+s38w/uxzMrPzYS5CtzObq4HSoWF6bP9t3v09oTKs7v6+YEzKexRZeQnxRNMtSZYRRzWna
dn+44xueswvQ7i6oO49UE858HabFX7EABMXFTStJYd6M1aDTwNPyPPn5oIlJO/7cCGWg7X2SNouD
5rOMHRewWukE/FcJ9sdQeFXUgSkM/bc0E80flzHkHXS4etUzzNOjjrCM1w35iednakTIR3h97vOq
2/38cwH49S0yYhpa8pkrgirSzHYuRr6MDM+tSzDbbbWrpTtxely8TRlhUDzk2jhw3oNrc/2crplO
nFjzLB1jPjXN+62CJMkQPCc3X2OrCSfb1Uz8w6qmeguGLjVbkLsg/4KnfxHDuGLAEqqda009r9ya
UcBS/UlaqD+ErmaEeCHJV4uIGFjjPqPuWc0/RVZKUbEgE4ritVcJ1auXG6PovzJR6QhMc2FL2lta
AiDOqeILm+YPJoL3GJyyjrB4JfvXBUYMgdY/fS8ayOsd+Gm4le9y6xEPsmuTRGKaFEDbS1+h4dnW
dmn+4VPtNBKBT4ZYvyA1nJ4SFfpx75tU+uMiXVSVMgQ6YnZ5ttgCvz08a7pX8QNw++5INNq1inJY
PDsGnLycVmtfZT2EKK8tq3vAAjWgqiPeOO2QigtC9m8ZaAYhtWT//Amd1bhlmQq8ZoS/UsUVucOv
QpljKqXWzLMJ7xH6pJrjYfBcdwvxeHCyIHK4OTdk7zVJ8bkgdJz0mduGx4MJaCpRZo/DN6Uspv5B
3kR2XuARMqIBjjwnwzPVl/pTh5lHxHRpT7Hz4lwbPZAjHUGPJGUauevmH76o5wYSk1Rn72PEv8Pm
1FyEOImuDOuqUcsWTj5HPzN6vY0HHtRuYZej6/miU3dbMmXwrMw5Lci38lDavvsmR3cqQKAvAl+k
2y0jvZ9XPP9tGkfJc6TkmFB8znCsd0L9oHnVLFENKTYSpeyGRbj2uRoVXrFKVvHnHfsvuBdFxwpZ
lvpLN3FCErcNYgdLYuKkFg8zbhSU26DADWJXL9eX4JhO5Hjtm2eUKUnGLNF43f0POYTox7zIUj5c
Bd+zDWo14sWNC6fIY2b4DssOwEYWCEvxqy8bBw0GxXS/yTFo547ZkXGWroMyKr+VJWWxQyXkbSbi
/2eDocXoF/FVhiQzuxSCOcBBBUpCqKK96Xj1v8ljcqtiVce8H+xYzhO5dVZWvkelH9+bFK5MH0ts
or0MwoMuz5DCxXDPQka4hJ3hJ/MKjy1OdwlDcyVCqtaWI/Sg4/CA6LHw3uLsyn02fkLl3orct/g3
2qGJIxIH+8pqccTJj5iw4MRn3Cdn0rXJbzvgOtEukRGSMNNDG3d9pMGvnJPu9VZl1Zl9kfnzD8ve
iH5yyZJ1GFFT1Gvd7jlEwQORONKeU7Fip9WFFQZF/AfwrjM+qr+3zTT1sDEFOKMkhr1BZKYT22qp
DqVY+z2/zXlMdQNq3rF0CADgjs1dIOjnH/TOfTTINfAl9W5kSQdr51EiUbnDp5W7wnUrUmIitbGk
vwUrG2+HVr6TarJJT1wM6T/U6I5bm52kZVs21YhIje7dHKq2VbKbABeLNLPRKkMiffi/2ejCSowJ
tIAFVDmlcSP0kRUME9aYU03LgURjFHvKEljBwuLk3uEh+rdsO6RDrbdMYdJ2I6LC1LroY9hm1Syp
78WgtG5TlY3fH+agsvz10p+0ZYFyD4MV1cyAdPidGJuba7hEgk2QcPZqnJ1W7HrRe0VB9Bhchm7E
0Gq4CrX9UTq9/wMl+/8a0vl1tfxxEZuTP/1RUE3FqZjBSueL6CcgbCod3xO/fYydvrfgzujb05lS
DVnckX2BtVnzIrYzXzSMC8zH6R7TUWuf9M5eTQROmGM46CwoNKAUWExxayoChGINWSrTmkz4d2fi
0joJPTUmSjAG4zIgo4p9wzDK0lQbXexdgBYwG9YBDVR8SS/+m2J+CBEPlguiAz38X3YTqLHUrS2C
c19a/ZB88lK2rbL2hBeBjyFkIrOER2XCzB2S0JNIZYgvNvuzLnEo/Hd3v6SieCPVzV+A03R/75PK
1pTSnAZP5ar3v4xeuvyqcdlJnPaT1rsoyk2SE6Ixpm5NXTcmAxA8P1n5a6ptxKuEoBLPN39KTu0Y
2YsMOPkY368xsVplA19iXl1MmF+4UV7PxiS7wn0D+KjVisk8E/JhFgcE/d5yzMEqq05bR7w42EkE
88O7iASLubX/LMDberMT5PL+YigV/FZRniamKaoYPvB9Wiim2Dah0H1MrmtGiEf1OrTLXOUqQJ4P
gwlLzTPVfBIIz8KJTJvyoToWfCynswu3L2efVw4JRopFOEOh/CzTfb1ft1BTCcH0G8PCOO9gZtnB
kpZhMXJe5xg8oq/lhyeWmBpcMQMCzOjsnANPBuzCmxyWP6h+F08buCkwYVb8iy3b+e6Gk2+5KKmn
bt+tK4JTmRWQ8Zf1CRL/8jb+hHGWTS99pG6539QFvpCDeJ0u4UTwD5qNegbMg/cHYJ+VUx6Ifi87
pZAUACtgwcnh44UNAIgQPwA5hwlh31OoFF2G+gnD6UIetcdMmuLxZqPszrBavqSDJiVT5kb1c6YF
ws/FeQOZ9jI6ntbmgNFkQaFKi5bK00MywX5DM8cxDHnmAx7HHEuX44Z5gn+AMmbfpK+gM2sKfdZ+
LsstmqckN+fQN9qls4ZigjtIdU6xRuhh2Gu0YvFn1LMp6ZiwSJJ4EaLW9KMWNfGktyIDT3jkzeMR
n4ld01pQSI3Kpqak1yjCcKEn5CB785dbsOBTxXC0sbjHV+/ny3eOlLGqbwQwMEDmd28r39cSofn+
fYro5gDQ2qdYQ3cw5mFlBfdOLt/y/kc/uZqnEcZT1RCG32WPDtaLPtWKg6s6q+OGKZpkraHKSNi9
6ho4RsrC/6bvo3oND9OdCm4IX1PThzt6VK8knwG/zoJRlpuupp0fRHQvYqsECbskTGWk/zThWxFU
OhD/8kiTQJraDFseSRn+heeAkNU5UTHtWSfyh7qZ+g2dLjn/Zs1ZUOnAxvmZlJPf5FKdBWpEvMbR
bNKbPdZxmK1t/KphHvAwbCLzOhLtmZof8GM8uwYB+x4cjf8RwAedPlopQxVdjJhYUBOE29fKceEE
tONzgH9gRzQ+/1sRocGY1j1PXf2KFejllbVOpDSTpubgZJttCXUlRtnY+IDKh/s/PgNlLKnrSdhL
8tqaLjkofgbasaZqIv8vTkXs28ys5jTDqf+WDP0zbkYzPeJZ8+bk0KnVaTpcg06X/X9VzVIPh6EK
VFWMJ5WL2v/CCVLG77eoB2S9QZ3Yzocih0dt9qAsJiPJSwphGB31f19W4eL+hy8DIcyyl7IYzkyB
IDewBZtrDBRHcQSU1rX9aaHDDkpVAVDikkA8p9rvOPx6JlnFd9dhdn4cyvBe6QRX7YEoehIcT7zR
4RiZm2+CzdQw/ybj0cBXeWT0q3hIN7zo9nzhPnXWYwxXNZOjlqhBrUgIScP+u70rINXNITo0rGfG
fCzBUhDyf0ypWssZDqbBaiqshgjRh0pVRTQx2TF55NTF44rT2eHqYppbil2ecQoUaz0IZmFxv7x3
XGkmMLM94WwnKCbk2vWbY3WhdkTyZMs5oE+XKb3b82LtgKkAzOW6Xlh1J56QehtCO30OdfCC0Tk5
ordhCoAd7ZgUXnd7ME6OPAnNouAk8N8Ghs7AvGYxqOyu/GvIit4Vuy8uBzkgeoqLmq9usfX859pi
9hTCYavy5zC3eCghNImzuqcexWTVcVVL+dPJPUD8xJMOf2mcF7uzqJzf1Lecvw6wsBD3ElcgJV0R
hP1wLNjeDZeUxsfFupb48ctoA4zXxDdgpl/ZKhFLxOXG1iMb+ch/odcuh4Sifx3gpUj7hA1nqyc5
lTsybpJhqK6oakPOEayt5oxdU31D+xwuohhsFQNb1Jq2yYINuM3yPNjfzddGXaaZEX1Zz7BzkWxv
ZsF6uP2Gr2x9kcBJZW9drlDO3TJE9zgQWKos+/ePBWX17YPZvS5BhAzZpaR05PqS90OXtEAH38wW
8YRyN+XF/uTzfyCNxySp2osmfdpWbt74zlPz9yk+nNbKH/BYxpR1GzQTnJ0+EF3GE4QDoIGvYf0J
ujLpHPt4PXoo/dQLD7bew+zL7QPKrHVLnez8TyysvCBtt5quHLRWnian1r6S3HcNgagfrRU4wrhB
bBFUctRbTBFYmFhJ0PnrGmfyNJPw6rCJafREEDrAAR/TtbRTxKo62ghL+5vX7OZa8a2rqSDLcZry
6lvd9TTGlGQfpCU1QcNIiiT8AFw86oe1Aci9AgUJ/VhBnTkegddq93HXHNgNo1XsFud3Bpz/hZ8j
bUk0sR6GysIie75TO9W7ygxhz2v+E9iWkTxGI+jLdrpZ/3eAIDx7EOeqzRUjTQEcSYlNpimIRj85
6Tz2kMpurlXXLFPJmx+IcXQeoUeKSjUr3e4j7UP0t7lsTSr1+tca7UAelSdPsUNNDLy2VIPdpyPl
QzOU3JHVjA6I1sC5ke5s25vR/HBrcrrZMOtfvLp7E4kjPhOjDr5MshZ6YY6yPuO6MYS8X8MCAGvN
oJKHwckbI1JsXsqiDEjTAnN8L8GTaqS+Sol0Kzn9U29uapAAJG+CS8qO6G3yCetnHaUG4E/G5uRo
O3YxCQs2VuxJdqSutTn/TZSLAITO9+LE2iwf7hyjPtZMiIAabUGq6ycUNv23L6gcXBXZsL8/RxfW
8lkGMLHUjbFOPd9KFpc/O5TK+wq30kcLIYVAIbDBIOQvJ7+N2V6EAGCwxklKZWYLx53YIoeJvOfh
6ZHmbnhi9W3QnbZzQ9Gv6QItqYOONJ5tKjlVo1H0OpPBi/XRpfG0fwHIvrl3P0D5d5rjt+fHM8QU
tWxwEHPel/thEfWoDXbskMk7RGmJQ84yus6FxbVcNWMKuwR2irzPiw1p9xu8dj58f4KZXCBaqN1Y
yubHSfAYfyiqyV8H2SQo8qZCMU2OzecP9qWjam5QpW9+sLrQwtV4riwSOSHWdYaxkis06w2BifiE
BRX2HidiI3hKVmATj83q0auj8dgCQm5RIiw266NfmtxFh9grT/NdeyPBOZOr+yc9r5+TaUionM/1
k0rIg6XL0gqNN7bq5OX5iPINttimsBth85xztTY912VvivbTbR8Y0/XZnRCxHRP01BPVjH47dY/l
sh9JkoYJ7t75v/w5blwEhY9QRJlgg9qc1K/zKQkoYw/0rpoPCqR2PU0zS6DZOpzkIr5U5spB6RV2
FyEFlN6KF29Zwa/YoOz9u68CRVd34GS0Aq6lHZxV6fOOE4MOjNAgbjn7T5NjfpQLfRAAigcdsHnL
RPXGhkCIfiVuEwUAl3d6hDM6n50ZVNnwAcH46cQLqq92IA2JTTOidl2d0K2aWA3e7zaG3AVyGJhF
RY8VHIEHzgy9zf1zlQjPy11amBIae8/nNZYNY3tkScWe7xj8nU6uXVNZhmK4q0YLatjk888y/4pj
UIDwuDtr3Ckci058HQeO1qHwy7hSzv4Sd6K9r4UIees3bn5Zd+cEqaiIcXj7ioT6le8ymXTykIZ6
gTGnQqoC5MGKXtdAbbewxM+sP+iT7sgcn/UkAEOcLxhFFJt0JD4sNs7YEuI+BGR1e759vxS14QWN
NNfS6bOegMrgrYyh2Cz+wSsyAilyjzeWDQods4QcMegRsVT/qJfBuPPO4OTMBGqhjlRnm/FHHolM
uZd1Uogo+7bUYtlgx1k+Njz9YyVS/oIhTt6zLm0cureSnqDBdF9G+663zG5csEqiJC1hBRlQtO/w
Mg/SGAbX36v6cboEeZtXsRV3BawRo9zGg2LB2LDB/dquCxMCEjVVjb9pRo+nuF8Yk8jB+dqn12C7
znbZKt+SA5hdLuLHnA9aw63kZJt58XYI04/xvdV4/XrfjvqkQak0t9oKXfWfUCFf4smp8aGexW1P
9z0lGlLgAphMuLmo+1y90GraLwBzwIdHaaY/ySgEzhRTxwlzMxmLipNse30jgYsoPqk1Pys+YXYl
F5hDnmFNC2ActFlkDI4LAd11iHxbBxuQ1ze8U78xKHl3Slf6uKCy4wE8AgHOf/SeKCO2YNgbCkur
kkwD5D6QCvaep/figBPlygWUjm5VRYnkMhcMvsH/Kmx81PKgWvpmvHM+6vs6vX/95AISadRswDW/
1pajHtL5/AV50jA80HwnlHgZYJ8lRdu9C+3fIun/J7+Co6+iu532X6Rg4km3c9ZQa8T87X6qsaLP
3ztGLzVUCpdVo3qpENr+hVsz1YfiGjexROE8u1gcZUWqn48Z7Jlcxro471aDyEWpuK6l+3hT0Ejp
wf6joHcRVYESuNZm4hqhXBtbbOVnN0MveWCUnSpAKlRmPdn7/m8L0CzNR7uBn0PCJmvhQDkEK/OK
TiQoC8nDuDBJnNFfZzBfl7C7/+ZsZXvnKxefDLij0G4zIzDNcmJnk6+7Id3rKQNV6xq8Nr24ON0o
BqYndSucfGVezS/2Ci3YLnABPDqLGX3nkwMyt9PGNR6VbmFnrn+WNtI+9vf29ERKHiman0yoRj6C
Qcm+JKtZkxZg0IuAO+0zyqSRf65l4F0gzQYWnmJmSI2RStWRkbdj4Ao0UBeOgACIb41uJt3TybhF
0zrZW94ANXe5n5nd6wz4dotuDY+vW6FcM6edAYmz9E/TwnKvGWaUJ644ghu1NCWiEK7rPyTvhhPg
GwDgilp1UWP9EVLOl0JX5tHKAdzyvy8vEiSHH8N1qKNqO+i+fRlj68XQ22alkCo8IG6gEBZiMAWO
h7D0IaLlOC7m6bH9zv65VKHyPp5aRRJd6hPoRhN6fyUZV+4h/LCzBGA57td8nfeXc/4YDGLlIozp
rRbc/bJ/y/8lGARx8PmBf/J8/4rVHkKlktXEeSxMHzoR/kJKFG86xRLFMhUZ9BPtnKN2o5IwVUYc
eQiyLJwqD68VnHbw2drp/y2rf1Thnx5bmPgHL1t4sfiVBBzbbitQcEpvHMlrx8G7LlUCfJFmVUm0
FsIgANBRdcL91DCgsoJDqPNr9laWNF0QWiFyTiqQcJRb4x0ECY+zWVrdEWjkKemh0XG3jDhP4FKC
IsSoGSs/5DQ2bJMHIiG6qWk0byN4k5Z1KfBgEsaYpxkl+i3LU1uLQC4y5nz9sT8hZajWy5M4MqDu
yxm7R843q/SoteylolxQiQABZqQsX4yApkHR/8JSe5vq6HkRTOIN2GGPW/GwqRQHnHTDpea5PwWt
5kbXj9Uy0Xo/40i6S+kPOPtJB4xECA2XsDPtjhfG8vy7JXhVJDcjcB59xQIs890nwl+YOs5190In
4qFAxUSi5A4HQpXehMOApnfGGkSZtzqqTK6YIU0NJ8OuBGBKOVkLZsh0viPIRc3oRnNiVGIzECZi
tnHNR/UggT0j+uQsFgItpMaCwrhOKAimqjMx8v7SCWaZKe+cyS8Hl6VuT/mcifgYConmIbTrPUYq
vL1OtnjygiRUNHYX3rx3Nbe6ZSDd2Z1QoVdBeqglic1Y9qtZa0g2oZE+kr/gP0qyywqlJx0eVdkU
VMJZw/KfZ1EVS+s3Ut9gbiINlk6+iqN/3Bgi1uqDYZOL8WzLjUPwUYBFOnL3MdOT1UK3IDnbULFO
VYUZVwVCnwOqr8xT6meRfGy9FkIzSlQY7HIheJEajSwEkS3qIvhagF4LVvAkJgqObXqEWPeoz5im
2N5a1XS6P3+Hh49ufMkCnybcJ4m70ssyTxM5Nhn2NI8WhX94qqoN+Z9C/wg6luOIuMnb7FiBdOqx
hIo9bQvshV9Rw8atCs0p4UyrzmYNMHSKkM+32sJieJGdgGWBq45gaYmAsVbu4IDfTBsNFWGHneSk
taLtCRKgIIzTywgSF+NR/H2Xbp+SarinK8JMU5QSrBv798L1WcVtzRlnjMpIZ6blxll0X6JvS7gP
qyciER+FyOrw/Eigykba8illLDaU7f8KXpy1DJ0oH/omrV/Fh4gUtLvDQaVwzsiLeNU07sZ9RhPz
jHuLS+daNk1jwmJWLuKKrjkni9/WhHT3fFz4XeRMC8QKhsIfyfqDk3l3wnrr44YZULNv6m56dad0
m9rSV9mLUOoYL5HSsX3loorS1bd+Fz/WHhvim4c+OwdxRbhExivJLZOne03A7ApcuWrO02z97jim
5UPI3Z7pQ0LuT4CyLE2tK5KG5PIFsV7sNLw24ofouLlm8PP4NiqJBnIR0doK4pVe6seMToWXy8zm
Li8TisrOknhVcUWMY0Esg+jPGWpswyT2ADkf0GbJ68VvpUUJfqgykxQWeNQ9jNszvQvmETcxNkrv
JZZRYIQA7KEQ489+peQCWYOAu797JXETTkL9xFddtPAV0q2ykMPsctrUoGTDzefCi2Y7zoIFY6vZ
4h9xzvohYD3amWzNQpSFThGymNN9xBWYSto96BSojzHzqN6+3Gd+6yxSwUuaCHVGmfrTWkU4eOct
kJWwvPSRih1GHOIH60ALq1w+iC4FvVjC/5v1vTeafeBBRdCZSV0Xe3zHcclZ2uE/wohYCSu6OlHH
jsT9KuvxMhGXZaxQ0F4wFiAlY0KHL86KyqCq57IsAbDm/hnzN0L2c1Ia53lSAKKRZZO3mqNmx0lj
LKZ8Wr2Dhzcb+sB/LpEU+VlL95NB+WH2rsqgAnbPtFAHM4oA6ViNy0I1xZ8UAKlClSWj6sKR5ATB
KAAETHHN4HdOo66961ScP9nCv8MQdIL37jGVOe9gvZ9tDx9l0SgLNP+amsBrJB/E2LnXpZZfz+Sc
HFqse8x6PUVWasGCr2jLiH6jKeXQCmrfDWPkr87XN5ikTCQFMbW3zdPgRieu0lSsT/zs3Lrud1KP
P7e/gTehuVVXHXgm6t2zjIW+MNuvRdvz4bD/QzFfk1aRBzzyFFBaO71/8HqVAr4Rp7QH93hRHooy
qMlyCkFlRXjuAqXjb6KQy/2RReO+Xb9Uesm0lAwTlxQiRedXmJ4W/0ot+ZZ64lDoX0GO9GBwsFFF
le3VzjVIfhb9RpN91HAr2FmWe3tpr0+RapxAfaUBbjkFQAhavepdfYJ8fv0JrJ2J3HD2J15DBnYx
qVBX1dsrUxTx0TtChHYEAtOzcMQhkMrq5qUdJx13T7DwklQohVN0/fvWqL6Y7P1kTUc0K+7thxtq
m+iK9ZcwAcIxPR35kR2Nci0FUCJdcdDbvGzStLNoxYb74CwHfTVV2VYa9+x4be+TI9fDzYNqlslz
OwIEArZsnbEwKCzSj5JEuCw6+hvqEXg+zsRx3iLk89ACBde969EGSJ+4NKZKALgi9rGeqgLJPtEL
NNf85tTv3m4WSHfb34bdBAhvqwHgppZMHG0UTg7+fUe+6kmbhjVZ8PEWbUXWvTNV80G9esgVsqoa
fAB9q9YleaiiOfbh0OcQLvVlVhbeRMzKzLLFQTqNyHhVPmrP3Vf+AVuaPPXMMDGKGbcWhwQAjg/L
j19BoCiDH/N64VqyVLYKp9Rue01hSv68CCxO8snG4KtT2Qe/RDA++as1Zp1E/NzGzgYDDHMqIFhT
kOnruxyGy9g7LH3L0IRFi6ZfaJGjFtQhY5ePHIbs1kRcvZKdoUW6iINTG8Hz63enfiUeNu112b/z
Y4v96c6Fddsd9ohagHL2DjktmzBCHQy7gUOBvceeUfPSi4hj+stDp4iz68gbq81l9IXdsmZcjheN
5QuntHiMFJZAGyysR0GnZ663pj+uf+/heBCblCY3cRYTNKcFuxMzFjtv4LGqt47bSw1J9F91BV0S
yypd7sJI+zVFuiCnB2sKQhqqhShY1GKDVPvfIKs5952VPvp/UFMWLjR50y7iv3CKe/TTqdc7CW0a
IQ/UD1m7RvzLCleqxnc1uVQc/V1fvH08bRw0g28WnH18IdFJNhr62EstS7qRB6NCj4dcBSTlPdeM
4NS9jJO0+4fe3ySqr3q0WkXXIfw2Nxs0KSoGkrHUQa9XEfBzs94prLg39Gtz96lYg3T0s0GmhP3V
5Up6y45/4dOc5IN96ZFE0uaXzkfVsseOLs/VzMc2m6dgvKVg5oP+1IxXd6dfBRwUwqjr3aHBpyC7
Z6byVl7ghdzte11gjX6RoxydSBFO/lnQYtyDXQDlLcOqnwwMh0sHQdChnM5ucQ0T8wyihPC5phD3
QqOaYDxOxlu05FmSG0a3u2V4B2ZCBTGOpJ91BAmELDVq8SX3NrS06My3L/eZi5G+qU7LcuP7N//o
Wgjeb2J4aKXsVRI4bZfgEVY9sYF9W7hi39Kti3FovTJdLbyGAHaYSI60Aha4vUqKfJDK8W1FrFW8
6KWB6HMtBmS3TfpTwxS3Qoo5eeoFwKRH2trXRIMHhstr/Hoig5X1EG5xcvD8oVGmjxI113tkUoAa
zy2WRbm6/VfnPCAMq+fX47ie5m3BcTVuE5nq2hQLBCJDqT4Ol6H3L9kPy0TnsP7LmzhUsGDkXQlU
P7m5bL+prRB4UQhyXo40vQZUiRm+6ZpuTV7Xg/KLNFFEcVTg7bSsD/jHF0nk+DfA/uGtuxqBSD33
77Un7c9MS3UipRdtE7lSEOt1j8477XwzH9EJ+nTo1dJ/gVY4kZKkVA+JnMhunt0Pc5thAAFX7j0+
6MDbP/K77D3dZV4+TXZtL6WrFXVaNoOXVKhSRL3SBLADBHyCwzJg8NA31hRdh0nPqfWT2RQo/E47
UJBWeHy1ivlMYBmDZxi3svG1SCimidl2RUfTCgUCjhHGldMfXqk8UxgBwpLAfruofnpV1JEmVFaQ
3HkV1MI0z2kfjhmztd52l5Y0QPM+Y1FoTPiy68Sgc01YoMX6b3Rnhk2b5ll6srin88o5RWdhWVH3
YzgDfcR3NU/VkvHmuV/CgAG1BtIeqSO++n4o63ZxzVXnJ1JvRX6wyiVvEXRnkyg2NVtKlFoa+51C
k8EYVKg5NiMv+0sQ5zzOiMtxic9LzbawUkehpt8pHTM21r2Z3uxFit0wmOgr6YCx8vCxOV5rRRx/
AkiBCYI9fWWOC0YIoguwBcKc/cyIj1k61bvTBYg6MBIkRv2oKdTgixbiUmZMFW0h6cnprPG0kGnc
2WPQhmzTXFQUdlteu2GRa0DXoSefID9+kEMGI9BePAD90Cy8JikethduxNONF6te3ox4Bdqw5X65
zTutZ1UMhZl2C/vSfbPHcigkkk3MhZQC5GCHlJsDH87luU0CCBJt/6cDp86yblxNaXRPriJ3gcpM
Bgcv6vVpgl6bjvDzH3kuRt/ocXYkwhXzvKc7i2KuPfGHSrBi4tPGX1SsAlwLADhji2PCE+u4vfh5
79qUQZ4H77Qu5l9+mGm4PMtlBUXxtyCjsXTvD95eofP8s5XGnL4GbEWliJZhYyez5GokElAEbipv
0F+Z5b0R97mPvVY4VXspCoL8TX3aJ69xTpY8ZkcZQsHFXFr1zv9RxwMnkglA73KIitNR0P7EFaGE
77Z7B4iU76T+A78x2iY7w2SW9cjJT3Z/wq9u20znrgT6+3XtZ3H0adRKsqmfoG7UeF3f49CHFB7c
nS2c9B6Xac729bOGN4RMF1hJo/i5oct1hVNpwFI0IL187/sFrmfXFzmJgCJkAwKn2PK/hDkSyoCd
oGlj/6Z9CTbGPtUbsYjONw2B39eh6rAa6o2i+rr/zWOYR+wuxe908zfdkmwKdhk9bKJmeg06jeNz
gH+DxSDsMZf2qLzE4u+Vcqg637mxBs2EPFzLl4MQ0hSRhosvsowFlZieGLUZcN8i87h+F1qbUb/g
Bs4Sh3bLBPrFu+TZA9ZKYK406F3nIhyW05e858b2q0nJMGRbdwkkJz+cc52bMIlamxle1Qcsky4S
h7WO8VQdCYMxjGHDcQJ+6qdoxePm3U4vVoyoyxxvEIY+AcKL2+BjAoNhWE0rC+e88xf6+CBDdNA/
JbXXl2j0L80OZFli/7GyEPtXEd0009qxH95Hhd4/aAJp0AfX0/txx67WwsJQ5ad4DgSA8o7obFd7
SkqvGdqHpW4DKf+QTIkvmG83O394IIypMGa9E/vf8cMtFbqAlgz1yaG5c/6e9X1rfVeB44cOnIdw
kZ9oYC4jQ06pKznDMoxqBjKQqKwuo5BbFndhHITGFm/5G/vY/Snj0mc3nJDwsgxhvwBoKR2Qyz89
DRMFjd9JAymYTbmr9AgNTuEOhpExg+v4dF+lQIaWWcNgHgO/BAxv/BlPBrAShUnzLKbyUfNlUdNW
cx1tvKlVBx+nMlhCSQaxaq+8YG0HdvzchFybaHkKI75XRgRIJltjRcdE/mZkNfYP7/IEwX+FtPzi
R8NT9ESSkKSH2lpCLxKcHsfKLcopGyXZgKGNcsJ3qHOj9rPFm3zCIxB6t63pN27TUiLdELmi4AFg
eWvIddLYQDtPzNm3+EEoqRyE37lESrXtVzHLsQwIFBP3DmC42WyYm3qInhHQS49gQkK8cQFfD8vH
7A7FYY0d9il/fztIAbbOCATkZDR0VDTiB5TA+zn5BId8HW4zXMA/a3cx9VFmavxdDDbWKK1qYMMT
SDs2Q1eVXGnr+1ozCq7opLjKq+Zrl/i4UeCmvg8Rl5b+0w8MrqTNtoIs2OStDAHntNHDQzwun4c+
XAU0i64JP/jXcSntyfAQXMqJZVGuAoAbJr3isQxvY/20yS06fRkubZ4Po6PJgAf3K1r8rbIZFBdu
/y+ghz+tmotwnA5kWPXlbipqaz1EZDbo2XA1MtgZXn5ScrWIeOWKQVcaOW3+ppXjPVsYxeFfDIK1
WevKrxkAIM+ZPlrAJ1h9FmPkPO2rs7UujjRrLdzhTHJpy+0fn1bInkSEfxAqfqDgRA1cX7U7aDwR
vQebGQxQWkmxih2YNTgVhCW+z11EI9jXJzz4p8wveNLI9077Ziu+m+J/mc+m7pfxcZj85JqHztjJ
EAHeY8daSmLgUCkK8FJkcDoO8Z85L2NZcrQi2gd9rrOXfmhg2ixXn5DA2ir0PeQ8Jq25Wt5IyVGq
KaDN271f63Z5o5SCWdX3jct6TfOvKcfuzB5uBrPhz612BavgRhZqEPcpQltkYNZlhrdMYgUTspNi
IzMzJ8r7UIfVNMeFqB0zGOFXSR5AJo6zzin47a0TfI97eWXIwM0s+6PhkSbDQ07/QD/L+2FyRuGt
eSqNsZXOyeBv8FbqRHxLNOMghTUse9K+RHNFE97dyIuw0Npl2ZLXWSjtswSY0towV54qkpe8f2PW
rWKtOGnIGdpAcd/Ueuu3wMpo/jOMViJfEzYRixOLox8Jb6acgbaDv5L5Fyisg364VWwaSpsBElNo
3O+emHlsyCDMj1T4oMHzDKYa4uWPYrp8pYKCUS4AOBLeDNgl8yrKU4QqQZ7SogHej8tKq8lv0s/H
WKUy9yOnMwUM3Ys8Ve+/j2G97dnK7Nv65M1hLXnsiC688BbavY3uiQTSkZjo+WA5FToDqFvn961q
DU96fpXRxFZvNH8QH0GnxEtIlNc0cXwjR4phoXi4UsZMUEm+89VpdHpJ9EEJ0t1A9vTRGlV5Esvt
9MZLuwPBiu98Ku0nQ84Ma0668ujUY4PAjaWAYLeh1zoymX0VX5ZxhMZ6BX7+Qix+j6IhUckKRAB9
pFGP6eTxgChK55WMwm9NNEPwBitL3kbwJAQykB8jDyzKevN7yU/bBOn5GBERDWXAw4ji67hbWWCG
CGOxncEtpCO4UBEh/h421NYZQ/AQHVtF2ZsZLkC5QYhFsRgNuqWokNU1Dwpk2gorlzHGQmnOurzn
2EyMjW8McEdVgrfDWzZc2dVsU4+zSogbiBSIU5BYPqSlG9qcvhT/D8aAJPDtRiqZUqZnbWOcKS7A
U+AQZaz4V2lvHpZSsYdzAjdaJiBgnQl+jjfAQLrm8ufihv9HSLQtsKtha3KEMysu9oxV1dGBZxGW
mti7cJrf1vEw799ig5FqJzW+fCkne1wsq4oE+5OGjqCLwXU9o/67HXASdiNuECkDmf9vPvjZFXyy
msOi/l6O7VHoMo3vNGtHkBrRbbKBxDPHJgJckI9+X1kUclUA4czX94fYWF5cf7ntSuIeOlwIc1sT
lkLzYfvF48y20ghfnRTx6p2u/xipoAVJEIxwSm3DHNIfPM1pkYFkI5BPZCBsH7VMV0U6oHcNYWNd
eIFBIjNcIPougJOCL+o2dYAvTd3KM3jnu4l8Mhk9QdBaz85nDF+akD2KXQW9hg3Z1GYLJkVsxZ8Z
8ojcelZZjbMzFJQB3q/b32EikCGE+ilFwviNiZKJswXQXUW7edE1CS/TKoTBWUZPG0Kd2/g5QCeH
yjagftfgX69IRKtdHJQn6ZqVvMOSw9yNsVrNAXLJ/OxqTJdbr9zpw+zDUW3l2RG92ku5ITKHcSLM
Ro6hUaRyktT5QIw8a2XYtp4z0bC+0cKrUjTu6DI9lGAzLP+q08D36GZoknacf6KIL+tDhQGj58Ct
bmi64dzODLAMBPVopgKeeQWLzcBk5ns0mHg/nMTiJ2mvAMs7YYrXwCMs1SfdaPg5K8/I2vVzPWRF
cABo2hvBa/MfdV0jPFqYgSXRjlngmz5tTPQ8nCmwngay3Ebz06s7eAoH+RyZjRQrBwDxvbQx5d8b
XtixY+b6stej6loPL0PO7NMwEJ3F3+C45QulI4Xr3pU7aaj8aJ8sh3a/jQW9GSBoZrTCsFMuWEn6
BPscHwb8q4908S0Pitg604JEFfIJZcbdoTcyEaLoy9eP3jWws+E4vhCcV1mT0ItQQWQP6TTWIwOW
YmrgWvfrpOsTFu18VcbHJ4VGUpLmZI42UUKPwmtYnfh8Oc3Kh23VWctNOcTBJ6JZB8HxFNjrTAys
4oky5RRHLAtigY8hcRQLcQ6rUywdiwwmZBi6E5QDH/yx1HzG17ERw9L9yRatujn6I2YpEJNEH+O0
+fDXzITh+FOHuWBPx5N4EX7KmEaqfPSes7NLSQykJt7NaP+B94PZN6HzVQN1yjcV6sUR4gTy9haV
lu2lLSEKP2LZrpJgK4K99me/9P2tK50HxX/lUzImGlIJIChvwU/U1gb8nZ3sYfOTk/tuL7JROCmv
LfNIdTGbmmiMCW56djaKE4ceMEG7YmfSqnnlQtLFcmWcubLVCCVcBxECbB76afj2OKUsudi+IBHs
9EPTnqeaO0/1NYtxajYC+nxfqEkCezPu7Y180eqNvkpvZmZNxJaXA/iF8cLFIXhBAFOjNHtwNlaC
Y7dMx7rsF2DQoP/ObjYJUfxqq+UIEWZ9Du6+k72uCGrCzkzV0ae53Q+S3cXO2xabGaxAiI45ejSa
C6HR2npCcV7PhAuJeL9SVxWH3D3Z3ELZldG8/SaWnNvdFnfuAKIKuq9JNSwM+6Z4XaHRw0HnOfgT
7ut4dLEGKKexskruh+btuG+BQ/LmhGm0gtAuqGCahYTn8IJyvZngrFVwB3cHoLhHk2ztRcgE9K9H
ElJs2+4od4QXA8eJX0BapyIheYh0JKkkdLVgbX7Fym5BegqTXnBIcL+MgYwk/9DhS+mDcdwYEWOt
v6Akheid2wDc8rcUmBi9O4mLbYPYjEK2L2ZbO3GRZiTblKCCAIxFJcRo0GGUu7L2cdYduk6Ogz/4
6A+sD1sb5npwN0+EFz4P4ta6L+XY8TyKQh67Knm3EfLopqbNYg6Ro/5Pe5v28Gskj+W2iUNoVqPf
y1nYjxvINZsgVUcbk9uEMmO7Oy75NIP1zZfY20vz98fC5m/yXyhxzL/aYZd8EYCVl9XmXQmRENec
XUcjg2aG12H2vPokNPLIaFFcu8HUyDzc8fYzwCfsFYhKrgTnyyzPWApnZKyfpAf3EmQzIb77aT8C
rVj9s2n+uw5IObQaoNPM9mpsqsCji4u7M9TYa5YyKM3/ZKwUAnPd8ApyWhn6rvaAWi4kPhmlTAya
mRPKSct1c0fiCOaFohY+PRrewC9V7CQcsm70gmf+T8jDY65W8KGcGstqt+wfpyGWlUY5vrMG8DlZ
eqcu0nF4ZE4Sj4egEw3H9JV25MKbj4gTw0tKN7o1XYL6ZY5kPojxqv6/6EgsHBDcQivOXBAOBGK4
MLO6Akd+eTqJ/U5sKlf9H7oX3YY5dHNs3hs6m+44AI22wFx+hayuNqmlBQJ/zDUCJ6ueKuVRDyUu
cc51kH8Nje9N+8r2zATebFcoDwuLoRtNd7H4v9CV5WYU52wLXwD4V27vaV8ITCJKVg3Vwy+zsFDA
IVYbAd1a0kvGLrcLw4iRKVoS5e+Kt2G94o+FidzK14QhD1xpwUonnksayhHKI6g5oAm/+kq9Ly/k
rfb8Sd+H0yO9RlROdpwgZyyvM5mHCNy8OGoia3E6asbaKGrLEA0crD4/OywQs82PtkoSYLCDLGSR
jODnaNF2gvmNtsPezD9/StbM8wKMpHQpQunt1JsWOGgZcUbGQricPuNISSLp2xJLNAzliK8U377+
qWP61/N665vC2DAgvU8kUrIoJAYDtUPOTQlRXyLn+vjHV9sM6QWRqLBsw56m88g69f5QaQ26/8OL
6okKdppzJCyNBZvHGcMJYtHsc/n4h4+YxB2Pglt0jk10KJUd2LmjONIUvnaxrro7tpc110AQEWp4
g+z/gOSdSyYE4lqMBnVlqetMAHgThcaHZUWb/zJe1bsN/lye1QmOGCRch0Ji3x4HM0QfT1FGo5Ft
iIvRXk6kz3Ix8a8coLEU57utv75eaXrAnsJz5bd8tv69GqT75P2sQAOIZnlHhvE8oJIMRsn3ToL8
yvzF6zOHGt2xq0o1hagq1pLO3PL2qPMuOwbE+88o4VzngvvcI90MMqf5o1HWxvTzANUJ95cxGNCd
XvYU5p+I7eEjY1g3XQYgGAwSDxS32H7Czm7GkswENLDW9dyhpC5b3/aR2aL3Hsj87peRnc00Pb7z
HxziGGUeEtIqWsFAd75ikPa1hg141oMEBE62VSukQXlZn2cOwVZbus4v73+YczpwWt1VEF211TEd
sTO3PLq0qXP+xw71JsePsQl0jtecna3XNZKpDpRFdlpiHjIpJFrVUxw8aJnfIGwNo77+Mk0oSXC8
XeLIEdtZlCn91aHc6B4mA4uC5sDM00BQFQzw8p4Bq5hGx3i3+ZkdOd9ByG35mLaZ5I+LSLn9jbjK
qc9Nge4bfdbnGWNFfjHyWeAfiGtNqOYFwRsi0MSHVvo5TIjKi8/W3bjO9uWaz8YHefnCK8yoUMU5
alT9gkjskfGiotXFFPs/DQDHuwec4YuMIMImlI5B7IReADfZFuf9aXshnJ6JboyIeWWNHSGaTt3d
aICdjYtWOZJBjLL6AbeXygd9wNY7gjeavpk8BltJcRCBdtb8NGmoZJn+ipL5eviI2S3LWAUeO6uh
DJ7u05tl+UuxnEFuxt606+YdobDfYQgFXUCPOk2WrEDnTw5fQj1Lcn3kQsvQLKZSiTZ1D+1GS9ob
DFCNt0TC5ISTiHpTJDu5TgB8OjbNwDEiWe/U1cTRQp2HbkX55EXB+KiOz871d5jBo9h2DH93aOGr
o7eh48sg7NlMWcBn4UQZHHcVt4aHahyVo8WYopbH2JihVAHB89WJpTiOxlOg5xtWMIuB4+SgAalO
hhUSp8nICOnHW5c4oVfWXeSf8dH1kIfqMo6ZIOeBiIak3Xj+iohDzAiAq15BU9aT5CWHysKC04G7
PBYBS5Ow74XGLgVXtmRF+j/jRfEFH64OAIwBIVX3KIMgeHjm8X8Sx9eifbrzslWvKHGXU6sFJyGw
kRTSQEQ0p+YF2hXcDu5BDThXKaBDLV96HYIcohC0EUBGq6bZu+Iku9CYkU4LQ69MSNwP+hWT7mMh
u678TDJBv3cExxmuahgyIbtlXDAFBY8NT6dT0yRQFZodFpE/al5+SKf/QqCZPVmIznWWHZtUTCsn
R+a2rwn7Xcx19K1klrnu5MEV4nC50FYnQza96Z+ulW2oINTepHmZlURr4DN4RizyZtT0fkB/DhoA
jbxUXnEk4yxDATzoOGsmRR/gcBpAwqwQVyvbFpfCMfL5eDee2rZpgGQtaGNNX8Z8oVASmAwPm+tT
Ud3oNM5Sl5qWfM4o8hMaerX8QpTnCv3BYcO3R6SyAxi/bn869EtHUz9m/MOtOaZX55MZBtCQ5vnL
whXhequhNkmohWtq+UvpTP3KfxhFm5ReO8/ukJCDaQtmArTRy8BHZjiPvY+1+noYyNPEpwInh/Tf
jdW3UISrauwtS4AacbSVV7eOnIfUvnlFx2xQQHUv61D0uagGjdAjvkfMpNyQPiXk6cvxdqcMe3z5
XOfGuorD2aD+lZeZW+AO+jEdqi3mGCDmAKX7X5WE8WzwiEizIQoE+f6XOZw1CLG7OxKyYcx1DiI5
VR6zVLzr6iI84LSJUOt0N5yZ7uMX3xLkRytJTy3Svj0SqCecNqOqiS3Q9RbWEuwKJR3OShFsU73x
Y34/3Kk6/LuTVmHQnRa1oFKgbk+aVu/dBZ5k31jl/habSOH0SQKe/T5gJgvcxAhOVeAQwv44ERGC
INDzdjxzPN2k6DqbNsjUgeEz2n1VpPTEy7271uOGn4PWoWzaq+uA+zlV6SCmQFrIzkTzQGXxZ+s4
esIhI83UVxMTcVsdA+i9e3wlQN5yF35cbGSvaMixtrz/E27C2o/DYh36w7GQ9Bmjj9+/ZcQDKgda
sE2BpDQZGP8fejFpae0SyfnwSV4hxQu057FqAjU/viSna9LKGStpp7hm5a5SlbREbH36Iqu+1YSz
YFuqYjFUjbZQUEN8rfYvp+eNdT1YPNiD0lqmcqf1ONYg9EQ347bkdGTuvxWSqmJ4xBtLC+bQAIKD
L9hEv9HUkIpwmKoOdsVHrrDigDHhamkt1BLpSPm8KwE4StVcK3qT/Vk1E1OYTOBHj4kQORT4Lqci
9vlgzKkpTkfqHW6d+5x/yKSaF7iWNFscAlMjOY/Oo+ta+ba6kEDHhh8H4r6qb3hjMPMrMqkD/ODw
PEJeKqNiyMpgWXx8JoOZ7njCmCty3IEz56yYP/4h3nYH+4kwCAdj8k+mmnlC/0OXVTS4QMlx7i5T
j8ISZ1VRTRGrB441bw2L+ErHWaTID4SiuWDPzDzeZdmtWlPzUW4ojlJ7nUSQ1lIUAo8FMo6Cqa0c
NPpJNo41B4kYEsMm6+c8t4jmBWjA0+h8Iei7+EZr9EmSRTwWS5uHd3/fMn4I6vqo6R6UyztGV2m+
yOxKcP1EXe14gpm5ydSDOZmNy5SEm4S6UIwpYg95NSFPIIAGrEjjCaBfmB97JPPOVEbbKaJYF6lr
oY6LcAulxvGoUKRw845nHkUtr4/5jiBGXgNKQZ4yBxqO2hhREe2Yf9S86ipx0D18viwIiWtCNhgH
+t+KhyON+fLrqckYEgzwWcTbNOLt8JJzHa7gicUGRE7hL2JvYAQXblDk2uA393pU2yLZnC/6OZc5
0uxgJyxUd41HUUbI0zu20nOlwvKO9nE3lrXHaCVNJr1I/EYuS4W99KC8CvIu9pevpYGQtxPK9V5m
m1jk1Z4Q6RwExq83A1YNIZQ+fdg61dv4ybSkipFgWW2FSdD8xcUcsLby3PEI5R0V56bE6v+eGpk1
KRs5884sdfKr+emi7OaUGi+z9oCODVjnThEmzq3aiID1+B3En1I7zFgYXMx46R1H4mWi9aNlColY
/uqX2osxVtfcvRA/aS6v7C+z6cf5KYWEiBTgTsTWXMws+xu7b891YmZ2M3AHdzlN6Xa0scY7MXW5
g6c3kt8JpMXuUeW6W/adrl8o16sn1D0TLG6FcqW6qlgYxkZ9am4utz6hwoOR4UCywNNNqgUrEnPU
11HedB8KKvwCDJToABc6tb5qN7Ioq9HjZvvupDEAaAxkRLaSgp8D03z73AtUkPSmc7TiUbUliv0l
jGxI6T+9KEpBlSBcGgyuyB3J+wH0QP60hWweMZ9/M4pWdu5ByX4PvA1618c+QVv8SKrZ2bIhwq78
uKS2bPz70UE3G4oeI/ZDoDLMsyJIla/+jDEJmXiUWvgtOKed/qqftkR2SK5AlEBvJDcz0KlFGdiG
yUoj6Pp1QeQUMisqKCahSdIjOWx5/gWylk/mSxhjHTLhN7ks1txvQija8wWgeeEBmR+2CUMQst3m
s8llDMnSqGtKGHR2DudzyeQp+aFHDe63osMVSK5rlbU4ZUjzDVldLJjMtduDqRDcw3/JWADfQ9GO
vn0615IDNdp8TZjisCDQk/WqC/Cvq43mvAyqLSv73HeqmmMb1Lf0jOT2q2eBiDBcGHjdpeCJrLHC
ne1n3WUEcmuSGRcXuVTwo7dZk/UljlGDbJjAymoDBE4tIJE6auByMotkCEdppkMZ7t9VTo3BesbE
Qjm18J/co8o8aeSlKhZGfa+MF59kKEWNSAR7UzCJywhWBNeFHfisyxACRnB3729UkRqVormUuzoj
MC08AKfnWN29y+gS1moAQrfUi5QahuyD5eGUrEJC4+iGgMbrGD3vvL2h7S9tEfCS3vbS9YUxTtb4
k29BU/7Ex7ZcEtNo4W0NFMW17U9JAl96Kri415F8nA7KIyVdFJvDQ1JPwD+n4JYMs49Ey1+AQNyR
FdJmk1QnAd06imoNvDKQlGgH+O3rRevBSPmvDbv5DGaFf28Jv8db+fX2MyXQU1h1ivLFf/8Lxyl4
vgMRJNL9BWJIkEywvViT+U4KxARslstgXot0FBbL0KauLZFfTz7sH8AxQRvBCCFFvbHqpQPZ9j2i
Cn2VP4y9SY4KGqTX1M5NLMxHjnSxesl5BJcetcjMuOGTmLkzaYgfKhZjg6tO9+nH2zcMg983IHW7
c5LlUyNZGO89Sx1N2lWbkyR8039AssK/4xPBb+BEoaMr7KMN/Yo4Zzr2vcBqMmEA81Yo6UNu6OV7
WzyKrCaixyqewNv95yrN1j7OdQPVPuuNp5T+7LVDWllpUTY1SaApUs3/fHkrnU8NXB0NemOX457S
7LCKGIxxcy9refOeFIVdmFVakEZWOUqW3roCdoB880IXbqePZt4CiLo5Zvg3hP+tTWLKbNJgYbyO
T3M4+S44FLdrNlqAKbjfoHsqrepsQ7X4BC5v7DiDLI8UnKkO7Dv2fDaXQc403IGNE/xfXQKPLFOn
abt8edZwA9NlYZnyLpHbEmc9tYfwY2aD+O68aMM5Qk9j3tKrV8DTNeQhJOjYMZeQEGAgSgO2sF/O
8n2+erYB1cXqnKMJ2kgCIimjg6/MFx2UNnvRHED8x7qIAoLFw43rLkuTItEfacaqj6OWmAwVryau
VsBGClmZqNMEw/2AL0uPibjDbz3woiSdPLZimog9qMInvftjklNxuNHqnhM5mDZQGF98DnHRaogD
kid3DbdTxoeBJTtjKsPSqG3vCWxMcFUr2/HB7TG0NQoQkpTpFlV7MBghLdSJZS3InEuO218zWAi4
pHDwZxai1lRWvXqQqPJcTzPBd75EtFWgy/7Rqju+KzJOGu3bjq4d5XXyn6ZJq35+M34c3Ypxse62
r+fL8kORghx6nyLF4zEmDyqAFrD3mbgdazUFnyu8hlz0mJjNfto8LBaoynOXQaWPmaFYFVXiDk3N
F6yycNuWyF5fcDD0wxbUHZ8LjTpb6A2wF5MUZZ973bNVSP3J9SLb2oSWj+y3C0os5QQI1UyrY5iZ
b9WxikT/yYfROd39USNPYzPQ6HrXGA4it0x+7gNnd3xEOIYNosjNlcH5/TwFPKEWThV7bMQ4ZjpZ
FsREtxnCXXMsRNY3M7Br95fQiyqM2oWS0YyLtBgWRxiId9C3BZazWA4ILV0UbkLJR3u8+rMDmK9s
WTUbk5LygEC4rPQxu1PFoyZbr3X/zcorX1b9+zLiq4Vs2Jp2d9obZ9SD0BgGOohYWMLFL22MZjbl
ckwv0cM+IJVBxERGPeZK4aMccfSnMTCPJrpW3nwKbuxaPa/KCJKK7wi03b01uw2Tg4aMrYgaMEVm
xo1/G39d7lINaMLYoXKUQoXRYZ6YeWYqVdi4aEmPWa5lDYSSYHt3W0meYwwF3GgRO7SYC9WbGtEe
raQzXhWF5NK4SDYdaFeLxKM8q8tJxzfd0gf2cSP9Vnmg6HSBtD/vCySgaHChCtcA+Y1rMpDuSBnm
qDY9PMWKdWYJ068CiABRV4RmMr1Cwp+fEmNGsXcgsRY+8/Durq72knMMcQZwex9O6CHvPw9w7FJO
UqnuLopdiA1ZXSBftAoPZSegYETvsDXq4mx1GW84lU4jddwbp7+vuypAJUrN7eClghzE4Vt18z7I
wlNkkF/inoqEl3oo5DtbstSelVCsDHkQvRu1DWbfDu1+4iQrVCMIS0ZYJoG918EpkKa6fuNfgvZO
XsBNQfuH3FhWG/4C/A/JzCHjzfZW5xltgpgKiM2h7tTIdFejDU/GW0GEgXYy0KQjIqRqlr974qWl
3hCVBDt+MpDQCgAzmZ/wjrdXqxJYEhy0cdalHNSugS2jFk+RHnG9FNEYrEFA5mxVDzmWF+xDI0Iv
NeaLksrUehbq26bvdneBYzZNouq/2zVxSYRTQkS633mbVpseEVDS3i/wbrTqC+M/QIcvybgv6ykm
ptbjb2acp7kdVmWXe7XSNz79Kn4ly3SeqBvAR5kbEMqxGK98FDbYbK7nShCvVsZFIiw5AAyou7je
WSUEMo6c8TI3cc45FZxJGr2jZJQYdtzneYXnSoQ4CNluFTsinddTGjpELc41JO0UeC6UgG4N38as
Yad3SGC37R/l7vYIJ8b9OHJg5IdYt7sbgihQoqfMz1ZJdszsDDFkbV/yE4nPYFExzR/1FD7TxdDJ
8iHwKxqfe4rdn2m+2LicoXr8I5B+YXZU6B/CwcTR21rhl8bJdwgtdV5LwwCCtHlQI7ucf5coEHgB
zn6NSuv/dPxpDsMCVSXVftGL5EUclhgQPZbrkOxX8VuQJjP+Z3nk7DCinmdzASRGKo/65c+Y4/BS
Q0I4e4Ru4/jzqI8KMHDYHATAl7hB9VYjRp2RXAViHTXl3uzvZqsr1rIexhF3RqEiFQT2tU3EkanH
twwNmjRV45FDIT8JJJCtH0Vhyci3zM4Kz4lhLkrbBXy2Ftk2pcXtHUNNONa7Ae96fTeTfNFFkRKL
PYNrS9PU7aNprIA5lp1kwOBNPtuw9+2vwMepqhQXBgnoQHH9QYXvQsJlwnldA/dkP0hFHd5VHMTR
c3rrxLTi4+haZh5fdFXVlOUtDmqyHTcim9T1wB0Lw3hG9fh2K59cuGBVQiEuS8nsRCZiBmDw4lGr
RCqacnNaG+VRjM+vWZHYykvoLkFDijcb3dXuXpLmYFGOsw8VTPpmtFNURCQ9yVSYDwNaMeLAkTYR
1TVTFAennvqukDCojt2wdtbSvRAY3BIB3/K7BxhqL88p9oa7KZOzlGVUxg3nUypP/gRND0dQiTFK
zD8WKN8kLoLGZIy2VjqgEjVV1mVzyr6UrxsntndSlxChMF6xzq7UvUIImDCPY+ETDwOHlvwT0g7X
73Qgn2WcaFIR4uY86BCTK0QqUGjO7uFZ0Bb8ecX5wmwFRwqCnqtnuwm1X2pSZVgeH1PTKxoadmqz
AiRcozlPtZGIgKBh505OuqWrAgiwM4twxOsNMHWYtFDEjiMIQopWAsBmd3Mc779MeHdWHRHpwY80
EK3gmABZmnM+q8nZeJj7Z6oqzUrVVY8xc1BQ0A1jMy6CoplmBKhp5mp3iTfl7rjlmfqQ58sI5Cn3
hJEgBqiiZyTWUKRW0Pik3ZVA7MQLkW7CKH5Kl2C2UIJoItngqZMRwcLTk/vRG3jcfaVZmtPUtDVJ
nhY4ul0Zh/DQxjG51OBEFS7VL6OGiB/CTIqsl795qPTpQ6XKhyi5f7jikufQjnS5fARdQjrXlEdO
Hk3VwRh/7vl7rzST/y5vMaAFhEuWqSiKkKWbRRZJYzz92gUGTOFeRIZWKBtgXTV9QWxaP9+qn5kd
H3TR4m0wEXlXduFAe+qRBlZ5+qIu2L3WKCatoGmoT2hfPjdSdOOrpzATaB0PMYVtItxZN2Lkl8gr
RoyJebO3cgqbebXlJtpbf2zCOjR3TcMqMXozr8UjNbjuCATEy/QY7EJdWEs4aP/jnhmf+QrB8RWh
3M9H4wk7MQTcflRObs3DIkgdhCejauGj5XPbnYy0gGQFqOSQQMhlGNj0t8zZku28O/sWa/sBRjda
5iqnCxasBmMOccGznrsg/cLQZYQZx7LItwdwaBZeiCwuBMIigXwRh14l5249pBQ0+5W2p56DKaWg
5onbsNE2Wn6BCq7zTdjfG7fojuoLJeXAGBzgx4gQPDu6fkpxNQhdKUQRX+Oxw2vgK7GM/eRFtyah
zVNzMKmhGmJAOhmbllfWehOcmQdpc9oaW1ueFHz/zNA12L8FwkOj/kUXxGNwZtsnhsm88ETCBHiN
hF2YA3vAlvAZ2s0b8uHZGxKm0/R7V0z60Y8Mb8lnAAJpHI3k7AzQvdfxl+8H6oX+FvwNz06FSiKS
MQM6etuwzTK5jjKJ8pUd6355US+VB4FcLNG3dx8hHeSSSwZeswfPjsw0Nb5lW11l+rKIgT058UtR
7R8aRA9vxCTzFn910aWiyO3/dZ8C9xWODJ3Nl2U42g9gzQod6aHfqnhopW4q7z2RqAmsVtbvgYDO
Du1a8nT/oZvoj0Slxgc2bLbw3mFrElz0mGTK7ANNdvIC5oiROT4BYkaOJI0GEKuG8gahoDHQ3blr
F8mHbw4I3zAUmubsblf9n4M+5U/wS8fkJCOpT3flESohOUMt9V7ScD7RymbO/K3cwpoVRyTup6K2
ZxLkBNWxfXE8pEpbUJbJr8AeFawUtZIltqALTXtbWVRdP1SgLqXnMqPoySfhirUMrvU45bnrelGh
Aq4gAcVvvP5shO3C7LuVM9H47SxWqkO9JLtyjz44+hOkM81qQU3VVL2kQhL8YtUBr39fGLUAIrCg
36NSiDKz099Mwxg53+XkymP2i+eKQMnRvujXBdG5N8iaUqGnnE32/PJvgDsCHcAzXlQ1mN+AU11I
v7z3x/desD23qNvTcoKv3EEsn8yC/dACFvdmGTa6s576p+m2JlEW2bgABZebSjs7M3xETMOT2xJU
CF2ESer2D2qphXEjJybBna1rc0AzdjH79MiEp0xvrIDRs6mKEqMfEMqoKNnO2SJ6sN9C7uGtBZoL
BPywk/1X8yeCgAkxtsIgJJLSGXbfqNjnz6efLho9PmcUUh10tiJEdwMdWSlvr3Q9T6VyXTIiWLHm
K9F8JnkW/HYZDR4Nd8nViOGTHA6ttC/OaVdoYzBDLH/+lBSQBgTDgWVmLT0s4j55yTFqTF1K/RIc
ahh4i1kGAUKkem6MmyAK8vpDffPeSAuMLBWoQQYiFmH4grvysLsUhJzpztzYaFdJcEWfwaGz4N3H
Q0cz20/wSkZYuhxOpF4asIq70UuIbcsfrFZG3QWcB/Q3KwbUpbfDTLoHVF590wJvc4Yd9TpHMQ+o
j64+g0GGwEuBaOMTeNjrdcm7k9pjR/sGatOPbK0GwbLFUwj5eEOODEeBbJObl2zr2lwAhDG2oELO
4ulNm1HfygOzCfbCMdbZAxpp1ORL/eWvJj8qjKo3sbyK3LazCnXnP/jYZgJ6xX5nf9N2IJPndmUw
ze0ER3ymjuX7ppmfoS0ecabbrpts5PMPJtYjdrlbDV1ktwVAJ/PsVnnKEnaQ4/X0xBFGcuAsrS8V
JLbIxYJ48LKAfpb1gjzhMKrc0TYp+2XjCbVh4ESf3K4ZiY0MVHRpPgSk+8PTsJTkQYaqez1TIkxT
6ioVsoCLHHA0VxRDYvXfAsomoXMf606Xe6av7UB0cbMDLVp5A3EZkMZA5AYoGtaQDs017bdDBxNu
nwZgZyep84w85XlHaqqc1lrpGkXF/EHCu4flBQUsLQTzJs4ms/cCDGyP7v+SD49GhLKt+gDzm2vT
SCv5/DAGv9RMjnOfcS1ue9yjn+2wwKtsoavTQgVbiv9uCk5XyRHczGNt6xgkv+zWhWQYRAdZb5a+
Rc3kUFStRXbz35Y1A05Cw0MYcV3u+2F5XNnHeg+bfcKhcCM+toXdnaeAhfUflwaBhFAJ3a1zE150
33K+8WeIVuHesfDnJRBMxes0BfjKGyT2uKev2USobY8c9O16dVyGGokudz6Av29v60d6r1L+iEdT
UTVL45GThk9O+c8dma5uPP29IoBIdQ1j4+ZaOKiuKQCPfq10CsYHFg+3aW7Zd+q5LqnjdTLiP4r5
LmD4WLA5t+YdXs6/3v9lAXaMF0npYvB007psfBQttvgqZskrw8pMAFIF3WzB4A99iuLkN8toEbGr
qBDfDs/HGIicdiOOxOj5xP1I1aW07+k6nW9SgDiMdChNNngBzNX35fa78jpCzyZiukjOfs8pt/n+
/2HRPiyvUDbQOfbGwsT2X1qu/LATtlNoieDm7fTcTqbJ43Kwqz54Le5qdp8+KM0NT9mhUzyP/q94
6JspPbwEVa3hhI4JDNj5y28EQ4kNe3jkDWMYOmdvDZjhamZHlvl0uJ+lX34KpcwLK8DjfJf6Jj9x
DCfm6dj4mVTQ9AtQYUnLmavNLJH1yZGtxbM2nodX2bnNhYk9j4gQtE7CwsjGPWjHzX3ENe/iddqM
YG0+9g0jW6JBMUXgB20Z+ALGrh62+TDdoTZ9+LDZNLrc3Yyr8dGYobXZntqZo8JWVmrXBZ8RNll+
rPMpcrHkbT1GAflensqKiqg4fSEAqS6qWmJSDkDb2nALGqe9xi6VxZyC/Yfd8nRACkvsV51quKVD
vemXqwYjnv+WgW4CxZpzXRh+HUNzywnBnYt089EUVWOStkWlt+FJ1kGvz4hMx3AC9OklRUvdH2X5
+FxsVXJ5pxiotyj44RL7BIyHNkxV37aGdZUo1zMoqnOx/pY/X9BFOnyBXlByUHX0GtX+Gsboyvmz
WcnhXq+Zxjlk6iFW0GUSKTL0IuRE0R2LE6i53ZXNkD6J4AF634fJop0KEFyRaWci+YXiSh0LP68O
4+g7Fw+l3lyUw6ZM1gyi14HfVA1paxnM+SrHUDhFQyQmNXhDAMCsJRcXEO/ToU78wwV00rsSCggU
XY0lr6ZeYnmcwq8mzElkL3CsQ51VaZ029ELNnwOoWgsAvL5hHUK1xnfEKf1atHVkDDxcuPMhbrQS
sL2E34jVXg+qtBQO2uqG/2X6OI5L7nL0oMRLSB9UtQGK1EI6ZSmyiynvGvZcGdckTJJq7G2+f0M4
rxMw2llZvmi+y2qMST8xQC6Sc5bk7MZ7U+Dy2pKy8MUmF93wXW5Q1RqrrQ3FfM+e8sOVA5owR8+7
+nVVUum+TEUUc9WQ23YI2U3KlEmdg1vOFMJK+n5YV5Wiyi3KtNomurnDUWmk1c8sxF5QemRaGzfz
9fAXlwMWivE4Jlx5yr8CRFIf/AcmchBIoDgsoB45Hks5jhsYAGTXVQjEW3hSf2w0Q40/AhmSz2bA
RMiBMJTrjkFmON6+IH5E0zNUBnRG/FDbEqNWQKKXgkojMJ2Hu9BI0Rek678vL8XLogUfG071dYyA
7TM+IYHH95qpeFeuRHieoTY3mO62JvHCDtSn9Qy/3AWRuOK2Jae8ojmJB95/BBeX27ZV7aavIZg5
KIcpPClwV2mD/yP2+3gtbPh2FurkF+/uc+iQv97j283Ky7D3P0vMC4qDCZSDWrBg/M+5hcRgnIZB
Pk4bEKhp7MtwzM98Zo6eeuGO1dn0nMbHZvrVKtHIRxWjqS8e19vZR234+IJkG/xaXjuvFOofoO77
/1rmGQ0VBsTPkJIeYOkHCN0T/p12vWjHw5fFqQMrnNd1ZSExSPUdCi39gPMNXWimbJbBm/OGFPHt
6pCBw1P2vFGMZI68hIdISsyiRxNcPJxqn6Pld1RPhZh5gaM4s/eiYp0rAg/SzSORONkjPmaem/du
TrIgYSabkQ0jZimP7tFk0eZMFx7eC9i80YTcUZYxbJM1UpfWnvp+VIbpnWvaWiOKg120tXMRJFNk
cszTZOTL6kATbaxi6XoF11+Q6pJz3tL3sc7478hyvy4/CKsO2AbFEp8GvAx6yJ81UDpyOi9FTEgI
hm0Clv8HzFYExVzMPj1ZzdyDYNM6GCYKwpcU4+s0fDV6yVBqajeSn/Uz9HHpWK41pTc6oBfdVYuS
CyUisEI8suwDBNH9sMhNzAArUS25WYdCHit0YIIjk66nbodLOuu4KVRHI226tFgDE/lj12KnT09h
wXwW1s6ct3pQ1oRZHqlmDHguWat8T2rwWqfGmEOgyJy/WL3euSg0ghHaOmo8u3p9to+jZAoM9k8n
d6SwzTiaROci3DccQ8gU064aAwIXODh92lAGjrCASLptyR5e+QKaxULISlg4QOOCe0f6coBk60MF
94CCFcSvvLguUV/UWIMiSkA18Gz2CruGyB1XTgiBeV7NJWKVu4mKBHzB+4yrnpdF2Mabiyzhz+Bk
yFCvGSUNO5yXU46z9vDK1yvgbUBtsBk12NSgfdQrScbnSlAuJgwq3HvAq4zz17QlQa/65Y3XHwCr
p4/1iXmp/OeeQotY7dM0MyGuu5AO7zTezZltmiUP8MUHUQkM99JdWIds3IZ9x7QvJw/hzX33VPJ8
KMFJDJkC0+ZKDCmKxjdTUOTqgFizr3jG/MUpK1g1co1wMlWOvKqBBpzvOUfopbH6hoPCop5Z4sUc
/XNGQ5VCT/JwEHBTNCduLG7DAX30YuHX3q3Of+fISFbZJ1fujw+Y4n2LPnru14gIQmviOJ7BQ3H0
8iB7rsjdH4y1a6+L2ZzfHgFx0qNJwMwl0wPBoqPmMlBB0/AJavLzOmY9tk942xuB/Z51hBlDMwKk
A7nBabR3M7MozMSMFYbbKW24I29JV0FmeWxiWUnD4b8hxzuf0ZoAzb0ApDb+rhNR8j2QLbdWNTpE
Y9p74muithyUk49BcW1xKWAAZS8QeDSZEIJRCqjK2k8sR5ArWCVOkO0IoE1XEVN33cwaZc6kSEGB
oFi7L+wlPh7aT6B8gb8GW4XhzOlAgrvBZdy5vtEhWA9DTPKIGTJIeBodtjA7aM9Ny1kYRdYd4HOa
1dMlDBlpjKjnMLSV/vunrovwAtuuvIf5gHZ6hwsxkGAUNE8EO0iLJDjguuRqpHs0aDGQKMA2IH08
c7Hfj8QeUcGvltWVGS3LoJ2OyQkip7w18Fi9gQI1RkVatCUTrVo6AbgrepgSXL5Mtw60LP8FXZwc
FR8C7mRTWLgsc1mkea5UFNcy9hrjWElekEjgfJGjpoI49Wl+ZnbC1CXof7oqhBiz5gqV7s28Hv79
IDGWAR8M97tlcCOOXFXlVOge8X+w0WTwceAcyvepBLavnfHWI7VPVKCNrY28HbSZ68F4lh1G0OFq
tkuVe5dRwlFjia57J8rwv2o5k94IovCjvrGcEfLWdV1X9yaCq8pdNLVWY1kwRarZ6Qw9DuvM7OQa
on786dpDx8grtsvMWiD7+sWABO0VLjeNiXYTvmYF2ZWi/8He8z21ogGi7dPVp8htaNWJKoGwCO9+
F2GKYuTY3INIJ1VR4tp2LIDS3F54tOqdtneIVGo31GUNBUb9jS1bxIdK94SdQOGpzl9UaNB81YrC
kXIFepkUF40UROlhEnSzSVYIRT6HGN/6SGh4FietZIsb68d/o0Cq1nqb/Ld3ajqhr+rTB85ki7Jh
Xyx4xCVbPZoqUP4V2pUoWLtYqieZKpYMZiDEybfjik1OVHil7HMXvxaQDm382DlbLSV7DDlF1kOt
MzCV1sR9b+yEdoiHtQN/iWwZqc2sPGMGf14ZmIgKu58N1z/6XFxUUzs89iHBfVcAhCJToS4dDNnu
mEPQxU0g6aiQ3NbbbrAq+FcF0IUBxzytVWHwrtxn+QywbZ7/ylrBf4GvjFv0poo1mBXFsO/HkCAX
vPf7GQ04XMeAnuIdzU2p9DVTg2QV6k9kYDs6R01IBb39RNG9DH78NvfMt6EHEylfmtwnjleYTnci
8eXrsWPgSAnuj9PzRQuGgHl1h7mIvNsAtshKAr3SG5B+6n7jlcQvcmoTNzohziUmiNzJ5Uyv9ycD
ilxj9x90U12CpGmn47O7qkwGeW+ZiemWG48GX4SJOQC4pnfeVkZkVIGyNBKOqHh9ULg8pPzP1dMR
HYsttWGHQF7LFgLespsMG9fOpfleofN8coshpJprZ80JjzSO6KBao4aC1fJASFkDzUCuEVAWoFMy
3qirhMF5an0YRn3KZSu/X5MMHy3xMBHi4u3s93AK/h4Bl3HDReWaUiTtvr+kBToXcXPDWn9A0dBg
9AJTLS2n4W/y72qH4ly2KxYA751XaRI3TFcNRoj+rYPGUDcKzespsjVkCYuJOXDk7o2za+3eKNIt
2AtCZieDE7QNFbtGCRNFcNtk4VjNtRhyEGfreg7dQuqvYrcws5/oCx84CZLt9Rx5Mpn8AD8lpcPP
vG9p/+pYyFsa1dBGrLkMVQW7CnwMs5yP3quCCuk0WiKbmZXrGPIm8DgcupBm6Y9FeqCX/AyvZxdD
KKI4zvp5g2bnInGXo5jU2ZFJR2ghjgftkYFC5ZBjw1ulrt2EvSfpW1nHBCRAcvdvNDCQYWqxweVw
yVAZ3svjtulH4nAioZjYYw99l2bqr0q6V4GZBc9IX3L8txboyG6KLpSrKCKk6xa4eSndniCgF9bu
l+DS221/Y3uJQ/KKpnicxNnkjLQ4WZRu9fhOUgIaOn7GyoAf9nbzjmM59on27zJyHrTkR42kjhya
ODvZNgAHvwpS/vWtCzAzTKkybpA0QgGVUQWun0OfsuoPj4AtYGZI7PJCQYzK9/s/qzHF8Wod8tpA
nBfAS+QojGZN1xd6Ik1YnEH9MwL9GzyUoZVZ1w9xSe02Q7x05MbuONwGfYoVuDcmQ0QQgXgky38Z
wE5uteh4//VduKS+geIU92UYEO22MXX/bOPwrmcFvI7zI+ky4qk/uvL4uiwJ5v3F4c65IrRnt9co
iRK5qqQpTzj8KEBisMYlyXgmQn7T0KbP7H2YsGBmylKSZ7KCru8k5a3qmADcWg5PRwmj2/CkDR+I
oL7CFnnJUc0dr06sPj4HJ5b1a6X/+tBQVsWrnNe5ZuHr2FHex3jBAQ28fRMLwQicWba1vkdirqWm
g/2cdIL3H+c6F4f1Ig+rKt7Cg2vBVS66zWAFztnq/MVvPISBVYTLyiX1NTxHo3ie1iVbv+K/I5Jk
GpBHKH/iMw9Z1HOKWeI/ErjadpkPxeXHuONLcupVTtair6HwxDSOZhJXdrMWU5nEVxfBMcpp6C6F
Bj9bVLbvt3FxAtYk4kZATT7ulVRCk1bfiym4OqR3mdD9svXb83XAFsWk17R/I83HC1PUIIHL3frK
Z1pXiwhgjfhAjdf1qHFehE1PTfHnVSsLJugNFOF506/nMCDeFM3M4mOBpBAsU8OVNo/+nzGKMawY
lREtFd7DPLQWhOuuAw6JH/E7F8PwGzThL5mJkamhdHvFi4A41MhIumBzP5MEZoR434rIT6aUZGjk
7X+K+95HZOEaLWakB30We4ZI9akChTRaytuEMw0O/pfN2g/kZHJJaFoLINeKtGItu6DTCvLCDWjS
6z58yBb/W88XDvsmVMEyaGy8SdqlIPWenb6gb7y4dB1wW35w1SQ7O/G7nsQawqctcUCHowkNWvAO
tl+01kXcCxsyiq8k0KU4uynPOw+rZEoqsje9oQ3/BoL3honPHvTulebFvH3Tsca29y+Db6kY+BKx
Aqc3P8EcrpQmD4IeQiSSFz0xF33nAJ30rDH66u4kGSjyV206NPnYunQFOWQC4poiXXcM37CWLwZN
YGOLTiof6igDnoXt/O8CxHJ+An7RFKWL0CCS792HjayZbjd8bdOXd4TmotQ2sPwa543uWMtfE45l
1opMPUPgxpPsu6md+RbEZ2kXXswsV/w6JWwcQUPhjrYa+cmhhBz2+b0yP2hiJq54eMeMtPudX02e
qIG1gGFAzwTuq8tHzjcFTklDfBwchQ3Ulr128DOPpcg87gYF6fYhwMy8SxA8FsCvT5WpK8442V3U
JyTt7Qj+7ZPUJol4/L1q87SmHKbF9Vyj/znNWIh6rooxtfF9USFW9IEX7M+VMaCqGhakFdDzahkQ
q/h4V+zA4ZG9GQYfFJVvntyoxisVlWUcMh6HTcD9WFy1lfBXv+LO8okPg+o/koIduPL5Og1XQqm4
tVNI4whU89OtZ2QIk1otKj8QC4UW5sGTgr2H80u/JTeNwG+/y8HMltG/R3RjyFcsTNja7nuI9wV8
heihkASeFfGNfOdqC8y2z9CtqPjEU7hmL0XI22qZCjTqhudxGTWFKdTqC+MU2EV0HmDIyp8+CBSm
nlpnS+96RieB2lZRmNln+ownOpR/5eoIdWIoTx2WVUKfNwQWWqG0L/mCmqxvB41g6OtEDAU2HvVb
b/5yWEdrHA3EnGbJTqTbES7hkgcvazKqbj7PVUupnttTWGDOZ1uTMBPodIX+FF9woofhEzw3LjIP
gN4tqJayngzozz6dT0Qq5QrhU76qhz+e3orvwtW78z5OvmWWMvEWvrdnE+jslCoYETP57ZL8kXAY
s+e+rc+59xYcOf3MCfZv4d0OzzcwOgxS3zHyjmcQlWqicOrb+tglx+BRJAOmifSiisyjIGX949BM
QK0zlxJc5Dn9lt9hrGfMZBTRxESQFhR3P/ZDshRv2WNRifDdnvVUhXyJJmvvwSRv0CDoJHgb2HjP
urQGixcTvdtK2MZOjHObiCLjZwTonv7hhNN57KUr3Bxa+gWu11/ED4RjoaQV8YfoQWld7YJYSgkv
48Kp3935wrxpEpavg1I+FRa+QwaJja2dx82Hca+XjEsSWxVf3Vg3UgHixM8kJ4X7YF4lz04gXRf5
hhKZi6yThM2jLWbffnBqnxEeg8dkEjB65P6WMb/XGbKlavncT/PAUXBo9hYXO4WjVPmWNTc+M3Ks
0fzX3sjtbN2Ib6k2FGAFGyEEC7G/CrSupKM43ZuE21sCCJReqgE/0u/sPoWyIoYyva67qlz3f8Kb
qUYHaWc3AkP7xk8KrmTssthRPqvlWV1mfEzB1k+UjLPbGByXSbqyCutefoHbm5KxcuDIPbAqHTul
Vxuy/inFYA+4j0v8TgXRabZQavZE3aYlEWP9i5JzwhMuJsjGXnZxZKpSHAweqnWZ7rKXDc0Sfro0
Uc/wLMXR/P36j7FgAEPRCDWV+YZMfDVitY0zJxUoqq8lVFMxtTVEGgok93tLQL/kntGYLeGI+Fjx
yoDAfyOKVKwg5fR8pXGvu/pPbo4HrK2yEdl/eFroYTZFVSz7QS5FYi+OO5c8hEAguy17O0+SLQYF
2LIkRqDBmBlpB5ENrkx0pjLDpphTM4lvupmSGMXJoxKrHQgAq8RISCWV0tqI2OTOHyqluIez1jOM
hJ/yiKKMMscfQ3dgbl4QUPA4l2dQrLqw0ZMr1cFm2F2kTogxVVnyjMt4OanT91zXEQaoot+fwNNc
mbMLH2aeCs5p4S4wg0/OQe86uMQRrN45sofcspkraSVx/1dnlamh2cTr7Eq41diVNFQLb4KnsYZ/
pABpV4T3K2cXB8onW8y8dey64HwvtQXBvDsdmM+4KJqSfiIWvY9hnJ1FMni4jkq4KYVl/ohzheJP
8hBKh5riTEnllVebuqteQCvsyPU6PYBv/pDit8iUmHaBjpElJlmGN0ULy3x9DgQNZfQzZBztV/I4
FDZrl3TZ+qm/6oIDZIMF0uceiYxN0DEL+17gwoaWuG6hM2iDy8u3f7tbOmxYlKX8L2vDRf3sORfy
sQKdpbTFv60ymOYi2IueeEtsNxtgc/vw/PMBV1UM8IcOiF798wl74kVz/ICoScrI2GZLpSDQLvaR
w6LJsH59daIsyD/2LHAVqAkE58YauRkCS+8Lk83fj07mc9o6cw3vjZVAKWpNwJHr4nGjYJDEZuYE
quaIyKxEKl1FL1RMafqX0Btps/lN+JZ7+UmZekT0hiw37cbz9jKuVtyVQAhAQNxVsQKsjznXPH6S
1TTw8m7Ifzf91IpXHgOf9MhyRsKdp0zRmg2/jOG0pc4mOFh3O9EANPNIpTWcGt7XVXgMGjMZmqgA
oUqGP0jpOyLc9MrLMtVQowjPv8YoaMn2clY7vsbuHgV3cNNjkyp0yQtctHEIRZmCmS+oQ4fU26tU
4zVDAtqa9LlwwFL5fsBvqCH0eLgpKMxHlh6/e8vLP/AfWTJwWcQzZ4NMhUm58poDuG/hWoY0E6BC
0esW9PfI9w3WzFoFekpusYbPnlVEjEgit3LJPqf5Qc1TazkEpE5R7j3pp+nm5m9dX4SVrrrIKAaw
tXpCy4HfLizdf6tRG3rFzz4OUca8zWVVyIVLFVka/Gg5aqXihl3GArg6DInDkTWYChvZ/aSE0EMG
eY1WniIb/Vcslhfr4RCHLaTci6DR1vCL/vF2bAQQzSiHNA49YD+8xacohB2X1w5jpcJh63XpBTkv
RWmrQngtgE9+cAOPhwxEyTkUwhTeqSf8cKn1cOnd4m74K9vc4Z2MhPHI6Y7Y7hXCEMgo7yNDWakZ
B4bvAFc+obGoAN+PBHKJ+eVh69Ld4/Zw49OLq7o4FqS2nwCYabwsTBVDuZWc8iU7WCeR5Sz/C9vA
jT3AH60FwKMYDjTZPKiw58uqTa0m5TXZ0+2hoaCrJws0jOdOzkTqQNGpYMTID/fIXQXqVeLD9jH9
CbHT6Uo4RRSkHvjCmwfmHDS9tQZNfLHJMdfsLfDUgbfvEkG/YFrP7mQjNT9u73XKWjlWAF1HTlVn
pw0dasoradgrAkKQYQaS+Pr5iv4eXS+wm2bhMJ6SL94BiqXXseDZm2UgzMZn/px5oFUtC3LEGqol
U1eJ2L8rWDoSnS4lWcNzc9uILogVlqf6p+fg0nIPe6/RrGV8rs8YyRg0ks2kXYLjK02zxLCYz1ur
ghhyroaXEq5z6Ys93TpOGlQgiR8U7/gsT0gMeq+ff85fggqiIJ/+DnxbKAQpdvz2N8lht2DtL7V/
62oml0AgyfA74MoUxT123CzYVrZtSz9awA2/cOg8L5eXinWBxrhppyvvOqZLHwBxoIjUEggIr3t+
eUDTGKNGkUYVtzZ9vsHM60QhtUQu/PAPFu4RQcezHOwHFGjpVeM3GfaSZL33mZPXdQ3J0OWHDZBd
b6c1qjvN9ca1kjt+nX9xtJ6ukah6ltoszFmXn4m2o9ER3vAGEFLh2C+UGaV84s0Td/QWX6BJBfr3
nUpQeL9/PS8oU/y8IN5hcqUsRm7PjlV1+LnM3X8wuiLE2mZXfdgWtN93qbgvaeC542gVS+QvKbrp
/jj89rwERmrU2nGBoZaW9eWPqF/BVbpXgqqCveA/dqg2d1xCroLUqmdi9wWqNJsx8YX15Pcpvk8K
FpwtfRcDFwmqjlM9wqMfP9I0eEhqGLex0sM+I3trpKeZ/4FOvImJIXdR8J4kQyKqh4twky7ChxQ7
qsa1MxF97EFAhcgEIPgqG/0i1JjLoVLDJxiuB84rSxP5BpUtrlqx5Ruva4PXTVl9QOsZjCvaXQk3
dEqKfYH0aW5P9E+9NKTmKYtSOhI2OQwgWLJEIqCJxyIS/yibVPembMHgHP2tgSAMpdYDSmhpMpEz
OYrK6z3Wnw8PYb3zXbI7mPsON45Dt4REwXZwOFW4FZtSMDSLUf8NOS+xEEpVRn7nLVvlETNB1YGm
L1vO1km1zQwNiwptYNNWMN+t3SqJRZmEZyC2JsF0IPed/Rn3FmQ5KWPvfMRZXjg1DPuJACdlzaEb
YUWnrtNpon9QDoOTfeN+a8s8XSE1jARL4sF+sJdQ3ERUsp18YKFT8tBk6FtF5NqqH1afhxNNWKPp
IlJ3xVWVt7GqPoZo8wE/cTjw+Ouin69B7aDwqg9BhR7+XeEwN2IRbBQ+fDAhziiO5b28IUPVrLDt
xbvF+Th0Dx0sqroC9WBKK2dUcAiPwKx6IzLXNEuY94hiP7hbW+72h7Ues0xa8fTi4fY1AzjDUF5a
pfEEA3Dk6rSaYAcePjjO1nRab7lwKEMVu1OzQDV6R5L//b1e2SBX4rhymzQM1HGQ4lCmx4kJ9MUd
woXJK39C8RlpPhnFnCgr3fZDFrvIGI8bF3t73CgvmlT/GY9FcPWwR87QiWdS98xXy2Li3YXKbdCR
GNmGsXKaHb4ePsSCkWKe5rtmz3OEfrlryTMdrFkTtudxa8U8u6U1o3BqaewLjfWHwxZuqRSpZo5b
jLY4rqBDBEX/K/lSqG5j0GC7hINOTHXRiYqZ+KISe3DwjcQRAFkB/1foJ48AfWTIRI+C1EYPlMJP
KoTqaEeUJDsRXCICSTq+Juhn+Wl0bNXnPlz+0wMhJUlKx9PnCxTq0EirK9584/9KnftICg4yOJOi
w5IXZu0cUBNw5U4wCGKbCWWtkum7mi4MERVENaaXsd5+sUutdvwtodmY1Lfpp5ZQc6DIZDxN08KS
l49p7DqSihzBwC8NA0HKLFJ1WWHZSJvmTWKKgwVeNFaYihGQHP5j0kMUK/KxTl7wVLJcSdWlLx2S
AKHJJImIU+jRwlwMW9T/+13zgi6m3mUGonKP5hWr9M8Seaa1KLxn4NPLr1njOMLEYg50Cbuj72Y1
0HzarWCR2T4cDdhEUgSDZwS8B9QdspYERrUSHtRavNP9GnWxXh/tshsPhj0IN84Uk7HnA2AkPk7Q
qT5x4KpcBBFrVilLihnFAEQ6cIm7LLh9I0BrmjM822ImzJ02LBqwtw69knQeE/rwRY5pgnGBlttx
RRaXaRwBRjBTvZ/ji+oRuDGXlG5U2aK7+jiz04GGttUweQXRu7QtBTP15IyGh5BA7fkOejJ27uo8
k6lrBGgJYdt6q6Lrdo4hHT+EQ/nnph+cgkSDBiKORzRUbvTAdc0ojgjETk0aQV+mVFH4b4J2LjdM
1AI25CRILM7t88RgGzVTg5LJs7xSfp/rNy54xZ2EtkbOCacfyTcBLo9yuvPsTVw+aG7TlcaAk+IL
YjxTt2Nu/iMFUcrwLwGN6nQovXJ1c+/cGGAg/ZJ2djnnFP8NGfE8z/bQLNEmDsfY9VXyhGhclsEF
4rnoyetVd1vuS//wfDkB0n2zdO5iU+t42316s+6TKHhPHGIY4XcKFxM3qfIcW/RRk80dxgOPNoX+
hAJO/xBteSGSx3N7xWSXaa8z2z3F05PppB3+sAer0mJXL80b9KWMG5/ZzStTRJhLFqg9KyGUiOtM
uVCODoJpeHY55+FCEYzGTxD7iP1tYEug2hKnW9wU9NbW/r0wF3da2ZRe91+kPMo5ZzFfChwTa8iy
7b2HMQfn/pj5jBw2UitmU5lL9cDzQC6b1gIM9YFhhhJaiogUNrv8LB8z75X8QWVsxr6mbs8Fu8cL
KZ6RPLgUmm0enQN87Pebz+qe4z9unsZjHHLgrRwa9kxMawTDhySmI7upDnDGKzoLOzf/ZPvj+6Kq
fc1axP5aPx5kihVNYyh88o76d6jHWdzNnctVvP1E2LXfQxGyfrVZ3gDR5jkkkLP5M3wkeH13khU5
Z/w/oPuS2dW7+CH6ahQMbJaibbqr6uINR9JmDasgS+wXFk8WTLq8mELMJ9SPqZOI+zwIjbPuVwOg
zodq6d7jxCPlFwu4w9BMn5nB7CmdHF+szUcadx9VwBm16AOV/dawpm+stp9ExlpfG/CFIcca8p4j
iklLH4FT5cVaAQ2LxPSkt6gG0e2lr5CqehcUM1ReCLKytgIIWmdx25QrzY+USDM2DS++N+oCzvm0
kqU9x9A7XwEsVUVO/1JYN5YEvuyTi7AUzHSsImDmpb50J60nJcbyYUEAq8AF7LS6If9vWM1yYEqb
BZw3JXUKjHf+gEv6dkhgr2wt3tRQLjztgPdgeo01FL6LWAeCtC8/vH6ppZ4yTdnvNi2PAJuLYsDq
dhhasxEEkn7vqq1tYyaOVwjPQoL7TuGis+D+Qv5spa23osBQkj9WRgE3Xa69M2XTuhTssjUwrGIm
vR2Rs4qnpMNY/9EVNvS8P6f7K0dFHEmEQpZ9TR0H7upOyjQx1b3l2VprnLBG91yr8OgJdU2BG2oz
PNtUKlvptuhLPK975djAz5TiRUFnRL/bzxluaqhF/B0k1u+gLE/WtMBR3vgo6I4EPsPV6BwdzYqJ
+zf0YGf9pEqcTZE98GHleM9Ni/kpqpaQJ884l5UnyecmAqYVf/CNLLysLGPpBV50RMgMoxfxW3xb
uv9tOnra9PpdGWkSOD9mekOKsQewOEHQipcDOLRvbQLSinaeEGlOdEquZOQTxwkcd12PGjdmeZLH
g+XEHivdMdToVCgPtTqX+ryxl1TgZeNxhCNamaoeVdigf0YZ2YItqwox+62jv5EOMTgpkJ3cOEJI
LoOFV7v7mkqzcHbdwBsuxETGj3TiYv2qvtWIp94TDrUyAs1hgcpCxwcAFpfN++cDHozqvwuWWenv
y6wqV4vDXJUpHUQXUPIZmHUXuKq9vm+bxL1M28JBFVuaQGb/Jpivbz8zu0wwnmS0GGZ4HOWWtHPe
QPzNwYfwg5AMbG5eig496oJm0Uho717Q3G9tpUJAU/V1V773mIfuMZYVhL6SFxneB6W3sKGlj+VQ
/wdCNfh0tqnhuj/eEswGjmkJBAmmk37iAtiU9g3xQpfANyjBEj7UoDDK+D8tcvtfk+QfaU/GYz3w
AbgfEjcVEPB9hyJSD8xX2Lji7JmMyAKDsNPIpMHhcj+JMQe7ESwCqGOSanEKABDX0GMa46ACbBUF
wI5topCOtUWAQ42wmSqBpdjH9OHHixjSk6kl3NZiTti1XoTROW7mG+SsmALJgeYfhWeCi5PRiTrx
0Dmashu6UNaqSd77tXL2gSYqc2GZ1QvcBW0dZ9NELxQKJJ1N1wM8wHmaTkQDH/cT7ehPGGE9DQ3s
bX5rXwyO3RhpFbVkRFUyItK/gW+wTPyMgyvjbCxd/q+qAkUHESjZRaItmx6ebagN+Omp3BoMjcAW
K9awUGCsgKzgmuhX3/XqXeZ5ak9XpujQ66E+srMPuV+EHRNYzeQCydFUB0bG9Oz20AYnLkOYRhW1
2co9VL7fjUFrma6uogKsmpXsa+sYKJc8jJ+wcyaPC/InGimcmJKH1gcBtZZJJW7VIGMD6N+KO0eQ
7mq72FnaaXQ5BTU1DQTud0KdRVbLNKXA31HqsezeOk+KH/k+hsNsyDn1KgfAqI35Gr1bsWMxPnsr
UmA6l3gjl9LAI/dxQEDJt+ELr1Icn4fZW2iD/RUUIZ1qT8I+XMzaWlrcXuUpvlYt4hxtjoYZTDoV
y7t0dsCnPf8UQAgSzMNU+U3ljNm2zGUYh1YQo/No6VABndMFIRclbYU0A5zWuZGvsb1qk6E6H1vf
FWZETXYEnauRWwnDzK+BXK+yiG3dWOwnpmHauX/ls9DjiJss2rtMqNffihDLPSuFH/l9qVmSj/AI
BPRkcXaqAezxapwaINeiHQZSYlPnUUWnLLmLeMv2o11Mm1x0vHM3m8c+FuH7BmrP2kiHL9nW3W50
9TaHLCwUCH6WBUZJZWcTebUsJh5wH4X8aptxP7Jn9KqmufmoQQwBw600FemHRdLW4b8Fio7gLPl+
vZoXeItjXFlpnvZq5mJrLyxdxHLmNcfJv734m0ACu75hmRtOMQIctVssQwDV6XOU49PqQJDpfivT
NHxmIHALpiviC1Ya7zOP/BfOh7lekX3HaTfT1UyqbdmpqNOwQ0vY+s9kaR+UWQAivJh0bk3lDkdH
P0gf94n5+T/yK32i55Pr/JBHGRFvLGfhjyF1zFdHA3TzHIaDUJMdvQXobphQkixPynS2J1hYgpQS
R3N6mW0sag5PKduQ3u1VK45R5wU0clE14rP46t+ZOmiAexHOGZ+M1q9fAcQhuZx44pZXwqj8cBzC
0IjiilwvSSZB/0lJPgGhrKhrSK2GcOHYPsGZy+fFHDtWG95fJ+4O9l4oc2hrFS0A30mUyJ/teDHk
fo5UY0wX8n2Z1WVlJxz4SVRfHR/4TZVnpDmUCcbkgFdpW+fzzf15OJZYv9fz8kxDUZizZ6uergc7
kq51AzD4S/LU9FQdbQ6AejzABlpWggEANDklG6xhtHPCT9kJAEThkvPRYGZ47S0O+h08uO6xE7m1
QLXqdsOrr8h3WHMivlNKj6At9jGEi5/tdbU/kB6Lz5f6qYVFgQy4Db4yYcwSj9DVQXZAqF2i0w+/
sRTkbI38xuxGBvHWiPZNyzjhEl8g5gbTnU23fUqO12nx5T3Ffnr3G2fQKicSiilTdMSx87S2afes
514Roxmf5S/KCO+qeYDIBOKdSK3pKBCO8CYCI2AB0ZzIPONoPNGbycL/tx4GJqV7v4hPEWJN/fk2
ud9lKXlO6TtejXPpqHYEfNSYijc0aqZgUO+ZkKUi0War1WGiX5c4EUGPFcturwlWMFdQK9JLVOfz
hfhuBUUVEJyIGcJp+uukrKwbKSgKUwF+wwloiYYEA5lSB8rqAEFqHvMWxKQ6JJuwr/54ph9ftjGa
bAg4zBIlQxy9RC7LknOacSLnQQuN1coEcw+2IRloyqi8TobgS+7zF7Jb2ibDIrk16qPwpu2/tfUn
4i7nsD6GqU+gz5JeA71e9r5ER8L77Du8iaD19coaRwfpVYTzQiCmMIkgkNyXACxJmTWK9Xr0TUmi
FZm6303ppJl3kGp35qprTezrwYmtev1s7MkOHNmxr5SppwxyG6dKk2gVf2OyH3qxScJ5AvcMS6Ih
GK1DBWUEZ1OKtOOSQpFLC2mJKRTrRCZVGO2kaWqZ06ng5FCojIjwjfLI5iqDhg5x9xARjRk5pPDJ
XsNm+7ugERHdKG+jS8plEU1nFjc15My/VaLkVVixf2a13n6968iEMfvTO8w6ccxeqnNcFAtv8C8r
u2Wi1eN4KDd9hUehkhLTxRk1qoMvtw5//mx9IpZtYWMQtz9+mlijb0t9jjHR6haHtdMg1Wbikee3
umFjWzwsE0E7bufqRU21y7y/VXUiNzCZB1xL/kCnZJCrO6121J580im/Tbdev9CZoQaRDq8i8HNA
UfcuIAHHwTbjZ8Cnbm/C4MIF10O90BFBQou33BsCjXSFgt7RvrDovDxyo2TUru3CzPC2ZMM8THyU
+wFDAI0gY8r6WX2vY8QsegZlk+A77shJSEGhifmsDMvYnOfMSJKujPE9woYQNVC+uYc8Oz/Fi4Qn
OMDaM21AiZRISGdCsaNtOHDV+bH6pI7+UL/dwhBs+eFT3+2tv8A3j5uYdcrQnrGqWVAbckcgYz9T
G0Y8/8pPXBtQ1p4nKxW1Hb3+zkWe0W5H+haa+5kzB83VB5kApOR7sCWEhKoSgS018WDZWeBmXKiO
ObyXmLXl9mCPHKH4Yez/M+pougiJDVKLf/CQ9UcTEg1lS7O+sysmSNTJ4YD9YRK+TIdg1/EO29li
t37Sdhy0Jtjp9vn9/TzYM9rFH4B8u6dB1H2PJ9RcmFvmMx2uPj5IiQm+hQBrqTd5W9LySMAAOITo
VFQM2bZZFNuCKlqWhZZeVeY9hnEMmK6OUTQqtXcap0d01cHsFtNbnT0wqkr7xUqwmzKYgF+EAnZz
2vQpn3yiFzElp7gFZziB6gVFLCCm6h8u3k98WxS+eJaehW0kBCTExXJ6NYFpwIyi7cElO1TpHF40
ARfwFQv8IjFDH9spnwQuYHX/MA/Stv9ZHNJory1jIPVVgPJ3+wsJ50lL7b9sL5WUuTFLLE6yyD8a
StjuUK+tTRiJ6UKAOViTl8JoHP3EeQGAzHboY23NZGXXAbWDGtrDy3VoRSpxaECmvzsS5X0kSEsn
fbPKO7clwwXqRHB7p3SyfAT8nC3uYTzht7s2oHiTts77WCPcaaaERlBm0F5XcRcekS8VhL8hdvNH
F6wbw4RJ5s6MrVtcDGQFb+v0zG308jFMYYh9GrFr+gEC/NNucWtBlX0XY//txOg6hijf7XHEPaUp
DgtkRb6Znx3kqkYVhievLO9yKHitBC/dizuu2iJVOTOD/oOgekMjT1f0vAYT+Qk4poG+ejAfTeP+
L4njuVINLtEu95bd3p+WzjyScTkd6FK6LnAObRsYmqMPTKNuBAYQVU1/UmkkTDbVWdPqdKK/eWVh
36mpTOC3jRbAZR2ZgagWTouzZrKJJy3oLFoMRCpa03WOsR5HAxoj9RlK+1CbcenWKIRzJ4sXOOT2
/RVzUZXyjz4hhdnLznf4dQxq49J7MFM46l6uYP2cKC66AAIhsHeZCd/PucvSZ5yKKOhkJ2Iamts3
kFDXAEvmm6R4NDzKpuriYdyE69vP3DmbRBOJJG6+wlFONLJyrS8xnyDBIZ5jd3ta54cfcL2jo+hm
F5eOFJGgiSD3UHN/4wvVY5FS1W6FgJHu8qEC8tQsW7m7rklX1WJvCIw/95X6Z89xxbjdmIYaxfmm
zRuXPeI81t/LKuC4L9ewkW768Kx/PAUEqUhD1HmETYsVAYdRvU9rB6qZNP10hnR40QFuzjUIUdUM
AzLidOkzTHH74DveRwO+aMXw6t9NFGA9y2hn1u11I2IPeHIHi+981v7970h0zvcl+5gEP2vSx19u
N7TLPpDshs9yDV7KaTEHrNRjyv+2aaSk4JChA5hHcggV5w1jIO1ULnwOtUp+Ew2j24H8aT5a3Yll
bjB1Yp5B++gUuSVWoqrlnauS8zTiraR9USqexqb2EctsMwrazdVAG4sqNYc6MW7zaQbTUZbK4e4q
4hHr3CkSlRErTxphLfQTvEWz9fgRVLr3rGmDe7JMVkM3ka8yCDXksQb26d1JgVEHJg1wwsSMjGh8
CFg0nzt1c0B7u7V5lf/wzn2dM+wGLSc+XorJzSgJOJtQ8vYjeqxHKOqF4Ox19sXZ+ljXNN1sSRwQ
gTg/eXSQ4zWHmjunThv2Z6GWzFG+RN33vRSSuYiwMJQlGIzzqCIEJinB4R/vGIZ5+qZ7xlezWuoc
MVcjRDciqaD9fNF7veTiJRpU7fyKIkEDbHB5tGC8/ksjPC98fHvs1vV5PRFHdbIAJ+Atda2MAzU1
tWQmyAy3YqxcqxvQMy93td1KSgzjlRcfmELxA4nRB7cDffw0M843CnUpYh/Sm9fwiLF4btiIDVuy
m0Fj7jGrRCYOV5lj5VhdSRzr+9Q/ZQCmsr7dJUSNl7b271FekogeIxCl3d55dD+uMAXRFW5NRd32
1Ptl2ycgke4MXdOiQnUNnSKXcwEXDKRm4i5q2x8KuM5eqpodOcs2wPc8XUpEAk8T14RPyYbCRnB0
qQ+NhMir/B/KtiZDwFR3Auw7bFXQDILhdOhCzmyvb9ZhOCEpW92VbXtFW23xBDHvEubbbOef0mG4
GZp/9483bdldmCLfjiJ+687pMA5w8dw3XrnnmkMX9MTtBt9ZaZuPJEQE5EchO03BjlWkOD7mYXiu
FUBQ2yZWpIwwJCkqBSobJ7AbQXfSx8k0DVEjGTTm7VLyDtp07EUlwR9KbuJ3hj+JVVxWfQEkwlh7
hAQKkIs0dTkhjc/bw5JQbZTyNYne1/nOMKysV7+84nCz4lzxsrFJpxIMHKhFieoiY6BMQTDfQRmI
KtwIDx1akGh5q3YwdheJ57cynpnsaGxTF/sqzG9uLOf542CGZY4IyYZTArHwN1i6Sp8fsq9aouf5
S4BpaVSUtfi4CkRkDXEtty5O+VM/p/Hyy0uD6t4j/OJBNxxLdmtysmcs2UmHS7w0+J+Nm7xSNKDE
nuKgvRZu0lnSOC3MMRACIsajg41ahwitj/b/BPSZ4nova/Gznq7H+yhziZK0yfK4kZ/CB7fR7ygY
LaSGey4wWDNWxoqFa9dRw8DB/OP3GOGLcPlBG7uq0DB7oF583RBz43pd4fTPzY0NKxPOunuqGAhq
wvvibXJGg09jDQQnvEOD61MckZ1B8rcpBnzVnWTr8wPqAn/4jkP70/pa02KeqSVZq7eietc+I3gu
T9ZcFnkHKj9CWLzA/Ngym6oeOFJav9/xsOf1IhAhcZqIsyp33SSbWq1p/EX1Johso9eq+xxAwbAw
dopmCuaBNhc9KQO8ELs9yjiXZ5JoF060yioRQ8no4l29uJpL/CP5pdyOBRhNkdrRvDhcNfCnvhvT
1YFr+AFBBdZ3o4bVcdD9g54muTLWyiyJqK9NgY/yHupmiDENYuPN/hEpyLP+f9cEJsxX9UxC9fLN
bg4YUQJiJsTdFmksYq6MaUkthAzt9T8PCLV0+8VQKX2KyLGzACTwvAPSndAAcpfMSximCkeQ7rS9
9OgfwKvq7y3NvU93sdIlhZxho4c3ZFKI8UpWN/ueFwvphBWAR0BlG69dBi4T/SloA7O0tqazN9xM
mcLOJxisM3eL9YhGbhbz46syz1UIUBSKS2vBLk+Nz0tgczNyV2UkFD2lC+DIKSIOXoJ+uNJnNdDs
Y6IOJ3V07ybUP5Il80kR14BMESC+wUWnYDhOTsUK0qaMZhXhkZ6THY10w6ZdXTJGvuXERFjfwKuq
pEqTdBr+fw7DqC3OUQxjp860jiHKi0rWUZ7rJyiJJEVKv1Znuv4ggqDQ/sGCftGihIQZKGPqgIs/
u7UYaQRB+YM8Bu2vfC5Y7uY5Nrc12pxGmWP4RZxs0cNWOure1trx3V6i/TOWKlAwbo7K5RBa5SFS
7dJxE0Vk/tWXEp1uaxy+uYUd3RPXUjCAU2ZxvT5MtPtnAL5HemyNELIdY/ex0TOu8YmSg3Y/h4b/
lZ3kEucqGVmLG5mNI/T/+Y4vHKXeqXJ+/PH3AIEHWBcJ5UsuzqX60WSRmB8P4IOMYdOuA88vrsBc
2F+hC6kfUsN8sNQfNGVEdHc++fPUF3U96+dkdkQpSYJFZqnD8zZn+cmD2nMjKHKViApRfBioj2tF
c9bEtZD1SM7oEbDa/pAw/h6py7tRralKH03tX1XFlkvXAIn8dGWLhpdYcRd+vnrYp4YRuWyAfuJM
ItC8lY3GGzaygAjftrQ67z3gSwNPQrblCs3Cs6qcKDh+xuuiYbl9YZXthaZxKLMAq6XOVrXFVJOE
bq27xuHbp6dcGuYsws2Bx99RGpNRimBXNamLgx6mMLfYAI6PPseoMAVYlYgukktSwEZZ0Nj/IN8v
01jAcCjATOxprx2Ehix2iykE8wOmvWkkTV484QG/Wp631of2KBogJNSjqahGhOuWGgJ1QJdXqhGN
ZB09uBWFg5szHeDw/rCtWB1pJUbre93nGAG+4iihG1VuLUiAS/odJ/QafthhILcKeooMvz8jcnZ8
vtjES0WpqOcBBwIP/Tqs4M+asOd58/enSSmEjwqOVx3oz2PpK4JUTwikEwPXf4ySvI7OHeUYgmTx
oNzLwGxMVThp2FbqwlmU4eUn2IwvlnoAhW8IREaA+Z1x+WXLTMSINNhi/NfqP27q11YmsMfpdMu5
q9ymq0kGAc5oOrLXHpobszMNUlArhloDfSwnxaMeJ+2GbzAj+naiRoR142520zuycMZ55xLsuwB/
0SeCWFzT5QSZR9Zkdr8+4e3NkZIboR7N8K0prOTpn8Nl5Wu8h0FQ1SDc/Wg849ElSktqATKtVD85
NCT7SoxbnNCDPsKVL6og0TZv0r7LetZwMdP6MPhHKrGIuOUY/UkqUVVQSz0AD+kfw3nyBDzs8cq/
RIRqnGfD/U8tiWVo1ChsENC96phbf57WzA8+mQn+Pa1Tmjm7dNnsXa3gb+A1GglgN3t4G3a7j90W
4tp8bliP0cDWgJovJ27ZrGwVsy7KlZ3SazfRVHXbatVX8uNBDLYhIjtBcAi+C7PxyRx9wiwVrsky
VndOxXnk0lj5Z4ZkKzY3yU57HDo2Uq1Y8NcfVTfsmWDjyB+NlSwvk0SZq6YL3YZlCsJB51OJOWSj
WLObFgC5kZY2X9J8ICSmS3Ya/psHKHpdWIfaIwl8vQ3F6D5gZYmocUCJaA8tXwYrRA6DCsOs8UMb
9LBC3avysBMuPtOsfwURwYS9aFmQ3B4d81W1RH/tkM7TWg/i3OEnB56HdjslwW7gcnIE1HZlWCfj
NyTKkCmvsvPpANmextuYKkKK9sKhVFhFGHYISRpIe+LGZfQnv3FUqQHZiy+/worjx0ApX/M3jeOu
AiiCbBNAH3nSBmpt73Q0BgnJi76guS9dyk4rJ15QWYKZdVMC1ttoDhlavUj7tQSneSXVw22ofW6p
0PoNQFdYhcOXQnDnZRpu+nelq+zGlNtr+Ydl4QKNYV6J3G7DLAutoFiU3ZZxdXENPJR2A0sUBU1p
MRn8+BHl6r/26d5r3Z6r1oZGIwGl/DAuHq8cN+xsHD/HYBF7SM9WZLr4j1LD5qO0uA+KpDa+yCmZ
+sgb+ewbKhU7pPSKrHdiuunOOjQgat7wSD4sBeeA0vlm49aCIpQL4tQd2vSb1baQ4ZrsENX3NTQl
uhJURMuchV+qLyT5SixVA/EZkG5AHSxev1JYXVhinFUHZ8nzCf9n3iHM/hYRBNv/tD9z6LsCy9RC
ohl8ndfhGpWBic5qj8StZlG+ep4J3j16MSD8wokA5efZaJp9V1xxf6D3InnDDHQzwjLvBdSlztqk
QKA7my/MjvU9s3B0hoU6+XlGKh08emW+xX6hoRbL9NpPWBh1iYPnQ8u7DXeNQOeu9faBwoslUD4K
kE2itYKOlbucVIzIog1caNM4DvHUMaPKceoBQM3L1q+485ixhPtxCQDK5noXIyVW86+WtzR/gw+4
tnMpITbKg+ln0WHk5hYbE9MOV3sKrwt7FTt6w2FDveHGD6khFr5EJ27QnQMg2jVkijnk4Q/zEuxr
SjkpDtPytDZko98qcA2h3wXdQm1okZbC0Ml2W58DVhJ6nN8QpsLQJoZBtD0XNcaaNSsMkS877MOd
VlUFevLpyzDMc3IUH+1It7W7IaglIj/xJy7CfUeaHR8FMRTNEfvC/YSCbqJ1hIJKVwG2yDCQI/QP
wASKqeeGFpW7uNx5xBVd+1duHNgI+6jKv6JRSUQwwBfAM+nir8czTzAarSD9qFKMDipClsp3K2/x
KVChefQxgz1DsekHxeFlz+b/QQDtJXKISiE+1QQSVYqM6o09E7aDj+Cxi7YobWiT5KCKO9B506M7
nclHrh9t9HkzkEkb5vJXftyktRiBgsW8oBwlo2RR1Kxx4knd7cX8FjRCwd1BDRpierguZpOZNm7B
8Yk48IoxL4B3obpQb6LXPXAEyD3hNWLFas6K9VIT/1rEb1gH9AXnTA1n2SOHAZBX/EMxUBjMw2zI
3xI27ntGaH79zoc4gX9noiCC0AHqwRVTGFY/gWUUPD6ENC7l4mqHLxGGb17xztkqSZS4XAjzUkJw
rkOaJoXh12nBsCUaBEBUDZXfrlOsJBovFT4O5XHsyVIrB8GVAqii+CqCmEbf5RPr+ky3jmEv9HZY
aFq1E8iYnUK1iSukgdDYYUmr3DioQHNDoe93iAnG5jMFNZSfp5P2/LSp7SFXpUnXscDPzmmoRF+i
5V0r2+2CT7hhP/PnhU7J4uSp1g1YcRHI1oz+aefCRBpb7neNp4ET/WdMaevAEFfmYwWzGQXLFJ+v
OI3rnnMGBzuoTBDxlcgZmFHAn/mJ4cknSkGMbEwyHnZ5btI/otpo0U8B5FpKlPt3hYKBWbK1z67t
WBP3nKM9ocn4nVM91XBGGOSKGQZJOaXAjlRkComJcxcRZQtNZkMUGKBzmjIFhDtVBT8RchLGNqRL
RDXs5RF+Cd9EyPZcQw15q3tStI6FBgoGI8JyBQuPe0en7x/925+ESwMRjmjSOv13jVo+idiDlMiz
HGIaaK0bWj93QoEpREXLTico6Tuu2/J6YlShZ/wqz0/y//fVy4eVdmzHmG15Pj2RWuSzxLRIGEBT
LweEUutIsWdHF6ff3s2gz+EGrcDFMaGdpm3JQCVx+k6OP00++MBHjm8EUYWOw2YWo+/3UD/TpWBq
z1NrQsBIHMzASv5YbuIkeAZm5VQns6GAdLlOgdrrxhMzO9lJQgJoFp7K79/KxHduysRWO2dbuCWf
kUtrE1oD6rUwo8/5ZzMhvSMB/hcL1x3oPMDaBxH0M7WfMrm3eyu2wVAuQOSc7/bZH0TCCUd0O/p6
lpbYSGb3HZQjXAf4g5FeN4L6mAaZqhnLlb5Umyp4y5/r97BpaCN6l3fqedXgQQgBJ1dKAEAfCcJ5
834VKGvpEZG2C6MJkuFHbfE4LXI5fpHB9yieLIBevtEdwHYVi29Xzx9pI/o4IgD1CtmtAu74ANSP
uvP09r7nzWZ40QAbiDDm2BUxnAewdC52JQpDJoE4a2zkfE0bwleqO92dOApzGAmyDSSWd3fYcTXq
bcd6URLp8gxU/zlLQ/opQ0iacu5S5H3L6F2qGSWsGhzU0cPOsYE7y1x4dIKP00ksGCQthhP7Vcwc
5GX5cyu3pHvF2rR/CNMbt4sYkSn39Kt1JsrSo0y8wjpsrPZ+JqBpTMkyW/2QpTtr9Nb4DmDESIht
bKxbub2/SP6WXKqVdNkawmTXDo8xVKZvCO35NhlQTaErW3l13+pvEljnvYpBUK+3KIkdEXeT5ZY8
aNhKGXrPIDWQK+WdnckmhTIFiYGDbjYc0sJ2lHcmzYYPn8J/mDz/E8e3yNShG+wUTkiIZx+ugn2Y
00WQPPhBYxrgaErQsNkVrPtVGvbbIfHbw7uykuxLOoe9m/PI6E7sGzjeX/gakwKJfkbetnf7p3gV
qLPVdLwvizPrPtGsRIkiWy0tdkdOQeejONE81ex2ia4Fu4wLIQFiOS3534gKkW03ihjQ1Pj0LP7M
RipavOcywtcJgcgwyemNMgTn6u/Xs/lU6ciOZdIelkouUZPHw5lwc9CQEUuL4B3tG/hT+SmdwJB/
jUtQqo8T0Q52QCCOSJLo06TGq154dVDUnkf/FbuUJ1Nv22+o+2PHjVbUn1bX/0IX2po6ho3hn5Vo
7stNbWTPoK/6z1k7rfVoyPwGmJ/UFg44dUOiS+5tbBfXEtQzFMc/1l6Kq+5IyIm3S8HJEXDqqdXU
7kU/nNF3gwjztO6pYzBaLVf2dOPcac9tFEmfT/Mc97KSyglF8C7lEFtlbn0HKCN7Ll6NTQX5KM/e
3cwhQHD1lVta/weINAbh23bQ5ZSnzKKeETaYktYPYVFoOOjc7JkBn5oAHJ9ICGo3izTmpu3w0QxK
WSLet5sPD91oMUghU0xgqEg9vS0ev59pAgGOmS7yy/6Ar6cV/GE5V5pwOg2UWLSlre/xPzitqzKN
zaE6OEiPce2iIv204tkXu6c1NCzNWPuFEJ0vBa9tMEWxlZgVunFCe6uSOtjiHYL0sM6OYWLYdmcl
0oR+6JXoOQKFWgXlsLPY7CT9XoxFUwJHkFqcBbQFCCO6/lC2gWpweX2lKnI1sGJJgq8GLpjfhEuf
xIgMbdnKLESd0S3twGFf6kDnZ0MDTTtMkRu2ln8j+UQkrMDs+g1Sw8Zai9OeQ88vscKLCd6d7BR8
kb1YfkZFqB+eVm/WlCuEMSpn4v7Uk3jwgm3+KQary+ICv9TAZ0ZQW4o07Jqdp48wDghwQYtfVMya
uJH8BwqQK22kqUDPMIZ+OyNMXB+/OEEmzifFLyJBULJpCzwnBrPI2MTZh2aBBzc5EQwF7J6fev/n
Au9XE+4ugHdcUyA0mTq8eNIpl1wz5saLYc89b4efAbAzGvpJqYdczKsHVKgjNQGG1x7oW6QI2NkM
2u/aO61RZONvHMd0UJ7Xt+BoONYHtMdedm+8+YL1fce0HOPzKI/4o5g8R+rqqIzRN1KsYVRNXL/Y
PweREznsOagC6V6BlASphsj+4MycFvtPpmbPoJYBS6aRjfjHiocXHIHlrkQ/8TtQj+P2MF7TJwrz
nsLSmpEIMaF1LVkAXGhcp8fPccr7rQfaezlqFtJm34dFGjeJKdPHKMpfI5Nush2HTQSoMk6377Cb
H7z5f7VQF838AqYWg6J/SFa5VKGjfoG8R0pvmyFQtW97S6vcsdeP1ZGm2ChxIKTNNadsz439ocqf
Bl4h7XSkzKmbuVJ732py9X+ln50eAzbleqIokd3wv4FcFdY6qOmKW2/FG+SI5gQxBwbMBGVdCSHJ
IMMAgG3wQtZz/EQOs2nwycZFRP0D325SV/gSz85awrwF9ujakZggtF/N8I64foCkBbHgz+tq9pcC
ufcs6YupWxnS35GoFUCd32HTrnXDOAyqkeIHGNAr8AeVnMqdLY0moR/s9PDrjvcOEyZlNAGi+rVR
5cOmtj4s/i/E1MF86Puqwdb47fl83Md5wxsosNowsPhOlyW7FUw/ncm5RdJNpyp4xV+lI9n7pgHq
EvKvth98OuAAo3lZ3YOQbrkHi2OLp5k22UN4pYGngAlOszSi2ogJEOfe4AbdE6A25+EcpKdUwDaZ
mHj1d5ZePUNlGkGlFWYHXTKD+ba8kAKJXmV3Qx7d3WhMr9674HKnPiLUZ3teFp0WLenkaI1CXQFi
IPwynscGlY/rUNlJSEa0v1XbZq9TsNF4Btpv8rF4yKmTLhE/jD0hImA/a4mxOHy8/PSiXPBRV/Rk
PKAql6UtzShnbgI8G1zXlM8bykRi9J1RAWYzF9exe41jrvb8VX/46rAEglbRfJe+2GGMiFO7T1T+
jO+J++m6NzTrfWLVKNsAXZ0/DXiteDsYnYrXsonXQXIlHoixDj0RJDcdQi6xkMktevLJ9rZUGwlw
p9bxLB1Lxae0EqDl17V0QO/ti3fkgTRQOG+eB9mdu9pUu17lmrT95jvxGlADGdH14vPD4cDC6E0q
HhZ/yPSr7Zz6cxN7a8iJRUmGkGyW8K40U/Wh7Abj5D2lVfDX9fuhjFaP9t+UzNxA77cS4rQxnx+H
06qIcDKjv52cKccEP0lh6ao8lByRcYdX+obbn9yLsn2Ikb0oXu87YTaZvzh7F0JzfMonFOi/NTow
y6UPxaEbzRJSjxRx7Fo8842R74E6SsaWsgZFBYI2w6XtmmPpn7brein04fEm07fsxXk/B6HEfkxl
d9NNRISXknUFzlxaLvypyih1uHR3GUfoLUV8LTwNt8JdJBs5mWFWiQ8t8525d2fEtSXxLOyp8hFi
WxsnsQ7mDL4bkqRo7hk6srJERQ69Ejh17zxzva/EzqD8yDLkTQXUR/QuzbbRfZnnTST7vOESmxbr
9x3QcxD7imvJJm7QjKeg2jCFWl5fJqEHhHcpQKC2MXyIQBNlq84wQp0YGZhQU2ygiEDRATuPDWCb
61x31UQZ3g867jKWkzL7AbWpWU6rknW8phqEZO6ahPbkseDMYVz9S4YGOlv86QV4bF7aUq5ZA0wD
OuhI/tO8wT9HTX7xEvOGPc0GIITNidnvRl+HEEA//BlcUg9M3UuiJU6F1DiwHZBXNoVwAbTKSLWi
Rn8ecsl9o7PDHh+xE4ZeMQvhWpKRvjmQE9S4RDVFZr5WLKlux9Ti8asipNVCGkNYNonHQ4j2Mgkw
G1aTCPz8ZNl0NS/PeI/iIL2D8+RuMbXUELCl5K0HB/IxcQPe3PcD9gOMqw9oJZg9Z+91wP930fOl
ASxn70o1TNnjTVvGXoyph49E/TjzcBFi19jjeqmAKEvFuNdXW+xWn2jx7A5vveu8xZGAl+0FOQzQ
A19dM/tL8D2UPg7Ziek1pW+6Ozw9f5Mpog8f+ZA5jTkwObImmgB5Amf5ozzozoqf+VEewf48bW3W
1AXhkdM6xjmJg9tZq1xIIHXbm/V8YFUv/nLL05kznsy6gl7b3t+Y/9i+Wz9J9DXet5fX1rAu8XUY
KK+V7FoNveEeIiSRVaWMpPn/sY7Az0cVQ//MOpbrIZJqEfkv8TkPMneaCRb7zVd2iARd8rEgqToJ
xmI4S9LbVHllrJjay5EmwVH55cpmAVGEbZOlF7ahkcUfFAsTCSGIt90pWs/oYl31XPswnobyLgpA
dJ8XdTJzXH/41KHAJQQPnC94K+IPnoS0X61bxBPKsygJXbnbg9zDfsdeMvuOzt/hxQxhhB/5Pn2X
rcK0LVDz+G24/chn6oVLTZpMiiYcPdqyMWr2dBd0ywNicaCShx2Qn8P5kxiIS581KRVQsxpXCcYt
YjnkLbG1tpwE0Txs0s2asXxGIT6NNH3v2FCQntuRGvl0JFZjwWkLrgdOUfv7vyMtYs+l3OeqH9om
5TPiY45LJN9dc+KGWNZONjdFhdWfHBkNe79zFrwra0bHdc9G/EEGcJSF1Y/z33h0bGwDSGcZU15g
AYcba4zI1/hddPpdgygLiRly5PR/7kOkeqA29UWEAze7C9BmsHd8mR6kiAmgVYL91z4jXb0EEU60
8r+3qQnvJcjduzNHd/obxyfyyKd1YzC+ASER9Pxwuxfle7hgivwcArMydz30mCLrya95Q2EWAbUI
Da8dL8rJEnWwcmzRC4u7ta/plHUey0vYV0jBCCrpXbT3NYbPmeP7W+DkLdP6BTBIQv1wXS1On6Ns
+8hV+iezNea/jVyzNHXB5sLQ+huBo25H7ZMdJuq9PRCIqR3Obs2j4yuya/LaL5yz7G2fbRdWld4D
KzjbCwGLh4+QnZEOjXiMSr3cUcpa+pF1b1PCOIrYoypT01ntmSNFoQtiSnMpgiPcqBQTqEf4qbZ9
VyOtcOR6XTifHSQr5b7XBhBNNEpSUAob5pBUtR0wAYBh3qhbSbbJL/3229oJ7vdT/iBbOE11obHY
qO6LFpb+dprkVLi4nSHWIoLdZv995d3eLpeycgSqwLi+bSLhnSa9Q1R08zVElrxbM7zJxFJ95Fuf
uAjXnI11oEmSmB37v6O5D2QFveeHZ9NK8ORLZHmXgiW2Mv/TOIpmzK5LUQ1IxSmsU+nC6ZYui4Jj
vVXPqRweZtE930UCCIks7xXqL4ADadhs+dozW3ZwZo+YjVLACL0m+r8m8PKYdBnvnT5qGAVn6fZI
5Padi1bhDUryyncsZiYXF9N0S5KGxmaFC1NR1z0CUdMPQ+H6ACgEcvIjFqPqCw+u3R0mhrl5QFD1
6qlfYgrd8lYwagnUiR7mrfsYGwI8cIS9TGApQ71dHa7qCvoBnQ51usHmiuQGGghmflsLXByKuEl4
TuRuuvMVyDSLdX4cgzSC6vJQ9B5+J8OMbqN9Rnlozb1cxzLySTJgSMOm+cVnoQEWWGarThpDT5Yj
ErtZePzB0go3DYDKlGuE19jMwBSRqumLCA81zFtKe8bFfauzuGGVaOSwZXYASLDpGwCJPSkpqi/0
EmC7iknDcDHqDWGl2yowuvI2kStNFi/TIJCxgkluvhjIGgdv+yatNk2CkFf0zGHYcXTUrfgyRZWk
+e+8W6A70cIzeTfa9rK7rrvMM5jb4fqK6KF7zKgChej08tEddFbeak/fXSI8P/JggNz/KwhcMsFJ
JuG0GFNQ6wUkrZTQnrhyYEV7bOjwceyNPcNbNJuTfDFjKr3mtrR1/HZFahOu8mumX5GRkIz9SpTI
hbWyDEYrhpGWdF3JRa3LmkAxVUVuBVdEHJlJB2V3aDT2q6Vdkjue4X0/TtmhwhHnn1+nxhXaY1Mt
+BwpoH5w+4FRBUORW/wWYZa75NWW0GJbvD8XK2aG96kOvnj+o7JavqIr6TTgcbMs7wr0YJq5GZ+k
iaJk6rSXuuaubfDh1r8bc6p/IR5RNiO1lfP/a3spc3EMgH1l5+QKUqHXJOxd5zyTPa9iBBtpkeA7
BL8Eec6XiVkwxxkTjbe8mFc6Qwn4Uvl8T10j+EdhA2EO5RxEMSlVO/Qj9tN7WA5pDqXpOtEAW65f
/C8itiK6OWjcuhkdYfEvYrlou2ySk24q/LeCliSVL87Z4AtZnJ+SS+LZxSdY4LwWbXmwvLTUfF1P
wFe/aqlmzI+tMt0XSy1M9h7scThMartdOOSb9GJokk7/q+uoRVLWhrLKFoqBoB7/B8Y8oXHdeBjw
iHI2dLEtfHaBV8c7lMiKlNqT2ngZjczW1Pa9D6UU50Y2YSWb4EOhvjbhp8MzRVk1tgq5ZZ0GseBw
5MjEr3IbziFGs8ZvNaiNdX3rmMG5Nc9yRFvVk7uwwGQ4Nc8FDqJSD4PFtb5tC1eicCnHIFbOriLe
K+8rM3I3dMKMJkMHOMk746xdiGNiGxn87zDZNBE2C/RAKZVagpBuM3Qa2uGP8AOzyY7Utb4BFWK+
HBbzL1cb2Tv9TyR1TaJvHKVeWO7zGkPodbUQQVEL+OYKvceTCVWGuepbOYXrZGujq9siWyvsh54I
ks1E8+YgNiLdtnU6apEZPkm+sedXQOkogX1H+EKqkepQM4m+yz8I/u8YHlzWDKnc3ZIYZQr0thtO
qcFu8+uB+JfGwIoJ3AifDGgGng3DOSPcLGse7ptIAWiioP2h/J2DK7CZzuZ5kPkG5L26rckhdKW6
50Vo8R2KzTKf/xc1rX06jCEXDvc+3kF0bZrzTJsuEd1K9+E6ln80brUDelZ3O7aS2UYjl7kBz+57
jJsNzd+kXmIdUiPKYYyi67+MUvu7/rhu9zQp6//9I3PyVXbKiKkRYq9t9kJ+u/ShnNCvIUwRKb9+
3Y0gXSc2oD3OpSHy+AHRYt4CeZZJn3Sowen+DvMz2VhsKOf5ZCBseYnaQ8GdXW7CAAosFJgc/j9m
vdyba8OcgESoVj/yqCAnsuNriHLG98Ww8FLZ9lsN8loADQPPLb8S5bdUjmrbAwlY3fK/jaTdnSCU
2Z0cxnkEAm/Qx3vDBT/iPgCC5SWk1rQ4/oYbYSZL2OjVJQ4D5vx1651mFIW9HUiKfdiBSyPJgcZU
xoT3iYnRU+SwoOhzrLTMmv5yj3tyg3XwW0H1WJ9MPoKI0dy3ZGeo0nC8nlWWPZWTo7DhjuEEkN+V
mmRrsVYLJ3ZADBkCl2Kea8h7sgLSpYgZqYxHWB4GKWcdxJ9hOHZSmAHaysp4XHj079tuH58s3BGg
i0hVb5lavtFWKGEL7PoHIyJv+QoYmAcweS2oLfMBou24OaKWxXPNH8P7cVfsqhNFbwnoGUUq2qu5
osAf7B8Ei0zPiVKL2PCaNd+G1Y25SsMBy/mdvi+737Cw5hkVcq6wZ4oUvWPF7soQVxsOBNCuJq/v
/b8x2rap0PJh2tlGeYVu+Sbzfq460GN6DXhNW65ePncdVlBz90xdgBegIvLoUTgX0YnGC0709tgh
NUrjfhSRBHzxvSKbFWwXNEkmAmn8+RTdTtVKs/p5S1tBWMxYcvs6SnJcSKzx8Kk+r+VXY1Wx3Lb6
CvA/L3yOA6dvyRHQ7kz5V8tI9wTE44b4d9GlrjUcBCrbbXYqTm/6D2+SmNXunuSJgk+hF56CkiWO
u9ec6hW5c9Nb9wKTRRmFblgW4c1Q7cxwSh3m0l2TB1BV4iCKvpKJ+IA7AQ5IUo6cUEI7kycxyV9X
U8n+t2SpRMpaBKQmKOEL1bO3q9BL7aWjB5UqwN+t0mD1oxeCexR4q12EOdc8/Zzi4cFBMDQCm1Lb
SAAm4XTXOjlo3RgZCwhWqvfm3gAPS/PV1xOG7Nu5EhXq+itzMKcae69xednnQY9YXMhkkdVIFYB8
EeLh2hyrRshSSIeRArUsAwIHUzieaEgoN4wosbUy5lcZohn96MEiU16e7O5YD6BzY65MRUcjNrW7
kniwzdE6MBzSw6aPcy7VwuaW/pxwwJYpCVCDXGlho6DFjHj7NdWb6xh+nLaV7pojtTc0LxOSsRKs
WEsas9tHKwcPuc18akzv/elxU0poKR6X5E9VDRLvNa2xyRj+zNnD5x2TaDkgDhh2V25Bjjmv3t9F
bGr0Mpsxj+Y+gQ+3klCkOjqnRMR9BhPFyTYwUMx7eQYrQbJKJyRsmN5joxKeNHzr93u4UHJWrFb7
rqYCUA9OkgW3cqcXa0zWwGui63GSk1/WhzoOubhKI/ITAoEp3QW3XjtnBn6EMh/NXWC8aOiH2ft6
Q5X3Ib7qCHTfCl3CDkoAvkcABFVX2p2ibBW3PtiY59AZlZJ7sA+WxY/fBbJn5UNW8IwKo9M2dLV9
nXk4fD6RkFA5+eSn8krPMVfeXttEOvlC7e0Ewsxgp92guO9dvHSV1fUGA01YJjPUegvb7I9ZkFT1
sXkNZBKR8jGTX/Ers2G/SZWukwAfL34fp6CiRgm5b4fbqbQWyscqbPUB2ytkBJuo8c/URVbg9T/l
q5R7n1s6j7VBZ5OQGkeFDxIiXd6hkn+OGbg2RwtJJ4QJeD89NXYkU2bstjy0kKfOVYBTInjukpOC
L5mrwWBR6L6Zj5b+OzwGO9/Dmsq0PG8AxS96BM0qXTGmvJRMH3dHzyuwy4qjStfBAcufvMDIqfzS
yo3UPK3AbS3o0w+7jpE/r/DAg9rGFsnUemmfosXFufTdwis11l3b3H+RAUwT+m8EDRkq5r153IQY
D27oLfOlF7qKu6mFYIUp8Q+1xBMb7CJ4CWyJIo+VyNgsA7pAtii6rfWMJESlGcYvCIlOAaKs8Mjc
Wt02Eg5kOcH0rW3nfwgUzSgXdgLUPlZnd/3dmuObO+Pb5Mepz+635hWMHqXPZRco5rbwC9EF4sLG
kx1rKhWrypeUjfUyHu1ZrjE88rkgL3TW0rb8IhfyE2ZjhQkD8n2QAjKVZWRJDYPMC/ie8MM8n3S7
cBEzqJsyWU8vqyJbDg4erk8h5vSmqX8tscsIAVlnuVrdRvdfHAN3ncOms7UN+MUXbKMA+pTDqS4m
NrhoutTYYKYaB7maHBDAW2IWd+WRNFh1IZNsI4+QFXm3McygKv/MacWsjs0Cx17ELp5BZqnJTUtX
uR6rPeW92luvNjRB/11T43UBbvWDUpHs/LeH11bqFQ96dwqbPfP+kkrBZ9Up+4hHksEKVJXCQq8v
ItRM3fRZtunYGicv55t+iXeaXaVokVn65xw/m5yaBX+u1NRb2nXdRO30VSwcbMaJu65G226s7n2D
EAMQsif/+jtGlu+4R2KVUoftXancsGHRwEiY3QEIoKF4sSysvlAkek0aKXDgYp7FON7ieIA9/YZw
uTcC7ZdSZQ8Mq0u3Bowb3g5BCf9P/x0h2lWqdA+ZZfw/SOBYFk7CG09RxJRMyNByZOszLUyyqbbs
l67+RMlerkFLNtzJz60ujxWWVSweuCF0khU478DojwzAJdD+yBdoUCCJkW9+gQOnQRhNl8T/wR2M
GDT5S2wDDtMp2PfPSFWZT50oKKcW51/yCNYM7H0xFC+fye6QpiEKrtEj8VGFV2B1/yzw0jKH5Kq+
t7FWavKU31SI+KD/bk9gCn8p7zpziGhghKNwku7oOVSEACjybO9kZEo8ZYSwZln5W4WTlRFincBO
IPR128/KfRgGDgirxwmE6ICJJ1h7VtYCKd80q5g3EP3MwqKl7bqdi38XSjkjVjHV5IfQZDKkqjao
87Qt9Rx+GIEmk1jE3iI8SzX7UY2pMYE0/mMRLbAb2vXSKdtl0rFql6Nh5SmnJgEB7/hoJzflJOXi
RKJb405YvJtsLc8InqB35k+G0Z3mFTITNSaHaSX88BOCY9XVCinJCge/XqtzQuVrhMzsTKZCMm5P
zkBZegfu/gYexvzxhk/oTCewalpA1bznl9LkG0y5YCgYfr0fqu4cRpmhzWSZR/Jns5JyDDhQqSg9
eUXhwR7LcP2AXMhAVzO6fr9ZiTH/Il85IQFvVV4ODsE7cCcWq48TIAYnrhdsNHSfeT7hIOknB6WO
gRvDovW6LekrhH8kBPoVIYfbKOmIPeDzeDOcK73eGtirTG8A/j7ZOp3a4Qm2f3akK+34goei/4mm
6imT1hg0PIFb8iqKVCb8o45kFtPOXNfKbXsN3eYNKzDDR+/XTjvRr1yUiypggDZsSuGF7AzGEea2
jCTYMivuCA4qzU2gl/FB6E1ugoAJoxHtToYitoANkg+a9yQF5nhRxDX5xtXuY153YoWSg8EyXweW
d5IMjdEdGh43e2W/RaCCnPIssRkMqw3bMmcScLXRKiCGXDNdLRss+eZ0AZ7R7Zi6sGtWwse9vDEm
kbQdKseeDE+nA1fTLBuLhShNbC8D1ZIzmhiqFEZOjBmIDkolyi2i2a91uAzOxtMe6Ueo+ZCHiaQH
IoJq43LoYMUdSUB0Vu++hwd8xLx1lZSs+FAm9Alr44ur/XkAaLpC4vBac4IpkUxy/VIyDvK8Qoc5
J5/DAfv1cbTOSFtCZkOfSZrQowUIRtIUbExev/MUzeXTViJlgqlugJFka35VnWkBNxOGyXNfMQIM
1A2mwDQNxi1JntTh1DHgDb5Y3Kej3JT8JxeCNiRILjK1IadPecfXuGckv3wz33a+x7Hhtu75q1Q2
UcpEa/aUeKPSayWHeTmZcGlaBRenJml60sGwduDlduh2DF1oCkQSdY56JIlWzy0cZX65OlQepqbK
wnyIqPtVrXUJgndi+I3N7mOklF/sTZsE1pk127oxilLmyY4nVHbBErowg/rpzj0DpjYJq3LHc/rX
9PiSK7alWkgrQrAQFtArfY/Mp5om+N5SUfbC5DoDvs0fG0PKyU1Y/bwkRiqHM/MN/dRPUqokFMCX
m8nxlxWVItp5xa0YCT6EHlneEzk22utERAc89NA+KV8tDn3+0FLvhLfWo6n7vFGCUZl8cZAOkO+u
q9ZNH9gSOij/meDvP+kdq3qOcllucbpB+CNHP55LQt7Z4UF3hvy9zmCqM1M08b8unyk3WARG9avx
t/BJg4To2Lc3WYRNYpzZKLKfxPViXtEypKyToQS9GUBTfxrzM43bG/Mo3rY74r+xE/60+3MkFSbr
84l4Qn4kWO3gJfbBP7sQvQZlyOwWfId2OyohRmhuXAHfrpqHU0KYhrI3Azto/t6TvkNXvPwBCf/n
t3NKjeacD4WhIOMJPvTwlOreLvGP3xDuJET1mKiQLE2MVAe7VmwU/MVe7DvOpOLTgA863YpR+tOV
mqx4Tkx6O/WTvOxfMtWCOVFOcd9JDhvT2cVMKDbsmtNAUm6IbxOUgOOL1SGG/KoKDiKV7CZV1+Nl
SDxYc3JrS2aci/pnNIrX+wpoUlZcyReZTmiX30wtzfyauXSJLSv+tz/difwjZWpmXoA9n9NIBVP4
oI1tNR3PHEYJcD/8OIeaGuY/56buT1mWw5+3fIF/ZTk07c4USC+uGb0BgcgQzxIaRCExeVnQw4sF
yYvI2fR/2I1aZxn+PPseKG/JysKbIYTpk+gY3X9WOtc+QWk2EgO+PYLdjyKYZ8P5NVcT7jCeRDUL
D/hInQ/N9I0E6ZtDZTxn0GkzmXcwKcxwtYTB2THsY+ZQ9KEFB3EePGWLOBZUotx/YeSkLc7Rfj9w
ZFpzHo7BHlepBC/4Jzs6NCazOVOXblt1zKm+VHi6T2yyApOXadCIVUSYl14+Gm4cJu8Yqbh4yhAQ
PkA/VtQH8JVIZ4oG+chCSnWuw9RwN3347wfK3BKMMEhZHVNMbEbuZqTVpx1mCr4f2Bbvr0ifovsL
HC8GIlqVIdTEWeshvP9Ha3Zn9pe8jiRmbJ2oszWOU2ElHmmYZNiEBdnMX7K/FLVFF2Pcb3D1292b
vX108Djick8LWeig1Ca7nGLUxgomDsMWQbzzRCB/Zap+cskGCjSv0IFQhschOrynlWIITSLi8Tes
CSzwKbD8UkzIHF/t1DTm+KOTEDGv7JsRBnvyNlFTeLx3IEnohn9NFH3yo7NiVquzQ7OWBdAZbnNQ
z2jEwecLkJWm/E19juzBDEszgtftrys+TH6+2An6upAx9maydqWuN/ciZ+bXXa0GTLWtFPhwV8XL
jaOd2OtvB1qzEdjGd/iyFTehOqdxuG6AmcQocqk/BxJAoKKBxS9e0EgLFCq1z3epdcTOEmHAHxnm
QaEaxz1EV6pCQMS0Wd5u3zld63SxVj0pUZk6Btfy41QX3IdCqMPS6OuY955cJOgVWvmof351lZ52
NV5HTlhydxxE1QvDtYKw5FERco2oTFo+EuYaGXJmnGTRr5XXmqNvYG9XftnebFgtM2hAMjQhdd3h
pg8Ora+ANgAdyjQmk6GN+gR+i+h+xThV/heuu5nzQ+JHoOpyGAi6N4B3Yl1hJHywKnGoL1ttJp6j
8kIHDtHK5SEfHDI/OddqSE6oAA0r0+GTCl/lmgrEhRBPEKH325E3o5DeXn7Lds987aA9qwWpMyQ4
lcYkYNsEcTc/vbr+v3kfw6p0yID5okWppxhI3k3NU6y+Xpq5/wyqT3gMt7SCShl26sLQvHyTSWwO
FKuftPGUsCoNm8OOOhzLgaIFSdGA1bpBppjhd8QZ0z4e9Ht23aud17h9cWWbUqDsmDMlUnGdEcO8
v9i2UwSBO851s4jTLQRNTB6bUhTBUoqxLjML0N83DtZRm8ouXmYt8Oh0U+c3lhyCKXzbz/N6/yTe
AjJ7OphTznUsuVPvgJB5pfsS3v2mTubAJoJj7ko6ZlCgZczzlR63qT0tAu01y4mXjpfag/7/5kRL
8q//OPT2gwP3R8TpWHli+kvlX9leoEpdp15TaX4VZqJmd8Jth6b69SAgVFhh40BT33Ph4gGJ3TOQ
byR7zOD/3PMjo8ifKJdxixwnnr9BOwvkI0MhSkZv/Qm/LwlSrDZzCJ3sAmwAvshXBY9FSLrNfRMI
8lkh/UWHrk9+LNijbWHODIIG26h0IaC/7p5leGrXPwkY31hdXKIznS36LKs4k7fregjxlaqephkB
w9gvLplO8CEZMiJlsDNZvBQJJhvckcQ49E6oE668jF2o3DqgPhvXd0WALnh7uESOjNKgLBCsdO9j
XB6Y2BszLA22wt34g+E9gA33GX8En0Ql1lq25MaX94hOphSlPvOwHFuLg5I/X7eUci8SAQc/itY0
MpuOcA/4gO+MTNgoVQvX2OScKMflPWus6QBuFuntBbscmp2FGED7N7ENwTyNH8xT/o04QVMdg9tT
ucgyksBl5hCOUI6ibniJEPKYNciAqfutVzGGR6EzNq60599E6lasxRi3fZVdejqQVychSFbnZZ9i
ejQAIIEOtSHUQCpVfpvZQjXQXl0tMDs8+Ax9/vgh5p9Jn8M3y/ueMayKvjB4pfbG3Cvk5j00jUok
P9VQgcJV9/D5T8p/fAQckquJtASFhEa93RhFgz20M/tJxxppnFCMsiL6ey59Y0DHfZcSQhvYkX3x
9ZCrauKz6uxQzurFMFtljg2dxg9ULbtJMYVov6737tqvCgcHLMJo6G5TA6sF/M6sIZGSzn3cQwm7
mqvSJFYZ6PakkWcFKb/MDuV0dyQOcihaLBGcD7TCXV1FpctKJpfeSGgA+3oJV8UagwAVQXk+6dqF
Ky6Y2+QpC5mbr+dEnyxASLGo7gOsftKfhljNedsOfdPzoUAnx0fzt3cgUFKbT0Uuwh5sspN16Ujt
Am40mOvzvqBgtUXC+ygtiGe20ztBqXRffAPPaj+BmtHrVorFzLZBpbjS+iKVKxZto5o5/dVXdSxB
DmVqRMog/fgj/UqoZ/DDOJTnUp80klNQFqNtJEZvVIbUbmcWF70Fb/bdOt3bwQ7DJVetDT/GjCL9
mMv6TaX9EAkQRGGSUUboeElJGrA6GPQF7hMJARhlEosO2N4Bmqn3qvDYoi6cEO/segJzeKBEkI77
QPIAnF3LaY4WBSkiT7jAbQ80lFnq8vOq9d+MJkqhSxjK3ueFt68t4wA6EWguTfVTXp8eSVOCIai6
4tI5FTO7qx7c5Vjw8iwZ2YjWyr675E/e3Vqntnao4CV2BEdYrzWUk5K1Htz6a1S1aBgbAhvSK1E5
oaNY8g85UtBCenQaZQfb2JjENKYQxq48SHgxVG24sXmSP4txTn+4yRcqqxLG3/drV33PNdNOQLhv
Yqm7VJe+ZXOBycp9op5m8AoDwN8o1UKxonrx+siYnlMq32yHf/Nyi0LAXvCqyJ6YRuItJ3sS750L
NQQhWQV2nGFxbZ/4ylSgZc3HurhjNA3WN8TZKD+flo9Ovb92TmjJ8ixk5x8/7PSIcLGwipK9+iUI
bmShy3Swz/cNC9sUC/gEMnu8/5ozQcKrkvRZxETMQo7WKD3XrDwC+VwIJe40iSRUWg8qFjGWtWYF
9dgHB8SPyXADsDe6LP3gTfmnWsBA28sa+4zEwvLaCQzymvEqrCWtikJ4QIwOM2pzGY/iMFvjHJbn
GdFuP/iE71pVWpNnic8Oj6eUgF4nC8rHVcpSCCz0VjuUiFoiUpXm1MvIomjWw7jRikCjR3kLYuxv
OTSAA42ufQ2t3nwBrvtDlLx+E94/DXo7ZoYGSQxpUkP1Y+ZaHQi6Cd0zr8VTuWmhhB/60giUtv31
jAqY4hovnPSXrYKkdZ8M5P0RFu32Lup8MEGV3PIPhBuCl2p+OnyI4hXE8iNrBkM+tUpAAVn5O2sh
2y0r2/V1mq/ENbrLQ4snf1QqKM85p4QzMNZz9U6xiP+jYpHgpL6NgzSG+8T/L2/Wda3DnM8nnj8K
xM5oUdAJdRoqtjalUqvU7mGR3A+jZJSo9aLRSwrf0UTBNlPKziO8SgMM7D6/0pXMsc2TJXZiViqB
rYSMCqsJacEGY34ESGWoOdIlzRszLIjfYWodKoIu5K8VfjAh9H6wKnXsaIAvh5o44lw/RwjCdInk
GcZookdaRInPxZ8JqrknErQkA+iXqsN0H7ikDkawvXIqx1CV9IaglowAWWG7bti5g/Dqf4lTgQkF
0oxXfUXvlLBy8B2I/aBL9vQffkLjHflbcQ4AtL9hASHUmwwaHbeM1Pn/5MsXh6IXMbN4Bwuwdlg2
iu6qMDluvrzRoY6SL4gcx3VFX3ynr03n4o/ygpw207v934670Kifq/ysnR81NDFYMRAQ3QaQKFrP
74TKU4R/hA5hD5sU/1YBxbNydQw2lc6fNMjdYTnsABmXy5eBMzNNXmhuQrIsxI1nkvWTqF0btJg5
Rkutzt+1q3Fnu7q11K4R2jcjg2Uan+ZQT67g8K7PRGgAw+HnKI0eIEgXjKcI+SblPjgLFbCbO53J
guqfcAgP5/K4tX58SQYOYpLM/NY7UzH677BFQl38uu7lUkYrX4Yco1vn0Nod8ICDpEXaeC3d/WoU
AjVcYsiqHIg9wN4Yz+NSqRXmALdgon/M+AzCCl60C8vskZB323Hi9LbOhQtHmRQm0thjP2jl6dCb
aIgGl12BLN4sFaB9aRT5w9WFQ4N1tHiGfmbmPI3ZD+P/9GFUZYVLV1VsiNNwq7dFwBRCxf/q3JU4
CX1yY9jLkXdzDHGqPX9EJpYwao8fn/a15aofh42sTX7tKQ6rk4dQD57sL2K7vE70RzlvnWyiCkgI
2bTK+1DHSHk+FMHcuq8ZyWSlkC4W7MXSuOZS6WmA1NDyvOpqlGYSQcc/5ar1AxWaunoynEjQy2en
iuvqmHwrNAZgjdJfYIdiGTcMVbzw1N1UHdpAHPfuChz/U89lZZloVgXIPlOXXR4gkkWy/wK4nZEG
6lKOZTBKt1b6fS7Z0xgbqEfijrw0ObQXQhIDsr7etP9kI0I9jhBFjU53KrzuWjY1F793OOXiJhOQ
hy2P7f7OZi1CICCPfYLmBgsNySTy9a5HtlelI0By18aTjIJ0jPCyxUnTPYuiU6SJ2aY25LHY2uHD
5Sh/JxYo07F4j/AnGSBAzgJXZSVfyts/p/j2u8Vxxqp05OtaEab2rDohBNhrGUgUhvyq/s8lmtgy
dAWmXgTOzuxMCSif7Xd/CGdjWKzSGxLSlOsWMmEyw6j2dv2d/aRgXqAQHkFMeImGlRCjGKCc9Zsa
/8gIW7TMRML+9Okok53TdgqOUljEQwV+h8h7DtY/y2ql6SYoJ+SgDZJ20RvE/rfEhFgA4LNCuSkH
Ir7ycC6LDPihEgX+jf3sTyK4fDu9EZ5Id4oOUhfTCetMqaXuQYQ4iW13vLSp+/kFF0EKMdHsnnFR
hHZucvomuEW7kB6BvJuM9l301wzHPIPkfh8vIg3oNiyxXRr0zpOgt02Hsp+yAVOS4Z56zD1YA3Ez
7ONBBHhSlJQn9T4U0Q9KlH/8JluRGUWZ1rua/cxRdwNjEIXTI5qafZDdaMDtMPxqhwtsmJj4NgSY
nM7170bAEfG1SHxHWU0BJFRIBjRx3nxvuss+lz0ujygauqGAiE19RI/kgc6ayuSScE5ZxORw7WOm
/tjQ/8PQjxE4+85Fh+iDSR713LAY5JG7taEveGs0KCXSeYrRzDyEWnXSf3vNsjab3Cm6YEHDgDSm
KEWJQJzk2Xo3TPfvtcqtBl05WM/zgawLsN9jpqICxGSRuv4bSKxJucbMU0dagJVeX/Hiu2FB+51b
Kel/4Ou564m3Rh544+nvZvZESowUGxS8s/JIkvx0y6cY5G6iTYjlK2rSWN1gfLWtTN4fv5vZK0mO
th9s0WX9zEQgkfxnlrkLZh0Y4yOP4nRn0O9E5r7Fx20Aq2BvRY2okzadSRNmCz4PE96Xp2ujTW1r
sRUWIlcg8H5nXp7f5z82/YpVCqEYEG7OLngo+Kmpg6atzKZAee5ViyRyf+W+xdbC2gagSKDw6U1K
/vnekFZf27kQjeX4a9f965y+DuCPWSHP5mQ9xD/WXBqLqBxw5/CHF+N1j6qDAWgrzoBWAX/n0mj1
bJvflydT0WOsUYLIuj6J/irrBaamLqwwq52zG+lE0H780hwFdpbaH/tAUt84VS44e1lw/ELWodkf
9JO1NLEZR3378MKcpY6Gr5pyHyy85B+09MbwK84xCP6sGacU9Tm+du87rt7D9kwDYLisp0oGpUVz
7QWGEjxPbqnMpkjg7CZU9jcGdzbXGoBq+yUcBs2LxJIqDNhE9YmEp7m2ndNYmIpfzficiYCeA1oa
umdNiPm2O/v/McRrZ/af3td5CJrM0H90COQdI//IWKSR9OIJu9PPpVmA9ZhtATY1uGthBZJVOyrd
+i8DrHamdRguAcaLV5aCe2648DvR0TPYg01rF50ATeeOoEMlcMOtgiKqWVwbzFWMYGfCxwhfEk86
ZgFOwIHBXss+7CHoalyXJx/W/nsPXJ2xaSJZNXmT6TX7rA+nhwt4tuHv+Xc8hsIuh138hOOYiA+T
VwENkuy0l0o4yIbNS4hGUrehBRH/iyVJpBetAJUHaPOl3kUND+856QsQdsonsXdKxCT3WB9cE2rk
EerAgR1eht1dnnxiYMvVFA0FFvk7GlIvNtTnXd8xDm5sEKfmGgo8owx4q9em2WYitgNvunh46GiE
4nK+Qz+s/qvrB5rZNdI1KK6t1nDfEfYsyJrAcBLRMvssNQlwKZov4Kbw+/mx1v91Cf8D/vKCVxTa
ZqAqfzzhkgPQZIiqE/mywh53RrXRNxQSNv9ElkinI7246ZNXiIQNVeApofJ7Ljf1XF1YtIn7Ofc7
HncuqJ111Rqgxb5YnMV7MN2DiXiM8BwMJWtmOAgMtuzBis0rTtk0YB11LjuerJC4nJ2DGrc8f4OS
yhp9qDwR4Oa+tFiyehgaJXYAA3Og36OlXTy/LKKWSebK6Q0KYkwLMM7u0B1+6DzgjguLZNlCPrUR
xd2pLvAo3kUt5EsMRVw8YwqiGG9wvw7wYOq7V46l3yl1QOwq8tv3c+FFqCzI6Qamq8GZbHrbaq9n
Pb575GOBNKr6yEw4UJiK4WCwSxBTY0jMLtxOry3Bg21q3Q1Ur/9uP/SUEME98nQUUkDQup9Rl70Z
as9efYOLjwnqX953+9VYXg5E+c1RmNR2wcm+UeshWzEmDiey7nu7VlgkUKwPQM80R/Ua7bw4ey+q
bSCOjD1utcHiUKKB9Lf+Vuy3JewEv8v72YBM0DqdVBHOggmx8ftPuu06lKYSK+ExHOIF6/cnzUPF
Gp3vJhEsSZZOt/jVAMFl+e4lf6WxbqhDdjjkes50XNBKZROQIehre9+wLo4Z0mWy7zU3S7zUKMi9
7zXld0VmLVxuAg4GW86yn7N4dNdbCfQiBOn5CxPfuc/lT5D/9xjz+rdMq7o8bTT301z4WXsrahM6
8DgVDt4whpGbx2QCyVv9ld/dNJ8EewJFrMg0crn5tnCzLO5S63a/YSTn+MiofLrXVMp0KQaS1RNb
5YK7dpGM22hB9d9ZrRwPHmR1McTiE4g2m8b9NwMJlnlAPADvabkrfkI68UMC2vDDz3cN/uIYynVN
2qFfY2bDqemh3BX4wSPo5uLj1vq6RoMGAf3H/LWPZSEHTJlAA9RPcC60JEbtCu3BUHQEjewZ8HuJ
p62B1jcxm35+L48VSYpA1Emvo3LN23uXWeLRy6R+eKuJHXsFv1oJ7g1VpDVDiThONIxovOKqhFZX
fRGbwDJyMFT+wXZL4+3gSFiRXSwBBQxVRKoEUdcm/edlwvwom4SM8WMxcrVGCUCxedApPEXt73Qu
QLz8OqV2AZAPYl2ral4fzq+U09W9gkGfZtM9RB7RnPJ9AisAWx7HIk+UHDij433YUzkM7SgG99JY
IFfYgr51EcVNkP+lZ/htO44Yj61oiaDsOIk3PVAjwq36BIih+rZ887z2tfuNWLMuOVCrZ38mBJsM
DT8IX6MzGTzvhvwxH+DiJLhfyo44zjW5lW7eWa+ZxyTIy9e7HZ+VpdUq2/YIEfolqTQRnQyUnasQ
NP8kmQJkjPga8zp5VX6o0GaOTxEVuPRNCLCxQuKi332RqEE+dvn1QEBW1CeBrIZPmUrEXmUndsHI
UpOaFaO3+7Om9aHw4C8pUikNns317jSiGIf66eQiTqr0ED7zrWpxsUNJh/jlJKmLm83YzEsqSvyk
3luPGBod0oAkhyzw5YqLrkDMXNACaPVKLfcpBZQsrARoq/TGeCFLxff2JfSTUszY4mgqCtlhbIOe
PH7Ie5kTB6BnEFkIL5AKJToKPg2MT0BHjdiBTeWYHrJUf2wW102l7bEYEsD7Yo94XMY7ZpnNnAxu
TOcvI0QwDsJwQQSpLjaYb7RN+4CBOUThNtjYoCRWylh9fPa1lmqqIDz+ut2hxiqIrcmM/abWdhFM
xvIoqYI78wyrH5f5uF6WduNWK6q0TzhIP2fddYtQUrmcUPICk7ItMMrEXqBgo4tj4ojWRIqNcG0S
R8SWJtSgmSJFuBS7K+BlkLteksVzkXD9k/vHpzLzpIAy+HEA4GN0bSMK/GgWsKub19UPL0OM8gnp
LtOjvmE4gax6LsSZuafBfPvaC0SSnB+wkyctgw2BGNo6Y66hMdqX28FwAZ9fu/nYLXnCk9J5Bhhi
bhgbJQ31qWOcErMYElURflsJUS5lbylUoQWCkxWtgh1JDfZYvpoCjV7asrEZZrsaFat1wH30Tlhz
D6kgfwWfoY80RSGChvJuvoBJ5v56WayEvLVTUQWEQgGgXosNFQVnB8+2u5GIkpUhvSSoKt3H5xC8
CpXkrCKxSWqT7pMmQoz69a5N/i8rc9s/jLvCpXqMb/AM5Swcbx/g83CB3EoWSqQ3zuOD8gOzqc62
5BYwOBevhZqsLQzjnWCypKrdxSc48Gw+GqxFyVl3EsSYTm24FjOpT0ToeYKH3XGaoU0U1nF7Imgz
cNf/VXSh7fUQjNDd7KGUuV2calJ20Kf9T7XM+gxEIOeRVJT+pR4yJQGb4GhVr3MybgEtDxRITzMX
gz/gL6YdpLMdJU4yH6IWxktLeL1c2LH8uLd7A3HVuTBJgVRNjBBXq8mLFmwYikSsaavSwjC/HFoW
p+06WW01Ap6ZEK2EkTbrwdeRQolGO18w/3IVsnAS/e+eMH4nl3G/Bx5/kkp48dSNLXCxKoXi874S
VwVED19rryQMUjTAhrO099KSo7M4API67Wc1j3g8pAXLMmdjilRtHwJV9Yg35YjvRAAFeF1dZLz7
HEzrD8JdTwrvbKDsCappwDKwZiW1KSsb6MDGV9Wd2xcXdE72aDp8tXVIda9klB8yzrTSsbjaX2mG
O1W0ATi9CjeeGpwMndUPZ49XuYUIMkbXzCTXpzPLtTTYofdZ+ZwTyyDRLWSNaMxqTrFSRHfdZoBd
EEeAg71eU+o9nborRyA153AtVT8LtZTYWIATIYBucjwuaQXPucJGW5Kt0YejZ+ZwtNhQLfELLs81
233vAuLikeApWIZ4Gz1nQrvqo91vSA0rVYqxJKaccnvq8KPrdDJt/0ASVZ0wnwPvjHYWXm87P4/I
urcYmOKEX1HUXYJ84EbieaegJXuAEvSCyKrm8NQXh7eMbNyV4BKKErXE0Vf8zLxCbvnZ7W+QfWI+
Jze4nJgLa8tbGDKEw/oc6si1za4oyJMBzy3Pjft3nNJzdwjm/RvWvJh/X7sm7KhaOzAbMSq/auNm
RhYiECTfM6RW+0X7pwQRMBTVftRr+McWE4MebIKjmL4JfcJVlBJaFExM1/K0tdYzcEVdcRLHWCL/
NrUZ8AFasDhY/tNq/ax1eL+STnoh3Jdts9/pPTtzmUG5EIPBzQpw5sLTyAaFkvXdmE+qHBrw3LZc
nStqQcq6os/DkMYKb5vSVYP+SyXDYqqUDDoa1o79mB1I7tZFS5ikMSpEYz+KQD7YZbghyTbwqVRw
tCBInvDSMV6ZDocEDP0j1qqt+5vpfQqPhDYOkq9TpIWmr4ZiPGs21WSXFxpyCM52jpUSKeXzSicC
bdSzi4jA6WjV79KWjIK27P5z6LCoGImnoQTY/5hKis/DkirUmPOcKIlVekihKXzbFiINcWgyy+3+
tGN8hbKseNxnRA1xuvA+xw0xsTFaXj88TD7jFM5vfSoxEiD9k5GIypJ2UVtzEkg9E0utnTEeuSZ6
Jif7Z6WAkkS+y0kelWP1njkNdfhSiVf75c+KPFNlxHQt5qDE/QiEcOv0mQThLlPaKwrQ3otWf5jQ
DefdDnxCt67DQObkXIl5yNRhCFHxGqg2a4Us4QWrs2oM3vRkQEMaDTegsNgInvTHq+HgvwzU3UN3
t78XJdnpqLZNHT2hksC1cGd1cATCm76VNCUmfPKM/W1YQ01ccALq6s4ryzcfpyL/iQkuRhMyLju5
+qrtLlg6XygIiJM1dfHP5bFr5AmWfXk1xEwQUaNw4cX79PBGwMFP2EjltT1lIuwgRCeygDTU+fw/
tLPbobobRtlThBZiFl2Okf9KNY/f7NMFWfpkZPypxMTn1dgpqG+RK+dYwYiCXc5opgm0nWSj+y+Q
dIFiYSXP73NJdVjnuKbD+6rdIirltFFmIlHkq4tjmJnAl04bjL4wj/f2R5de00BLsERKEwbKB8j/
FAxwCIm30RSvYwsiAu7jd9Ilifws0qCx6abnkNDFXxSd9mC+dgG2vqUWm709nYxLSuvWE/MuZp0/
mBs7nwf1b9miA8VnJb1HP0xbcVIB5Ly06SwRWZkz8g9jfUfxYlNYY/upeuPBkPj6d+3qydllhSsy
v+Tja43imo7m8v8/1z+kvIuPpgyTd9BM2ukffTiS4HlNLaBGSrslqgL/jBFuX0EktMS84vE2arFN
C+WDRKQmJ0UV2lJkcf2tfYPgwSSEHOU8OoNuk8k0DzP0vGUr2DRy0rsxt78xXh6cfn5Mar19EZ6B
NPRPB9/aSDyxWsVclTlWISkQSBiQcnS6FkPp6pxEhtLK6yfnj1eRLEABxy8YEttx07UkBfc6aMBj
K8S3f4+CNw7lF907QnXJ4nFp0UWXXp1hse3AD9IyznCuMG20uK3Bi/oZp7bgtc48NfqQaxu9VUVK
FU33xRERopSScTS4NGNe0VVEIoUkTsBakOt4fMkBgpwsU0VwTmvVhix5OerAqZTMKeUAsOLCJFtI
vjQDWZb4JQ4ISHpNFk6xe3Vls5sXoeR8t9lpWbjyzdpkinmTQvNensCDkjaruMYpCn2mYycNYfyK
LmZsj176UVxUjElOcmCCvhp6OsltFSwwjlc71IS2wOYv6O252OKnTH6OC4zMR8yCOrUCurR1tA/q
FVtiNlumNksW7NiBOVKihAlGt9dDySEhnc6Sf5N1iYrkdrdu2ZFROpMNtPkxfUNHegunCvp2pNJC
m/u468aFpe0Av8jC3TCXn09VqUO+l8hbn1LPs1PANqAgZF+niwu+PxE97UHG8AC86fmrUkmOpGa1
nQPLEairlCX9kMNT+06Zf1Z7lKY8vHxwpZxhVzZmk2lUBYnLRiYOj8FoDZXEEChqh1mmVQXrO5tf
lYQDTFK0XD3NClqs7HvtLfd+aq/wrR+HycUrrbJxhoCqXcdTgM/GOu7PBCVgg/xgrjEXydK5+pNn
0r+dsvc9m/cejQt8OdwBXlAUhnCuGge6qsBaKYQXiSLrVQLJ7Rkz0hWW516jwl5IE97WAJv1H5+B
4tvdcQKtqrL4mFNbgc7NRHhcIehDVcP5g9E4KojwULTYbZyRl4Ov411wtdN4ATB+s8l78Tw42W54
+qvcogt/loQX6wVjePSLThWaBKKskzx+8oer9R15dLnft8rzm+UQ3giW0e6cYQ6oTNV6muEa+c2w
//iSzLfKCPTukqNEVM9zG2E0tseyOkRf7dSPTEpZI92kkQj4yf/3CDH7n6TdHwV9ehbepxlVCYjL
LmD6jfLxAiDzKuHv9zXc7TVpNnzQtSXf8e7g1vW0JptMDXB1xjRW2wSh8E01FYRSeWCqcrNuhCTH
9Jxm9ORPrCZ+Ua1NTL0mIuYGJnog2pPrCgwahJIexwrwkDnxzT0lpaXe8bUCyXt9O7JYLJB3NYdL
X6xk54e4EOJoMapvCOto5t+hWcS+0VPyWXPX8jVogEePbh8wxFVZe6x/MDFGXJjdDxrAclAtNzk8
oMNRrxzZp7PbOk0wnpcJGj6OkXVik08QDOQQ2luKVt1CYbCmu6EAlYpz4FxYF0ggk5NBgWj5MEhW
di/0cQyUnZF8UqW6lYNSRoXqW/Ucf9fAUwAcFhIftnIj6QNN6QEFvg0K6gzBKSN9KV2BD9Ao3Da3
mNlTS932h2zQsFXbnCi4aLAQHYmWxE2pSog0jslxpw5KEj9HDegt1FR/kVHwIHH75LrsRZq6uaLU
6XSli1SxDf0I4f5Fp9V9QEw4hVa3hLhrDr5wpudm6rzejZkmXxhWhDnegMXf/wp6R+RJjSnW3+er
1h6xVquWE6Dbm/7oix4KVuM5vg5FKw7TgRSa54SZk95OMAkLRfDaPKPxBaApaGXm9joUspSKYU8v
xwwWoNwhrY5kftO4s5Y8tSHtUbrbCtCQlC7tLGQ79MoW+a5gweJN2GVXN4/jY2oNmFyQ4pmhWZt3
cdONTHP/sgzzRTLsPBRt51oAHZ2pjk4c+AferxZh71UeRCfYAsybsiRvhrCXWdzIY3U3AJmlnM1y
jOFkTz9C+GYFdsYNG5woB8qHoC+WpfMdOh18LXEv+lFH2mSMbG/AMoIaYmi8CFWQGgOMMGYXHZev
eE45PYog/0eM7mQlM0MmS6FQgJOv4LVHSZfC+DH9QpEAT89FxjJKi5qXnfwBfNSSb18VB6NoIwOl
Dnx7lyIluOGFkfuU/JlzkOgN18Pc40oxilu/bg7+fuOOFtCDhxr5Icu6HuITRiAy3ne7qHxyUCeg
nTf3HwZ/iP4Xhi8HT0dK+UJzXZ5sW6kZsrLWSke3YCQW1o1JoUbwi1DPH0OoIjCEc8d5L+ZB+/bQ
5ar42e/RJpqVBA/whJmk/0m46ihAx0gDRQ5DH3lIrfkGsfk+rpkCiedvfs7azkDnLqX3rkoxn5g7
tNHUAIB40ImLw+ReQOCl3ngMjyuMzrZxNEYepKdAxTq/j3DdeFDQEPyg0mCzWK6XEaorEZuZalie
dlW9R/gEA8mRNS5rVHTuAPwiNbGBt5vEF8yyKxibJDU8gCFyueQHTFrAxFHIwEuf0HPI/a9l9BB5
3pW6adENCv/DQGoUjARjmYMI69KAEP7ZfARHtkUlgMhFWH/OTuXEuR2HEsnthOFGSE/NRKoafdgz
52JUup5w9chhRKCeYflBY6lHxshAxuD1G66k884CCc5zPYM7ho+R9eJVDQisdWNDuT+SKUQYxaYe
oPJxAXDoBa1WCZfuS1dqY/jfzBKNezzW0xUxV8TipXyV9p04xrFYkaUFeb3nVSNE1nRQnZQKe61C
HNyPtVlzHVro8pBn/qfKWvJHD2o1CGN4YOWQjp1FCyLGUyfoOi7yDYy8n7v+OnZvWKBeNI2ccugZ
S03yqkutcdaKNSl9fDZuk5UDul1+HFWlJ0cXyxwmRL6FoCTcSvx3ti0h6UrFqDuz2L/n7Komsp/W
m2vNXsL+YsVPQ4u0sLGw5kiORYv4FvOzQtTriA5BlXOKlNflT2arn1Wz1Nq0LaGiOHk06SKeEZEy
J1eiu18onwPA3bTeJ2ZGyjAjWZxsxC/ZYuv55Tu9iBV8AknxwEVX61ulrqSL7Cgvj8ynVEceVMTm
AcyqXXCxviPsvJKaT35MgJ8rGW6dfoMbboedG503mJi7NkNcrtmri3zSBEXRpbuxwa773CRmRjGL
eqiL6bMx6oAnkSVLpLT/OZE29E5oMr9vEjgjQmnEjVWzWJuTpyFiM0cSnCxLnPI5FZ8Y6MOF9n+N
xzVTsYID4EUCGQp3gTYSfa5iYgSEHdr1oZnZsCMgArBtVI+kDJuwZ5DxqT3fIDIA0u7MoBxnB9Ah
yWNeto13nfXm4NIsmPhwb5M98Zoz+eX0GgDFq0HIa81LIT1gi64vnPnDz/5RMa0KqmSF7HjaZk9R
Y7NRoGp3SgxVSfa006pGlu7dEx/ZTXOXT+QZbStB1rTFjBbW0WMuDznR8ArtNgha/g0XMYq8GCd8
4M8i9DWXvwcNYcQho/tWkuk01JkBSd3Ht7IBGy8I8gyARWpXTBbIDW/f9/+PPe+Uk9l4jtNOmklj
fAWYBVPDdc0mYzOvRE2Op2MoavJG9R3AdyhisgC3Dqe2qMdUURKWr4a+v28COTrYX01Ht7WhZvHy
AnQybqSYw49pIcAcevUd8leA5FEs/4/M3ykCFYOdYsjW04sBNmMPq9h3TsEmAR3HuPqTPUHgLCjj
/pbfDCBnt3Me3XRhQJBlNbOQWJTax7LWSllBNvZ6n/O65jqOzG7BqEzE4647ncNylXGurG98f5zx
lAfuaK1dxzFgTDESsAYJYyABWWNNUN5LQTsxe3A+L/XlWoZZ0OEFD6mAZlfGPvAvJdaCeA5PJZUN
ezWIs/Gm5na0DRxXjANuGM0S/+dGbdn4gPb+U4oXzaN7boiNFvduATDzLEt6ohle0H34Wadc1KIO
A1bHAdn8BjJ/yyhYABgLwnN4r5PHO9CxdjuHCaImBF5FLkkDs61ql/n+vic1Ljj1VNEhHFVbEvM7
84J1AlVMBMfApQRHf4qXx0MdWP0dNEgG2mY5LOfbJVhA+f4hw6ZteXluLjTR67j5vqdn4ka0zCoR
9Qkh4Qx5OV1SbPoE0LrfCpkdnkq51cFXuRtYsliRfl6Wy8IV5Frlf0WB1Jei/UjI8tOPEGgBbhjH
cVUj1Cu5Uj0SjTK5tV41wtnqE0xQItQufXMHbJIjRnl7skxyiO9Cd6Wjf6uM7H/cHcA3hP3fZ5MF
F8V3DNVZIVYxCnJ0d4//wQQPzC9sSQVkvLyjiylG8rLsWonp/ZRPzhGBb1caiIeCmIlOnHbXEtV8
VctMGTF0eX/HDiUqTu8F9nTVdGk176khN6ze4DWvpDeynJmr4cOBZMlX6Owbsc25PCajKxCI5eZC
j7TSRCyEuHtOMv3s/EfrQzOF0rmzBqcXGtTJbynvxReLC6eqk6966S3c+hhItTVAs1dDUmaITpDj
VrIi5bc6EHp+YiU/tERCq23Ym+nnB2dNkWk+QWpFce/FTnwl4lbROo7l/Yf7WTE5N+ndW9bgBH7F
25RXMPav0024tdhNOZlU2SCIYlOXF0JS1+h8bBjVDYdk1Sn4xVkG4oiiL/HS4tJfFvMHd02nngPm
VMFR6ICxT66yktRc2yV0lgFDXhWO+WmdKWodQ29eIqLOdhmSjKBkqTq88t7Uw8cfDpiDZum2Kkg7
s10gwE0AQfycQVQzu0t3G5ICi8LtYWQcO/jqd9ufqDFw3QN16Cb+Ga1VJkHCLg/TPrXRK/jl7APH
gpmzTXNL7eNYvUbJPgPCvuClJ6Uv6cY8k2cH3eB3+hbf4LFFiZhJ0cgLGw7N2G5Q0WsquVob8UW3
SBQbdqm8U7BksaV0lSN5c0R3DQ78JdJcO4UhtgcduuY2F6pddAKqg0q9Hwn4OK1PZ7Q4xmaP6X+A
Eg5GcQqz2DC/oS6ykmwH4jKvRWPDe1xoTuw4DIGYVeGi97U3pm1kdyJB+mZ7FDM2AXGDDuqr/n6H
3yfLPgTPilifVd2k/FJTInerOo5xa9W8+CWBCzy5GDg0x/ewFZ6TWXpgbnNpk2EjQy3Z2Omba5qK
OyuYCPe0OirLcY4ZbYv33TEi+SCTC/EBm8PrjsCsGwmJBZJfIZIy9loMx9kBRPOyM2VBMoCF45c7
WrZbZAavj3Fs5WaKyuONiT8Yri/HnoLTiNMgLx/i+9/JRacUfSpX2S7px+vcWIQvME16KlVXvQku
hJKXerhx7Yc6HkfonRNpl3A3csJIY3cv0yaLIoySRHFWqsoKv3dVLTQYvEY4f1msA5fzCJX1HCHM
XilEwliQLmtZLEsg2hMCbwU+B3VegG65NFqiL6g/vXIobiyk9DU/0kcOEz85t1bxMwA44/YLS+TB
MfBF22wamDP5+YuSn0vJmV38yf8U5vwwQRJK6H6ScI6t//ZTkhYcaP1xSe5NQDtCYPQGK19Fcp+m
peWU5IA1K0PUxQIcQdYNBTKM+Agdry8F6TvL7qEeQlzMi/+I2LVoR17HkMjic7vWhgknM1fMPCe7
+bsto6pqDMwCHUNe5rNvlMTklpdkmgjUG8deCYAdE4GTPzHFoEwaQqpzV0GFsTywZkHOJXzlZDFL
4GUMMFwgRXnxH17i3n2NqgdIJEO9fjBt/oW+9OQpA2f84ptJQaFBg/dpJ6AzmJ4ryl6mCb/hMJQv
loMHN/OSsnkpCBTpwcI4u2ryHw8Ezp5BGgvbHwPu7bswrhGYZrv0lYba5ySYDRV+4CLvr6Rzhp5d
cziychhgWdaXCvfjbrFeGpxZkfQhi+LNhM0oWI/Jon7A00tRHwhm5rv9skpl7lWXQbIQdeXBnCuN
+YTzpIvXh0OwVci0UmnUFO3Ilnl3S5VScr3j3M7fkzaa22bO1Sy+La5cMuwXcc2o13usBbkg8LYW
9nnH31w4+8MKhL7FcD6Dso76hACxGyyFRKUxzyO0B1nyTJNk4v9dSoaLCfRWAhLM1vS99Ky3VFpH
qpxaJFB0Fi9axRV7iUdZCtFOKzGS1SX5JfGB0IyRxyYnJPQ348ydr5aXeEKkSe2sW5hziKrAVd1A
W6InqkzRddStmXDBkfbR0ZDUm+dDXhAylLPhMZlHitYsIF/J0oVKQwo5p2IycFlQ5yOh84yKfDQ8
OBXazBSfCJ99NbSm5le8lQBTVtBg1OJA7Ie1Foy1XigBAGjYD2+bIAnPw81w2UuO+v1TWVi64KY3
4f7m3VVPI7b5ub7i2jaZd3idfXwlWP9QKLEMYjttUKdnaIZP02SIdKAFrTPl9WsWDT3AXvn6o2on
Px9MQvkwz8AaGrsMeQB21k3K5/PbuNU3ImajiBD0MCPi6oWdUJqqk8DQDuTJXeZP1mcVEiX9Idup
KUdIYhaSRXIa4iPCoRkRzqXu/JL75MyTlvXgUfverJubNjPaJizI2oMAfg4ltCl/Sr3yyNtCneUy
4+NfYxggPJS1AwJSQHUVB6ZGgoxX6WdkvfoW+KY9qxwcPRIcZ3Fyctv9b+eW7CCNTLRKEleYa7sC
s657bzma9ZWUPTRYvq94QskiAQBJfd75bw9f8GsPAL08WseItaQDdf2I1OQyjPxreIi9BMAddtwX
qIeqXLPrbKyZ2Kk/PHiRnKEt7SJ53HwKLSMHR5e4YlVpqFCfUYJAfV4tu86bUXAS1nMg/g8rAeWF
IsMo6kzNm7G3PIH08qcfIHBVqWjhKEGZM0taysvLNe7i5wP3jzz4Htu/UFeoDac4mLjpO8b3u1nB
+B5XlstNfSEaUnyEZogdSEsBwZizAJZc8sHvO2ewLr6xyfLziN5T1LGrJjgBYT6F40chX0IXbFB6
elzXeLyt2F3ZkrrVfIM6eTapdP1MSBcnRGkOrozGeqGNPk6+LjMv+CBh2vEio/MgmF+Elo65vov8
BQtxM1MkBPhz4l7NqRWZRSBnDzzmXOGHPQKyCrYgQ/JglS8aR/SZki/yKAUJxMbfTsv4F4QN+IMN
i256KWiT0hhoDsISVDp9+/eZn/fzepiUTsQTUZj/Ix8l3/Drp++xugh4l//7PBnV5JUldCUjVMr6
yxjLeQug4fXsHclCLdzZnx+KPBucP6bKRrLzeznrtONBB2hDiCItPXTz6EvDmPQiVjmyA4saK0Si
o2VfrDdPXXmI0wyPan/7gqAdhUYsHf6BcDWyGlL30gkK47bJ15VK0FosqMyZWLLHuTIg9zDYSqzM
zGMPda/0iHuvSI6S53/a79HiHqDP9GjU8UtvLqI/NOY9GOXtGUaGM/QBm5LrpxTqsdqsX0UlThPA
3pQRhw7YmQyZkuilnuUXnrWqgxSc9XU2vFbgDWe/PtYBuuaV1GMtXZ8DExs/wwIQzKzlCO0x/nF1
8h0x1m8a5dv3nRdSa0KqbCtJtelkZ8TSsBNIIZWH6NDKwvPGnp0S+yQrfi8CV6F8kTLJeSoD+Z8B
9crPUCr0B7gOSVbSfXJ90i1Z8v6DXh2y329AtgguMz374xAJd7olEhR0ZubSwIpgEWTCv7Uk6d3d
qWRTDaEWCaBivkitqyOTWuKFYtz5y/gTo6Suu2Ot5eeVfF7DNdCa9ki+OCaZaN7KkIcEmZXZCa8J
GfsMULsmjkUOOJz9p/P0cc+lL1hl3LhUCbMWE8U2YALkmIA9v5sX2skLQsiHUHtqILcb1aA2fiJ6
LyUMfLk2K3sheYG7zh5mRY/VWdK20fYPCOgP4Wil4CFKBBCyaqdxEYxAfXQlpx5Qt5UrUJIX453X
qLSjR1z1M7Ekkf3hIgJY2uV7cSQEj5urdd2uuMsMGCGkSf4R/v4987rOQq4KZTykx2qH7GoMQOWg
HzQC+s+HXL4tMLx0cFYqU6aJes6iRaSv94Kb6WdYKtDvmW9MKlylB4MsoccBgwfpdbSvWeaLjBuB
8HomM0Hh+VwrvrlL3OgXwLIenI6htGRqpu4d5UR/I/lXwhjE+NCD7Uc8bmbV1Av6WWd4I0Y6YIzR
ZGe3V7OFJcL5VwtViqKfIeHwsZyHUuJWysfloHCA9bGw6NzvH1hHCexzdj0s6HJBFjMMdD70Hd6X
HBPijUrMHUpDorcj+RytLjgN8EXx3xnDKsPduEe84FU9s5SHJyOBXRyT2BmbF7EXnnYu5FPPx/z1
w4pYfYLzcocvOXPEMnmXfa6H3qRV5rkwZB0TIuT5rt3DLavybD0EhrBkEubDezQHQpiti1r8ZIOE
YPx8W67bp+rbXJ3v5cVydqjOcFMI+wBMa1NweML1fmps1H7S7gbhF3xqnIMBCMaCswb49ukcnU+r
1eu5LytZ2BOwMxckZCKiRr3Y2FhUgDPtAhYf3D2B6f+PNH+FqnK9f3OThFseqY2rq+R0iQWFsOlQ
zJVA4GzO42ZD5WXkhr4XpVVjXgaJMJ/+SrYGnfuQJq2P6pbcsUPmuxIcmY2hFPqNurpdp7JiFUml
b6tfIQA2/nS0ZPMUW2IKuvZya2tP4pyuBmE3cObl589l58caBuKk32pylGvm+lTTuvjC8UI7Bhsv
y5Pg9ZG8HRMEzE1yPLt9zJguLMXuP995X2MW8uxQxjdWIRW0DwfT2uXekhVW7msNkCi11s0CEKX7
DtBBbcQ5MKcTKz11DKRPuIiTmN/n9lXedP7OUNb4aHB6eQ08Ck0RGMlcGBgi7z4dNFeKsd1elszC
fMhaaN7ZWgbk6DMo+ZFgaE3+262QEK/sqgjQJLQ59muqoVpDW7yzwfHVWlnt6UvYLaNuDKrF/Zzy
j4M5NbCN+YNKFttaU8JZRZgfwN3bn/zE9yU7Gq8K7w6TLCVvbn7fau/knOkpaKzRVW9lTwqqsrhp
h45REi8pX8k8TxjewNHNd6TSeLk6COagFFf5CtOyyl03fnBffDFG36IxBb0WbDXP+3Na3ENcAz/f
ac5V1TICpUh+ETl7zswiOPobjSUS+ZwIdGr33FI/cZodvq8UIcYL4HvW+bG/5qs9CRUS4yTj+l49
+A4zMDO3/fLtFgfROYxEL0h4ITKO/4VAG/wRpKlHfTfoYGBvTUaRtCV9pC4kS/RKHmv6p+yaId9V
zcF+igaMe6M6lyZbAqvENwGmqjCqMaiCwpkU2vupmnkAUYK4tUPXlAl8KZ7yXOJTCjBCjQFs8gSB
PepCSJzrWtpZ4axvNHr3hcB1WCwtWnJm2cAYiL+Ik7EiX2egauTZKAiNCIP0uMftnoPyysEvHEU9
fefIfiAvK+t2OO+r5IsMHJauTLVbxKd8YAL/X+NmFRfNEOHpPAB86dylH6amt9t1kvLKfzm/mEwU
OCRqvfjvfQhW2Of9DBIWsWMo/b2lYiurwesndj1CTDTfiN3DwkFZXLRMTEHQ5kB3M/lSdBca6vsl
5qgJ0DgTnusFi7naUDOitvu6CAGD0XCaP2XzL4coD87ziDzDUYgaAZamanHDrYaahYDSOI61zFwV
daF2NPJSv24NMCJ+7Id9pHLHCYEJN9CKrnk0xbWIbgfOfrPm9iqoIakuwN4Rp+DfUUz70jLnFENk
J3POv9tx39fhEixuTNlrW230nQiPfMiLPZTRxZJrHgn47LtznRa6MHbSsr103Mf4J2+tPACC+83I
xCWvRCkUFPH8m5AljsSfcs/OyeNSp2oTy1rmiELCtUcojQcHSrj7si/AtkQdyBHS0UoQQ+2ghu6K
FwQ1OTj4h61mYb7NCWIkh7OQ2SnvOPPLIfqoU/cEPegiWFn1VwpMmrvhSau7UBCA/t0zOALUD7KI
Q84VBZY15W11nu/jEi+m9uJwjeXcWw+t/oCWWGmAA0GXeJru4pUnZ/RLCRrmlEn0x8DAhCohtRL+
rSmPHbD0T2zFTINhIywB196hKefq6mxBuE4/I5kNaozMd/dMt6xGAOAjJRuFD+7h1uI8r/vupWCb
xHq9XF+9XloA9vO/TbUE1GIN+n11DGawPikCG6AgmCPCCb5JpOB5EgRXQa8GnHAzf7rezD4Hu8bG
sgmARurG5AJXyRoSel2sw3AksuZ13Qg/fn8XaaKODkpPgJ1anQYlLZDoIFI7uZELec0troL3+DgO
hyuCAoatDBtqSa15payVJXX70UFO5na2SD7SkaLntIJV3oOkDkIjdQRCxWXpj3C7ZHdFHe89YYqJ
c+lBKjKrVi0ZofyN3eSEqIrH2AUeJr2slGZ0uUv/p3JeHB2Ydfk7en510d+lJxL3aLT2yUbeg5mL
kMn54m+hnCeEmeIgj+J0FUFgHe4pgnJm11Y+6Z/xDHnTv3XyNeMMbe2nbFwPwLIVrTrk1q8W3W68
YjV0dRTqbzd9C/wEM2rVYwlX0cbzqq4wrprBlnK6QCKuQK6a0g/8+4Ns2562DBzENsnEhQ8/2LUK
bSqGw4Jyup+db52houFb7pRez3FOak3cOx2H/cgNRz0UAgj9+b49h8gtNLXEussV/KTvMykVZimA
TbA9XYSpdSI35SNb/fn4RzNLnMo5eYnYIrpJrScoYNAcZNQ3h/btwsPLmHLGW6tS1jXPuO3qQBgH
7oqNPuLsefE2fPiNqk8MLSWtaCvT0WgaGYYsi7xvykssXCXmqRQo7zAjnBZqREJdKuTHV1c5kbOb
Ag4b4JFYarRo4C9DlIDKAeWaayB4BcPR9bfD2XF5bN3PTW3eoUvn6qnaC1+xrGwFs1/Dp0e/3Bq2
3cE1s/TELYeMzQD643QYIx7KVdCQHz53mMW7bcDDooGYyZaJoG+JBMVVbzndEHQl8k//KGqL2J2S
qqHNwF590jCAamNy4wLSRIwk/9YJPycFxFU0qyk2/k3/RQpsKv6hr3JYepp0Mexigf+t31Iu856Q
RFtAeiY0samPySXqZm6gZpN53DNFhUS+8d4t3yKWPOhO79b987ZtWZ9BY7LzfClP1mA6QNkpu+vi
huceuxRDlrzmWE9fsL+REFqzcUqGEcZIwyKxpiWP8BBJgDNqUFghR34awl++GBO5O5dD560u1yab
0DTkeG9phF+dVzmIVFxsj2TcUdmiM+EGheyg91B+YZ5/7FHTiY+zRJn34DOby3uAyOBlQgqpng9S
EbERR3rm3AaMl25bYtiDB3bd3vvU/PcmAtKf8z41gr+hPi9kFaKHVr/Sc3egLILHUQcXsApH1zMN
2VrnBoDSiuZlVsNb8NoPUQsfCMO8J0imbMP3YkjV9Mp324QnCXcr0ho7eVn8KGTc5zlXWC5G+aMi
5xGAH5myABT3/Z82jJL1oLuE+/+uFVsQuwgDOIJXrFlVFMO83fAjELAugOONQv+rX4ZJAGBXbzwn
2RO8iSQE/Z2K/5z1dgoPJ1vjkXC7gNEvMdbrxpOZHra6fyC321oNQHh2YVJ20nxteWjUqsYnIasp
3+KDqNGA27dRARQAVO7AH4bC2jaiiQA02k37GE/ctpamC1ZXIxQzpYUxVR+fW7tSIfxhbBeqicV1
yqS7UgSFqbxZykQ7BQnKprSIDtZYY+9iMGjxUEjqoqIelKySR5H4evNNLsGo9czUftItllqsl/hB
Pk9Df+qnmFvGwNcsfFSLlUCNG1FGkc5oycS8ErZKz35T7hk4jh8TYAXtCjgcl0q6wVeSYm70jnrm
D4DaNcmd8e6Td6b6LC+87miP8VtgI7gcQNwj75f0qY+OYDY5jFGkYw1morhaEcVNFq2YgJ06Lfl2
seTArW9uhBDKBmPPOCZC0iOq178JLXQ0hplPryOZvCbCoOSgQt+2qKSx4sJK/Z1hUYfr3bAbSCSK
Vszfxa2lQVqcLY/SP6Ph018c4K2SrhLFJzKl/rDdkxd5JP71k5NaCjy6f1dmKEkefcsNN+W/v2mo
bN3IirsMWSwlgsnNplR5a3INKoG+Hahx7lz95Qf1pDwseSGfqBXoKhndCYYyg3VCjtuMXpO5McvJ
EHvyWY2/9AAbHhGUCb4xRIbT0CL3JKIzdH10WK1RBtZfCxoyRqQNPXUPwF2+ud328fV00yUpbodD
Db33EJVcQjgMCvET1/BinWg7/AjSdRSsCXO6wSQyzTbwl2WrUzE/aSYijn3+EFzMkj/ZuIbCFp/X
89ElfGMuPudsEr8Ht5rR06Tcy4hxQpKTJqIkreeiXA3sDCaIMvYvXWu8s6d4VX6S7yv4UWNDZ+IO
UqwuQ7jx0a8Stb+wXFdFOHilj2FDNJ56gPY5SeihlYDBUOGJbFqp1lUHfgyCJmELOQhdgHjHy4S9
MU3i1fbJG37z7+UOGx/DjzMFxQh3DDBVIOTTuX3TfgZpHH4hdToWbQqco3YdhPktMexNBD9g0Uny
iEuoJb5GXNISN1i5ut/Sp/5qeax/flQUCigdi4TnnCeV6kbYbwuxgW8WMeLHx/g+zzSX7alCuK6E
Aa6cn9sANSEd4J80jYlZy+Ze6cmsE9VbVnpz3NLprNrAmjMruPGBzAn7cKEocv6NrDw+QsUJZrWo
uu3nUNBDs6RjQXHhK11oaw89BUBAm2FwPC70XCL+7hdCJxwTOftdfit9IROEnfCMm0OcqO/oDd/Q
qkv2zEvTsmgIqVuix7PoCBsoxwuRcawi/civUGWvPo5RLLqcUa4lpDNzIRibVsjB0qUDaQfn5Eq6
3FZFyeyhwm4EQCNUo543bMYEJUDzwD4SDlx9N9ZX+yuSWOyHAN12idihgGqluTKE4wD75E3BqEYx
BuYxZg5/TUY/+XcWhNcC6xUXEyHsOGomH6YbZFVNw+il7QhRluu90dZHah1Wt3r7rnA+62P15yut
NiWkYnmjpDfo22a/k0sCCpCGTI+I7KRw5Hz1aiSVZXqwKTlMGBQ0ye8mpJgMk09dl97BJWRSnFvZ
NNmN0zVRwH7dA1eTmTOnEuwxJBvLv4LQqP7wjmODPs0nDS6mJp9d2z4SHDANkxa7wLvj87Nu1FSI
4pHS/001vgURtWFAmeQlbaDlO+/RZ17W/w5yZD0nAwD98kkCTywqRZIOMYz0Sn8aLiXY5ycBU1zo
U+FMVq21d1oT7IBCk+HRT7kUar3Yrt+y7JcbqO62Ukr6fiQ9Cn77fWo5ORYwIAadiMA4xFAz22Qj
bB+BQJLfa8Q9LB6b7fFUcNG8UEaciCQr//+HGpeEdWfUttoy0SC+qngKJnVv2XJlH+GPnYfBEZy8
aCi1VqfdzKV0culIKvzSS7T/r6w7ZaQQSZpdDcrVrq6hp6gfEM8vRbaJ0dG819518qzD/6Czu5On
duHaRJ9Pz7GnXE/Pm+NRZzvNA6sC272AWQpy0gPysWvTm0YssBub+LB4YlliZ/HzS05wCpJIwmNC
Jd4Yf3OMQjUuPdIP0UiNEZ7Lrt2Sr1Btpy0OvqfD1EPXhAN6R2KJ3cER+x6kminpnguAJEWWoTAN
2K3Fqsn+333xDgCyveGq0JAb0h2rXi1xh+ffC8qKbx6qoJVkxxXVSNgdDA+xa37UjZC9QLHSRGfC
6CQ1CeOVbUa34hyJfTmcBT9rJFZl6hs4qtuXFEGBnJBxiZyeYq2hbwSoUZVQVb2Qn6OxLtuHSByJ
4vI0Dh0HgPT8K4mlPJV7AfAl0pvZ/+kR2vbkj8v5HyoTPS+bwOUL+/ofsi1DuD9UowUvzEMnkeWj
jd8pq0Hsf7KYQfVjaYjnB3dxjLp8WqAExFVNAa1Tf5rGRxP26CtKap55g2KMWFfPNnY5knJqTIIK
RvdBOqaWltpFg9lSQAIAYJeXpzXMOwAx87qk89XLDXif5xEp8aU76x/bIDdz+h3FC+D7w3Kc1eWC
uzOAuyx+vJyxZk+g8RivSLALi6H98fwu85A6kVzB2NtraU40YF9ou1zS0f54A33xVtBrIVCAWQuK
sX+XvGNH15wy+pZWRDVRVZtGjeGevTl+agWRSAD6Mam1iR0jrz7c2RwHo3vIYFPEGr7iqHm/Zw+L
LQoB3b+iOicrbRuDZ/9gLcExEKR3ZxbhBk4vnFhNyP/7KuQuId/oq42iGicwLU8LLUZi8L8edkW7
QTgtjXOA76OY6dNXtpXg712Dklc5HjyGDlUQOJ1XeMEmWZe3HhMOdDQfwMg78LqS0XyN1VPR3I62
XXjvf9+RzNaawmNXWXLJncOSJouhq1UNgv9JYL26CTNjsfE5Bj2MM8fIpqNI4v0WVP9pgevlSOOp
QYgiYVnpfIxHucqqQ3af1hTCzGyrYZmwytR+eqGOc+7xYO5mT6sJTF3AAWZd/LOp8vBe98zJSaT+
wHqOYjdRpghFM/jt/86zP4m1hUWh9YbjfKfpYbHiREkph8QbVrrYnvTMyjvAuxG8lSZcVcERjbOT
tw8Vz2r1aOcqS3w6bSk+00gYw+V9C0L+57NUvMkFrxO9qx2GoMnX03Fk9/o10G18yby7NjDEAzie
IMuL8qsYrb+vt+fcy9X1dKyoZl9W0Q1KQ0hexoZ/eA5oD0iYSqEXYYgqUxApYuAkWGfjGeHCw7u/
qbhdwa3+v5+6QiLNYG4LvPFwGQ2jrKVWx7p0iZTL4XcVezzwjwJj0G+ndJU7AkyMwdRMbKmd65i3
1f7TLnf3ZXdx5jRkf3UekyRaZJYD/tvqr3/WinzCaW+JQhLL16TnisrYcTzpw4mbDGvuJBUBjGFT
XWCBM+6jZhnkv/3avZWuBQjX3qDe35GXfVHVUZHA0Mgi3Fx/dJY2LqHWoQglf6E6weBTaUgu7N/Q
fpxFv3fIcADaVSQxOvYyD5VToo/MMOlZ4iD5mU4f45sTypAKeYtXfcaKZZ3VpF9E4BTDnbG6gjgI
QAZHi3wgxjcXrjaZg5K2fTyq+Ui3n4LpIDDElfTEcl0bU3FC2FAa8VuHmMWYI2euOKDqYF1IyCCw
A6cHJgunFZCjI2WiqZ8gtofPMyf3Cha1KjqlvkoiQedtWR/rDIko9pGek+mDhTd3IiSuLhXj1NkE
Af2Ml2ATj3du0DPOsiA79veUhqXpJuEV8LH/KdSE9QL4Iug9BB9ZJvY2u6Oehz1Mu6GJXQi9wbU7
qk0tN12/gZbTEC7P3oZiGovxFwDu2zDA1xhTZe2FBx9wUAfs7B9otqAu1Xn1q0AoJ9PnljDZ5cX/
S/934dekmcDmoAqfrGWAZgVBbe/fROHTZ0EsvoupLItKGo+X6Sor/ibdcuaCmWOO/Tw/NloLyPVe
BRxxqpfrYHd89gzhmzL44+bj1viVYLiR+TEmVjIU609Ow6yUKP/98Jny6KyBo5T+zjDSBnCsEd7X
OD88soFWWrKNsMuKNWpYMH7EJ+xygJYwlcmwbItNH0lQrcspoiRWlNpIsbCa9ABELDiKM8pQcVVd
69gwjVc8Vt7CEAbxzAro/z9UOO9vmkV5fonwFxU6mEkDgsrAUagrRAzV+8y89R7+5UE7Cx2SLiO0
P/qP4FcJyPgyxfgabGAFGr0a/CadNJBsWWO8Afrp8ijgOGLA7Pc01SRW6Va0tCFqG3j5QQNwb678
Q1E5hXF/qommjSVwEdFBUvKZRZGXEsAzTMD21Zd6W0Fu66UAITuNZDug3/gzAXfCf0SeWtv0tAKp
9RmJmQ4IWWHAGnTIjKUu6DNTVUVGckvvqAo7pndnbXdquQEW3WSKmTK+FWvaWb6YIIp8VPJEe0Nu
eDnlnJpMf3WtgNvOBihHTg6RIRVpmGsw0Lv4yy1rrNO9r0GvMUetfZ0oLdO+yrWNjkI2cweC1JFV
AmAeXN3vq7LtN33hW5gonumxEDAKuQtIHcUq3hJ1kO0k3A4+FScVn+gTPU1CWgAREebjOvNZ6osJ
snORTAGRlXDDY11phT3XlUjWMw7k8AWplCr3pg0lD8t8bARVjIqEW4K5BhY4bbVjFAdDZQklTVlY
vhOl9N3t6EhYd6hpr5rQiBfYQTr2Gvqm9tgJqPp4Piy3JBcnO6XBkM/FI9DytquIrqnqzzeWsb2W
JfBZXiAPq2cHQV8l+G7FmveeBQdcHMf/Q74TQIcMQKz2WmX882JoLjEBlpgzKjryz/wiT9tI8cHy
eZU080VcFRY5M6nLmNYgQ343QFkK+VPavkg5l7sTX7sg1keX67MTs9Sq+OWEny2xvOAa/y5fh20W
tiKHxTzlW2xY1yGrEQQceVV8dfwVqY7zTvJoCNGJre4Y9bHvmScYFXRTGAT+NelJ3ZKEPeLQdRYM
eDgwe3y4bRiyF2+Y/Ng2biPGPQMds8CXQrdcjH8SsoD5md1Dklw1oHflbU7/qyLxlx6APvZlNTdM
P1TgLBEGTlZWmUdzpz4v2Q7UugJN/v/STpO1SwqRsiJGPR84wHN7QCmtT/08XsnDvcJU387uW2/+
lpV4/zkh9u6oL5EtZUznwXwz8s9oBRbT98+5+9JdQjmhbJX94bqnmScifwu0TQA2I7QGvWLPfdre
dSS5dY/pb8DjBZW+VkHK50RM39HMDx9HUTseZWgeqcoxmuzBBM/WMrUF7gLwt31HsRpVczycjngE
aBhao0tZai6rAVwNQ2T6LPvd13WOYaNxzJjLTK3qEd93GXH6+nj9rR9yvFQxMHeQSJYixL1NEFqa
pCQHWAq+TD06ihvsZbMugEYbOlLPP90z6XEB8dgw02iTOcsN0/AjOSeHW8YJ0H12pULRxPIKQayW
+RVN0t7Um0GOy2ceM8xVo+0KelK/ASRT5kdV8zVt1/5qBc0k2V53Vran5AZ5JdobTBQqKKBRtsvQ
U/MGWimGaNtw/rb6oAWCbiZMWSgSoKa34a9CPjsRjaK5L4N5gMmo2+RD2YF1Ns6/Kj97Fii3rcBh
ZSVS5nSLWXKse9Esab4liT1k7GpmgpcUAp4VQur0SK5X/bPbZS8dliAb4WDT9Tfef1fq4/ZLfaa/
/Nxvb8KuCmrZYbwdzD/cCLgMK8eBJPQ0ai+VZUwan0uWjVIs2M2rSRHuJmMlS5OVzxEY5bwYSlqw
1MypQyiQ+Tj8LW6k0r6QS/c9W/jiJt1ZGq7BFYj/IrZsfPyjlWGsCDagaTVVm9dhzqPziSPfr3Dk
Kau0SO/yxaUhRlEfhpsh8WQ+tfL/0gZ+kpLwGJehcbQgfVoNEeZyAbARkswgp4LruNsWkB+SH0cj
pCg+faKUq96mFolw/8zys6x676NaCnEcILCFs5N1kT+YgHtdapk7cbbWiPCVkjD5ctc1kP9kI7pt
XK0QumSkj4Vpducg7zno0PL8qHvxWf3mXdDr3JN1IMsluliwXxbcJlwae/s49e70LBfwEAtV6Oi1
aPWtzj0XMQ0OCHU3KyNZxvPVZVtp3WW+061Dadu4FECdSLg4Mp3G+ehqRv+eqIcsAw2w1uszVPoN
IpRR+ly6vkWHin33C8H3WYjlwq2nqk+/h86V0XuaBc7Aj1A2mqu4iRJiAH7qNcqCaqpAQrhPyJqw
/OJLDnbqDTOkGoJljHqFGyolKXOLzRxnXMV+YzfQTu3BEQv21UDVVqnJ+egaCsZR5lKur3LL8TMg
pisAiNRnrfCEF6gk1UdwaW/5ObHePha+GC2a3fxL6q+E+liTNehNFiIwoW8u1qPAqL5pWqugONyD
2p/LNgLJY43YaahYoAfdfAh3ggWHZ7jJbUhdSHghHFCxAdQ418aiK+/NmuuvLwWw3m/zB4jcxIaq
B3x2AozCLmwXMd6ncDgqLgLDRwnev29rx8JxhpiNnkvCCB7QNHz5wg91lc7J/W8fJ0ZMUNZ4rR/t
CTJywcyfXSxHanpwDonuZSAHnr9HQssVNNok2kYWa0riwLDh/4b8GcRRBjb7BriNt7jADtlafvce
t/ewbzGPuIlX9wOyG8oO6zYpAUozfTfI0nwaN0PvYL+bYfEg9kFuM9sFyMAxv2+pztuMywOVLXVC
ZNNyLBhjBVmcUOnfzSNP3X+SrUQoG0WgxfMqTXI18mLWoT3MDcFnersHobDbufXD9NeGODZc4jOJ
mTT+lCHi5jJcb8R5aDmawpP7uITfAGphE5dCB4yJqFV2gIhZUusvr7bKpP9xXdl5qoAcD8Xq0/W/
c+QQJNbCautvHxtRjva1PhKGQ36QE78sPiIkdJCsL9/dxSYHcMD9HWP+XQD6oyCFZ9W6tYbBhVR0
y4eaRgKed+Ir4ZxLmY6KLJJi2Dsh1VyCtPt5ORHoqgxpqePf+1tXbT7DVTwdHRtoA+JeaC8rsiPy
y1ssb5UpZ0auuUKOdqRHqTHHVCffJ1txdJ7VwoWDPGpTaa3ASgMG5Uct4fJMPsi6O7wJUj7v6M/q
LJT8GAgTjZ77Foxd01r88ksnaZqLgzxeMNmch2CxDz6ldYOPDQQYd10nWG2AiYZqi7YgKSy4TcaH
KB8AQbpo+1a7NqNwADo7tCWf3KrktvOAf3E3xMRfIk1F6cj4KEMKqpUwdwAvKQmPeCkIEbq2lCeB
m2/wBaFSqcjyXAAJ1GEqfnm5AmClIrS5si4etyfOGP68jx7tjJI6ox07RdKm9VAYxX3Hy4OtlwUK
1f0u/HYt1dHC7r6db6WjKKAxXzflKhSS15pgcJ5X2vpQHyLrtYhITdFAQctTA7NiT6gb6Fft4FML
6xp3RpCHa6CCv6uH5igKF/VFHvKsgpRn38WxVVf3MgKS01ItuYvK4WUSHkhc+y52mJpGhA1SwG8f
r2egjmq4bppGwbr2WhBFld9K+p8iMWwBamSaLqu1rdyJ1swI0VIdxXBwIuK8XGz8Z/0dYXXcJPgl
7Ha6n61+7HseDf7DJEs1+dTBXwNM3xvbbySL06BBT9Jw4hmigHLQ1AKxKXLyMfWyEjLdve6DyTV7
9KxEByfuDn8nCS/tzeXfPvvFhnHLVfvkkKo1DsOjZnL0OiiBBpsIfG3tqMS9oH7bFBENxUi7Dj+Z
F/XyNXIGjLyiUl8K4WmODqJJHF6pq2eJBNEOt4vss9hVFYXbV5AmPs7z19G0/I3pQz0dN45QXKBn
GJC47MSitSMfN4kMXswqKFG+SM0rm0iRrep8iyIpjUp7RZ1mZYV/Kbp5qnQQ7CQ/uXnZkRUNwfyd
UKPTgD9zFKihv1JJTvW0kWi9CWq4Gnot7pGNz17JMM/7XRpe79g1gq1c2QWig/9yppVcp/o8arwn
3x7ucyCtY+Uui2SQnRh6Z0xf84Unadmv1/M5PNllG/0UcbK7YAJFz2q+uxiL6Yj2ePGoJm8Lx//h
O0TmUb8AhgLuDqRl5cEUF160iCS460e1FE9xDy0wUoD+KKLK3IJe7xVLTF4VfdcrzGTxBUqwbAB4
JTcTh7Qb9Merci18NH7I52fgYAe73qoNdcrtjN52Oqa+kIMHjWrzcyb++IUkngGn1DPHDlX1iAWt
Kz393kbfVGvTRXrIXX82PkGa656/tpWwZ8F0eGfM0szD25y/vQDA7ARaiAq3Xb3FrARvUMTEtbed
4oIJHdHlxbwN8LRa8HvRwXI54pVk3TpVI/13XpsVSNZYMXFH4/0e1P9GnSRdm38Var9L1XMu5J77
Bv7qw8dgP0VxiCDfH3mxBGv+kmrdZTxw+UeCvJtFhIE6ixBrZG7v97OUZMLrReDhOOBgec7juDsY
D0s39hKRHeaTg/qbi9brfJUR9ygz3FMDJn75UYAPf3I/qYU7zQUOD/BMV5BcXzrJ0QQkzX5qdH9d
1qdsy7g+ODJF8PHamA2vMSJylDn5ZHGjhFXo5aQHUEGBxbkf51r1aYiTRV0TgpoYYy+HFFfHuonw
bmGuNTyla20JvUdPeqTHALshNB7gAvpW3mRCb/zA3V+mjlP0+wNkQxpSw5ZIKJNtq/GAq8MsEgoe
YEmaW3o3u3412NZpjILNtPxyVa/MZ/td6l4GcJpOz7+Kgjzq2f/78BcSyu1ndc5ab5N3+OMf6Vpb
rOK3eh+/joh58EoV/q1FRLZCI9AbUdgoTLh0C4eTwJxSNOQk4Zbmr3/sZ1lBzafLi6LTDqm9EWDn
3eOV0gOEhWyIPq5wIwQkvHSwdJARn936JC8jUEEXDklz9PaPYgCYVtvU/Ndm/sWYF+WH0x6gfLvP
QkoM6+xax+kjAvN+K25dvPBKErqjzSEqCMUJS7xBqLtVBjCJDtIWQJSFeJ/XkqcFoJbFag1ujK+V
LMYhnHO9UGd0VJnHVlJ/e7LBMu66w2EpI73ZJArITzPB1n1yex4BO3QF9ZIiFRzWKc65DYNNFrag
NOEtHt9vFY4uNaFwd63SiCEJNp/OqEZJh9X+96Mq74VO1rESX7Y6ESptQXpZmZK5WeCAFi54C0OY
ie23iu47r2qDTrVLJ2jc+0TmHSNvSKvBfm2kM6ZA1AZ/6rnBaVIFPwcph8AG4LyFng91cnDrlBhr
6objXJacM7JjXRaIF3rX/1VaSipP3mUQdTZFBrZl66HczmgJ3aVkYq3bTvUQFS9XLf8nNb4Q/kPv
scIImZ/0csWBoABmf2F7XBG3EWI0F1SipSASTfGo95lUaG0TfEPatb800o3RkuSsEDa4IoyYh2+p
kjOe7FDK31MyezoSJg6aOO/kk+Zx2heyVSTi+kpYFbfl5yBkj3jbJ5U9GYcg/C6QmjfxqyFRgjHp
TqG2nAe0FJ+ck6pjam3j2vn/ZARVv1jB0088/kVZh1ZB5H1cJgd0BNCsxjBBNOr08f71N9ZwDkjR
OnlnjU5PMxfo8Gmr2J99LCGsROxRCUIQ13doat8HrRUvin97r56wwrWZPMTnrrrXxUJHUJettZ/D
zkMaZS4raKVay/P5Dtr0fdRw9zOuo1OMKvYHpAcSlNbzebLPwy5z4U/6iK87+9V22xW6vJAzBVow
w6yo/DgEcsPD2jt5FDDEr7iLOhOGUNaX2/j4k7n4XETioG4fRl/uGpU5A0p+0RT2vCKHZWKs591O
GinR6UqTkD/2MFnY+GADMSWeTVdUZBpHBjeoU4RvE+cr1N1s2h2BQcufoCvtm9XSVYqXzzJZGw6S
7Vl01EHbO25YrEFLEiowaMN0oqFuhCZOriPlF1ZElkjTU779/bVehWCuYsA52+i45JXH7t9sATvI
23Gzw8+qSSF7f2viV2rLGjR03j+yCKkbJ6dwv3enS9Q9xzb2N075jHkHd6McoxdnxmJdwzvLYRQM
icax8XwvbgwqJiGoxl94M06Q3jkr0cg5jxxHgiePHsVzN9rycvzLPZJrMMf/N+QNqj4TRDkGZvrQ
CieQsQccQuPIS4gPPQhBIp4lWQ1uguOyB9QU3fnMnx7zCkBWbRlST0mJpxanB6mtA9LYMDABnERW
hF3lBv8a1Ub9VaGoy2+Xck5FxrYK7pOECMzX0ab0+d1XhzV7uNWf1cgyMe8V/wujmUb9wdAl2PnT
MoYR6BY+8lzKSofTpM+w0ExGdZ9MgKCvn9RVJHHpzTFCWMQ50+9hg6icuQ4CUemGqZrTkJQaGf2c
sknkfjjkJToRtoh/sweLLrseDRdEr2KkNsF0QLGfWbADz/UdwlDXFynzgs12BJmS/sAAc8hQHu4H
WBmzqGOIJ5AgOS/LhEJ7eLSCxS2uC1Mm2Hlixlldoqk9iNB42Pr3ShJ0OaV6rvWYFvGJbBFw3CwC
NG239HUeDHqr1X1pASNMqkpUFpa3kNduL76mULBYJvC2vbzXIDQDLR3NPKn7Oxndqsz/P/lZa8qO
NVwgDAQNR0Abl1xW9nyuHyO8LhBBEdfi/zi11Ibg7E43vpTHC65/infjPcSSa8ztSPGERTaFf+cV
5ZcL6tcsNyaqwR2bZPlL1s9x9lrGNFp7OeznE0Wc7aFSvwgtHR3Gl2unWIgbOHjxQ9bOKZW6EUO4
mydie4f0V7PB31fX4GM42jzip/KLm371R3CxehG4jnngwVT44JV+k47NUHkwtXSQanjJf/lqN838
WujdcpAvv5JfEtGHN/EBI/PqqJHUJDe0GhksZB0PZ66I/thI02K1fpLKNyByb/J0MbYgsIM13jHi
jS0PHa2URCjQdogB5P/lbp8Gc64BbP3yXaf6NiRTOzA6TpIMmZB7ZmF1e5MvkBdhCICFys7VDfww
g0EKm+hcOCmPObbB6TQZjnKUurW9QOxr2wIIjv3TBYi+7G++ofjkGUoGVQbmjFJY2IGksj+HIHnb
LjoAsIJYEb31Kjg1thqIOcRH+gs62ttfpnCnDSSypSiQlgsJ6FiltXB+X26P3P+eKMrJUKu+XW4n
rmTs2J8kcbRNCsgmQcoi6NY/4BTBXEZhcZoYT5NvKCDRsE8uoIra5a0+Uai+rKB4lTVVOJKOQ7Iq
fCeM7HHjBYmdUy4VgDoeol7PS0CAuOmODJtBZPq/UKPHLHadisfkipUyXABSCtQUz/dXSswYYB5N
6UgfuTkz62fNw+kcrGq8x23/L4q35ObTAw7Z6TMLKy1dSzp1gsMRH2uz0ea8Oaa9DGQ7ACf1y1An
AYMFz3GFRC8XIqHoBkMgBgZ+ingtcYlIqK7E+QdM3QWWLjuMF+wj6FYBjN6LuSKfRyDrON7ZFUVn
IzEq/wMomNXj8kJ66xEWQnb0yGWKW5KrKAw9EhyrLJDbM8LJDvKeUFp893z0AyNkw+w23Nra3Am4
Iay33jMfIXY3hcD/NALiBMxCHO6dEGwIEbU/10GQaymngYMRDn+5euWgoXHdKFUiSNNOpkAzKX8F
VwCTEfnpC+6F/xHddrsxGN8ygNBOXZlYTKZatdnpaXRRZZE8fH5kqN3zYrAnuEV5aHVar3jg64IH
og8c3kSsKRk0A/iYmnJI2zfkabEVDmgt0ZhOuaRw4TM1Ozb/DWCFdoCiBc33UCKtf+Id51IBp4Yc
reVMpzUSHIswmyYjeIwnKqYENEbCi3d9B45fVZ8+SJd6kkqLRat9EVQeIp6om0JpxCwEv35PIfKT
FSPaZu0VjN3Fd42rYUQEgarU0jzQChPT7ryxFKHfcyVAYSN0KKxDrG/o7utFEPIslArifkG0lRzP
rtrPs4FvFJ9LQWfVK53PfHi8PJLufGyFgz9mMV1preyOIBF5cWD8o0Tv7qEwgmKBMk26OlNLsKhE
JiW+9HjCmqVwqxln+K1zxkgx+ZxHNZmR7zePNk/96mSlf/mBjNAmxZ08Xzu/5VgPXugXdHSHc4/n
Slj6ybTiEfQhFMIWk4tPG7m5l0q292mh1c8/DQd8gaFakRz813xFM1De4U/10onFUYRZYKxOVpmk
FSWpgv3zBblkE0tH5jo/JCIicMXTKHcux2nAD4siR0bFv4eECfP/FLqlsbXL68nt3o5xsitLV+mk
F7UTvPH/Yi0y8v6SfuOgJXzS51sc2BGu9FTLHKuTGqHBJpeaSJIdbjnmL2GPLHzT72eBoGsC4KpE
Rwn2scI0LmkBT+e/CDg752nudwON/X62BK3QcAc/NdIU1Gzs+g/t8ryVR1/kOMphiz0ah34qgdLK
5p3uOwXFDWwh+L3pHroozA/4Orup9HGnWbm0NmPH9BTG14aPxzzn4Ru207TlmlR98jfnFfFlOM1v
BzQPbI9Re7gtSwe5Y9RsIBpY3geJVWrsxfSGnQ9CzCktyvZy7eQUbZgL7A0mBUQhrVJxdNJYyCxq
TDYvORY0dgWUwg0xu8cKZpNZCucrltw3L0aD6JfZEHdG0EcUCbKsNB/xFFZJ7rlb63UPzG6QUroZ
UbefMy8rbpSfpMwKq03tmBvV+XE2GpqOsCzvqjfJ359SXASylMCaS2Gwcw4mu8LxdZl+EsbpeZH7
u/LsnI57+poijvkF+WvDD/ONtGt02EKKUAm+fXLtVET8Sb7bNsMopvlDBlVaBSY4Z8JeaSdyYv6Q
SYLHQa8EWwO7db8nqC8n0d+uEoVUmTiATWofOVD+2NjmwC18nCBpaEe7XiIz1E1+TrKz0IP2a8u7
QR7UHyUhSrVjDBiNyg3fLHv7inCCI926qLTh+NIEz1gHaXtFdRzLm8Bip4jPq0+kUoQRqxxPjGTs
45TWvS+xidlnaB5NP+h1bFZTE547TGzzlpCzq0yfk/RjtWH/z+K4u78R5MveaxnUdL/ceuoqK0zs
pvuPFKNs/UlkYq+2hveO3Lhq/AFZLGUzOBjWgUD1w54Oa9DUBjd4RDuDjM9XuHeU29M2bIQLiqy2
F+x6sx5pghgGYy1QFzvWJVeFSwBiiDzTTCv7pymcvcSHqVt19vDKkShvQAv73aJCuWqTEE4znUu7
A56zAV/v3BRpgPwEsov0xljT3JgJ4vo9Q9fx/CbcFnFHA6UJ8IcA2UiJHYYcZNqTulZlwbGBKKsN
4SEsMDPDfAw1I9MGO/V1FOS/gGvuH4BDBLsTvaYiR/maR6sAc0hSFnWzuK+CaUmKqCrTCbwAY21v
y9jfSjoqaifo0WVoVTr91nmXyCic6k25c5+jOX9+MV+asdh1l/GDthhh1dQhKGZjBrRMp2RPsHE2
Qbip6h/87W8mE9bL6LCOEV+SCa+XqnSwkCArsfj58JUwAclOEQWMnnWP0Dqd2AWlVXW2c4/SKayA
rpuQKhNb5vzd6bbin+QTXI2gsEJ0SUxsK8MQ2pb4VyaP3QZs1Ca0CYu9SK0GLBAp8M9zpstD2K8l
o+N/IfxRR2i5SUYHGT6akfYQ4kbokNLAvboOhbXB3t1siauObRdIW/LQYOAkCdzt0lhQdkjwCsNu
bPKomglFkK5YXK9x+d0wKjLRH0QaiR8yFBbXb0ArXpQwqa6Te3PPWclHsDb45lChwuxGSo6sP+m0
AkolAS4WrW6ROQ+n7J4ct80dC8fVsXf17LYOPUN/ZnLTdimL3VAbAYHSxQgDqvOYOTdW7c4kRWJk
wT6sghXIGG7Xz4zn4afhQVL5MrTa4bKze2HJyAwYLr9ulkhseCG0pT5RWUlU/TrgfWsTY4qyNQkX
nko7hdT41LWOejl+0G0nj3xy9Ax98+It4f38grLCrweXbBWRrbMBS3z52x2/fBK7MPqjsLxhUbSN
Ek0DSKlGYtPoki7zx+GAqcahpFQdGZe5XpM4UDHUjzF+NlrrUk2nDze28XZFSyndnkHdPn8aUsTY
dZuzsxcPxxvylFR8j/2LV7UH3OdWxVVeH6BsfAiM0qxHSsrwJjHMmSdAUkD2wIw613Ln6KWPgjzI
/oM0l8nG5aBE+XW31Zlkpw1iVigZIIiSK/9SECBFQSIqU+0Y1LqwPVnniS56yG2rfrR1irg4m+u9
58EFDfLQHP0Flj+PwnbWYj9pKLZtMC2kEIQIFEGm2SeV9nHQxssHokVEcheT3OUTNZF0NbBbHerf
m+AWeB8/1hPLb78Tsuy95NwHJVUjcW8H6CGyqJOHLxut15QFdFclMtR4M3XYMg6iqeSz8s3/v1hz
sJH9bL9ivIzVRIXGyvDyXjCwbSnob8RqEt1jdMLp9xesqCzGfLCeRUGyPYLA6PeEB15hiXYyBvuD
FZ4Mppk/qabCd5QL872ltAeNLQYwFAP9PEqBQ3fDzx8U2Zk27Y2CBGdoz9t5oGxzENvZNWgJ4P92
NyU18x50iVBUM8y3sBjnlcrpU0KIg4C4dfB54bMt+ZTxs+hWJMqxiv45gnbWa+wuG2YpMwcg1yqf
At3n8FHnT+Um/Vv9kqA8tkAVyoB7+M6P+caDMg2NoF5qTqAZHaxFZMKqzpbf5Of6DLKb7M+BE9eH
85iq2PpOx3JlhFSVHPePh3jWkc6qhI4uF1UxvW8hgALFfhF67stxcE5zIDloieUH5MR3O8Fdnuad
VWpQqnlnqUiJCUzWjAnRi33kH/1K4WRRpzbwaqlpGqxPWIFP7F4pxpm8opnDlwp4NrPGH9V93YMP
bC4xYoAublgm/WAop/P6Z5N8QrnWwNByXVUtsX4cCy3SHDfJS/FfflX4nX4X0GB3F9ESTO6nQjt5
4rZyFfSTWo2XvpEZCyasUfCQolWDue5Q7gdbBMaAYRBAxpWxJywMbpsLr/gXyim/scAzjuxSAnZG
zishvplN9eRkoUwZBTKZKkwgtX+swSB+YxciS8VNQTYU+5+6zSB/pR8l5gRrq6YjZOA784pD4kCI
nIwANqsmuyRl66TBl0b+9wMKBn7xNzo6bmQWXvv7x/noTkQc4iT+uYWpdoMI2W8oNXDglmlsWiOB
q8WEPWicKNhyKOiS1OWcKYVj9objhAJqjrTc+vjM7wqYU/TA/KrLbwhwaSXzxAvWI1MgqA8wwBXp
vQeMpg+qGJDbBxaieAft5EgMv9z6u+Yy+NKOEPghBwrs8iTaGEqgl9N7MfARBzaA4aEaWLKurvGn
8HnP5ew8Mp0C9r/GAuydjfqcG/oD6+89ZXBtjHyvaKmkXBPE+brqbeFWrzjFhWDu1Nj3avg6uIxS
5+Yb/C35OGTZeKkP/nW6lavNU/7omeNGa2h1qjM8DTmcwKA1/oH4iTNXAWk/XA1idP/s3+N5Hl1v
cEeU27d31mv3fojz1piKj0slJuDd5Tnl/J2Dgxm0e6Ejzh5qgMUAKbUSfRZIaU130j3lO/k3RxZU
JW//aBoiKBc+GmKbKH1rznmNoqxKjwEoF+tGMTYYIk4q2oX0flmgZR3XYdVVqykUuPxwLpbZQM0L
qGXEghNW2Glyv3x/fQWmijb2SJyHeIjqQsZ+Qb1jNYVJ3YkxQfG6qrWPvK63Fs2MDE2rjPgeN2Jm
RsxTsQvXcjY/fbZXdH287PR/KtZx37OtvP8zNIsUNal7/VESfEv98zhkJpK/aaAXrvGlQqdEq89x
IV5RL2FnFsH1at19mbHzOwfcXMcxL0pIqZgmRaslzTH7x0dZEAISsjwy2wW2os/qWv02FNMf6s9k
ADJzdMkp1cRYpZGSqq729xJKh0wKD4/cauCtCm0E3ri1pZfVpwtLs+8zWXIbK6JI0KZJkqOoi40i
ja9dDVznSn1DxDSDa01+xPCT8U0UnBox1aS7ahTIGyTaztOTkqC51+eYbb1meLr2zccUHxf5K8q+
fTvDXjMl0z61hplmaMVmd0ChNAooiI6CzbCE+64vcZj7Z8rb3WvhQBlHsHyzqEEf1pavo9WuxNl+
RRkCG7m1z5g6oWXxKvbAaW3mEquTRo659x2aiD8TS+WpXzDWM+H7z56fbQbdz+HTpcOMi9p5kw+x
ZTm+i8zKlPLro4wuJCtuE4qwyA0tK6LEwxELIe1o4TFbei2AFvHtldM8lmx1NXF3cJYsrNvGfLoQ
64sVmuQZm0xlIX465o6MVVy9sZ79JXJB0NdZSBLWfDFxHtrG5EfYrbjxTpDNpyPcrdfTZFkBAxiM
tKsTuoL8dClZmmM7hGJqX13XmAsmpFUomJ5x2CF7CZM7KOP9q7IbEQOcK5kSNWIKsdKCc6GkkQcE
slDVYlkmbEQdz0h8LyfNqR1mwLp8/oOFEqIlaWlJYGifeguN/zK7eqYoWm1+mb6ISCe+6Cfvumvi
A87v0N174v49+JhRvNw/MVX5TRi6L/a6uXLCtN0TjwkJD6/+oheauK9Bo4Pp3YG7RIcUvAu48MrG
3uLq54g8eS3y0lMbKniCOxAUCVYVoj1jaJWy05B2IcXMbU15K+22D2mASLJxQsbQhC5TSe/jkIhN
OEv/FxvAjqu2Bb+ZgARv1miNuFlzIMLd0zlR34yQVxkc0vT4tD7usIQJYigBcOH2o5U0bLuXTWjV
YorUziuz1/X2RRgbY74jY3JNJ2p2Z5STEsneHtbwe2QFn9ldkM6WUlyfMnoQcO/EDEoBantVSOuk
z4Mw0unZNb4c5AUHbrmnAEuhuJninM+T0xkyQQecg3gJEGKre94ZEqzLao2tNjEzPopWv6bffQW8
xsSsO162uwmYRwFjWFAcVABhIZd5+1wleIuY/C11Lp3Bti+WfOR4s7ZF9Zo4tuKM5STLLYbErbVp
J1EmdntGVW6ruW4BWZSf7DDpm3ZP2VzcXmxuo7rmEYENssed7yU1pVhCZ6lypw7sv3dsLvBHTkNh
q9GKqwcjFaSHIDnbVvB/BZG5ZLw/quR+WFrkwqGcdTNd1I1UNEyZSnCmCyyyJQLOOS/b0XQAwjI1
mnuNfIAF2jPO39QGP2ofC55QqZBA5Mdt6i+0qIhsB2eyrGQvcFg4P2Swf2EofnOULbyoUnEAOm6+
OI11AG0XHTivdSlB2EASiJXlzCm6qUCHoaN1uhdkV4KHcCSG4V7SRDqcYBduVd0f5fzzX1YKCpSA
a4Au4xPdYUU1qVWQ+nLT7OkzmyBtLVIsH6Al6Cbn0zItLw+Mn91RiBNL5/qsGytJAtZHnxNUT8ID
pW7Sld7VBoiAR5Nnwn6boT6YZWwEp7pSK3u0Bl34myOoVSmYrbIR/71RdjdRiMjCee8Rt/H+pzE9
ciE1knwYWEMi7+A2gIdmpk9cEdqP5eNKNb4Gu+bExk+W5cGzteakELhLp7VTnZ+PPG2u+18JGNha
eGzwDf8+0Ok//uZngs1w1T1lrCxn0K/f1H6o+Q8chiAfr5UA8UxRbig2/G4ya0ZHcJDS+9JetbkO
yCFWtqeeZhgtqyBjRvCqvC4/w1YkIXo4FzOO2f1ikpqbZuhf0cm0CVzqELLoSjNrWBDFVANNLwTL
PbJQ2IalrlWehN1cSMTfjt70SXuch2nuly9hw0cXJunL8r0Js/Ya3J2GXa6Vshhgoq82LYEe1Km4
BhQJLDGeSfzTnfigK8PC8axbrKrhWQEPEJEW2F+b7VhhSpXR6JksNeg+S8+r1lOBjg+K46UdRLfq
EreoiStsd+zEER/WYWK+tcLeXOBOnDSfkT9FsM3pfZxmfF52B+aS16a8c+991sNh6r5sAnMM7+pT
bfWMmshl0sKtX3oj45X0xhTnB0qLBA//j2hhUkXt5qGKV3iIOj8qJYW0tyP4ZMw1/jstRmrO0ZYC
f5W4j/VMHmWme4iDfo2bPkhAX3M4Czl3yoio1ZW+9B+9Hij/hFKqrunNbBFEgeW3R4sIhCUnhr/0
RzTpGuMYByweAHC0kzleDAa80PwL3r5vrGeUM7P4rQMjoHnSgIWu35fZRnBtJX7DJZ6L0SrKrztf
Vf3BmGOoikoRpyFHOxfbKcTR7VmnJLYA2DI4em7M/oAbtZxomFSgj1js7k3SqiJwuVGlhQhunQ0W
Fdirp3Ba5wfNRD5gUD3+vVVmy5501MH47O+4QlYoDNeQAzXh9R16vQWqt937LOmIqF0qTG/6pUED
/xIdzprJQrY3Gyk+9g77CIWxH+D/yripaaByfqGfJtuqAGMJ1CTUtXITHYHA+bzW0YiS8HHtBGnZ
TpY2KtqoxmeFF6wEFMQjqLfhr6WepBGxXfhWSz02mWzJzFq9Cxk4mnYttr2KVdqP96B6wCMcRSCj
r73eqzH1pPTG2uDM+BRHlQqoHuXNFeJPZAd7bjyRzX2flu3YYpRr/pZcKxjHFptD3TH8vl9vKSkZ
Vm1YpjDp6GBhRJGCVJCEwuJMWCUplQ37fMX4Gz/ci2feT9TWS92u5fhDzPXywiMGzXkPZNdPlY9z
pHbAmygmml1ncztw+pPi0KrLytyYe7OHy604HxgOdCnCrM1cZiCAC8KA2uZzsqT9gjqUzN+2UkbR
l9hLyhgncZRgyQBm5QzfMR+ZCeKb680l5QDFsiPo2Gy+FiLb1TGftZ7PlcgQUh8NfHLykhIIMNG+
JhE5AzzMR9F+kK2jg3eSWvtwoZONSMHOwAOZxqqU18EbEE0eRh7JKLp+jaqsFz9iYy2pW8e9vevX
77DJIkFVAIl+bnvViCwGLz/tzTp9bhkFy7LUgyaMnSiwTi+nSoe9w+co7Ekg4UYYwyMerYojpTTY
JjwZMh5Bet64CRBg0GTrohkFK1YySbJ+ReG4m7lbSEmb7dTq7vrA3Q7cCYy6HThi+7lJEbdCVemQ
K1UQQoiidWWy45zfOgbc3fbM3QTfx8w7HI1zFuYVBA8wqCV+5iMdTZRfmfn5xKKG18lUeTCxVxS6
6VXcUpM5wq0A8dfTGTrM1wC8lRTYfUSwhVo1abRoxdMBB31pMJo3Ij/BUIYbGXk9ebhlMjqpAbEM
R3Xj1Judmz43Y/TRbxjIHwkEMSZvAImBnBmBEYVxTED6fgwiivfpiPy+Vm6utHQmEN2zZQbqqVnc
xQlpXV2IomGdnxozvLBv+uJdCMgKfFFbznsPUMxe7PsNcyPUejtAIUh1KBghzvj/bwwIzsWqLSJV
SENTdRklZql2sZsy3xBaoKClJDH6ujvw67EfqpW1i5UiNDZ2Vj5Hu2JERNSAnSsvU/a8CnFesyHo
RhPJmYPTZ6BWe8p3puRh2koiGwaHxyF5Vkc/JsYP+JiTMjRDqv5JOtwgywddR07ctTr5ztkrIAIR
8oKgMyP7OvuDSluYtilbjq8MQU2Deo/ZdVEJbraKK7FJ9qiGIYUzoigkFroxb9DFt146DYXOFhTC
KgU6El5Qur6eYdnoblIRrO7OLxleUK7YS/12coQstprwoxHDVcqrpxjaai3tPXSyMKFBLgdFT1/P
SgwFwy9bj3D438578YPl3vlzsbkBKfbmJ9l7/gmxlK4eytQGtnmf2Rey4+XVc1gLgbJafmUv6nbt
z4aTo0PGg88InErezc4v6ytfQdM/TaBYqdC2W1NbDBziPtsmmYxoCuNdnPfBTRD3PZEY4c6eU6wj
D3Gq8zF8a/J9IN8eL+cBGKIEz1np7ukxiFKNvYyvNL7pDjDEs+gfkZw2/aZTzJZwC4qiPSvvBm6Y
TM4PgGmgmnuyZpQCZ2J04g60P8GNEFwZI16UWT7rQWL192pUYcNZB0W/2uixcLtDGPb0OmEk2Jtf
Qg9KpbFziP7SfnROHcBYxf0EISCPYEpnXVFfTJPBGX3V7077cSCS5vBT0nqM9Vu0C7A4hNiKNAAf
sPDSmlCLChNSVmi6FsBa4WIH0uouTGUOfxKyt4YCevo17pOv8l5UB9NNhAAIy0oDEBG3l1b1WvAQ
WQNE9LwAx/qHMpAmZ3mHnyoi6dSuoQDJ0hcsOhLvBu/SXKExVurZ/dnkciGFVxe/n4FnChIJB5RG
SOtFjTTL0G6x+7Rfn7t4kCQYTPVI9l8rx5CdjtmNPmA+8zjqzMYIsjXRp5sJRGPNlxegIjGwrNyp
8pKMU4t/5/oQ49y9eZXCozZ3szJMeGHvbL4DEH/BRwCCRaz1T3ONbw5nuh7FUse7/mdQvjxLYDxZ
lFAOgtow6Gbyto3C5RD7CtUhr8KB/WLv92rPH/HDsaFy7SXHpKWOBl9Bed+wFLJwbdkm5oyoHed7
TVmnFq9vJO7l79N3x/xmLwXtpVoxSMKeL4grjlJIJG0/svpjGGxUe5zCxZpzxTstB6eXTbJi48Ji
uptiFLeWt659XGcpIAkIxIuL6rTA04CxZcevHybPQoxZoJ/mRZCfPMTHhdfLIZjOZVlpSYUldxHh
uIwMkc/QQR/zw9MNzRWEGLjkjJZ+VSbm4+84cc5/qhZWVAZ0YRO5+kyzR4VOgJZ7yIemq7IRE4p+
DCuLxjEfn8VaNtOqzpSMyY4IT09rfMhdTiCnGEqKEhf9C6WAhZceGpzB+vHqn6SPyMlSC4qwrWAV
wlwAFC4CcVGPFZ9zycDmlTA00QcUszvNiIa74A4DrjUqRfwsNaB/6AwlIxKpz2OVvF46fyc+Ib9f
HjVzjr0m2YNub2x7mHvO1ZIwb/1aoJ3zxLlx9Sr+PmVOZz2D6s+Y+OKZiNcgFPVY3kBOxaihdAaZ
BM9AYndCpc1bYgoTwL+KdV1fDaP+tHY8S/aYJiz3L1J2iONkLFguHvecHIf3DoWp1vDScA3XNanU
uGefpeVUKO0RA7WCfZcFt/D3hA7vkyS7Zn3WdZhg3WTjoNDdS+lzZtBcVJAYGGCO5emiwcBxJhXr
6c9MkxBLZHLTl68QMVAwyhWymsFUhwcmOVK6TRB0eKg61NDaHX4l7vz4MgSZN4wbqL9qRrJN5F56
2zFiKfGA0Mh1NL/Qmntn5eal2qOFdjHtN5u046PsrC3rtepC9V+l1QAW4t9nfBUiNfaj/Nj3V4Pp
QC9c5Xx0fZew/AaEsiGUNCDzmeLY3z7MtujK/nhwYlWWisJ3YyuTII8PdBxMNYi9AePXC8WsoVf3
hXqe+XVHxwN0pkbZgXrDih5xFoliP7cL6puu4baj6rLWxHRqkH0Sx1Q/4Ric13d1sfubMdYi9N5W
09cAwYxnMMAmGOxtq9XOZWZF8lC1d30n8uXXxIiSyNH66Pv6pch+wG8DlVqlxDiXe1k8sjLdCI63
BhXCryFhqUE6dGej1WZe4wOD5nI4WcMBVrsKtimHJErOxuMbk7C+aFpPMxHM7c+AzKPO40ziUKtk
RJ8FipX88Ay0W3883FTBls1zsnFapruwb8xQKemYgU9bZUIudqq4OuPUjWkhF3GGi22qqPdfI4MX
FI9M88+b4bDGZ47mSsEF/XCV76z6AgqSA3h4skO04XsEf0ngD/HgT89gvdhZDyC/8nMVRLXmj9be
erqRLGOI2QWe/LFEcBRlYvSFNEeBONl3AJ6BB2bz24S+nQltJcLhZGQmsXPawVBdBlIWUlAxrF6N
6yHi1csRjpj7WhHNa2ffIkHobZyHz06lMs9cDTVD/74Y7lKgu4m1mXUNOwy+msm/tKPIIP2tpI28
aXL9ZICUC05xVHDDslgFjxvE/KTpTzhrlacDJqlM83DEGL6lXmDlIPjTjtzR48+bmVRUwYynqlMT
VOFVoehh/krPnKExD4K+grLFLx5DIcKiDFTEHw/FHbTX34y2Ux7xvVMjdakESB+eRcaw0QnAXGZi
FY30xCLlsMuIlAihcd94B4y3U4JxKEWUb6bNwUXxIWwap0b1QGC780xwKj7RK54kwsoVMnzFGn30
fbrfRWA51lgKFHA5EKbs/dn+5VfenFpsUqUJVbcCJkcjprVkOttH1I8pkLIHqItx/4FqWwHFMnkp
ctM1dODgAZnetqtKLAB1t7UauqCioSorkMrbv90VZWk7ri+jJIcOyxjSeVpsjgupmA57+bTE6rTc
BWRn4yrel0hFCJRh++LPobmCnX5J6+PEq49CnO0iOXBDTsgCfHzBkBHqFDvUk0jo4VfxK0n8pb1F
3zdUoK5js+WXRG5S3Mv3uSDRYS4DLkW08kAwLNXLl8UpvmsEtXwKNsuwCPWHzHV4AHQPucRvHe9n
XHb9CQlBzF2Zx72rUHR6EPS8KWBu55Jqa8ofoKWLE96Qncq+U78E2AKqq5sUXy9IbFnE3QNcEnko
xT/UgK0HN4pE71XVkCNMH3yoGwHE0pdr6cvWWGdMQ1huiNEu/k87JDAypTjPOKEkk7+amFK7hUdL
SC6n+nx03fODb5JlQpJlWuk9owqArrPe+JLrE/mrBnRVzelxRnouaEmuDefQnq3568QHtWlXxu3y
8YEme1+xHTowmAg/lK10CGT4We8p7AA0V6ZlEAm9B5ohk44B5lJB0F1JFgycSWX5Xq9Wlp3y0b5R
CnhjUZuD/tN9XbLoO0K9AWlRQoaKvGrOpAIjXxv/yz+zQOEBbfthIA9j+9lfI9XaPksNB/UL3Eso
FAM/Rs/jK6j2fSE9qfHH+fqUrKXDrQelHBI7gWsmt+azi4t3348Y412VsC2LNm6/td98JJ3mRriP
U96OKMVIPSsytwxRr43p08AoniSPNto8cK15IxGubPqnY8g0eOmQSoMjBY3oBfd2ibZRZ2egU0bP
9Q1EVsCuHV31yoKOLk+1WhMqWsz96YFtJ1W9MM3o2UsrnITWl55f250wT1DJ3sGQZLsBdQ8/svrh
aCXOrD6SvK8dtpE/9wAgBbMBl0eV1hJ9rgVQIXx+9ozEp3Jlq8nHFa4CITu8HJa1cWb7DThKEnGL
NgKJUWR5KVHmsUiaqbaYT6L8r70jD+U4ts8dGH6fgc1mgR4cwSfvVWNaFFtP5dxN8HOTo4P0hInB
f3ZLzUboCddVh/H7J7WCosCmpEi6n2Oy/YA90PLBlK0Doglu4ru0VswVMk95Av47+lx83QswNzE9
ZN3sPwY0WQLrR49LNA3XMO4/0Bz4717nktnCQWA6MDy6qUVH+ksZouIJ/1LRtZ/gPPx7K1sPzhJk
bm/21DyS5S/DSVC8xH12HcwMpuOhWVj+rJU4irVCaZlb9q2/xEHFBKjsPmGZTCDyTEKtsdCSyiAV
nGYLmjCWbT9QbH4pTZZqEHHV3PQ67mu+DdWJmbPP4TA65iGTl5CBSDpDvkkOBav3YKxSSFMg6ZaH
+1hwS0HqcGPk1CSFlHETZpjJ4/rZG2EEyV8WYNznWqNK9V9r8R8Qthd1Rcv+N4W+LJlrPQyvhrsH
4rXhrTB92SKXmUvHX/DqWVSZjU7vVq994mj8V7+KTVU7esngxHUMf8CFzEIuEigsLytN9+GCWlOs
4us1klZvVtoNAwdS4o3JZHdnw8mPBYEWG+5FITucXs/aMmPOlWaseoog9NGCKjCRB2V/L2Y5hfXz
hI10IJp0owghGs20jrEYW0qryyLNAfxXsb8r+U+qbLzDP39UdBFYaGKrxBb27Cp4iMbqugX/9iD1
QGXlw5LvJH9eIlsTkyCZVvx4jEOcWMK165zKd5jh2DFubJDADSfPWHGjZxYOytGaNUmp1FPr2CL0
AgoUp12mYKdejJS4JWphJxKVurK+s5NBQOGNWj0XDxwRo231W6PtKsJaxXJ4bfPBfCu+xixe6ucl
qLWxiHumWUxkAtateD0vQqijkJkLJRqlXBn52v/TDWtgeEPP276Tj5+99VOSkySjwbV7Vapqtz2i
Qe1aMoahlfe71bqBJ1lrJoWe7B7dngRCf9B9Xix4tX/p2F4Ztnuq5bxfkigdqph3AYudnyZtRCBt
cTmpDk99iB8E2xebP3ipmsAAtYABMmwZkzVQ92M1HpxJ8g0dHGMg1KU9klmzK9b1lox/FD+UiRgd
KSfXop1i4TVChQLi51AjT/plXUNxOKoYx5jc0RwzhmdycApYOYsX5gceXYuq1HwXZzPaOOptFA3h
1ZXne9yNubbJbvPrumShxIaPP6mGCw8xkXztulqPCiEtT3n+XrxqfHQ0txQf3Wfa+VBWa9nkT66W
wR3aGxEpJ1ubJec46TUfXQuDhEntJKDjJ/oCXm6r0vAM8sDFNYuf4I1jbMRFsK0K9BTjf54Q8o65
nd2KqRfP5v5EFF+ZngyQA4suVh0+ogrrVdsaRDuqbUVIm4v5ybTZjfk994ri4cfnNBlOajlCnQkG
um4vU3zmKERJpboFG6jmAe9ClTa7g4VQLj80chtQJEDoda69bd5ugWCzGb1sf14W3jxHytQPHIbL
jGIdBa0HL6tZLff39d+12D/AIZMEGzMAsMdRW83X1EKJGRJG66zQDhndd36zJ5lO+HWQXeO6kNwA
k59UrFGncfAenK0FIfgbW+OuPtfYXMHCGfWoRrsqjMmgwrAPgMebeUkPxvGBmxBNv9L5kE2FKQSf
AVrwo7Sy9/ZOADqCes3T6eNMxN+5z5z0KdjaljencMVBjn9X5XRiaz1OrYZme/XUNnPGtXV1lFhI
tHNUwtw89Y9Ycg+7AHWlyNxeWEnNcz4LuJ5ycx1ZOMSO9EUO7CyiWCazc3JPxdf1EYm4HZx0vxMy
HLxWX3xbkB7yB8rPyZkg3juuyleN48oDrHc1mmyjUoLt+zprI800VsJZAzlfX2E+gWNOm+U90f/a
QzDKbJNLQeNQt2v8jYSjhDhEZrGaXgtsWpYnj/s+INBRtlxC6SjGcsFhJZPil25/dq0bdCJBR+es
yPIxuUc2LzqmexC+DifC1NleOFCZVH2+OjaknTrCq0I+z2HImNhcaUYy72ratte9G4ADlsYsBpp9
LufmffDwm115cL7sgkRj0UIz4qyTvpQq8RQQ8aS9dGyzQcrZsA5WYcQFSwJuBlfNBObDcHzexj8K
YmUZFZT4Ed2zcQa8nLOB0PASVnbsM8+Wmtk4eHWznteAquh6PpkSTYvTcgnMGbN0+H4wH8RxMcKR
EZMK/TdfuMpr7e5BlT+j+d2qu/VZCwoDJQcsyJ6XnsUZF6wl+ZFUnG1kTsynymyeUOfA87+001My
nMWMYiHOkTrGExHpr17GkmXISVcSajuDxtCj86XpxslPl3UbPLseMUgrXyKy3SDrgKdl5oXsRZSH
+1t8j+pW2gvlj7mJ45tFZgSHQlmbuyOV/qmkdrV5WRgAFo50BA4BWdXC+Ics7k6yBCpbrNJQih+w
Minr+/soMmDaa/tSO+WP65kwq3u1oq33KHeFitqByXHe18zEUW+cXSqtj3DQ109JHSrCBYkIAVLv
HpYGqnmCy5ENlzgNeM/SYLALFW1ig/1T3Nrhq8obnOm4dGhm2bdL9qrdpnS7kQ+Fl6Yo5c+dS8eo
Ypz9GiXSWon7Vx9dQ9aNgaiYh1pHMW85O946N3/7uKXhkIR9PZ2WQikeM10iq9RBGEL8pmaQvjfi
po41MkWm2U+di3sZTtcOTjccVicFkznFDI1i+cKZSSB9kQydFxVUqU2C6VRMhO/praqJSysqnLhO
ewwGY5aEYUtZSJ5tV3Id/K7McULE1/3F4r7HR5LxGJYogzCiRtXS+gip2mHkMCiJXlq7CW4bJcMv
G38Mk/vcHmAG/LaqCFjGcqIW4qbobsgFjjBM9N1p0ijtetlzpaqmP4MK0eopwYI8Lgl8mrKhrNxt
8PF2X/15omlFFoWN8+MfnpXJS8Cg0ny0FVCvSwMEYzVgqgm41jUJafDOjPFYbhWU550kp1/nq/mK
Xcro0yJ4jRHVbbfZa/4JcpnkYPbvDZqvTwSGZU6AuXXAEbW9e07h0k1MyFbGHaIVEZ4OLYoArX4F
20zItfe1x5Q2QCgkl/ozEBPmE11AWh363q+MVoflpqnTiGyQQ8tMGIR+bLzVD/tJExPhBxLkMCVk
o2BTvdqnabhaa9R6tFvEADq8Wz/dFuA3d+3EETHpqzOI+L9sX1xwiwLSO9PXf1QDw3w5IXoXgdsj
7ekCPxxvD1xGABWrmwOsHU5GuS/fLwevcv4eSDnwy6q20WCcPap2KUx6OSxuCNvfZcp88xDYVAGt
obFfkCKF+YW1uzJUmFhfwWjiMrHXJSLADc80C2xD+B8HsRjg4SL1BNLTNhzYQy7jHAnkh1XURDGT
qwssIIHSBY3RamgDAXb3uT9/YPK88T+5xbuIymY/a8imMHxScHvc8WnLVz/nyz+6PTVQj6CRBfIp
7tY/2oJuRHaB7ihbuCJD3fhwGC/XasGBcYdqG6pgybruJMUeg+GfYYClYD2rUXUOB9OIWVHO4N6h
JQ2jSlB4K+VRup9ZYJofgUJ5Wn7OJji0kMyuUGKSzKLtdTTAQV5LN0+yKpbkN8x4pnnlLJmNkqjv
JO3yOAar/S7mDLZXqFLoL4NGPahEmXoFmxcS/y3EvbVq2FD+N7s9/Ro4uD2yCgZGjRAarYskGPI1
vzIlYzHOFy4wVAmvqU9kge4fCl5qEqZLEzC9K7QrfAA1vcuXnZeB+KCtA0o0n91bYoAqfYoXXk7q
lfzIn8bic82Oqc6I7EKxujdlhO/9gywiHnOVsn7793FLzoewxBOZ3S4Bc2fzYfErpoc5QsMCnZJn
q6JmUuYMF15PJWKVTzxzhGrx7sAm0wbv+X/x1qNSNmtaKHKjmnMUexqFG/DXOUv8Yd32BzLiknTY
XVHhDAH5eFyrnq9lpf/n0BOiw6nuLPj60pKKOkYcD5lpOVsNE7b9Ck77rgDRVgCPQ6++x7nLzzTg
y+T2t8L0R8ZB2RVRovpSj9POXMN01g56KgSvRcxeBEo8ZpXQCE8D6xRKtZUWHVe3tKi17jClbEFq
tQK4iTQX+8qNSYbPVeWw1x6QXqzLJhaB7FWa/dNI7kTkA2uCi9Wq9pKtz4IEcu4lyz0oMhbFQn6t
CI3YEi3arBBta2B1FTBUWII+MXGEAbvyYu68XmitrDeVZ5Z3lXp4GrpTLWF+pmGgTnkgd9JcoQo3
Vz7Soo9QqJCq0vkYfa+eBhkAfu/nmriTQkNKfCNKrYdxxNh/t4UQySeytXmmgfWnnRUwW36cheEE
oS0QlGYjleQcqGDPo8dboiAqoGIzdZeRUkLg5tnFzq+Rkt2HSeeqYTd4f5uYfXArNDijGZlh2jJ6
dXMiTML3RWH3jbA7fzybLh9mb38jvNhkypiCGqKqqQF5mEFcU0WUM0k/Z/nbeHtUehZH2C+GGbOr
w3IVg4gZ7DEzgfDvT0I11DzYC2vSkd6rzaQyQ87nbxLeA4ndD9OGRxkEhV1y48UIVicNUk4JeUsj
Ku+SnTooTYKRb6wnY4efv/HsIh0k95tyBZYsI24H4LcJaMOiwM/v+8zFFIWjfE8De+ZSTLtQhIsg
io3QneR4oewt+276ML2xrSGQYoks9BrUlzYnk0hZiW8KwgtH5AGTeBzMWO3Qu3Cqh+W2h5MmNonh
9xnRTwXVt1bRu3s9ODd5CLnHbIliouRGdR01I1wkrLYGZPXkvf2/41QDjC4kKmnr4W3CHOqLf4cx
gd+TVVSUmxmFBA80KyJfIRQxUSpey7Kb2ogHZAXJWguOiE2wPAv+t8FJpk48iJ4Dq4kiQKcMcbYz
gE0TqS7fxx7Ws58JbJs39DbTOtwptYvIveU6WSxF1dB8Lkx0MeXtT0vYVe2ucfb9F466r327kjhg
XXZ+e9UaDenchqNHQPWwAdRuWewdZzm2Y+iGTMvrmLHNx+FchU3C/2lZFxjP4WwEAcMKU8zKYMwV
x9CCpIEfwROyQrZOYnghbaBDHAt3l+vAIA4SUsqFc8hnf/V4hVhSUFU89tzuKr0VPn6z6R4fSxEH
ft821vXUkWvr173V7zEwYMiKLUumb1lC6vgc+Z0YrCd6hczP8eH0QtJMGUvelf+YQC8YEeaNEl+u
sf8pU7qp+ZV6Zoh+RrptKghq9EHqv1eHTItOKr4eO8xsxIgtGiOlwBMsImVr2x0wGNUeclhqIbRo
W1KJ3IMmXrx3CVzeN042TZfJGnzT338CqbqM+S6LQ8qDYxyvgb80cdeS5ssrZ9iJDDYvz6F+3MvK
uNc1MXeyHU8yEKs35ajCsYHN1d6bN5lrZyX3SkXqy8YXMpjYucx0k5b6e4mv9R0xEl3pzOlqE22J
j8MdgB1LL1WMgjtEsAAHsJ1fkdl3baBHIa1htKVEmHrVXV5KSFf5SEWSFS2FoNAHm2/dRBM+xO2x
v8fsOIQ+63IUAgkj7rJaE4e2PTF3R+a2ACEXgVVf5Y0bR69WRDYJAcxE8VSTA8HfKc/4jsNzy8gk
4m+iKbgkzIo9iU3On5XGQADG/3mlNiMNBXtOzA7KNNza+wxl6z49Vor00f2+FsHeYsVgy8es208H
NYzOD4JybQoOKMeBUGCVqVG1YLX1ikxrqjxCdeilPXCWJOocAsatUkTS8Q11aJ/tMe/wsecOgxSV
MNQG44tlrXMvMwBWIcgVKwbCwx8GV9UqUwetWsco/g1WbkqRQEllOpp7pBX0YkO+U5Wc+pI38pV1
pj8iLAki2cs0UBD+MHF2NmthiGomjKU+6BxAkHrWHL5L66NfmRLuPKDLLsMWp2tNvymrVO0XYbH3
ZPEdTN8mrzIEGj/M0/HyQzV7SN0QE9P2gVzXwobj9piqOmT9oOqE1scFJHOuZ+Yn6a+i1Tm8/H8Q
gP7W5BAMHN79ZAchtlDb96GEdh1cGzg36kI2rTewkKnPHDt2autxfSrWCsX/1rJS076weTP/AOmd
onaRPBZetOAQMT4z82mmDPO1luPmIT+gpmF5nppqs7HPg9ZkHwwG4SNWiNPPJqafzaZlBrP3IlPX
TmT6+1AkXrjdc3sQgOmxnnS2CTlHjgyfGdXnw6Vblljqc2A4rV2dBb65tDVvwbpAQvyDKyR7pgtY
nurbesLYNTYHJga3PnuJai9v6UPE1HOCe8G2kRp6eYzF6bWBVhC4gI0za8jRYfhuQ9U/Y0UvlGlA
DyKZWGHllDMVoTj6GpQB8SNuKDfbyG73wieT0TssctJuccfJFmTEEmvcWPPD3Eij60In4jBOtS/Z
OcPq+U9EZ/DVdG8vbo3g+e5Ft4RmmE65ZzUJc6K08Erbduv3doxVtP5uLiwPD+vMR/J188NszwX1
6MEbUrZ7aabX62RCIZI7RnQTuAg7liSHPrECBfcivsR/4GmBnijF2Rs5Ddk7jVDXR+65BtRoKr8v
Dku7abuOISvvaEYlN0KUA6mQi4QpykqBzhXo/tQleGDA8JO9CjdytGW6dqywkWV5l7AReHWkqKm/
c7SMVKSc55HqMCf7HohR53nuIYPFTh+N+49GcOfBivEMZKOxzLA0H2b9zv0q1zy4JgoCyQ0GoG9O
v9iENaNnJUkFs7Y1qSIMwgZUPL33Spw1kru2oZ1DmZsbVmizk7l++bUQvqW+gtcNv3o5j5o/dCCf
wbJQIC7rAZX0iAp52XU17Zwoc1tMLeiw2NHytfvqWLlmdqLDoaakKWoVbVTVljs4JA2G60B1oEUT
GLK52Ed8d7OvbSb/nlaxPzqQuLoVYwPpIJ71yP/CNXKt1vNoTEhI8y99HdyvKt5eGoDM/I2H8Mlk
iXrt0zLhHDnhMHVylyecRYePhjIpmcBvDibkacMXc9K+xoCkutcNBvNd+0Z3aF11yQ1G9e6jIAhU
XCNN+D20QfD7ZB773y5jfmGHW9cT2DfTdPZQrKv9uypvNEUJZAF5vEjqQXrv/NsXfV9903GWbWeU
0HOzPTNyqXJUUGVhaAX5TX3uGP0aqAlTdffMy2nEqYcVOZmNVEjGpz/CtMd17EMNIcHmXxsE2bAi
wPaejw+R6Yl7gRssSa6cOf2A5c3U2IG9rd6kNRN5q4W3WQXZpmwVQsi+TupaUHuvqaSPB4r4DzeI
/aKA09STy5cx0Lk/WlwMN85GEFfkv/dW596ytWRtZpOWddlSjGfWQ1DCxyYptIRkFfTIDRDxgSqe
CMCiXiwWv3eG37YUgEKGjqhaBRJoubMVqb46HzjZw+HKLJwkkNyhmpLpEYVT2zYHbiEBkCg6AKMf
5ZCHyBJuE5g8M3NuDVM7AFAKvg7iJJxa4UaAo8WTynhjm3axYk8SKvtvKkObXrFucIh7MFjqD9YQ
RjKaXZPiYNmhwWWoMuX3zpCVBRSuWxtGb7u1Fp3c0Cv0k69Q79kXAioAosV43f4YwmqQhDYYnCtA
8tEpEc471h3RNEp6ZLvMHSfnfQm0J6ZO2AjLed56wgTBURJfZitD0AR9oDQ7R1CDr3qh+ET9fawq
CO3eWKKga3eGCxD7MwsNJYdUHfJLzAGKjtbVMs4AboV1JxD2Q4l0AB5r2gRPPOMXUZBM7rNtXw/b
izXXIiitkQtJwiMFiQNnR5VPJrN78pV1mr5LKocOUrL4jRdKtKR1INJY+vQ8gEjp1G7vPU+EyGv3
nJ9wFuLsY1uPEDp9kbyfzvakSgX6iU7vP0cOlMTQ6GO0lsclqZK11ChqqDzQXplcfHTwY2kbbQOL
ZT5IbA0AiVzpCSEP08hUAyyrCWzVcV0Tz+9AyCXYkRVx8fn3IY7F2ulWOm/BB5LNNtmysF/6ssWe
VcejWwIZW+WKwzL1O+c02HiBXMeCC/VPWQV63XSCIzC+QPHKrlAQDVFwE8hIFBMlrn9SigQJ0BSv
IJxGo/6q2C1xzsK3FLHRhuTlZLHj9lvIRtHqeeV1ahtcResfFfsJA0MfC7FZN3nEzA/Zy/NOebNE
n1HFZyAmcQiO8tEXOCTJiw8XJm7h+Nud5gKQvjmclNZagoMQ77JR5NtHMrptUIQQNxmfsEljYupo
x4bjU3e61smpRnfA82QkubSbzk1NYYcsHBmp/Yhg6FWFmF8y333PLLytXg74KMIkQ70wDfKAm5Lk
XnAjx66v98Yf2ZUvb04cDacfUOQBqlDe3AKjyDJ5tg9ZaKXh1knt/eGsmPKJrQ9Sb9WRxlOT7Nl7
Tom/fWSES8Vm7TUsFQdublBPNc+atnjclJnBQy599ZqlPkXLlv6WoeeOxMlQTG115MS+2fBCsITU
PXX6wDeyQd2NwqqZY/E2QU7Q87ESdIGrlUOvioDb1F0XoGCvbXmpcpbKMHV3Wdienuy0RR7Kjxi1
k3RcZxF9j1nQzeMmNMKKt4EqoeXGAwYrxBz5HyQ4q1dj8sCUtfL/xVz16brqxV2hdCfm7Ama5pli
xb1m/6lBG4OHUQyY8uYTryEx6LHtc7Xip/TRcgx9jU8/oIANKqFuUUxJgbaLPIS7i3mictEBY8Lu
kpu17kzgyBVvHFaNm7/6O6iU1qANksBL212eHmCgNXtLUgCXuYtPMvzzpdf8QQpXaXaqZjce9m4u
ec8pvmY7RlLgTxchqtJv0giX9suHvYVj9rAJY8tGEBZDFXRft2WVVYXL1+5dLo7DfWlV2AaUIJb4
S872LxwRJ39iJQd7RacBe1DpGYCqiWzgWkUP67ZmlB1fGLgzOMvQyF2DSH2YyzRwzREWanGDfd/y
vWzGl/qksCrPk42KK6I/evtJNH1MIHNj2WWN55INj1aDJ/Os9aHBH+WQGQ4uPKPpwNpBtHXNe3Yf
aCoj4VWvNDVxrkQr98VA4HJ8ie6gUQ/Jxm6HfTTsv0AV8NpatAjVTxz1L7Qlny2O4xKoSiw+p+Mm
VgbfLJFiYiJL29hiKgMnZ7ZOLC8FPDe2RR3N2u59AZaWpC6KqRoiN/n0js+VjQE2qy3zojX/krrT
UD7unHC8ChXZpLGP6K0CTSmEZO7a4ClCiURBu+NG91WigJKshq9PK8wA9M4iMy6J5TmgDgDCn9lS
jHa2AZza1boBHDYFarcnC+fbEhjnl0x//iE8NAthtHcmK3LE5Tr4tm09H/ZZkvmzqE2xuIjze/8i
n58/zyKlzDgKccPH4d0/Qm5/2p1IZBvENShhT09ZpXDjtZHCAqTUG2O8t4U5Qiz9hAa4i8F7AACQ
pk8jOtekdi/5zL0hoMXZnyeVZkZPSoQWAUtzRGez2o++qeVYxXH1CruZGAg929dDwN0o7Y2/bwye
S5AWWvLbhWmG7t/jYl/0rHTfeIWsfaiAYoDJ0DS4r8BWGwbhsAU6zW7FYtYrQkCtm+suNEW+B5yd
Hxi8GMbvM7W9LMYxXIeKxqJQnAgWSTTL0o+BA4yTMjoia5hTx29Ujxp0gyuFewL+YdaAiIEtDQE+
wpmIERHmvOmsX5Y2OzmwfDIEhLdHfNhDeT7IksyqpM+YH2dmf8ZX0YqAzlJ9tHvDlm6MrAiIIGfo
wk2gE6/sIS9Gs5kWddPt1iqeqHVHLfy4qk+4zJipe1EOZGcuWBV1A9hGFQkfFlQMX6wCeyIMxcDe
MWaDeZPitmepPK5y0AwIgbM0X0g01Zvrbt/+vWNJqzX06CQV3T2qcBOPOSOk5s3JzKzkqczQqnXm
rpljxEpe5lTSj4E7fJXN8U6AMnumF+SGM417UiUCQdkrjW4gHXyXd2toMy5JQVv/PjolIKZuFx1E
lcakAHUNwar7cXCA0DT57Ef3kjeHu3X0tt6/EzUoJbdHFGpMMh2nF+8qo0rhqU6J1chcVyUyG55k
T+EwBQBDAr6ch0CUC/qLxt5UV1n2ZhqX+OMjzUr6yIkJ9FT/oYZVNmwL6O6Ib/ocGOSx+lvn82A0
CEzPqo/g8EdbrJIPKe7IK/VnPjEeNHjuwhqSNkt7KlvoJWtjGaecwimRrkrXx1s4g5wXsXs3oe62
G/z5xjuadmCJUybvsaAUSQYSQlguN4jIRHCqCFsnC9KEtMX6kPZggI7tqg6Acq3BDYtFQlu/+U8U
9dn1q3tWVJAo4tnZaaVheOr3dmFnvH1YIOixDbvxivQQcO4hCk77b3Mx3EXFTO+cAvjqa79q+agK
Ku8xOF3k2u5Ks9llnJEOm1Sdiw3DmGShUwK8+Pwin/SqS1Fc0e7L0D+ScaxlI9r+50aJYWE6p/so
dRLFg4APcFfgV7EWbwkPnRRCvmGp8Wu4Zita1mmcSld5OsBqN6MDy36P7DW4m3HnOh/hr3rsQttg
0QIIPoaoy+IgCtnNRUZSV2NvOfxseF99b6BQJhwCmWWX6OKpJh1TB4PmsAI+/5atP5WPe5WxoTQW
93X+vEUU3oEuCFx0oibLlFEtpYNSGBGtP+NKTE6KtDGSEpHlFNLDAGDG4/JbeQbptxbNN70dX91Y
nwpU+vyFg0B4/3Kh4Wke0UVvXw0TAUZfT9CaatNQ3a+ENZnnv6BKvmZYJ5hKiYSA2otpU8eN7t7F
o2UDFm438VVkB/jm3eeE1GAH2eIdlnyNh0q4p3X0YE8fR72miuB8lccsZcHCEb3mKzr+8fP105Xr
9rjvXgQGPiBFgw1OWpZu4B9JN0hnhYHX5Ohgp6sxEqAXCEB4lTrsNDeYBynnPTFBnSjKDQ3wJLHd
gCevpf4mUPqIn66G2dLKQkcXRdURvraQ4x1Y3OSc/dt6+widXqdwi1GyYoPZB3oD/LkvWeo3mxY3
bd6sY3AAcB5RjwstjFuTqFfvtm22HIpv74r/k/WvYc01Tur0kDYWPGSJzb40y4CrAgD0ktVV00YI
XWY82uDgzWKAeFaEw+MAuE9UD3+UDbriwCx26XXfNXBDcjmCbh+wP6l5CR61KaaTKgxJ+PHbVK1q
JQTY0XQc4vDvwslfUUraqJygAUuqAlHip9AimfiPhvIn6exSHumMzMBB1I15t/nSJpgXTGmjueOj
++NRRHWFAlkLj7D1tFC6ngwIbtXbiHIoEzBibqWSesxJNJ0IBR8Nggy4weZizqGMDcC0LhFJ+/4K
cETi2UZTppqjKfCpnqdHcuy1zwufDVnRfGobdlKKSeFs23rw9GQLpjw36VIiGav8fPObI/C6jIjM
uu/YPRBUB748qkpE3bghLj8lux/zQRESibhi9IKjJDD2qNQ78s6L+p+DAO39WBrnP0iH85SLWj31
txTYZ2x5oNhVunDVbKgvmd++MhcDhDnKwLfhWjoJFOwiIBVx+ecQee9iW8WXNfJ7k1xmWbwxWNxE
BpQrk30S0w3haiBOtn3wSyYhW2ZR09aSybzfUJbH3hfHylSJ+MCzW0dVp0goAq/cm1RSNvx0KTYP
O6E5RIACsmhIh8z7hXvxCQ1gyBwZYJsSWZGT51Yqcn26anZHdjLM8gDuvx9TObYGajcp1RE6E70x
ABckkfbEKssV32SnPpJMpdZ5cYADyiXYnO2dkj7m7KYbscfA14dpLL+5FnzzdfLkjNknYb/NLYHB
rQG0ppx66zRu2iWLQI5R4TQq6apKvHeSv46uZuaXgHfEr7zhbeGOnZsWXPOOQNa3XKfdoTDUxHtL
twHXTV73tjohLJcyA5TVF5TBa1+bBYmw1Esdv1zuLqauXF0Annts9jiD8blVvCn0339u3pUm9Lwp
GyMCJ8/3AYBZqvU2+pLUz4nIxHpRepBR9LX4noU6Kk4o+1iuGEbcik51KEN19E4+MiwdJwJX0tTR
FEj6+JpmeHqTQmakA1TFGt88/vrnHMvaW+LWCLxGb/KPZO28TVBRmirQhtCmsEwpK6p0ATeguxSE
tyP9EhesA0yinKNMw3uIgM3tjJMd4JlsxMycJu7MnfbmeJ2ZT+tr/CVtVPCC6ib1Vs+O4I+PtyJz
53yWxFBWgRmDovgdxff6f+H+VbhyrTG+MTrJWchu7j5xKMMH1TzYBPrfW09tcK5XnJJsdTYVi0Zz
IUjBHU6IZdoQfB++8e95NfFCd2xDFw8R0wYhXwI/Lvq+sXMg88L+nUs8t8377/U9oinPtUZ1kmUN
yyTx7wrgLPaXynVCPC5BwSL6SgIe/k9pUsLWzfiS+m2e7N1YTLw0vxuESRqhLbX4sMEgu93IwvsN
Y2NmXZkrIOYfpcL7RcoRk/WqOLn/8coZ+ipDiK0eI4lrOO4y6xzCo3tWVGm3VL/Lxawe/jnDTbh1
B8MTCIhjOfXLr2EvzRIIL5WdEuKjTfg/xiaXcKeaKUk37NC1c+ZtwT5BmoyVKvoNbCjwT80XttiC
65FVZ7Xko1fS39QRM/OjAUNWrwxqOMypex2/h2NCg6Chmgn1ZAxcfMTl5/zh8djUaLzu+HYAB7KX
ORhUl53QklnaOgVLDjpLJzKOj17nABefItnmfGzclS7O6qSglfm9a2+u9dBdWBPNiMZxUH2TZrg9
rSFqyO/+5tVaTNZILoqdOfqZe6I4dginsxOWQk8rAweuGDABYOyIZjy0ZKpi1K/yUqEN8K6gIUg4
5Dw+BeKz68Bxr5q4Yf8xFLcVCRruwrSoRVk+7FM9ClytTfj5IoJg9ZmFfnIb0GCgeZ45obKFbDTy
Uwl0DnszXv4tPOlsnK8XGBDSlW238J/+MqcPXnlmPttMDvMQyRxLv3ODgCjV0G9GOyfN24dF62YK
GLzXBDASmfclHg8nvW7SQGO6RM3Amkv0qYbYwhH7HWGJWzlP3g6kFuCo0V2O5d+clDMFlnFK02lG
oLgrOmpvwxmjCUQs/oswP2vakZY1WO/9o7yWFqNbktJdUPo752ON3/cAZpWB1kvnYIkyzRwoI8Z5
v4fu7bWxYmZfDVxFJn9Z38NSn/U7nBsnQ1g8hppVyk68XuSEBxwWHhYISIevUXgkL+nZUiZUjTxV
zQ+diRDVxYTA0y4mW4aEVyPJ/Oo/0Lm+JZuJwzgPPOOY3XywuQR5p9kw9ny72lvo9zyKot5+zZt7
Cg90WJ3Cg7IxLnCbffEhyO+OVOhv+cpTG9FGquGFxsJ2VQF+pUKbiaWIOYN52XkAMWzsvM3gPOZ5
T/UiHnvfExz6AmGbrR6a3318/e//dSaEmMHyefJewj6ky7aU88Qhn38j+Tw/5yQrNuz7Jx6QNij4
LZAwjxcpR/Jup1z2xz++m5LX0TgBSr1l+EvERn8TIZhnfhT4QGjARGZnZ6QAERRCXaGISrU0trch
Ki1A+3rXVOI6NXbspanbOhPLwWX8l7ZKT7iC7qpyt9+91p0Px01yu8w9agY1GYkWlQN3WNMZ2kXe
WEUnpasWoGTC48YaXzJkEAzVoqAMWNX4OKbG7Y+X/JQs8lJeD/fub2pqHVdi9IIdWyy5TzkU2Zu+
3ZaPb3y0EdvvhNoKX9zsmU3bqYZiDwOUX5x9e3FdSlfgXY5SxzNT+Z21ot/1fI6AFPd8qwNn1QHb
SO8MXrwNfbDRIhWzKL7Tw29BVxjo6k0WXlkTZZfUlbzgnblxK3o6jdcBZfU+mAmAx4VxFytn1A7k
0ehHdKwb77gJ94p9gNCY4AyvnDeVhJusLUZi1u11JtlBfAQk4a5uG9/RnMgz6Hd24bXGfNex3gFT
I55vEgF2I6SYYTc/rXceabtM+WOcLCpGEvCEPcXIuucxdBi9wmty+8ZQGrQ8HK9QvVYBxdAJstmm
qWgasjvKYhmEB0QUaABjxJ0gKr7rI9HuCHEgohsQES9+bXxFmLwD/hGMPRT4VXfYqw5DrFG/NG3S
5B3fOuiWCfWTZVXt9v2MDM6RP8fkFGb1LZzOGtGbyJfEF/DeZkSPW0LZQnLy/Hg8CWmQXeFVp7rd
iI3GGdIbSabGUOVhe9tmt12u3jqnlSCJEWG1mNhRdVrjAwc80X/3JFr2YfcWoHTXzdA7KwqCydzA
mmisS6V8f5ILjnSynmeWVMqlGw8aAU47lZ+xCRH3WxBipNP3tdJUhWvUX11/+rtHIz5r9XLg7VWL
Cd0ZHBCvTdpSxuWCIbbSax+Rd4Cist+1b+sK0OBZnwqf/RPyqTJmQel1Tn2WnNwtCCJAGXM+A4dJ
9oixrbqKXuxxW3YxpiaWoAecgIhtOnr84YzxVmrMIpF91m0B61maz4Xdr4QbGW3+LIobLO2xAIIX
IWEWO0X8pBdxrdD6mTSdCFNe0xeFZX90VIbnOLAimIqHB+JqkUydC7IZ394OxLvJEGLtwHDDDb0m
MfGdgtpCmUY2EJocvydoIAyDeO52DGrlx3+mcuzkUGNJOSd3WwTOafLzNI8XXs4A/tY1Ca+YaFxd
QsR6KEEiIPnecTfWJqy+zFQrerMFHH0rB0zOrZruyE8Da5o48x7feCX6nRNHrZR/EnlWSIikEz5l
4E6+sQ7/j5YCgHZY7kAkrwpu+np+0BY/8kfiUL1glLPq+W5TgWW3YyDvwkkfj1px5bL9+K6YGSVk
I9ohjbYlr3+H6FJniRvkh7ZqSXacZZ04GcgBO00DIqT1a4PK8tVahyxqAEp8u5Md5OQU3hRI8M/i
cBmq4By8KJhsfFJ7h47kFXZSM9rjFpI3qiAfbyQpfjNOFcCcrIPcVWNs2zKqI3rdRBFvtym1GqsP
V27f7MzjdPff9lEwPTCjTWYedRg1wSx5FzTttuTxQp2KVCgSEM7+U6hPbi9t5X1REoqZoJviU6Xy
9yjZGkK26PZBGdIKy0yjVGaI3Ffh9ujENoQ3w/xnOmdDSwh838jOrpzznQdMavPH/J5t+fKQCDik
adroDr3BKIIn5BP06EWi6TiR3FJa3HWo51VF4JQiBfIEUH5TPIfnVSUm1vZVgiaOB5FnszBAr27w
ABvlsDPDwlpygTYNDp0WDfJI4WaTLUvUnIvj9zKrMHpnt587JyomBw0TlXZoFMveK0mcS/DBVSfj
e9KvxuD+IZzN4QpyJsKlyT2gnn5kPgxmJ7UzopUdMkdF0+yz9J3b6hs6nBcDw3oHyhIWIzKhJVwb
XuX3pv3TdKvf7UEGcTP5b4r5Ir4INvFy5NIryOlP4GKV4VP8ehOwl83ZfjQkz6x0WxfMXH/GlvUv
D81W8+Tl3HbtiZxPqeNeDhi7ImYvTxM+TlkoApIWy4XmV901D5UK4I3VBG8WdTzZXc3M44V+dIj3
IaLlN/fcwSRrwGJQbFjWDlM5l9V2bf5SmO3jXhPZGX0BQWaABPiM87+EHxTSO4+A60Nv2JmSpz7k
21Q9Dd4r6uWBoY9fgYF+LqgSjzqzb9Qrc6CUj+K2pX0TuWQd71oZKb4cOhrQDSnnZ5fJT/lbdeCm
wvUieyV7V/8dF0vD0GVbza5/7JRI0lPSYYurWH1FZEPmtitJEJ8FJRmbVZyLT/0iPHmRJrLlRzf4
pefXuBU1d5Ztimrexy7HHImbFYRiQPQqgKUba0speG+B98dJEmrBlMQrRmozi7nCSTg1oFx3IgXK
cqFmWeGunuP9OV5rBb3ab4prXtXFEQVNhgIwjuFpyf2DHSYb6fdr1RfHCgaNX8Rq7i9L1Rv84pvN
p67HUsuBjAhYiI1waz5QwTFJ7Ait6sU0NZQ6ehy/IzYpSFesKWsETcjvmEYsLr59p0a9AkQNCHJ6
OqPp2bUmHHgFr1Rw0di+Zkz1BLTShFZ/kSHFO6GSrzPc+3mO2DqPFtth8qWrmyTmenHGnJZgEmF5
wpNsifIUEY1/OBcAd3TTg+C8F59tBOjSd4MFxSmJH6nY3D4rz9Y7cGBgqBlKDw6oIraEveNozG1U
ax941AO0xoibOdk9BwyctTxdBcrDugxc0taQNOpj/U0RVm9AAQKbXLt45EqqwT20SlR6c5SuT/rE
GeDwcLortBT4xaxMl/7d5kg65TSaVK/a7Y7er0CNoBGiHbmd9BIDrkupU8k0fQLquhpoq9uJvGl0
aa7ZRhZzU0YMnhBorGl+4c6dGsCk1Po7RqCCN1GB5cHOdy0ZoPSPx/sza8mhKXQ+TthSHzgEbz+X
5U6EahpMaXFwfZN4jCA/QywRj9Fqr+zrWQjJssRlKWRP6qPGURbR1bZCG4xptpRqcYS3ZHavHJue
hokZZHCe6CxpCojI04F5lJj6I9sV9zLF22DtGRFHqCPWxNamtGx0lMrdT+JwluT+ENLCtpW5k6MS
fOh2nrNa1ITXyZFipD6htlHIcgnA/97jzIvbpDGlIv/pcYeRXvtgFXGDTVcfJR+pFamX2garOTBr
wOunIIv++1b0Ly6EjUNoNEEnyYA8YfzkwW0+tZ7WldjGtRhNyKAx1t7ix9s3toZKt4aMpKdzNRTi
QoMxrWeld6IpBHqJi+nr9mJEZH+tOQsVR0Ocvyu4YWGr4YZTkXA04ywasM/YmkcEMgivT9qB2cC7
pnfnKZMBgqmC7OJNAdjY1OQQOjTP+Y9K3i0QV3924ufb3yyJdtppJ7/rqWb1qb6BzHpUgcUAR73A
Pb9hqiwu7vgtQEjP+BgWvOFLjy4bytoCzZAgasCyvdZSZVgh5fYTDdh5NtStmMQFpfLtHQgHeTUe
mbfQ7HcwFHxgTOxjc3qezvvSGLgHJ6RWl+0VoC3vi7anBqEb8YnLc8nMJMaZ2kQyHuknnzpi58HF
NrliwIh2xvuoMeF1esh4JoQpBW4Sb1bcnl87XRZ+20d68t5qkn23BoDCaJHrPg1dEdgYYMPNgsXV
/LKcVSLFF7ORNFhrMDutAr0ggscUzmnXjHwF5eTnkgcZlsBDzSOg/Xgk8mOF0aSCMGM4obMKbOQo
DTGiqM3gz0fALsGjqPzlqSH5An2bu9ttDZwulvT24/k7e5oWAp9ZGH3xtZR0syssPQotNA+Ve4mn
3VTUEe+ILxruGjt++0rkw7jwKsr6A5XPoWkxnz9HPBisva6OFcwKFMS5YHUwNdZomQPDKGdEh5hK
3+5b6G9h+pR3Xhhjp329LVUfmRVBagRTdd2IM664dcoP+MndX2zdr7KBvo4YUkpKvchNDWTYFbQ4
G3AYrSdy/5mYwPQmHWumxuDd/rA9e/aVbMFHBS8fC5SIVOCmqRRf3PHL4m3G79wFpi/BCV5v4A69
/wMQloDayts+SNszPJreMrVh6kViIZLrEusFBl56xyJwcV2Bdy3fbq/AJ1rL8hhoJV3d8HdZJt67
TIcTHq3m6s7MApWZMfOZLoBkaistgFf9OQSS0VlARsBKnDC/lSUZ6VSS1fdDtjkQYLd4AM+TXfhQ
KSyYgTHGQ8T2N0Lb9ZtmOVBLFv++NTRONIPYFKoZ/DitZoIhXgguEZfW+iPwlAikkocXhWGxDmJI
Fqgma33GeW5PE8V3zyGMr9A1QQZ9Q/kphWZO8XLpEh9jMPBlsEy1MHr55r+ccs0om42fFQYu+DDv
MltrofX8yxil2v02QIKUuqcgBCRlmSfujbYFKAv+vP4Yq1NHdDhm9XJOTydUA/naziqtlSjZ9494
nBipHJYdS1pPikgCWq21wbs5kZBv3nQr+EM6+lLdB0QW8IR/6CRu4oHnb4/Y6xMaGCX5Pqkw8GqD
8bRsNsj8F1urlVuryb40T24JBS4SM1sHWwco2Sj6irYVakL5lx0CAucaArSkm9V5A+BTKX/jMfbf
yctTS8D14dxompuHsQXq418/fltyeH0NLqfuJ9DAR8KfZYvz9bi3B5Nv9WBDIoBfgM6sUDfovHoa
MFGxpygyETqayWe1YqfH/WaPfPdGWbW/bGd4sc6eSpKuw1w2EYEgTBkeUhde0HUAab6rdYECJ6ja
1BbTMv1OBKtwN5eKjgK8IgpeJ3Q4gQt4OKBu7K0tR5PwfeNIyaDkIHu7WeQFy6ahjPuuzh4IlhAG
A1+o7b8xqcJue4N9anUJytFFXchc1mMckXSH+ylzGqno480sM0+T7GAMuGgSBJ0RW0UPJD/0b2aH
plBTBscvK4cB+bTbt69D/zOKTKWeEZsBLRHpjETMTVilEnSXuJBhcda48/zNzM1xG71IUmPWN4xC
q1cy+2D00bBzYt1OWZxO4xXSHQf/TxmUhl6/zH43BeqluSgkvklM2+AxtFYCkus982a1QOdR2ITH
I/3JVv4H0aARvye4OHrz0Tt/GpkQxLxIoKC9fW9ajIQwv4orJJgP9h+6P7vZ1KiAXoqkdyOXki1/
vgR2XhX63pkN9xB0ihgwXsWwz1BuJlcaJG7LEm+a9a0wA8H0Vycg07mmFKiqEgb/KVbrGrdchFsd
0hYoU+vhXySQiPTamQx6cwfUm9RZwhZVQLWvWLQ0/0mndB+ZPGsaRkLtHJrdh4DWa7Y5J96z9h0a
xeJjLyxwgWBLKKfDe2ERcZHBK+/wCG/4a1UE0xet/KGSVXg5SIZdEH7Is5QurfwGfUkBy/0BFgr5
STsnR6p3DZbfc/rSg2jIQCDGuiQQLy83joLbCD97AJKuSbs2oJ7eoS1AjKUz4oLb1XdU2N451p59
KwVXaZtPOhRXc8xPsih/QFSVkJkeASFgOJc+nJRSivqXneosvLeAXj7vW9FNqTQTO8e41hdOX5r2
m26rfFF3oeT8PqUOcEgPz3Jsuk/1FiNHnIfHuRm4uQbGvWfHn/oXaB8wESHLyX2E2VuEDALgv/qF
xv1got2BJTMyls0fcQzkzwkK9q9Tm0M4MhGDYZlNnVIUx1JzH8qsxyQcSj3Yb5k1pgQl2+cnPIQF
OT6elrWrg1Rd60r5s0vgqw2RlbH/gm1HqccBAzqj4MxPRxMJo+34rE69gkKkn09NDD5GZIsvTCBy
2L1xejcTqh0yJsH1tm2yZMyBIO6IvUIZn9DVnkAcd5cGaPvnoOwO1xL2UaRxNQrIxDpIrmpMJPur
hdzkgR4Z3BPAmTViXGi5McfILsRxzlOP9fxIQDWx95m/zf6z3hU7223qvtIpCDz7KuQ+j9DcE4jR
m42c72PrSLMgHXxYWfEoq+QBDkLLgBpC4Pjow3GRTJp4wC3ix2v1FMGff38IPVUcs5ybQ2RTyyhJ
5G289tHkMIskZ4+k+x/HGKbDKDJsvXsnJw0HbbKaNadiVTppnsw/ATa4wi9IYe32U+QFnxY1CwL6
r0ZpOsDFfD5NcrB3Yk5y9rQ34dNvYVUpP7/Jm6oWd2wO8J96mgfVVofbI8cLAu0G/hGbA3UZNFQk
3rVaClCpxMeT9rxJLGGmUmiXkjubnJwBEZWKt1qWG0s6kGl4pD2we9Rc8NeMEqiy+G9WfTVJbUdu
/mswYlajCWaoPvUhAqevEifND8O/IE4yGNkkCgZgWk71BEWFMbzXrEQP0Y8oifDdvJ2LL6f9kuOq
lHr/FghxbQL7sgAPzyanrY5yIt6KB/v/hSdJCod9Y9WCJW3gSBoN/vTv+3AlnDHyqfrrp7FO/MaL
riKvAk6tIhEvAuu2yXOPdwtFb1QeUui7K+EAXz3uUmJHEGamctJS5MiMsdC7IXcD5EJa15txkO25
K7lJIOXKOdabySIlAd8cyk8AMAygJ2CGvZsUWHyOq6N23eGGjAHjSt5JLYiq2hTkqvQXqvixBiQo
+49ZVBuiNLhyV0dHwYoyizx02f1GPQIAxwZC40e5SOH3srsRoIYvhD9Z3RYMGeru8ydmA79TMa4w
lYc/azXovaliMCmlGz0zI6TOgTGiGAqQQLCp1eaa743rAuTG5lgIdRw8P8Z/9D9jg8s9VAiR8knx
54Fgkt8+jYFKZbFvqbv/tWe2BhfVxSfVK+g0JeOGzUisIOL6a3I4ryxrzPK5+bf+7gya2uAPL2Wq
o+N4iifg6Tv3KL+0YlT+C0swIyJ44c2Ryx3cCwsiDM+5b5DTpg0dUd0m5PK08NDADQHKfx3MUqRe
an7KKglkXa20rV3IuAA/hwZGdC0JCVnloOM4bxerFXgn8X8ive5m0dWNOrauIdEO1eL6157oFfav
rDabk8MPbqFeAIjVxuCx59/+WMrNYpsPmMeevbYzI0lkolQuPoRba9ExlBYTwT+GDjUfkT9ihgSe
dSa6MjUBDnkSHMZLMuXJ50IP8dsmlyt6H7Cx6RiyDDZCaVWtNyr5ox0upUT+HCOWGGBjaVrdhkzn
kqi0hacQ6KtNXP5Tmtpjm3NjM3/ZdQHD7MFmS+Ag4wqWDY/rZfR3VN5/SBohksJBFc3Wa5B57wtR
ZK/GxG39xb7YHXIoc9xo01h70danXc5Vdp3lBDU9gozJNfIuL5i4ELqtbDskSK+ruJxN8GvBdSdn
34Gndqd6jWPiBppbz07EfL77LwkkqqZFwMiRNu2L1StjFlJPnJN4XSh+g3ufsql7ZEBns7n+fjWG
vxvpIZTzo1/wzIVq/Do99/wCV1FAmAxvRG3yDckmHhEjpS5gScjHqUwzbi64n/VPNJr0DgR2PpPS
xc576lP8ropDYxAqb1M4TrcNBUuLxOekBAkHvceiZFW8U1REZlkbZekAH9TbbAblTCEGOAxq/VQe
LRkJwOcP8xJaI97e4k6WMX6mTbn926DCVnPQ3xKATGcLohlOrVTxPBx4QsZmK91QCnF999+JNSjy
0gHmACy/uFmVubdzA2UzvLr2hjxeZDVAwb9RKu/l1CX0Qbyx/kMAldiVXYNzx4pmvSfrs7RaqsLg
Mp5d1R601cCx7OvzDI1ek73Z5BAzNEGjum3WpfS0chNF287I1si2EOCr5ss39vAlA8VMTZv0M3Hw
BNUkboyLxMILejtG4NmRuNUMfuy+yWyfrdwGs8Pmk6zIcT/OobynVXfdbL7jYE7BJCe3ZDQ5/7nu
4Q2Ut3IYut786LGCk8T1bKN1JU/+Ed6X+O2zNfqK5HsA6+uuaduplOxMNKgIDRq9ei1cbBb2BEcn
RAlMXOOUVJDtyJbNET/WA3nQdHJaURNvtqZpTFsC/v55YwqISIrY1TlFvC1mYaR5w1yMeN+3hVGu
OdOWY5U4l2l83w2CcsHOhpTUeXOe+uC0vSvymIOsY566vXqyOwbPawl0bJOZ8tVN5buUMsJTmol2
mxJ1o1ZVp1pdCeWaLsPTkLcD/z5ZRGNL+DV4ilc2MbCqTIyoXPfNaQZOK1BvnaXvY/Vpck7mAk9r
KAAqJDSkQHAaPPV3fEd55xLdyQUI8AnhRSrMDNcjpbI1EK71cizAu2QYmTfjPsESMIDcKsQ7isqt
uhoSnUoDPLBJA9mbWSgNZPM/JYGsrS4K5MM0D1AEee7BHCQzkRwnijv5LHMpWlUp5SuLHOjjDPne
J1WP2eLMWUu1WMvq+P7cUEPGhvKXn1oIVPCwGu0o8lb7lV7V6HqIp4wJ78fdMgod+4Uzd+TMqtiJ
1lXw/dMWq7AB3YCnJplNf4X6joToRqpWAXnp51T4b+WBlujapgCAJfwAitSRrLg02Vq6/yXF4wCk
HN0YB6vCmC4gLDpzMIMX4/f5qU70FLq8DLZ1D1uBOLtcfbFPJjC8AMqoLV3TntPI81eqkiU1surW
tDQP7RfbD/55IYZn3o24YyoxRE5VgGjwSX6x8rCWOfH8bciPKvj+95y2iRk694NwAEdlVcYDMLvY
XjPV8oLQUxG+3c5dbnbW/zXoLTGDyF+zhz7VdM3hAnQ7JMt//rLIo/I820x8YkplNcHVpvFRZMVJ
uTaZVj+6Ag7FwjenQ2qIdAZOoq49lMYxXcoamBUf/Brm1s5XEqjcPQH4Z7rHqygB4ESnSn2zx9AA
4jOtAXzz4KUAWd53fDNe+GDM+mbRsyP8RukrqofMq7p875zb/ImL/CGm5ZvH6rSGqrvc6ozrLr6X
a0NdpI+WAy0AriAWc1U/MqHIDPlWmjEYLyl421fmBTDNDy3/doRXObV4K2Ql2LLEy5pKLngbHmxc
yx2lTfgYy/96WLQbikoN+TkcS0zbRmzUA8KjbOMyYj2RQQuUt9OT4V8HWn8JQqvfG8YtkDMJwfj4
4MC62CYEizB0o1yuEe6MIQLnBOQR3jYmkIHkR7Xf2NGsX2/FcDcHLhyXPHD9vuvfU45xecizxMeM
fB+DGA3g4QGsez9xgwyDP5KXrXc7JDd5T5/RlhfQaG6AV3aNV6lbPx8t2fbzxLc22Xsf3mop3ejc
NbsUYP4qM1ecRuX5O+OgL24NPQbtovecBhrftcD0Pt7iD1z6vU+Y0hdUtWykHdNErBoJ81Fyxdfk
lOvwuWfqtpoee1iHB6g4p0+VK1bI1T616qcs3AEhokCnv5PpL6s+rKjihFSyyXQaI1cNZ2+RL2A/
cvVyQrAm8nqySC2XetP6w8gfdZVDRDhIgYps6e5kmW41L0YLTObxCG+eNdbWLjIv3aZm91yQeQWP
Fasy8uhOAP/s7r5BXpgKRcXFOgzqUhGV1Imvk7rWV6fo5FOQoxSpMQZPFAU4lx1qMeSaNuvomPR1
4Q7cPsNbu1/Q1e5dCO7WAOOSqc5P6BaWjoHQmdhzjbvjAUks2QZkLCXxeTwLrpj1nNFElWesJ3Lu
mHhVM6D4AGtf2NnHwFBW0sUDtiRGM7KZ6HBqNaYifYCkwf4NDeNDSKShIAuVuGB+6i1MsFspT2pJ
wLpI0AZivMGbqqxLnE+C93FmphIrPyetL2CIw83r0h17UR0/0PzCxKAdMOol22expP9ifqkTr/hj
xzUK4Bge3qI2sZEuwlQkIWoh6JA4JnlDKiXxVHsuJhkyN3iPrXra0VKb4fEz0Tw/1glNbVST5QJC
MTesIbWugD0t7WQXRaR3/8Cx/vo2XCG2N5x7skD9JWofVHliepK4bWUyip2LRNrsnNpDn7fupMYj
7o8eR3o26oGaAOzk4IY/OkPmt/hx6XfaXHX0S8FwSBrLqN3DS4Nl8Gk9ThEquHcBsnPK7LXsyM0m
OwVvJzNCRoVA1+cm3yyiydJ+dudw2WOciQWqxvHeYNud0rXF5Alz1VwxmoBRQnILbLRcmxs4WC0o
k1xBuz0ua/q17wgpVjf/W+hSNAQQKuPTQE3dLanBSYUgJFibhiDRlscOgSllYiArujGuAuYw+564
TDeKi8sBzlXpHMwPSs0RcHJPcWA7Mmr0aGQXTGaAyVOOOKMMYGU2JzXP9w2pZ7B+IcdG8HK/Vv9V
agRAhYrSLsyvlIveqP0XWl0BjotZ3ntf/su+c/dRZmtBhrykwxv0KFoQH+ABVMiEOfiMJiH8Qzgd
6zaiI+m911ixvCPu65peRd8eXT0WP4K7lVYr9iaHiXE+AKgnqRggAqkhM5Dk/nrjycHlqnwT6CWk
Ji1S01eyjrO+1+xe42T/F4564oYDYdzUfxWhIRgWqQkBaS5Mi4UzpfeBqxvF2pF5m6LNlsqPmS19
5+cErSEPcLyCH979meJP3Phqz04MWapZCKywfJI5MwsxfGL8MoS+BhxnaPnsWdxmHfwUvceE5bvi
Xxzs3SE/bXHZkdPXXy4VSz3imurZUGcg5bcgOOLq+rgl4aTjyrAZYMWTkGQkEYK+cSk8drfO6RrE
oTK+Ftnj3YWPv37IHy12ppwbYxHieirFCC2e3KbpSn1D5Sz6sg/GSAv1ubakpLSjWhGYEUjGjBWO
sWBdA4s/FL1F1cHY+bsHhVYCr5TZfnjrw3Wl5XoWXDEUOgEjOT4WMnGR5pQB6k15wsGWUEi481eZ
Lw3fdwfZvCmsYysJep6JWfsOO8PSLXuQCGytiHDQN0o26UmA2WP3qYgnj+Y1BGtHYk6wzKf7DAMD
p4agrYTQL/HXShoQ/BIvzCiti3JKuuR2MGDl8VSCAP/sNqoKAHAs6A6yMqoA/qJulshtWq84idq/
DZqXLOIDGOToMi77OQd3igTLsqY4vKCQ97Gw5L5txvreV/4+YGCODIO+5h/tfb2IuWZHbCNIXtmE
URvZKR/hKeaNu0mkuSNUpjeDPdTYzwc6AHEDn456jjR3GrrdP56Uc9yR2apcsQpu8yuqZj0vmMMO
w8bPBuYhWwmOieM/qn0S+c/Tt8c9Ants9VsU4rGEwlk5tEU9BdvpaLB8OuCO348jRCTq0sclG19j
H0T33VEDT1vIiHF4YW3LdNuFIbRzPlbFMRv8h4OaYC9Dlk4uZvh2madCJVupvuH1OgxiLYE4Qp5P
QT4jtM5gmCDOtuDnmX5DJk8UDCsEF1neT4D7d1Ya3iIUqSC3MsB6m3ENKbv7ZzYEoMZlTEV2DQDr
JWW1q4zmXvAoTtouy/jHckxcKiizRK/Ut7K4qcRF5G4OBu/omlk/GfBFVeI0szDczdnASJ//ds38
kJJYGmmIlVm27ICi9dnHJgllsB2UNJYZGnZ3XWCzlrdvIABTWCvuE1x6uO6G7QN6yD2WJgJkYTPf
p0Ms2e3fEICCmPpIgKqFOEY6cYhCv2j0/3AWla/Z9y3qFxNpBIxHxNDsswC5D3AinovNBFBvXGAZ
B2QKEBaRc7Ros2E/RehkZ255sRWI2O6ny5Hx2KzSvDHZXXnQqmCQKs4w/Mi5G/jujbLy6aDIcAUA
vkJEK138dozl03pU0JCmaVpVyO645pvbjEhUtctIYeFZeorxDH+BLR1Y0IR9aReV9g8tnRrw+Ivl
oZg9x7RDSL5oL6BbEkdfOST+odrFo7hQ4DjclgrAPDCgonNflWOA0hXrk1ZmNwObqY1WI30T0tUD
9CiEmPZEPTIcPXx9PUhr2XCXBWOL0/9NR5eobbzPuOt5s1RKA+x1vR0w2nDpxUamnTgLWm6ZZfh9
5t0dcSePi0IwzG9q7xwt382IjzL9yljORlSMwo7DKVDPz+dgZi84Jm7yNYlq7tlSfcodxFnXGNxj
/oE9ST2TaJNyCtnndjcR1Fy3ecr6RGS5WkAWFGBuDfq6CQpJfqM+82diQQJw81o1Kg6vLS6DcWaO
6DKrvkxoegiLDY5DKp4+XRtibIhVxfaG40l967MN7Db95OAAKuIGl+DlN3ZMHFANZVZE7fknK6Qz
UprF8cq3BSGI/GbeVUC0ejyZ9K4zHfV4RnXz8TFatPICv+dtcXEDMmHBqXzAtc6T+8La63k+U1fr
d2NzDMcoHc2YDJe313NtO4UHD1mW0aOL4AWs1z3qontadIp6K8KFoFQcgYDHSayRg4k8xxgd/EDC
bEnRyY4P0j978m7sUtfkjV1djS58eCcl5TPYh+VOVXG44NH37XOrTw5OnUZvhhHhugSiydJn1vwO
SqETJlVeZsQ8rBQJRp2YUj0CCh/Kx48J1uwyMbKdn1HJVadCKP9PBAz+38hx2UCjtESvBiXcH/pA
4zX36hwlL+o5jgiHIxy8Y2Dc69C4/DPq931o4dYiHk51iK3RIZgFQamUmZ1+IJm3rQY63CH0x1sB
zbyqtn+nlifqCvoEynTDQ0LgiHgb29EifmdizAmg37hR1hXe89wFnYdnE5VT5DdHgTxkGbTXNStW
hogbP4HuL8WnJ1mBITAIbPPnrl4g5SfYyUPhtBO8BN24V/eBft/vD75mBQwLUVIac+50dMR/2Knh
5ogJCgW0WBAOZzQS/VU+7IReluFrS1GovFJsgvepz3FSVyqM1Urss70g7F21dZWKcK6LhR+PbEAF
+K8k89UV3zoJfP3KLM8K3zmDlX1lbVusnOPBBNTn7beN7a0JStAGY5hhcOjfMYJwbWVA3XsK1s1M
UcKjFfbh1Ehic/6X/EcP+IXK4NxGDAn9/tG1jTKoHXLazqDmcYUbkOBKZQxpSRqjkD2FxFChTuT5
KSr4iN2cm4V6tSVzQUp5YCjWc5tfdcX/PLY4HuR8xgGWGiLZ3xzd46XZLlbRhTloQHsrc8yXtVYe
vD3irDcvCigDdMypGK7Iitjpik7IIkRkSym1ug/8Yw19+JrczBywyMM5+4ZAUcQHvuJ/Oeh5eL4F
4qRsNKTjJmAuLMLvKH5enQ4Hkz5ol826NV9aBV8rKeUlnaX+u0+k3ieXLubz3cxV7wucUBW5G91p
g77+9Xy+Cgv0sylLh/SN9XokU75qEyaHdBev7RwdS5AXhHeG6IAR/2tTTBgD/Th9t5zdM7V3BoOP
RqnMt8YylfkpL3+VvZmoxBH1WnuOabtElJ4yb42E24slB9DGYzC0MmSHQ/Gs5aheVXzygyTBWrwj
8c0xPvSHmHECfiQNVIfNTXrOC1JjNJHMEAZSXXZ9XdI+A0ieCPR/B8aCWpT512TC052yBrJz5jQK
n75KRtFJhhH0wkNh/bs0lPgM7VJgSYhiqqwiFMe25wEwMMiPWeVLzS0pbEraYDRIcyP+e/imkA28
zp4gDKh+OWwHJb1LRqYopaoDLa8Vq7dpa3Wxj9omRbMhw2zstd6h6o9dGkDK++v5c/97MKHWnsmT
0EqO1Vf4tibZw2NPNrm12gEuZoy/qyg9YMWMnIuqMBs0tUDDmoaWrB4JmbRIqU40ojDv0QvmQuaf
DuHNUyULJzWEmp5t1PXqR4YEXnSl4D4IA6WUxZhA6v3lacFOocDFWvkNQWh2DKzv+e3CG9A18pCj
qwJ3/qieHXg7ViBQk/ZvJCokmvtcRk3CkJoAtca5Q+IDZk/5iIJHoHwdSSa6zEhqpN0YMdQTq8Uf
bwTmolmxoTWjl42Vm0wUTB4orOobcNaHND0XF/DZCFDhHsyXW3RQZfhwk9VOvbCjRymdxUmpBcE+
mob7GsrBLtxgr1ug8i+DcRPLLkDtyFrAT+XGq2kA1O5ctfFlBdqOCFikLlDl071ck19L+ZCFbMqk
IbdY1YVrzQDJ0ponlJGxGHlDJ67XbCTIgARvn81VBBabMZPgkWQqoPJT34Rdw0j+1rIjCqMJ6L/Z
qGhX9XvIq2TkZ3Mayaol2y16Ryy+EhCoavp/JilMEhROg8bakcRCBwBpZQby2+kQ6Q/YRkWXhyRk
5KhG+zuNQoQh74z8AQobghbi5YwgBCSVvVpCekWZtoA/5+6AuhFXXu5U7VNrAIeFefT/Qd0QTUKI
6bDsNV8Sxs2tve2X7q61V3NO7TUaudoBW+Q997ldVpqwM4+dVgz3lWZUktJrecWdi7ReCsRJXn3p
nevRWbaUxWWVL9iX+FpEpir68ueoivuL4pyZARp7/bMXo5wjPd9uB24qwoUPFHds6wHGZt53JZYB
h0wNm/yvNTIw2tBMYQEx1BI/khZaoxb9U85NcKzG6Fe/SKfLr6mIrHfW5UsFrBogX614oCY2lSqA
wlDLL+BhPfbE2bDf0oR12ySNojU0W8+x/p0crGZRGwFUQzlV5BXD1TDpIb/hpfWDIrXJ5kBDuCaw
DuxsDrikOveS3UBPIjVbM9fDEmTmaDZJGjFHhICIYtK8qI6PAw7srnt0NHwSByycJfBmeKT0mzeJ
7PIiEeqEi8L1NFfJy0AenQfhPD0iV4D6G44SdieOEbQs6qq4IlOTppBmBUiPjE6Jo83QYTBqKZ5t
W1WjG8oNRB6Nhip0S5Ispvt2tCLIWkezwlZePa2yCgADe0wQ9YX3ZRHZSZfGb7zcM23EaCTeK/iQ
6TWaaFTXRivsRq9xY8+zAeMrzgj6dQo3x4PamJy/D8jnc34nCevUUfUAoWQxQrcHejsAxuBTjw7p
qjAk31eJGMhW6rQsmKsxYmfGWMIf5UEpnvM8XF1KbOOYhHaJvbdM8xkQCFUeSta9hBQEUYck6pwg
mSmpuGyYrxn2lxsJxI4Jy4+O5eTF2zHH7AazdiDAX3NqiK+gnRXxAgWHyGDIXLsfcSLuMyrZxrIS
7fVjM2Qofq/ANKeIyQmvVM5u58+d04l3capJ7t6DNH8H3ht9GY+JbnCiauSlRdBi/8vtsDOrsTN5
uUJCSjAZ+aTamoHjvWhV89TeDazvNPqIRQsYiwZ7+NppsIVDopTmadhSkTPNoe5CT4XnmIh6KWgD
2En7QxbBvgoSc/ofxE6bkNkSZk5Rl0scTbqkjrISqRwNGjrhGGpzeNwU2/NY/CRAwP7WZAaKQ6ne
gcnqPcz6z5YWz0I0kWThOapcomyvYTRe0swWqoeNojwuyLL6zUKLqzE7zn18CfcU1Q70AZ7+EJ2o
EimqKLOKAIfNh/85bJ+WGuY1FmznOF3vZN82ZAEFRCs2jKeFTdh7PwNnVWfIBC5VvtIdzKFl0mLG
QKyd5FmhHIVovqQnB3aeIriw5sWV9ON9W3LyrLozx4NJoyoJN8BzErrA6P8LghEPwvgfF/8N7NiM
kiQnwoBr9zlq/lL/JLAvFyVrUGimwsblFnjCcos/ZetqF3vGVe3mu8Vsmt6C9DXMaWfY3j15AeDo
vzCnIMYm6jycxt+ZHkgvKkCumwNNgF8+8FlzepdRWdzUt3QCKh6p+cyoyVliblPVDsQ4+m/AZBrf
0Wa+7PxYwg6qN+k01r1fBZ/0Php7Q91YQfcMDvnhIG8JS3yzLF5Zl6tDrzQP1jl8jXKiXYXfJuOO
wnQ+NNa3OFIRrhwKpgd+NiY8CKKQNlMTcMI6GxMb06II56aebjx2Y/4Pz2S96MvgWD5vZIyHJ4qy
Zy15RNZ8IC/lCkM5Uxq7UdTxgg7KRsrfuZYJnWJh4RRpyfTwYJz71+wf92Nve1NqcRvZpGXDRxGF
dR+35k7Xes+eoiUexSfT5j0LgTUIclQYSTF7YD2o9AwtdrUqB4Df0XChCUALvVtnKeSYeHOrCfS9
B1WzigkaUyIm8YL8l2PE7g8ZX3VhwWNC/xPd3hgmgvVKml9Hzs0hkwZhdk2l9lW2h9OkstegFPhr
pYeZhM+llLqnC1UyzPyslFKF8bT18X/rDhkU1NbnUnrMV4X1bJ8BeAE0FE24Y+JFJQutnwCOqDt8
NsSZVR+MC1sIWFJat7pzRUa0IiUZ0KiF19FPkIKNz/dkuJblb9vYzApY4AvndDCMmCVzkXd0ocB8
oX3YIJJtbXA8TDyWXjchzS9Q2Pxpq/s+jJafFHJ9hbUGwNmO/ErP7K2PpJRWifhamPu7bwr3Lbck
bNghiew+4aVWPySaSUTbRIXXr8sdtrNixGhI1TBWFKOaP1EANFwRHEvMij3l0hRXUm1SLS6f/3Ih
IZcmkmSEYC+aQ77+sU1CQ9nAWfd/+PfCDXwSMkLdaNyMyFW2poXRa2BQ1zNfHkNKw2CqmYAnVpHY
zyLJ0Z7f/rakwVbk/a67dcnr36QBSJxU/XQ7z/Jn2Do/CSs6VRj8qpn/pZpm5szmnQiMdegpT8rc
0qs496kHgEc4uGshXYiYud4RKdz5CCPLKIm4oNenIfktdp5jcdb4j1Won4ix6tdUN2ytrJX6Adtj
oQLS9DuqcbOE06uxyZxnbFChMrfmZbTxH4i1mmimIqk15eGG7oitakPNaYdnMRJy1aEys61MtvRR
KNy7xu8u8ud6pEgt+90CvhBmCYnAa36G9p7j5PU+zBOqUqYS9O4xbdvfFhQiyKMtj+gO149SnIqR
mvFgdeWG44Z7aVqfmfE/aSXVx4oEHtL7XnYUDWIuzePU33+axbZ5Ed8izu5pavyU4qR/bF70x/EQ
qXZfJw8qOeHGAXU1447vStkAMf4o8wfcFricBW6+eiWnppgczFpCab6q+Z3+hyJlBZjXphup1Rvx
z6TLSTOEnyFhTWA7PeONU52ZOd+Ipim8U9QuVbcMONIviV5vMDZ8+tBYwp+9b3YeE9+eCW5rR/vc
DYpZ87lICFUCbAkuGC7GQJyKysxKfH9jMjOqavnr1dHC+n0sOPx348Qiniv/QdQ9O/hjQ4meBWIp
saIB5rTlSF+yDV4g99qvPmj3KD6am2nBT+xOCrs/22S+3lg5JTCPahDSp2x88VwxY4nMwwN6+npv
PotPHk8DChsgYtelxTfjHYVvQL90/lvthGtF/Nz7H2nLrjgf0456pxhsCjYcllTlQG4NiCeLUTsU
5R3yQkEVmh2Gr1YwnQC6of/SHRnXb8CAi4hskzHKqSX5fTm8w0xDcv3yJqCiq8slnujaCT4xT21T
YdpRvD1MHJ8JnpZi1aNhVthel+w+wSXwl/TMM/03M5nN0LQzGJMc+SQKDQ/wCK58t/CRXGkpGDvu
49BGHl0RAKaw9xbIzISxQ6eaaPBsP8JcnygxW2uv889a49Vhyo6d+jdURVB+Ge2a0KGw/N/KAZAI
nxqgxz5lVUYlN/tPP3czuMen9cjTPwWsm3YVkiDXMjGTMBEjIO8eUkn1FfBvfpHwIUaTUb3K6eCu
a3El4kqK22ApAoBWlvDH7w4e/9oFdCwmTxxzVuOAvGSNQUDZD5d12AJULyEeEKyUmAhiGO691Gaw
6VCQ1FOjYTN5LG0DwdYIcaA82WyqhKi8NngUBzZQDO+AL0usVgxVoprg4eFHVSuW/tp1uvfG3h9I
Laho+3LadRiZpHw4cLy39tYgP39Do2ZpSg6az2ffPsq3RQ3GXMxa9BxnIFeVXj6mMoXECzpcAKFR
GSsh+UWqUYn4gEKCX0HqahPYeOzbPjeGPYkiszO8VUygByYrWAErQoTS6cfFiR16egpZ0nHHxeAz
w7WpBZcHXCcL4zmM6pUXNZA75Slz67IGNB4dpFmStdP//jzKwa3Rqvj489yYlRANOdjKpPJzgDJo
mNyqA1d3SDbDeuaIA8XXtifv2rutKuDUJKN+JxjBmh3AfUk3Ac5X7daKOegBnopX3uJywYbdyQ+x
QHJwWtltX6S2IVH5ydNKBWOlsn86drL/DQZj4kQN83pgVaYg4IkIqr9xUYhTpBSTu/ARZrm7nAWt
wM+Ptl+0CNNDRUIqY/FiM5d1mdIeoBrqaV/1+dsr7M0YjxJqCYZRvAEUHU/3JU2Rn1dIzBLvsvh4
xAJz5Vr1DvrmCJ8io1iyOe98wOJ6L4pqDSnfT03RsmL/N+jkisXKpVTzHrfpb2P/eHtOv0iONkZl
JuVVGK4T4nCeOmgxzFqtxJGR4G7HepVwMas8FIQY11O/ENYOU/bHi9xvUhSrKQx1xHvI6KnW0k8f
GsoebTgC6iZVeY2TX/KcG08LmwfrzF9pmzp5U1nEctuslq7bj4P3BqJSPHo4UuIkwAmQiI8LUEgk
HTKUkLP6awytRoVt4iLJ8J6wJwuo8wTx4S5v1XaGNDp3MSn2sKubsr+t+XM8/QSwrQM+zMbW+56F
VrwIymSj2Zuxn1sHDid3bsr5koVlpaodWT1CgJzAB7mZV5Cc9sj9fzmoRD88KOeg1QqnB2J1ugdc
t02+B/+7BDpWsDojr2Tb21OMVJpYeGlj2d6jMvIIgG1dBOo5yvNWmPiwvqPd2bnA295+ASiOak7/
01UtQwe25/QZW+m0hACZHzpf+aZfzArUbpF9Q5oj3LtlmfyOZxlDA5hM49uBVdmReHwdPxtEu9VV
1FclOx/oKQQdS8FaVCwUQKGhT7FtPXdawBkuZW6bD1Jhros4NW8oRUab/xCuOOee5d7G6XlQiupn
numfXmZcGPR+HcK62ZxK5wMTwnzcMuM3aEV9kvNR9r4VEFWCTxOhclq5CVnQTcvAOpkYK7I6d51T
H7DnHAE8AR0ca1EBhGoXJqvfV67O2LrP//q50SAKLGcI18d9+XLvkVRWVY6KIhcC6rwuK5dJkZkn
gUoH+tdKVH78FqDxbbijVelm8ns8ELawS1dOekOczmdI5jFt21Cm/UShRM/49taZ8nDI8oF4G9bc
r1MTYcZsZnXFruIfY64N4dlpT52qL8F16bN4kOMUhIoIGRdYAYxhxYJ4c31lrOZpdwPyPOLt4YRN
9QiU8o8qskAOOk+XA1PCJ8RaSoY1AHSK/x8eE6ffkoW/YqM72qKoHBU6D7zJZQRwRqNZ1JMb4tQJ
IGhYhbpxHubbNcQ2UccofpzUSsq4xTwkcIquWQMjIuCcuKtTrwuspGVEUol4FULKsNtMD5rV/zOl
3q6jnRnbZFdfmXLROrRS3DeyTyneNn9xpu+SAPeQdYOpx3HQDVmZhRBlGoIL5AuczlHb4YzI4xWW
oqHVaE4Sffiv3T3M3Ja03H3neeEgUjP17PcOmbLhtf/qh+c/SyXPh8+UsfI8ND+9P7Pwx9orOlbH
qJV8s1IxKUl2jdLASUHMhS/OPDBaWN9clIWqGZwNNcbiZrWNyEm05dXGETx3EAWr3WslRkHz+T1N
UYHde4mFOEJPoB7AHbMiBpc+KrLIYuqCsicSAJ3XmiZZfQvDaBrUk+RVyuuG98C84L7p/Ncszlz4
4okTYkjR26QB+Jp81ppKpCqgKLjKASbV/1VLmNGHgC9vuQIYzrsKAj+Q+LpaNK3Jsts+RWBXO7Wo
Kca9pOtWtlZztY46FZqqqoY+u9LXOjRKMVWav9ZI1tYKWkiP2u/bk6TjA9oaO/MvNQx7OzAwRlFG
kkFaMV4h4b/93q/sMqIVH9QjcS006dN/RjNqxoOPp3g5TS02LS632qOs+/OOvcDMfyfFCvB9NAmG
91OCBBTxo1lYbik4Gf5/K0kqWFHy2XTEijZLLytS6yWLXLJmc5Y17Ew8CcTildu98AVCsjYUVS7H
cgMV1djR8hManCFtDnxdjP8/yzP3jvOGPwGStA39jHThq7Klc67iZnI9yPQQxzmK9IP7vOhP5bRO
Stfb81DfZZu7gT+2b3bbSMPwu5bn4SBSZvNfwO8rSCeY9frPr9/4VY+tE1f/q36sKnPLG5zZIfYy
YGdD6HVO9hlYSnzBO0vf7qci3Einjbur28B7xReJDnUxiSIH2pCOM+eU55crZA9+NsXAZjCTKNrB
m5pU1RD4jVg2cj4Y3Rca+Ll2L9tFS7j0b1HmPuDoHh5vKVfETiBCohWNsbsUlvF5FbvOCU8baxqV
ODyGyPBwKGVZCSsR2vin+IB91fzEkSziO1h/dI4ACEzixSTQdPZFOIVDi7TmiQBMFvfGUPASAMp0
WNiZTPOLqDZZ+Cg4qxJ91nDwc7Aog7iqY72OQKFQ7zglwnO0ysmTj4PGOwlS3SR6kNY+/+wW60eB
UmCDjhLpRffnB6Doy8cJtsdYB0VfkPNLCGdetptcPUWfUdAsb+O23yrV5hkSXF8ybp5TKoYFRXGV
w50dCkGxrJU4xR8CSPXto0ib0/y2RJDYMN4EpuCwzSCxVR8bW4G1hxsbBrYreCSJXAetfAA/LuzX
A8H1PczMf8sWPTVwqhdtH9myJjPKEMYQdJTMtFKJ7HdnoWz45vcXEyXuWc/fMPs6CCVo7ph2se6l
GvR7E3o8i0nJTrYunJpG8Zd12NPmnbJPhzyGb+EKmV+aNmFeIYZCKburzoI1mrUR8qkyowuzzMUr
XInE+4hSXp0FfgOF1f8UruJi59KQWWJgH1/gonnLze3mD9s1+UInwVp6aGbPrOGAJF0xONhGVi7n
h+JBE7aTBQGe9BmobobCVjJKeHJ5Fi84V+hik8VN4uYIHrB/1OZNbXgms++GzioF/jmEOquvufL5
ymdzg/6dQs5Zo+9vE8VugC2XzjU17foH30wznq9+dvR1Qt5dUzRBzs532n2szdh9g/KJRFalcYFa
HzZrtK55MMP+sfUwwNjddTHhzC0DiRTzOoPvQDEkHPb90eVRgE7pGImkxOOtt/fV2q84CKTmUtbx
q7C9ACyTGJs+OFGmF97nd/htGa2tRvas3dPmzT+Q/iJxdkNuYNkSzbZFQYLDG6MqQ+EFwej8ugqR
CsLwwCPXKXF/fGqUYBXsKyDt9zI6HRkkvnpnKm1FI1YJ58xjTbHacBEZk93TloZtETfo0a2bHTu9
5XRZDzw7BXTqgx1Z6dZQwa10oOoDu7zMET4VXf7VukfV8OlBNvnOISagUdL2/eqzqnrxtqOfZws/
od7t2ey+9RDydwnPBK6/KEwTk+OHfBRGxkS6z9T1YMuXiiqYbYfI1fhycHYJQw6H7WYw0BDlGiFL
yojQDU2hmesi9UI25c+nDWp+o7TunqFczA2g0HrTkDTUuhqoDu81cSYqfLFqPnJxPEByY9S9nh2l
uHXtAoUbwM9HIssWYA+8+bmt30jK3IGK5v0axQAom7wANCXKUlskVACj1JLjQ370+Miu9CMctkn/
wCdt14NYzPLp0ctnotjyTRmqc0nkYknVn+3IufMHD4pMgzTUII+v1aZpA4jRWZ+Ftbkzt2IXTPqj
RNcoBJUv7V1sUkU9czfUiSP7zaRw9m/L28JQzpTxfDwt3oB1kDPw8Gi71jn6bd+VygsAOEzisnHy
Ya8ih6FUwaHnsm0MbNxCgXBr/S7fdjb4+g7xoGvIQEeVaC9NOzgvHv7tqKiSWgBOLX+5FweLktBu
L6FjkqziCf+eSqbMG3+fU5G5c2br5ZYNR6+GnUet1k+jZESGG0GwoQW1mppQOo/Ph6oz3ptCOR2h
u35V5AWc8XRiQR26B/D6gWlEbhvlepW11IgxerLX68uMx7KXRQCdiBMXYLKG5daum3oCCo+oTV77
t4kIhrRZ2G5ho4eo+QFcrpTNlcJpuRUQtYHibTYhTSDI2AgZqILUiFalsKh0/PiHP7TJEo84oVWx
Ts9bbYXiJn5KtCkDuLSFyDFiKRC5kKjuh6sv+CcvRk8hMwXBTYU+HZQqPzCGr8BbfRFg4ghpuifz
BUN2cddYhR87FSncIV0SXsCiMItjHZFJ03k1jkgh0b8nSlvAx1PoIoWR9AKnY1v5N0CHipNHjzeI
PMYAP4t89lZuirQaDAZZG4ePXZCmPv8gB3mixvHtmfPX9+jg6iKdaiWzYDHPCLryXiSOpr8sy0U6
vPpD60MobtntnsP1EcFxd2smird9LGL9LJJ1oV8N+loGe6koyCkqxi4+yykRDkslwV3ZQ0wfDEmq
+rQU10/SLcAP+G/rBc6iYRvJjo8HNw5bT7P2vD9JPR/Jpwy+nIEdQJIT8HyPljPAKvVFVMivTrFg
z3OsnynGs9NN4pehRadO663p2rtb9tZ84Du0b38ZbqNpA7uwNaFlLXLld1Z+FNVHlHNZE3NRgH65
ihTZDLoaUHE9JHiC2XKZHFGzd0Dfibzejl9ZG1rvMFTer+tzcSuN16/FN+Sg2lSQfNngFq41v5nY
byIdloXtmwZ+QlXQ02d6R6fBppqCqOu6pSw9+oIwv8OQW07oXNr1W+qS1KjguEwq/bLmU31HkyDD
OalHD8orTnKxBpI9rKt5DiyVNnqYP6JQL4AWETPhS76Z0MkFH+pj6uSlLY+wKz4mDg5xJpFeEilh
t7RzRBuhEuuxat1j/AMkBWg3zdSkwnOlRQMxfLcN5H1Q0LWGcZbFjEmLZw5ruc4AUJ3jyNPPTIz8
BrKB+Edj4+Cppj5NMuKi+S3+ANnT27e1Y8ECMq7W5QrGHpnsoGpcxCgNTHam94y/hxb8p2hZQPf7
Cit1OTC2tYe7H1yjPpbUXmk22qtNixjT3YGKablKVK7lCpH2x7nZZJZF/wGqDf7NyyqRlpNuWJqZ
ywj1MB2fa6B3CSmm9XeP8/8MFmCikR+NGFQcKzXDfJPxd2AiCGHaLz83C4uOsT8LuMgM68VJtMNP
QEkjFIe7XE3d6hG/JQXR04OnSBUmNDGZWdgFwlruk+pbmsm5oRiuhqPEscqieuKGxe+5MolfNz8u
a1vZ3+mpp9VcHpsh/LKamPAx4vLOHpRkRV/xYcYknp69J4/oU32vT/deYGD/TFBe0GzEWkU4xLfL
/iDbXwXNVfrS0uzqDjbBYH9XL9vAjtU8fqCmpVTxuktHYweecpflcGLGjRqcs2J/nxokfWFjnsfl
Mh9WZxucivDu1Da+v4p8mCjcRT07fZW5Qzt+O2kwrbLxK05EI++1tylPsaWjBWInUu1ZjEk6zCTR
prbtNItvl7CWUJ1sMnyh7ATpdcqt2jtvzV/6WX4cQX2mvvSXsdC5leoyQ1MDF/pWhbjveJOb9dsb
JZoly1nXY1SO3cCOHeULENJ7OWM1dMtz6UtjhVLwpdpP2zl+s4LCNROB6/f7epF1Q1jyc86JNoQw
6Q3JMhIkivhYh4pS6k3VBRO/Hrk04SZK9xvctFNlRmyPOf+TOC4ZLLFMxWFUvh4HRfJ0bEV1jGXv
WdpBDx1gL/reBFvt+aQSG6RqN9RYUCJIJd456YgTU2hxTZtts+tzLeBIlWuwjw2ATEEFFB6rxd6y
m5graJuMcjtyrmvYMUFZs0l6zuJaNm4V6mnmuZjLyOdXUxXrnqvTbag3zvTzbkifXhmX7qq6uMFO
8Oj9wbYPecf64bwkbrQ4A2Fr3breGfUWG2dALVd2Zh7wa5QWTG9BjVqHLWZTknb0hN8CzliY5zPW
fYHavUQ1/T9qU/1y+Umnk1N79Peqj6FqGBgsmvU008bukx++/0SAgzLiyxwHfwvI1uLzom0jJOm0
GGIlA1rR41O+MkoDAo8LKb1ODZINY/ZCO0Oz/4tvdyrt/Su/1WSEfPmchvDFrtxCePbO1ZOoBv7r
qi4td2zFOhHQk29TkJvIIZ1lgLFENOeDgmKurc5Pcfdtgdi/ecUgsG/rn9XIpkkoCQFy7UaFQFM6
0vp6zJNj5AKRNZDRUV3dGFLLNjImHu2ya0Xxex2y122mdD8sSiG7hyy9DtRaNOLAEoTm42lofILi
mA2lEZ+FSa3leIeWPz4KUeLu/GzSH9JqW2LHNGMEmchx0N1y1GY0qP2lqVsllvbLB+OCZlPGSQiX
zkObn1WPsN6uPgyOnp25iKtSGSI59pFCau6kj7cyM2pXqQSQppTL+bw0oDtmcFmMoMPOgYbONddG
0/4x+CQD1clXoSo+5S6egoVcVVIeaxTxoxf9Km5Mxenw73WoY9FX1dBXYM4wfLU5W0Sjn1+mXCj4
dSrWghYtCWjLZmvjkUIxSKw3y91KLw0mJrhF9Nbi+1sjUteqe0b8tiD6ngcDakuotTM8tJnxsoh/
E/V3Wy6457xTYvY/Z4EoRurte75njxute41w+z9jCQeNfFCjl+/aBGQUzG9jhc3iA2SuAMKz9eRU
+FELeTK5JVS5v4dt7LLV+GiObbmKCDT/yBcUettqZRN4VzOQNGxc2Bb6/fV8XSdA02MOSeo56gzX
1kO0vEcGFGecZbf+c/foH6kq4vgoWjgs8N9qWCGVof95TO8YkhvbpH3UMduEC18EkYELiK5TkGmB
AfZXdLm8XIJO8glDQy5T1VjnxibiqSuIZ1tuhTFXrqMoCHUuftiy72JDrVJhAZUka5XxvW1exFW9
GxP+dtp/suw/lD/y1YXRCMMi5dl4tQT9/sZzRj4Y7Yu864GZ9kLBL9Mk2IW1RDEToIoMZymWXncn
5yJzn8DcjCfFvkisW6oyLD7YZiT6ROgqbLj5SGGrrZ1sM4AUJXvgEj5DS3ysH2NWMoYm+x9cUCeb
GYsFtmXxoQJSsRPXzoR6ehNNcEQKTDGFMsRNiEup9ibyWMhyHpp59pWGlGUA6VclcTvH7hYtE1uL
9EdMeK7d4TkZk4SdwmZOmbGqvOXOqfOVtGZ66Rrs+ib4ilLpznMcrjkm55RRbwY+T8olMEsdxzrM
rsYO/P2VDQ3+8q5rKvACkP5EIEbcNOe9qwESUI9d+ozipOr6Zh71CMUXPMj6gXeZ+GCpqv6o2hlO
a96LpUhSVtF4vNq6xyuxRf2x6JCy4iAqCbUx2nroDZG3ueBFsH7OjEjec3N3BGol4VQJVCfExvzD
lTMRRUf8h2VlPYWW1Le6SiyYngQRTZycrbqR9LUYoqO+YEEE4Pz1AuSoj+XLIF7gKW+c/FNsxr8b
jTG+tFyurfLH75NfytL1HFU9PYMXXfPVUxEn2mJyZkjBWa+pho88iuvDo29OHWHjvk3liDqq3O42
FM3XhEJDULS5GHXXhMSB8hKZk9d2iPlhUkJutDHj0kaGfF6E1ffHBUTA6gLywzoFMSggBLDgIq5V
5Y5ijaCK0jb+Gn6EGx8bihVPPILnKCFhIgLjj6Yo/7EtJzJgE3DUonWZZ4vEdcv3i7MIxdkfNgak
tiy6cjGs6WmI4kYtIBDLNUqSU7zqGrKMXcgvsiJPc21EWtEFI1R5Yj9jYUVFVlwh4esFbQBJKdth
7LtvCSSOHpriSYDQO+aRBFU1S7XPsk5P1OlUQMchPDIjg7eXw8zO9z36twGzn8jkGrnFlfvzQesa
3+zqT0TAfqPdrA7Gx7eA746YYp0G7pAvcaXApQFfv0upJfyKqBqc4AtnuKXPToOV3ugax3F4YNT8
Z9JgCciXRV6OZ8PTtRkUjA31z3CjPjo+tsA8F4N44wYjAZnJfMPsdh+VbDKf/pzFEGyE7H/CkcLz
krhArSKDlAPfHX/5W8/9NggkkHLpyDIn42xDyF+I2DfRVACpFmieMXzrUnlaGqYOh3T853h5NhfN
aYLdmTj3g3YNSk0dBWSrjYUrbIL96v91aMiC3D5xVrtzfnCPWfB96zmFRD6gP4TcsPVRxKiwb1Pw
pv7ZGGBTkBMVdpC8WBBEvgEvGoexN0h++ZMs+pEgp9jXJPOiG6tGe3rtKkCcA6oDp/h+8Q2bgDio
A5lzSQLiXRFvlqeKBJ7nM1cpX3ZqkD4rrVHLcyAPF1TPvxJLKYeCvKY6KBlf7sF8EU58EvRZZ6bT
QRYM+G6LaasCXdukDJZ0u5Ga8F5avKLCA8uh5xgUaqZPv00qXAeGpFncEEuWKdR0QZm7dmsSuBVF
t+SP+bPeeGbrgoFp2/WrWbyiv3K758oUjxLuYGLPHoQuyaPFlKv2FoviZv5ULHeTOo7gaNnuLBMa
UoVMX/01n8xhEicVubVeS1aCChyfYW5N+0tDkNXkElMOon01jIhJrwMR9hWHtCYzi6g2uq/yF3nR
QvgIDHrEO6HaVqRYBr/aLJ3cDMHWFO2L9p8Zf0m+2D0w8qouiVVBHAR2lJ3A3gASXzbj52+8H1o2
8kt6/5QDNWGKXoEbZq9gM3Cvef3uPynyC43pAIpVvR3X4PHRpp5Nfw58c/Wye9C5T38g2cfgbBEi
RuUjZu6n9XWzpMhBXjx9YL7fuEBeLEW52HQN1W+Xwpj10u/6/lMbVPdb2fpZPMCNRJ7VoI8Pd6V5
8ACj7OEAvZI49TIlRylGMwnkY9sjauIvQFcpl0TkFnZ8QZAomSU8nFGzNQ/ShVQ9oC+4IUHjblSi
Xas0zT0Mg2d/e178jJc5pWM/fYdU460iIbZ9E1YIoPSahHV7DGVHieJCvdn+oM8T5XSFZkfKwb0c
jen7wBkR+MZ2p8NWK1beXbtQaWU6uYvLav1fR6SoUXoqKfvByXVjRx7PCsA2lVda3uMfvMzioR/P
TY1TzL1NKI13nNWlp809L6P2dmlNRREfICP2VzaE+Mc49wFqCHdxQGHmhpljw7HlgZfNrYdrTNQT
+lB9dG67M0cSSWDv1SzD0IPZosEIDfhzXZRmoswAJnDUa9e0eLCPoc7+5jiMWuvuiu0uTW0N5LKy
kodVuw7aRRZwsB4NPiau98/lipWsrmjSm2RzBQXQeTVUffYnm3Ej981043aAN2WEGwg0kSmPIxoo
o7vAAsb5BKNfkhTZd4WzJOgQ1vdZs6XjnvE0QZJOGXMFE++M+5oE7v/dtERjdJClAVZjI3UDG50V
S8lWFApIiVGVMfFvK+MhxxXIKprAv7JkGeFcoWEzhgn3iwQT8/iXctM2EYgy47nkuQNAYhODqDsi
W286ba1TDP3mScJE5ZmY7TtE8R2gCPgjqOZPjlSGRPnifmEVTnWx/Y19caS4t+75BUXMJEsnp9LM
whkWF6JiHHAzUTWtwE3VrhO+yuzAsaOMijdpe+sU+HFMA6QIFgW5nlAP5NJLfDkcVQ8WgtlSmuIN
9drRMvw9jM1s+NuPPdgYa0X/NATe8Y2eYljKWiCYfogDLTXMUVnCvhmdI/U8nDGqPH/WUtX5VjNt
zkVUDPjFKhnfGrFtCoXby3WDfb4xFza0K/8WGsGUqX/pkFDiiZI1AJDIIK6EwKqlWg8EOZHvd1cb
LHJ5uQMJGiU5c3MfR1qlvHakqzT8MJU7qldxMYCtMOgmpw4P6sK8sH+ruoWGOzjKkZZVA3r+r1aO
qKuLW2rbDTb3z5suF/iexFNuM36N1f4W1u7+t6yxizH6+26d+oSCBHf+MH7kxGcLkgemm6ooHRqQ
WqZBQWPU8mFPnbf7gdNXZdiz2p58h1uH3cVyiGDw96PbZNvbgGfLy9gnd+2lBJLlgjQSD7+z/tVx
2hdOSYoDoxWKXIZM+xjcpP1i1DPmVkqiIpT/ArjWCtmhEvqmo0Ozp5tUXpSdySXYMNXAvE7sxP0x
DP6AUxg1y1kh4NDHFevQxYMFdxgUYylKKHtFlJdGeaz3pFcGRhHPk80GljqJOxuZxA4glboJJjQf
cySLRhw7EzlJcbNKlrymRf1Tj54OqgBFrZwfAUxvJkbxYkk/JI2EjHhbiMmVsajBVBsabyMFq1tI
ol+rzwrXMXm9PbxcJaESN/49XRWqWWje3QGjOMOQkWe/HJZTg1oL0KivrQpLeTqkU24cDQpYTOXz
CSi5C17nnuzpLGvVnEDWvUkmPH8IPDa1mozGNUHcQSR0KpiVND7YXjr+XPJYjeVPVmjoiI+R6+8e
/UpzOl96Yf5AoteBgZ0dewRVrTBBzSqlfQ7dd5sk5mWjpi0v5W5Yd54GWfMOrPgwtAVnXtByQ9CU
roTw2fEZMKWnF4w79adqZp/2PCjEo/2dJmBadacYDJxy4VGg7qPOtm7qfCQ41TMzNo80lDHRZLQs
ImeGtHYt/Z2DHYbxzCQobcgf3fCtZcoGb41SuS38+bkKfgWgT6ZpGzYI/8D8ACtR/YlRErKHk6q5
BVGAsY/O9rx705Xw6MU4s4VMo1YfDVhn6f133byWBxCnIViMN1BXRVgX2c6R8qGxzrP5YwHI+aY3
8IIHJx7FhrkLwdAvPrRLWw9W9pkEwmv+6H0V3A5s+YbbJ8OpUczp0KaYCcQpiXpWDvpvf6Qv2dA0
4EtTtsjsEbcXRiPgQpH5IwjhUP/EHr6BBh/fpXifH3V8xsB+TbhnlmtSLdda8zpeyoOi8NkHC1L0
2qtjZaN/kuO3ZFf6hS9ENa9cGriq6uWBzO05JObvCjWxrnlA9b4+xqPAu+HEImgF1/sfyh5tRG9P
QPhDoCj9O6SURTv8SXv79XTS5fEEKIAyuLf6dZiAgpZUkKW3kZRZaZQxo4TRFHvr9kX9njyRrh4H
skIa+cAzOEuHmD7Trbsv8jTlH58TMgZ5u/KVFK/xPxpPIKC+oR3Z5cpKv10eY+6Q804YvMViiwmF
e2xwPfz+3LvTuVsEaexQ2zxNqIEq6CEffq3yvUK9xi02ncC4rSyG/A+a+W1fDIqLH3jrNHXeAtFh
NVZovbBwkY5VAil4xJHhBASI+vhKYW3x5AKreClTwO+b6RzeQ0dtPt8cXZidg7P520o54RPzVykR
I45Ly2So1A+aGwiyy+t9kYpPCOn+zkAA4ObbYQWNFtTATHkjQL/KaN+U1qSpBotCe9PLCMK7wgZT
dpLmJ6+aXxBNRxo37/1Ru9f1qtAP9YTlvziGt/JFABB28uzF3pieg/DRBEKaE0jOy+GUXx6HGg4M
tBtRpc1UdOdoi3gKeoZSfyWEOGPVbCDahapIPrtrS7mzDD5x95SjAAhzaT9cRewP2ppkz2K7qrt9
g1N8AyHMXJF5NuBMa/E3ZL1kmEmhY5fhp6P6/0DkkZKXnEy4cEhDZJGinjgXCjuKY9YMpsyJQ39b
cUevzn4tujK1rNPmzX3uIuyi/ineo1HThtaYLSUcbVKHxcsjDSMV2ChyGR+eVscXE2QlbthXXCd7
oCP19o8siz/A/ojwiumsy36HNxFre7O0Cj9vH4deyOlHjWrZ+jXagXETLHwT7gsLunaPPn8Oyo7/
O4IDXEYvZ/BmrCc2vPpBhtyQNwW4K4i680r9AS7e9S3S1gJGN6RWkpxyoe/bZ1KyMx6/VgXo/Lg6
3AJDs9t8CppT/EW5FVk2U9VJe6M0qVMZIS4f0dqBb8GWyO7vSuyWlOkmL0wlOzS90uvFw/qGFPb3
jyaIAPcIRP388ZiIAhW9PXh9PDHUUKBvC24ZtxwYPpDMmzSPO2XloNJ629c0FaJcNJTk8mnHHKVI
JLhmf3oXyI/gMtOZkhF8rPK4BLPKwgnGYqfhWik0Lv3JKM5GwNlrVEmmcv1OHV8Mwj673z9ay1zl
vOXNK/ULkceGO2AaTNIJ9O77Q0+Im9/r8zPEbMEr3oVVw5tLpPjzGsfMw4CaYj8x5KTXI1rUhd4d
T66OffP06AqdLw1eDU87qXD+kCMnLJeDPHrfeTlTjlWsHD1jRGYd/gG/S4b1kCET+6tOodxjW9dd
gSezDQc2zmUXofW82+wJ/kEk0cL2AxW2UvjMrbXPfPM1JDO1vUf8AIe+kh+rclKG4TpASxSMbSoN
TrAS6x/ER8aqvL8qhriJaeWUJP7dzPUTyVX5UzvHnhhPZKG+zf4UaWhC2zP7t+HVRzfggyBBH/u3
cscIyu3VQPrWMKC0/Y0lhS/odoEOdRADKIjhTVX2TBp162HdIU85Y928Oam/vf2PQLCvVx5vI0PL
gFg0G+qaq07KlaNoL+99iVjDyQJDjpBs8i4LlMD6uiBIftdsgtauUhghgxfx/2PYqs8Simf+j6Ir
gat0Eh8dwlRwakGtLD97L2FYuefUaWWKiY70oxmX5/TQ3wrStGq50O6dLFhH7Qkc76y8O1Uhs74O
AIDw34FHp0pJhYiFcfZb/ml1yIDmHaIdOIvDfQPMJ1qyXQrewyTImQcS23e2Lyymf/uFBJChyRCn
0UMIayStaBt35VlzESIgvdpC+vsHBOg07K+yeC1FvknRzVGZmd+gcBqEyNgEJFa3wVKtBz6NsAoT
AXnj5L5VyQ3BzoybAj4sNEKnq+ja6v42qk7mTRTDYLsWoXHUy4KzmkwohYu3+iZMTn2NfwIRO1Xl
grKyGFvlCO/Ib9lPMpusiftRIdpZaV5+HeZbqXFtp/LyWExBFO3OXHCOawBEWb6u1Ui5gdxjNNvX
GBVyps63g9sT5x8F4a7KwTyC0B2YpG6jXwVEkLccJZKyF9x1UlawJVI9KNmXnrgw8PSKq+BN4y+R
+W6++E0ZykZddV20pPopzBRU2BqYfs+zPCIjiTEDklQL0GasahyMFofaMrl5A7qiQm8oI8XGrX53
dtl7G6AwvEaYqEuvb1HZ0AWLi1GAuKkrX3reEn1CUqWqVjV5PTlTpeJzqo/h/w0i3hsBQ+WBUgS1
0gD/eSl4k6Zogox+5xWMO0pMO+w3uWtN4ynq4kgtRQOwRAwI5ZF6jOOPv7RqfxiR7+f7ZQ9z6mBn
mRz8Q1FxjhdausK1P0Z16Cafc9lFsg4mqXJM+ULstPDiSaqQP+2c0fNDXRmKeJUDQ+50XRq5n+ui
Fw849NPDDAWrstCzK3CzcGvYOhJ1u36nYEF3I0pwp1jTxNhdMgYcyvoOdObE36uoM37ru9+JnrII
hujIlViMcwb07UkBxKNZP/FY9gm0/28DoZVa3rLlx3g1HcLkTNsWvVocggGhFn4SPRCC/UscxoKQ
S1zYZlt1PYeCzTGTnKm735bZdj3JCgnKOten8MbJXPrij2dwf6EDM+PqXw5AXAoJ8tngTsJDFQU3
zcp0548H/Uh7M7bY3XRrivPMx4v/EtfW+qzpYD24HHvqeJBdkn87Fjr48hhF/F4VPH5NN6m7/OaR
IDHEMI277R+kXMWb7zBNTHXidWBZjx1Ar5fRclNFtys+wYmrifrUXBifsrqCs74ULk36B58tzE90
yslaYb6V9JWl4HNsI5xGSx8zTC6KLwzFghr0yOTCKU9d0ry7+rjUnop3JsP0eMqjAPug5RGJiUuM
iaswoEksGcp25iLk+0ESC2S0AzTOHoMQYY78lVfslfwh2iIGAJzxUwWT/gpj4c862w9giEhR/n5b
INPYIBJeW0H9fug+HPYIT+OPy+8oZuHdGtiny9UOYlUncvRR23BD5luXs/pnDCkT+kBLjjK64ZuW
9uPzcEGQ6xt0+K7lmWqnvWbO3tD4efJiHXVhBMhcHuTCoLgNI8AD1IVnNyWc0HZV4jLWEiQnI2w+
ua/bnhSXqUxhnFkAp9HX8JfkYdguDvWKILVMlMXugHqbxSSn16oAGwrfv1EQCRXfGlRdSvs9H1Z4
yQrrZuHFtefMVgkxpgtUqWehBdHgCayHylE/UhIl2XYWKb4i1JGgbaEBr1I32lRkdeDnqYQF/S8t
FhPJn7SQ4sI1I46VNmEFh96QuQ1tVZOoF0TYx0n/USCU376kzVlMAK1GsiXBrLvCsRmtyl02wGCg
/cBfznICi/uaXS0vj7wZouv1Ffw2tvGKGFyRAzDYyG06/ygHlzr2zBiBA0J5ChhcpAAw3EyrwCk9
WULxnDcepumO0NF6+BChUm62UY+GCckS8AjpVrbMQ3MAaXoIMYTL4fci+hxFgEbW57rlneJgNSX2
J120K7LBP0eP7ybgEXS6b8q1VDHeMmuX8lH+IQNCvb2MwDt/2P8ii7rt6PXeXemVtrt3ij8FVdCV
6L1jiQUvZXu2iOU58a+3AyXx4V47n5BckoWG/wJMUpKS/yirT2uE6RSd4U+TZUSHhDakskEa6uAM
FITqhBfE0lS6CqUFuDMGV2Q87xI+oT18vM1xdMoPwZhBaPNxN4rq6XFehKzSk2c1VeXt9ftOh0ta
6To68QMh516QKIaDjQd+TzjoI0UyNYUIqWl+1KtTOK8myA5GkO5TLihbVqBaiRlEpqybEI6DJ235
0zjWzv3bLG4Qq/tNTuAH8zn3QAf3jRjYtJeRKAcjOsBu6M2/zokuCl8fKroIyNiGr8A54p0+kKlP
13C4M6CWYZuZo8HMajeeJtESPfIfkitIpB0Bf/Vge5a5bTJVeQgizYJxhE4h5B9eE07l/KK7rCl9
seONCtqq+d08hYNVGnt+2yqlc9hNyFpDSZRtcx7mYlOUYKfCrh8EPDPZ6utnt+xL5E7KaTFcNB+g
CPdNcJXyxEfcHMW/RxtDjg2jyyNeRcgCEMoUj5aa5fEZXsPEIJIWenaiElYX2C0xS9Yqa0Mwhfe3
91em95IeymUwvxsjh/ujSTrxQlnL/6pIe/BzZCdAKkyhnvsD6Ge6Hv5QszTG5wYRjJwzFSEIwW0c
rpZ3YtbpH5x8u3JPFvJruA9MOgy42K51AyP/oSzPuqxKQd4IQVPbbQ+FLXMp1e9+CkYmmkZCZlzi
L1JIIKbOqA4VlWwKBNBTg1HmYf2jtX0uao8cbifjdZBsBk1PUoMlMr+6J8pTYAHvwuwo8Xl6nFKi
YIizuW8ZoCQcgI0pz57gEu1tcKI/WmckGow5qKdDLxRAL9nfqQ45dCiZQUcpUkgREWaiohHKCrED
ykaqe3F2CACgahAGKw8ryiYbqnx3wbwi4ZK4wD4Ubxk0jRfFOPLrgsRFp8uI7KpQw2ACwAcDQ3XD
OSJpjI222hs9arnJ2Cjrege3b1HtaN2BqSnujrann3vtt6y2kfQ0tr1OSw/8tBcAjHaCtL+ETb98
OSP7U/v3IuJuttHJ/BY2zLQC63hneYysXN4ohVz4UitVzM+NkYqqFa+gBFlUpJXNu4HNJPchO7M+
ADPrD78Tqo4B4YiEWyLhiWEwdPUpdED3zh249v1I/e44/A5cEGvvh9suzUIMw6bxEbdqIo3lN8lw
edGshOctq5cxpB6zxOFEQTmVcjLstqHIKI5MsgDp1i2v/NtCp8dQ/h0lLZfmleBIFavbaBJ4a68y
xlYx+kV7dHJsyyWStTj7e5aFo2sDCaOWUbXE4f8hLy5D5teFop0d3BSxgwCmrdckapTxn0NgNy9A
E4Gk+vQIN62WtfTsc7U/Azy7p4mQ3Mv8XuX6nYYtrD7fAmEuyY7BscQog4nFlAn4ITJhyxSSHmEV
0jJmU1UVKLC7r6YUNoU00Wok34SHS7+XJ7jtFmj9k2lQRhISdHeWOuYiqnOkfeVG3Qyv3t4kQT0a
NxQ+hfMrPk/foaBPgMAoXynNf8yRpmWG2rbLNSHkgri1FtdFYBcmdIXceZRMZQTu9Fs/mMK7wGqS
aZcWUzsDbi8NYZ3z0rO4c1KQx4cXoskGX0qYpjTX5E9MrvJ/vmm5+2BbajplBiOOoVKy5Prtie1g
11RHWtRRprxa1z/ov4rdLymCk++PwwrbuWZ/VgN8oXM3FjKrbcRdle7U0cJ9HYzxcq+Lz3tP6OUU
txOnkXSWAws35dUOnt/eBcCkeouaGeezDp5vobOipMaM39zsQbbZLiyj9PT4f8ha7savD1crk9cQ
QFG+U3fk8U29q3VfZMGdJFnbJVXaTAWc0/zmd9DiGBml+k+Eb+cx0rk4zuXoDoN9dAc244mw3sgf
eNijVO151xo0hCrY01g2whIwsRbtSqkryYfioEj1jSm04hVYKHPSzauj4KxfBoocMa1gKIM0n6z8
/cIj1nhtJX3bcLW414xcQenH2jPbHeJDwUS0qgp6xjjnXpXRtc7NnRTsQmmD8FVrZlj/B6vR2bdo
1D86GonvJtnjvTntOeNmrQwj6haKi9G1rct1w1AHeUnK00m7/+rO6/ZrXXvv+iPK7URsHwpN97Yy
pyZIuneg3y6IECosRMbuiAmmJuHEjtAQFebNQRUJviVLwSgOfH5IpmQJAauj4MFK77XER78fvfez
ACW/gb//T/h5AYdnJwDDNH6Pq/j6cwcVV25VH6JgSSkWtk23+xC4kGxMnklIWu9UJc91Qv0m1HtL
9f2tFUFIrOC3iBBdZJqcQvxNmWi8BpR71FyRGSfN5A5+dNm9OubgZ2i/w4lnca4lqUPc9AISWVXt
RH3FkGpXTvzoiI6n2gu6UK50Fz1mJtopxG/eWKnXrYPcOXzAyuVsW881Y8CjuXaw5L4/UevTKFVd
NZiXgC1nL5DKegMJagA0pRwST1lQ0Vf9g2tnVqXMlI/ilUmMtMlh4AuymuBajH4Rvg/j3Mq/R0y0
2IqIp+oZtqa+uRkxRX8TomPJV2PSbM62VX67A3rhxVqUBi3d6AqL8VoEZFhlUUaTUmxwHHLicOmI
p/VdPaUuU4PuP0/dTnycw8ctgMzCQE5zGk+3lhJ1NaEDbgpg4QvfKlyl6N17UidHpwJj6MEzNTVZ
UqSefGxhVohAhSgRIn0GVUZSQpLt6sxN93WQQJJJn7B9CHpeMhpGOyQ6zNZHhpm/Wm7eaoEItbZ9
S61D3ey48RfGdRrO1kANfRPt1uoDaDJZJWUgl0Q1xe85ZFRf4yQ96FSyIIpEaZmAS4/d9ejYp5Da
+F69W7OCWUqrhknelmnWIn7z+1Uw3cmMYG+9mMdQQ8/mPcW00Qa2L+o793sAqg+nkznpLyT8IzG/
/KTZ5Pk9abbzYt2ehnqXzmJu6j6M+vpMLYAefQ7ChMZsXAZe98eqs/aqlHHeQFarV93PtFt7pner
kjXfXN8ORylAqQK9RyoTnC7E7LZyhz3mjjpveW1LkPgctf3QZuHe+I75XbPbPdgXlHoVk+mKUcoi
IjCyzpKtldkieM4cRXT4oIJzlYoZ6f+6OcMQ/167EmH6r5ClZFpgoUxSr89XuZyYWX3eMC0EHpD5
B26gqvZeogp36X/vxJLyZ7mallX//t1MdZ8BtjUPByaICppCKv0pS2PILZCR+YANNYGVgaysPSrn
J02PiIUratuYf7HkygzUe/Y0PsFCa8dVHkOpJRmhQghNm1XWU/Nsw2m8vGTIK07VoAZdn+UdaESd
yuMc25fdyRCSmFkAi4fEs5fpdJ9quQkpB+4qUUuU9w3l5YlMu/eiIO7XbCzgJ51H1KUMuipJw+6w
9hT+FOGqhxbfMqUIne15GXCGLfOFVFWIadv3dgH5hE5gYsGSVJJAKqvJb6aWisNWbD3YaPpHMufW
cURWoGud3NViFUgQbcxwMOMKKlOOGxJplxRYeyx2y4QhVyUDjZIk8SRXinlQi/MBJFfJUfKSIGMZ
QbMi0R+QUIA1qohcHfOtQh/p1q41tEdHyE5DUzrxz3ikNju+Q+dboGuLlQAdJ8fwIYsM2zhzIWbJ
RwEZM6h15chOVpBbOVGXfgHi/QEE54ssxDBefwdDyDk0PoJhGm4sS6tIJQNuv9DVZ+r4FWrDrb2y
+0B90aNwY/r+u56QLRZOzkSm4/WYtwq9NnlqVjzV51kzmcKB8udOi5SNE3z7sac9DyzDtg/52xpD
nRbj/ETza//B2YZIlKq9sBEM8K4mci/LLzOfahM4rl1owUAtBMQKDQK0wjNjiu8vI13icD/wkafu
9KFtFR3CHSD+kK2f6WQUvfhLxS1TQ14tybvHGuviR4ALjeSk6V6EEw+GqWV4SaXDFSkqeoaHeAjF
cnmFKEbKV3DMe0D/ZkyyeBsZyLzAPfHFzC0gCAOPju7uD1zfQcxqHyvkavX4puzGyNPRFB7XtkEa
bJB9d4pKQS62QD7g7bRxWBZrg0oQrM+3VWtnFOVBHCw2W83e2X34jSrzAiT7JzAKTtZJCU3jRMup
A+qlbD8ksIm7zp4qd3h+pzT4A9TyugaVY7X36SdfQ/29q6zj9aUqDI2eeVJ3ZswCoLiLjPObkzzE
RKoajRaGKdGvdnXmV+asQ5JRotxKjmzynxiYL3D2A/bqFylWL5QbrMgIr5g2vmZncWMPzsxi5XDv
uAZiAI2KEHVdmNPoW1TBgFR4I/S2AAL6f/ehb8mdPLOXd+VP3HREo3xhMTE6eYEfGCmolWQLBj3H
X6Z8aKpgXn5FgSDp8a5NpyFcMLt6X9OeaqYSH4v0Y7Ml+xek1KCLXnEMRMOpQ37PA7/RmmQ7hc+x
OZZyY0xPqZ4XW2Y7n0/1n06Jq+wSaf3W/Tauhi6pHdEQYCf4lDUoU9g96bbO7n9mRUcope6IWOo4
w652P6EXeWczSiq8jb12Km4tChoh4FJM+V+ASvo32Z0Rrfb7cfbsgENZx+MbIyqepVwRmsHqjB+K
USJKmWQqVUPr83dVDdooMRV19ntRug01Om0k6ZgSUKcVbEbe3OJ8GesfWFVn3regyGd/TA3l/Oev
sYOYmeouaOmfZlGlrdlh0bsbolMeMKPQdwMJXsrjMdoAtr7LkaX9Z2DKX0Q7y7JjsmIX+L75PZal
NaQqvNCR7BnBJqxvq1UJ31SpzxEp1iERIoQ6IxfuJpuW6gX0KaLvh4VsbzUtA7c9Gqvk8+KgDMjw
lpPPeGlZqyOWDmlEplIQgx7VvmeB2Ri1ZQ8EGq0LTi2F631kaiqW4t9qOj0WUE8QQkxfbJVReP5o
W0TbTihSIMu/B1LpM66xd+lYYXDpqpdg9d+c/H+U5I5rmGBfS8tIJ+zHP8Aryq2/P2JnsUi0ulu6
bXHOxuiYzZaXRuETcwuSStHHDyHTaaZ6AIAohlLHFyBOcuKEmPbEjaDT9AORhkYLcnk9FiF0C1GX
xjgsPHQThU0CocayiMqpb3I6pq7fgczmBlwSJflqgEMk3IGQ2vmTnE++N75XyhmL7LjKTUD9uYrt
X/AXbavmPN/06tFzV4Dkm9de0mzMwTg5qeGrY7JSh8512bTNAxpW9pErNI5OeAemjE9iffJ1O8L3
PKQJJObQpdQQ+KeBsv4JN9dtbUYnrzdjAlcSGmVWi2713bf0kuhiQ/C/Vwx7B6MbsjZFu5k1eK8L
IDeGUHR9ACQB8jWTvlRJn8QLK4XouMN+tB4t8KrjetWVTQdOpfW5OAMUBHrVVIySu4E10sqRAye0
JaYrxDrvriH6np5UQ2ym+SBIdjr1c8N4wERYFlRpm58yBFyvdnfpKthPDsvxnN5JQejv9gn8ol6/
wJvEzXkr/7kqaerwRBI19QNyo7cal+HiWzlEm2xe3wJvexKyGGbttCzgZNZ721xg3tXh5IPpYuFh
oIm3nskklQ+EAn+NJVRv9PCQgyAtRz9X5yRsDgM3jdyuXRgZ646QEE7jSSXmsI67x//gkBhUnPGx
8Ya+9U5wEsVJaJSdUCNKK1xuf8vM4IgBUjfImPQs28rSCIlkz9qSx2Nwfl8s3K62TdKcoKfTuUjW
9bMNqcNbLgMbv0iUZKN5mfS/fAJYBZzVWOpI+BJJ6pXfwd7fWaV+TsRtGT3GUlOCIXSGwW2JFPkl
L1MwMBbPPG88UVSczXmwjkII9Sm8COeMMfYtvHbSaJ7kT83ohYzpm0V0iVFQi6Ew7dE5VePpX1iU
ZxqmTt66KWoLOaOPsqlPyEX/0Rn/6yBIoJaX5kRDad1udPX88JPJQOrvejt7ZFggiQzlieJGuIHS
UNN+NHtCcBYcvw8INgpvdGVrttXiCKNy2HA+A2HroJKo7yRgBNcaBj8ZsR8Z2MFBBgwpeZthwat4
HAoCs5g+F0E6ES3keQyoED6kurzcVLQfaXFbw2aUVFQvcvJsLkrpQb+B5/9/QYAJwqHan4VARyYC
QNJHVlpXQqA/Iiaph3mXke/6A7ldwNbyOoVRWWd+wAE4+LoD+T6UWrJhwMSIYvQoU9dEFSTYN700
iTFl5hACVjewEF3cuHmR6keEuhltf4oqjpq2zAbY/9Huqo8QUA2wRzzv7J8YnZK0VKd2cpTFhn4v
FRuzNOx7MkT4uuGzJlMlcf6dDWGVOGuDn50t3V214bznGXJNFcWEEjG4Dr7mJvO9k0UxK0mPX61h
ACXFihNgjvUCflHEVr/xGEYeo66K+pORb1reOigrZUuAx/+GkEZQ1Ino5ROmZIQbRVsWKDmLNdqq
jJqzX11k7acETpx1tqND27qoqXIowULn/lh0TVEUObdMRIndP3kvdlU7IC21doqHYfDesSbf497V
KKbPCXI85QKSZy0nHm7KFzOq/kkzwgkI9Ipwsje3BsgPxtrCGvaSFAZbA+aC8oO73rGYUPJCQU+O
sZk4umgMLVfkJWenufO4wYMUozvqGaHfSFgseyzW4f63/3KTFJTf2FX8ul4brvaxIlmxohIafi+c
56Hx3BS47eMxHthid7C1txZZKhoRrHJeg8hbv+QtNtwChPO+6+Tb/UwOXDzC4rDozyalB0sd85mP
E/MLf+5AZrABsKrR3CXjlgDu7edgHRnvB3RhTF5y8jYL6VnDL2hgqUpWSSVCEDlD+h45ItIhR4Eo
RD5FPtkdvAZROFF/Quh57uIaRqSb32TyThkgGV7V1NHonjg0eto8G7nNc055VQX1eWSJfPDkff26
yqcDyRwyzrACnq+9QuVHfUcan5kaumL731r2KgLRWdNhLWVu22of1cCNNgC0s00Lz02AzP2PmoF8
+IyE8DZqJq+BoRqTYtxFo47lFSEjTMFnOhmnpQYEM9daGANYI0/rXKJ0Pb2/6Fn/BQw5IwRX6jF3
fq89qZQaE7Y0qfjs1RzGwzkTBgaQG6Ux42u+5BexxRjYeLSs1aRqUiyf5iRsmCBymxZZ62mtGxYT
dg/OwVMZKUajWi+I2hp46GFeDQjpPQBoR/6jyY4vWxhm1mYLFUgO3/330APMhuZqQmfLld3ws8Nk
Ers2cEMY4EkGWA3j82GGmXbK2YPLni3yoih/37MSsum/onJiPGxpRJujK29HV6xiuTqRXJZq8+4f
ZM9wEMrT8LMGwJn4evBqCUGqxT6CJp2gJW7REmE7jTjI4Vum11npugCUO8yYZtiHlg8qv0iaCffa
27jcn05q23HU93K1mdiBOMNSN9+1m78JqT/80h+lT0nF9UC5FjH662pp/tM/NJTw1pvAfCpe7irr
61r6SgcZUhNJeeNxXbMmXWTo3vmmAA7ajH6DzZznsvNcRzSBklExrnWxa167nqkrIf64hfqxJqU/
fCLX7NEZVA3ilPm1ldc5m1qf/4Oq7ktviRZhEoSZlvXyp3kqDtHhNSUskva4hqngK74bN5rjpgf0
wj2P9iG8TaxkCq0HtcZKD0vRCx3vyky0/1132M+8RJJ1A7XuZZl7R3XDIiOUjHp7ID44VpsV0/L3
KGGnf4KIPYUCGXNEeWX23R8T5UVzULRp+93D2g/jz8kej9HCX1Zy7k0eDcayPrFq9lUnrTjS0W7X
kC+TUAax7hXTpFpMEnmGocspZVLhZtHfXtJqJBY+BzrDsJ5PsXvTybFfzWRDj7+oK1v27kvui2gg
T5d9F3UTglZNy/Bi+NRMCr9zyy1wCe5QS5OsxkHOyPRVrJEeooLgxwIbFmZEfkRV/QZLEww1jZAz
P+5Qxyczqj78DR3yz8YgiMz5LoNWx1838b46loQU018miQ68iciJUM2iioPOBKX/Tssg0C3Pzm26
pa68ZmyBz88V0V211GhBwCDVl2QG+GLEHIUIw/AKlAl04m9MuR0c3zmnmB/RS1L9E3pZ/2PzIR6W
0zGWIUemOMd6CtsTQntB7U0ITe4PNhC8tcvzyWQiAeqrcN1exEhXERrZFl2OtYHnn3rVSxpss94B
BSE/1nXjI5ryJ8b+NhkBSaJ+1D1CI/6PXTZXUwX18GyJ/P8wtFY1CsKeWvNz9xPZTIvFkwczyFHp
wV2G+ufyY+yM2eGkjR+RX5jSffj+DOjdz/MdBx7IyInEx5S+zZPsZPi6fzwpIEIIiST0Jr+Y0/2i
GpsG925SQVpyMcQRweMawZL+QqccKqOZB4y4j4vGePKVNL/1nbFaB5L+BZg109/jYqq+EnxQJ7rC
GiLAn6w5eEfWXfBJSVhrqJR6dIHN7KV6mXOH1jZzjoD7W/ziHwo5hPH3CBPrbxQjqzqD8bmDwHC4
FIcp1oUBICouJX7fwWALwI7D4E0E2N62GPteJegj6xuBMIZ6BmQNUBVf6R+AtWU+vAXG6lZRRDQW
YmGmiZfUrOz/dnbzkcT36D1Bhay9wXMZco+pjKlfMCfXR0eS+dWX0w7VPPLpFaISreLUtOSrgDLR
qyhI196MpQCIIywNzknohXm8kUhgZlN6e55kHsbW0WoD2vXyj9zOdOIh8NOx01hW45FNR1dRO9cl
AL/szJslfczRKO4Yk4F8oIdxKzb6xvr9g5PwiKArqNXLmTK9kvaTRjMWglnXOF76sr+rzQnm1zwo
1/KT1FMGjqmST5IkaJb3mI3S/u5ITFKaXEHtc6Zlo6yBQ28s1oCTBkvSkCU1I6fZkqJy+SjLC9Yc
VVD7giCib6mMiJxyFdRUyT1eVbB60yS6uczwZVTiJ95KSIcQh1M5meqegJBlaPmtzYX98PlvLLGi
lvyHDkFSoGVFA7BlnA+jR0S8DBjkXuRXt9h+D7ML2r744hCVByEh97cOaiHyuXIDpWE3egVLhxTp
g1XqXKB6GoLUn+xb9rlfIw/Mas48NJdyJ95vJi7b0ZkYJmAQ9xoNl7WfRdW6QAr057x0wV7f2Ae+
WHzDDDA/ircYzY1TeP7XzC7bcFPcjxRyTGwKH6R0asrdcYqDw25aldSW9UX9GwTaz+O9eBD69fez
VrIW8Nm9JE+lf4hfcYwrU3/dKzUQoNmKy5G0rF0QoYcWtX7DLGdU5NEQltCP/7fXfaVLY5j0dHqD
s6n6LWvru25i2nzdrWQqGy10arD4ALG5EVm2+jIf3KucNQ2UE5GUuzJlcT3Olz9LI57KsiOeVlEs
+ci0HQfPLvM9FWfJj1MYPrOlFVg8/MpYV1AsebTMUZyC+WFt/vVYog/z337vnCIWY8NDYSxnKPql
Y/h7jdWO0iX50d+PIhovYq05xjwfNvlqknDbKuK/hM7at859qQQLWIMQwmP+xBB0bnO/QuoHPPrn
gQjC+ISzxJHXXGEVgl8OwPF48P4L4FEEz3W+emGJT5iWVAAzaT+qTW/IxbOkRlOlE6VoMygh9jn2
Rcpa329rc0oQJWtohXuHBJRFLXmMVaZEmNJ09+ubBdh35V1Yu6V7CguYWc/OOFuqq0T4u+nZdgiG
CGM2ICT0McCvaQY/GvEZfmzqHWKxWWNCrGvLKWLloWFvWA6Lc9Nb6ngYZesU1RjXUp2qLGBHrJeP
lYEfeHCCYRCx3H0cIySH7nTYaz+lhMlx/K2v+Wjvs19bZNmbsW+qyo9K3r3oEpnlS2IMGVxYfEy6
o3Iog8ytk1bj0Q2h9pQULLMNm9NaLGz50Sva2oIoWSAXJaEhUAcyJhSrRrrQtWPMoJacpxpLhcCA
4G6KgPe10CaeKBsKQi4vuVMR8Y+2RC8kpnm7wef5ibZTY+Tlxmw8k31ZCwtdGEq2nvcGKHw96Gua
tnrGKBfkMqrnKwrVcqeAHNwF0f6XgpoeWqPnn4jDAtQzoumyYpWOEEary3qNkVUrW6hf5XW67QLI
hZWuOZvQZwCoS/spCV2/4Hvh/X81JH5GAwaZaWhmoBH1lTfC0TK+1W0UvUxNuMQf5u1to1suioZ2
uvdn4hRnAJqo14b4Wcfxp66BjDT24he/a1JlTzm5Mb32aOU3jSgXY6C1GfPADKsJSrut3o7tSq2N
U9AUMkkIjujLkawNtaCHtbdnhQObjrxS00/2OClDaOiM1BV0xS9iBUDCNN7nl9NtIcxFTzi6y9Tj
J4Bdi21CdiH50LmM2fiTcL3tUEXtOpCmr7ZXkR2o9gM5laSfqs4uXhG40DpJKQ34laxgTmLadA0h
aL6TIyiogEAJKAwmYP+lsPe+eA/1mW4eqKH+MfMIcHSgN2yTz1jjt1ifYnQ9f/pTp2Z6kUXcl7xi
dFEYtpiwikI4MiY4dieSEeVm4UohKqcZz+BJv9EiAMoCSNeSHOkl8jNJGcSoSK5qQv/Wu5s5al0+
/mRp/TIJwpfiN62M3x1KrdKxLQarEnfcX/RXjqBoxAI8LTzFJ7XuUG/4fnBLERHT4mlwst9otzkg
cvLTJwNXwJlXJuxXxHSMEhwvnh6jYDbwnZ2CyNELKgIpEGAu/mCC9+eZOdFof2dBYs6BiKs86+lr
ayf2OU2wjzG8iQDGlS2sEesDsUNrpKQgUBnR9i7rNeqPtAA6fkgWaQIKNXx7wosXXRFxuEE9BCYg
OIDyLV5MEtfLNEVGYGmQTStLYXhKnyc9ID8ukKl42kKEMe8rYq3iLKgfCTskbLd3CNHy22m8IsbR
nBFWr4d++cIEC+xjt1vNuasz+P7rc4oASHQ20wxbu9NOdX3tVfTg+0rrpMVmuSTJjwfj/WkdorND
5lASSk4e+cZ1ozKVT9cdzI+fVc94O9qGQlHjpWyGEkbCN6mYR0XTiIG0ORdquZ8AKTwLvf/1Ec7g
YPhcJUBgW5PEyzWU1NVQsFhHL6RV9Lm7fUpH9Qa0DN3PsYGiXQF00DK1ZANegj1Lchxlrs4EGw0P
DBBDqMtzXTALf8dI5JM96mZuO0rkNoQ2jYJMBDu+DAwKGPKF3x8JOOFmblza7SQcDgkXh4MXAM+h
ORqRWgx7RTaY1ZR+c9ZCOlkCPejRbwdFXWUTSppLe7Tfdn629MYHuewLk25mYyPxKlxdxtdH1e7r
zXvAwLC3ek7JANevQwHxttgfmFCmTQ5s5IM3FpAufCz9/QVdljUmXM/uDM+xFqFijbbHEw68KO4S
PdDShBwu0k/UylTEOqJl5crDcncvuI94zAnLpwpitBx4jrpujh6rL6Svh3Cf1v/pvJVvWqCklJtB
HwCSrv6HIOTXIiJv+Ve2ScDcwf/fMLjZlHfhL73Mzo9fKKt/1p064pDZ+DSeGY/coM8oAFyMddnp
3lePwJhjy/gu8QkmLEbWStAIfXu9Tkp98wwbhqSD6oms2F2Z6IMp2uCAWUELkX92IE9CNGdTnzhW
RNGsc1in/m5oohFajcZjFdU9F5FWmAoAxoPiB61MDLjcgGfNIHAxOcV7lgmKP8d1bQQIKxNlw0g/
F/3T37/DO9krdf4yeFPq7OtpoBqCrcUGkHvvuMWGbhfW1xBK25pznYJwfDtABEcHEII1pUbBic5k
lsuLoiqwVAFg613KpEY+rPE3x97SHXre03oAQxRUzjnl/l2FbwFKHrxlRkfELvt2SAgd4nbz0Dpq
7/ha6PEWt1YyPXDrKrXByrPvXsTYDgGKLxcjD701Pin7wlZ0D6JpIETK+dKj/Dr2aAMHzNVVwIuH
iLD7k3uzN6p1l8/YayHBkGNblE4nTdauSPRH7AOKyasUTe9/icCS9px78ABUR7nEERYixmmxySV/
dxTDm5AIcmqBOm+IgoXTmDt5uoTNg2rTUTfF8fs6zVELL8OsaPLatFq8uekQ+6ojaGmfdFNKMIPH
AWrgu4UDgpB0bAjzt/fex4c4SaqKGtmpdNT9uen8wvjlVRd1ygeS7W8/1v8vNLvLHk52sQdfpyKq
IKzQCffiHzvnY21EqLnJXhf53uu29H2WtxelvbUp1G5qAu9ijLopH5YJiVIgMtv1QmjUXnswGFdT
/gcG8qGvK+6DlQFk01VPlZA/rcGD+u44YTcNOb59mD+R3+c7crzEmH0aDmSOkAJLcJQii/Pedem2
Zaae6qlXbNqVdFuHi6gGwXE4zEs+BjniJ5y3Jd/W4dtkpKK/saPjMu06Zl+BvAMWr8nsHALRVh8I
KbWAOGy8ycgxBGukioTkC2p3oZghDhY183I0k1Dp+oKz6PrCWPOHBjV+YH7Q0i/aTI87/ESqIkHd
gB+R7UFDWAiVaJ2POb+YPsmvHxO/EscvxlHQksH/Sozs7P4X8T9huCZU9D4yu819e+kwptlckoqU
pTWfzM1QH63ypZZCcAESI0btc2MiGOyR/A1HQZ3oaMYnzL1l38DD1BHDRi9ztBFar4ZMUcPuc1ue
ero7tGNx+EB4Wh81r2IAwzppBC43bWjIzH6rD8ZvdvrImt2Zk57cbarXGJ3MUkpHw7zKxD4QX5y2
WG1a2wEXepG6xPTgd1BJ6BYGmeMbNXOh/+GlDNjpoSwJuWv9NqKS4USMtzPletrkMtWt6zyhlbiU
wd4F4Ngfowcl98f/HzLRy3SB4UpAexddiQ5Cvkut+6Y17Yis2If9jjE1tMLITgOfP7y0Q0u8yDWu
tMfS699Q/3wu/sN20/qfw2vsZdJTUqiQp5rUbm5zXVlRrg7vUtawcmrB9al6XYg1X1wc33WKd+4R
8N1qSc/XENr1IQS/CsI6cNLc76hV1xYmLzd+tnLedNk6+4qptQGJg/x39G4veVttD2n1osmwodBn
9jhgmaSOFKfzgcVJ/qZdJFGG14CAxA6KJXUG5oNxseDQqeK/5iCSkFO74akvKZDu9yRLTc+qRyna
h4yrIMJoNAQQLuaX7Toczq+EKpdZ4a4Mwy7s3kmPWwxokXvRX/mKQCuRxNpMwzNkrLMBlY6iboPT
eqUJQo0l2sih9+9TcYHJJuU6l6WAFI2Ak0msg1ZbfYjDI5BpbGnOIkPZNHOwpHn4YMiCVmeGPVJI
zFeRfFP1L2NLcOcwrjJlwLmTeYH9+N3BUlv/HDZNCG7G/z1jfGwjp+UcnJd/pENm1YQbGYTlck8J
Qts4BYjbz6dc0ktI9z9fI222Q3ibfHcb7Eueh7KYk41rlxs7HMe2ELiAiuwV/0SnkWN60Ynz0eZx
YVYzedZnqVGq4Ty4VNq+r7LQtQd+At1aMIt6V8ikr8pS0A4i9uz76dci58yrVtOfPT0gfCn5/v8r
lUDE2jbGfnJNn4P/1Vajs2s/qXlZoy9o26doN7NveAm0VJAE54pj3F14z2Q4ape5CASw30q+pdhX
ZedBBSC6wkalIBbXfB/8M3gSkY92La4p4ZfJsVds5ya/FxJt2a8WH0NB4yx97ib145ed6UI2ZuvZ
ND57wXkuzKL91T8JrbUjKp2GY8rPq9PuVopA9QIcSRhheVqYVpfLyOuSmRXIGCsi9U1XTzmJ4AE1
nOl+mUtVzQLsDVtHz32MTpv88yI7yzUVwvrGcIjjMemtC8QjDnRT3SrxGfemqMJami1zFk9Sh1qK
pRydvL6mIDggwvyf8ejAF99nd7Tf6vel1ZwWBaRrta5q099/j/f9236cY6lR1DOrcP/ECWk7CcRV
NbzMozLsak4E5bR5Zl3TifBvzDO4wCxUVmNAm15ArERdkBfPAqzMOh3VLBVSqdU4Vjev7g8e1lnG
Pf20bxghZwSODUD5AOP3Kro9CdrOvWwCJc/t/xb/dLt/kRZe6LWwLZ0kqQ3mopd29yDnnTg0YTE/
+sJ4vRkPHDmDQm+ntde/0iqsM14jwxLDEGoxksc4SosIrjI+OcVK9YNkPKLpHF+TiE5l6kKn/HIc
qT9RYMuIHJNu1Cc/4scx8DoqtJNZRHi4egvYw5uAk8bboJo6DgWe303LNV056cEOS0O6rpZDgIRH
zdliX4VVoIQvW2nRpNVR6KfsZLLfYx39FU0+xm1xKMt3PMgTxarO9eYeD+S6Jcmm72arUPbLOQZ4
Q8X02PPwxNwUslHtwr53ndgykn1JcNoNCGze8XmLEhphfM6gRnuh5hHJTLwyyVG9RCtwY+xLurKW
APxcviPfLpGm6LCVRymPQU2GlFtWzWs18qmwqvDdDvLBf9niuCOVFRG/lEqJpMquTbmE311eZg/K
PIsOzltYCkeUIDVueddWsyjCG/5HrbRcSocPxEwMU+Z+Eyp4V9fggJY9Tai/axknvcQLSPFuwJwu
mJeugl73qJVz8nDlgcDSZUP3qVuIBPm07gWYUrSHPYKNw6iqD40FfdWd/wNcEgD6taD8i9VvwQwi
uIlJbBLf1x8aPQp3Zr/XPaO0Jq5tVUDTY0K8l+ebp11hFnw+kd0aaBF7L5aqVqVU+ioVIIejQZM/
bEfvkX4PLXvrYNZ2/M14OnECG9yIqlNGv3czj7M2S/5s9MI91BKdL+Wmi5FC4XGjjNcOjzN+V/Lr
0tecHhFr2aC1lrnJ+SvNgV9sxr1sBb08ZxQd3iiLJLQn+3ewXyVprLCYjQx1vE2mVbWAB5sNYnMO
SHZa+w9Sl1bYAfIo9ykeTmbWriWTSEAcxJKqyvbYEcesgZL0544xlOafM2UJ3QB9Z/hjiL8uEbil
fKXcOUHFajw7e2twSN0t5o8w/ZQaEiSGe/tQmXLbJKNghyAAqdbri3vrYBVPxzJc58eO+c0GUXLA
GJd0jDDxGTzkqBpxQs9ZJ//7PNla8Iyh0k6KSg5GWTeFC5LRY2uw+YxIplPaGkLcB7w4+Ksazz2y
208YqOpxEmwbfk0Mj/mU8so9/imISVPgIKU+lYJdU6QIWnreQYt8t5H4zsDRdC0xMAfw1QWnT2H1
CmaT1ITtudCvwxheJsZjZ9So6djFLVZ5yCYufIqwx1KGr9eA/wSarWkdZmsYIj0PK2NQebyPwphE
FOHcTji5SYTxuF5pGIIva1d+CtqBT7hzRr4dTGV13u9wAxvp0ioLprtBABVb3s8qNjO+VXrAGCcI
rO/FL2jMfScZfrzY3ClKxE/6KKfEFHHieSARKqAexT6Api1YQ+d/TpOzmPTdWDmeU93ORnQP6HSZ
VMdFkk23xOKaw8WgiNUl+xu8PJXSAcnXlKjVgnR+VNsdESbNja6j9n1OdHtun8LdCPxl428zdc8Y
JWm9xZdSm9CJ8YDz6/cStfpxd5n2uA37RoaW2hRX3nY0iCk4DGWGYqJoX0mZjVrx9eHpSQ8+xNbN
TJU87ISsZWGZD7vDL2CNPs9nfbm1q44aXX29XI8W3a/UgnUL5pVG8BvBizeMm8Nr2cNaUo2Ja5YR
qhDSrg7AbF69AXeIU34a5h8psr97htU6nZQ3+OvG+YUKvrMeNDsGeiEwsWvj7fJbvwuEp5IuUAoY
3UPPuLDRRTr6GQyzqp0ggsOblJbfUuv/OTszUn2WFqlSc8++YHu1rdJ8lBYcUlXaJFkL72jt64v6
xaNNHbIR/FTbQdVbT78dfZ9i5pBcKiV/O1i+Gf7tZjV6RsPN9YzBclbpVC/ISeEpiXnGlDEn0p46
PRm/HMtTc7efHjoAiPHjCkVFsYzGtI6B/oMO6EwIfXqQfsejvyrNn89fKWDtQ3Uk4eptzZdFUJyh
pPQPbiFvun72Ae5MI/cr/jZUHn9bUyQaetUipQ17Z8CrMVO6/P3/lVJwaaQLVmnSDfCQkRh/3ei5
nIcU/TzRQUC6GzCXqE+yiAeTgm2o9xKRNKYxd+6zJrpFsxNMTvVwpbIOADeDPyAjpIUFI2/jFepv
llTHhmX9tju6SullRnUo3GHGryHTUcLgO2dP7I5BiAUwY8La3cdbqIjbLIBH4jWbU6a3EofStqNq
hr/xnaXODyXmIlmMxYOyE8IQPX2PQBApAVn3qEfjP/lJ9z6V61Lq2oRqMwJocYNL7U4Hp6EYkaJ+
YVeoyt6bdF1goVbrjF3QTXAh2QTMNZngwIF5scjUu0WE5AVRousPwr/9EcyDjKyohjw6Mv6xr+aH
BO4Zw+riurPM7UPI0wdZByzF0D+kLqanLfJZpnGX3AtZAf1CpR5NblvD0NYL348vQvueCXiZXMD2
oWjrEuhCbHzE661UZ1AloChreaxzTyk5O97pdpNIUD3NfM94FmMwCr3XNKT7qzExdLCpnSkVvWqy
1OXeEHbhTLWLbRUI7WBmjJrlqIn/rjlMQZTjiADWsAaNS04tb2eCMwdObHW8jasmrH6bEqRMggoW
M0VcxwMW+n9e0H+dWMGni76rJMv77LDsnhrX68scdvU6+qKb8TVWJdo25avvAGer7BarAwKmIKBK
4bi9wNRvzsmiWMOnsEhAER23ZTnB+MnfeHmkexw26lUkVKlpl7Y30alNecGBtowICBbyidfUG/XY
s17C9vujl2C0T6Vh4/jIJFHyrN5OfPdqel9bOqwKra2TUvIUdyj5UZ9LS7S4XjUZVQOHjS5b6ch3
zKkFokUQd1Ph0lT6jzxKyjuV7VU2Js8w1wPVi0Ru/yvOFIhdASdHa2sPviqfEHWtjGj7YfpzhXC+
d5c8XqblNGo701vyQTWDOFP8RXfo4/Xw8WjC4Hm2JZ5mLjE32K7uzUvGX+XUgdUSv3kuYwLo82iQ
u37DPso2iawoCKeZgJz9SP0Ivy9tqmmY3dMXkDfEYVFNmtpTWD9ctaJTLywwN+bKcULdRG/fUoS5
LaIgYEUdDugdX3eztYwdSHMjklNXKPGRc/RKaLEsNXliZkAEf/9b4ITI8Hotc770h2EmbcWIKUzd
NkoJGR/t6IBHI3NVLtaGSaZz3g8boiAt0HmTVURkc5NS6ZGEKoD+mKLu6oatKcWhyzJs24KABAYk
9QqZJDfe9H0hxcZL7Yh4N/oQtvk8xO0zorfSvguRJ4AZB1rzpoyuyP3XC/IIlbfZR9JjjnFvHXhx
EXWUuob4L+bLQz3xmw5XsJKAJqqzJP2rPkFIzBbQXWdKlLF4AzENOap/Uvm/KFgw4K7TGi0hTU8g
IK6TjDHOwRQTrZtRP834IL5dirKZuYRTzwje7TaikQ5ljB0/vK+aWJ87ZMWn56JyMifCWflwNilH
b8Fmk4Q6zA8OLVusDl6lE3fM0LaatQOzE56fSAuhcW/QZk7FcGmU6GDJ858d4A4KldJRVxdl3gnE
yxSjyMrI5ENOcgOcSTbpQ3dyUtNT/mBdntD4u1sFtAVDvIr7NqxGg0PPvfdPagbXlR0LuDJR3iRm
soJPMwFfYyxDCPHtekp3DZUcukH24kdGuHG/tpE+d1Vhj28VtF65KaTwazKFQYTNbMTSK5/cDpkQ
FyBpOxXlbMbRssnkI78TFnt5znXoSOv6+Da9mUnXcA45ZBOrcMF5IUJehOewHGuzj28eIChfvFdr
dyguokzYZmR16iAHGrmxZzofWx5L++JKaVIQ66sBJg/t6l7W+8HjXJSzl9ZIWS1XENGm0KFw+bjp
ULhi0p+g2in4mCCIu0CKdx3TL+nClcypbIVevxwDwDdlixiovAdcFM8a/CLErkJbdDE/rQCv4Lyc
MC/daYOXAbo+XxiAi5+sUnyMoKULiHSJ8w0pdI883svUpWXf+/yTA/lVXGbGJxFl6t8nEPO5d5XC
fQO1jvTU40Zec/bsYHK0gSmv2ZxEs1+32K7qEDUxJqQpfk51B4O+3BpYke8MMFdufCy4jKFnEb2Z
JgW+b5ztf24BI4mFm8lOlY531vlSZgu6tgJU56WAtJcjVIMVAHMclr8zmcDxyl5yyHhujdjbPQTw
NDw5h4YMoxWi8gFOhaOckA53uIixWFJKDf9RLzozPf3Af44f80Buk12CeRx/8CTqHXfnFxzrsxQB
FDcnh+PhJPUqUTqpaAFEv9ai7jNrC32FsnRn1yJ6045hVquUgZzoRNmbDTLPQ9D675hTGrmSMBVU
Z8qAMY0cEsvDLgpFPscMicRJtJ2+KiLYwIHAi2FzupE1+DY0w+VlksTyKEY0xyHsSZsD6pErzwk4
rLVwm4ZoXs7CZ0BLbDZaO6JwxnxflZm3P/wRa4wLOh9PsXIEs16aGQsZx9JmSi/rB/ZFLBAh9Hgv
64F6vKI3yhyYKhT+/hNQYXISvG6ez4NI/smipO+30TfVTyEpu+jLVokNDmQM/1meyOpd9uTVuDUN
SEUfbnJ61pxadX+dypkKvPjLVuRJJfRhlRMDI6S9n3cPYwJiYWMmKKBO+Zu73ib6TWRxfZi4SC3Z
uOsPVrEnQNdorgSl4w8+zBqC+VE/53wOoUutHrhJLWZFMTxP+09XyVr2CsLugJky9aNYb4x1ICzi
gCWhERewdb3mk0AUr7D0Y+msV3Q4OTf85VK5BlyzpS44YjJH8ZLvkIQGjvZaulNVyiWF05IwFH7w
OBlUroCkh+3YmrTJ7mAycJNKzY1h1AojpT2e1U4H3gdIgzYxpUA0MXKPFWIa8MMlnzxJFYKtchKa
keig1SWw4szhVfe8uJLEXskxeTXMnP1Wxu3jm1lYEJ4YTuBvST02Sj0oD/XIHzOnB86p7jeoCHDo
bccrSEO+WHjNWkPGRBzoKjk58ShTJ6v3Rv8vkiATWQe8ItmsNLGtLhNiX+EkOuXeV/jqhpuY+e19
5R24Lh73awQlyqH8fSK5NZtnas7IKf6qJuB4yNHsEgkAYsNDn3HW9RaF6FggIESG2kpyEKuEZx2y
eQ4ReE2WDpYI0b7hUM9r6xOfef9HLzo/3Po2v40MeDOkHBCZWS7VbQZFz1tgzKDdxogVSFROGC3u
yQl5um2/ZaRV/ryJVjGYS0vO7sMQV1mJCK/q3Bfx/a0dbkXJXZGmnWdS+feG8yshg3o9n4tvUFp1
hl5Ka72uK/ouhKJauBv4pdeovYh8EZ3Wjcvi7CYzgidADtBkYBYZ63EJZposTjJZCUr8mgRidTsW
5UoNqGToPuR493aNV+ZRADFnK16UjMf6ih+q0plr2v7eupn0HCMEVmFh4OThXMgi/5+zrgn+UXNy
qfSM2NGqGaU1ywwg+9bH/J3jldPoNn7gRL+HPM+xl2xxdh8haF1KoQo+aEFLunXHb5TOBspNMSB2
UvBARvQS0Ejb2Tfi+VKdTqFnvdM0sKTpVg8jO8fqkUsRIyLriHqmO5R7XUSe4u1QR5lMzb2+UTHH
UZcUdnVBvD9ivRcV96zzkj6m0GVfbWzAscjR5hZdn+W0QoraDLPm+CtlpfKJM2xIwcHuI26hhGmH
wVVBhgyfr2xQNXaeN5TFjn8nDsBnVYW+TNegRz8o4e9pHCYrkDnJV2IUcAmCQGAZn6Od7NTFcEW7
RTwC4Lt73qTPW1cTxd1u/pJHKNrSE2i7kMe357tqTYHGXnB0+XLQoOLHMZKFf3BpNo/9ZcJN/PW+
SN42PuF+7YNRGGCVaHXEqaKpvw3c7C/xZYv2mfeXq/b7QYR49jmQMqrkAIOeU8TvKYy7PF68xi2P
lfoQQiysIV3vpLiNz0rtXBrhzg41EXAs+SAXYXNNBKrLBSF/xkx4hqYtD2rGCAq4lCkuPu9ekQDB
EdGt4m3WLbtbtkjZUMQYxY6574VDXVcrqSN294/ARuaePEiBX43D1/PYYQvN5vlOvSbPMQFnFIcc
EcYzxn8NksZW9mLMBqfH1nX2zuOfiBB2IBhXG6pSVdSFxrghJiISQOinHyINJ/q0vvEHmjwIghf+
v0KCHHwEVboV31iSEwxIvy/akaUL+R5JIEZXYlApatSAPBtbW3PjaAOeZsOvcXMWoSar0M5CpkLp
9Ov/t92UOyHEzawmWbh+iH6tMgjaTqt/0qlDTtqCswrBR/MCG4kbrwWfIegB4QX3QL/YSR5nxv1b
+8k4Bs2BvXRBJxyaY5TmBsaUmMjBuvye7d3Fh4PKwy45JI+uhC/bbHLeFqSsaOzF5ePP4/tLDEP8
5EJOgDdqcTETCDF3F9JKRqzxjXHWshJi0H05TJOye/iFjjm5yM1eu/bEEKgvjjyD4RCfitjyZ8QS
dFfQ7yBCHKlejhavdanV5460VP3cu50ynIYVkDxRF14VKPFImfAFFKGTHHrr09qnEUpRtl8IEMWC
p1x1Lz90s+9IZdJNbA6TPctrzs28cvJrqGoUjAxLN9O/IN0zgFfvo+Mg4pupfCCb22ibcVYdfU7t
M4SCLwbwuPbn7r46KoXXyy67yhmvhWts5JkCPvSrbItpA/k6wn1lHSGrarARyPHmiDPYyTm0CA8j
Fm5L06hb3HoaOjZ4O/HytudPRlZS+3TB3i1Iy8p2BxfAFr1Z7r2C9azsurYIlCDrW7jhKgOOebD5
q2fT6K1tBITa79VdFj49GYw7gozfVkPG7PgYrZ1n9GWcllbwxTezGSytqX4yZT5UZkV+rgBwxn+N
ZzWLJDyLgw8+qLFuLq01pSiu8K1kPiXoemC/PhZGXCp/+JLc5ig8qKaTK6uXdT/YVoLTEn3FnPkI
K3qp/LeNqTl1/ZihknXUjVXeq0uBYFeRK6XcaMyu9zkChHsvmx5xrd5U4EQnye2qeTWGgWw5SUEi
VcId2ivJYF2nNMfQIjvta4X6IL3c+KGfJ+liE6Vnx1KucAAFbM/hxrC7GPwaIkOqn77wK26TsSJD
kicou3V9THgSfuL0Q4OHC3E93T3ujCjeDoIuFvUtUus+kPXvKFHJdVaRUcjXpO+fe6SSMMXFLjWJ
vr0FCrkuj27qq1XjjEsRUoHBw0h5ei2kfG+t5gtWA5+giaKGN1kG9a3nWYpySjVfrkUE1LSXocGY
7Z9Rq3kgc1V2M66Bge7PlqcZt3gSCTrgZx6Qj7Evt/ljtuGrON4NGJ51eEbWHDoJ+7QlJR8jpf4f
Wcqww4/DUWqrcOf/ULGlEY6MNkdX9N+a4aRzhvQiyeR4YMbUJXAKqBPKuhCM2jx2KyZXHRgbp40T
eaigEUNE2ygkuJ6CqQ8ygTC2ek956Wr1if4SLcEgBRDUDCYcIryQEHsCSAzI4rIR7pcWOfcTemhY
qAUo9WN2/O4Bg5xv0iewkx7xRX2W/WzxmFa/4qJ5ka7BT1LsZTz2AtX1IbdRYRYrTmFLxvu+faMs
TOoo/G5/7WxSrSs2tE+Wwk4R/Jd5ScSV834LbIVKQ5KvON5psJgF3x6lUUkOYtZZR/KE3YSKwMLF
1fJhft5YcgNbkwnGUg5CjMF3PxHZHVNAd3WLVyRw4x/a2v+xvNHb+4acA5wjij/3K3U6orJwTxVv
Lypr9/hLr58Qg1Km3EuV3m2pylUTNd+3K4SdF9ZYH5561N2yAVv3hoE6ib+KN1v9LJtAY22MKXee
mDzOwLPsqeaJCddcilwvifsduDP6bKgk8NMjc30EaYLy7bKimgfkJDtTiIYnZKORTf00qHnX3+nG
z+cDFJ2kH0i9b2PGzrErWaXHndySIIQoezkkuqdCiJiFNhUx+FmXVRvq59c535zuOlvKP7Oef6d/
P2+p58nIk02rXxOyC9jcnTRjNlk9Cd2LqTy3WdczX9xcreblBB7eNlf+BUEE2Eh2mRII7Qg6eNMe
apRtXyyMUb7VFJe0/wuWSUz2tRv8jR3Rj97i4OGG4ujfngYzMyNj6wkinuhllTHq9TXvIXwkBtBn
oShEwo96ZW8G/g60WXrq7p8bAwigV0tKCwXpS3dQC9AasWDpwGJ+9KsSElKqV38FLmeyOtWY6jF1
hhCWVGniVY3q7ynmJ3DwWuv/RbWC5MUO/rgQ+dKpaj/gYGaYokLlGIpPgMf8C8k2auJyHCMVtgSh
UQ3Y+OjRp1tt7KNycxbNnB+wXsHx/90bvpnw3bvtiJYKU5U2XrOEhZkHLLlDqUYPh1QUv4fS+EfB
dvilqWorLiVXso8a78iTY5mGsTGWgAB+ZCuWr22KhLWH86Im+alLAqfO/T8AQyvGTyNiCn1u5dxh
x2shaVdH2EOp6a0TOE66Nkd/jD/hYcfHqmFiJgdr6wyb+dbwVAwsfIKVEz37Xs7iasaYPBtHLRwg
7OzgUryFqDEdsHGucSGjoVC2uptI8fY7pUkCn/GdzUSiG43Hxl1rdSbregOHejPOXn1Vag6A++z/
ro99+43CHMdTGMUwTxyB1HFPUxmstgyS5v788LRPb8vuR7z6I+8qVG7v3aXBYNS706LnOJ0WO74S
fRmGsmLiYixj1mRaMzwTbAGXzX8OBGyjWwnefSqI3eUiAlBZAd8b0uVAEVus9nwX//1ZoTEaESMA
NiFkG374HCN+L0EuiECxug1aSZOSLPxMWejsDfKJlI0J73equvO0zLjUC4NjW/dwpozi6bwdJRY9
8Ik8VlzwRc2pe/PiG+bCrXMj7ovXawTCGqP/H6tyTL2D1Ce3BnwCLoLUIzYgReGIJeYyYkPul+rx
PqaTWDc+t3vtp8HGAQ4rod6wU+DInY2AnRMrcEMukfyEiH1ahMSo0PkmwlYDh2x+kGsttuXZ63Ra
PMJT5Ddl3jTuuAIUAGeVsQFYx3qesTPbG1snwWOuyjoQUdYqZfIRYzLJPPkKiec5wx7ZHpjwLzw+
CU4WwquHChuIf31YH9ZWrtk9Vcrf7v/RB5xw/A8f7wZDen10gXdquWvWkkEVspmDUKcLaflilhIu
UZsX4dYxMo78a5wZjlMRGswuJ29yHCd8b98EDf4pdecG6J+eNQ4M2JGHjI6RXkpglkpYjkME5cTg
YqC6XSOROGduMne2ggQMNN4Cq82a1HeiCZCRgzZK/Mm/qYLtG64S7DjPo8Nx8n4v5uaAE8wsWlsO
5Y6o29NyHDSIw5BoSXsB1ymqaYdnR2bbT0vxHcj2FoHfZMDNqrEXrt/tRoicZo1RL+M6YAlwckFR
xbYeT8eXXzw7YcyM3Q8dKCBs1TgIpfI1yCieyNJx2OwX76Nz74j/LdRe9gK6fvrxRMtHiaouaCbd
sQjya9frwm7Xcyhj3mW8TX++QPypRoPhVTex+MNSUOHFKec4ZMzrJlvVNg3lSd8jPrdfzEi5xTUi
y70JHZnBG5MWDb6+AW4BLhI2GLTXQ2O0oKZL4v+0bmFSHSMHmvu9AAfAOo1FkYu/GvaoFpY7spHa
DirgshdACZYuOh4HaPsvxja8VfJx4OnwEQusfL4JdeO3v+CXNKYQ5TND/WpwIhqqPGdbaJIMqqdt
JUats/AGCSI7IBL4tMYNFfDiUainahEqr36ELG28Cg67l/ZaI9xg2xGsb+WKQ0NJQ39L/YpdjcC0
7OA2oHvwUp093kPVQWIJ6owxdJGC+jXV236pAcf2zk5RKJPQktAYNE6cUmxzYhfNuo+D8XOVuVwq
afCP8A4DCJOV/VNaucusqpvzWIx+8OinKQg9dKvRfhbtQ3EafWwIaP5wLfQSf7YLkfnHDGhYggul
1dkNtPoqMCdNXMaCr65/VpwanF1yJIkQ6i4N7ES/lbg2OL8WvuUQArX5WkZFA0xQYLxBIEF4m+c4
7Bqq6Py5hwK5kEuqbnOXCYKDOJJj8fof1RWU3F1odUrxPpekr5wLK78tN/yUWcWrUyEpeoMBO2H6
1G3yY7F6IrFaiiNfDkIhL4ky8kdd9RKeuEYN8vVj81yYgH8Oa0WuP0p3WXK5b7MDDn3RuXiff9Ip
7O918RAOMpOcLniefJ9iyqe6ZUcqESjVXtgjuZMlPqqSiOJGkrI88neT/9HihgQMizTxOzyxPm4i
9Hzc70rN3rON+HM9bKdBovCa6Ng/UKYhOxbywETsSHykReVOpCKlgO2oNDMXJPtToVO3jCg9kRvg
3a8dKiEe3iZLWJd2+QYF1W960rLT9B9PPYnVwR2k0y7KffZj6rJgCZlFhvtnaQcTfEX+9+t32bPk
6pFTqHYrXKdQ10sfAakoO+Va2euxal8RGhhhbs027V+sTouCHBn7UTnt0nT/qkjrtt3W8mxPPf0/
UyFHnjR7ZhrC4mVotCE6LgnytVUsyvVZc/IMV+kDYQ9AApHxppa5BwX1Y7Yk1G8j/vEXFa8yGMJ+
xaOKjieiN7bdYjAp1RiCjzTdKeznO9BiTUOI6NRLHp4f/fJOhhHzM1VRP+fqW0uC27nkOgE0DXo7
5K8dA+PgU2nqDEZU4Qxt1lNg3J0Q0teU9tojJRON+9TYJZGiDQLw8/ki9wTcfmraisgfD3+NRUGr
5m8ct/AmBgcEHV/iXyFdZ9hk8+vE35RgD6iPkryU/bBH+BZ+hflmXQ3GG2kLHmL/AYSiO/zOAsT2
UNRKEPahT4CGbIi071qnxFE8wJA6TwPc6ANHywRsP9LXeHPT8EmyAVj+UxMI9l7/13KmrEbrTg0B
JUaD5lI5KbH02to7iwSeaY7LJSzRWNme6hOk/V0mGxPVWBgpFK9eDckK2vlgp1o1I790GbDyXD5s
YPGosgVd6vU5q0I+TjjdpN3gEdqdrS/ok3gFVD7wYZIsMB+Qi9PpurbY4DwYaLodGEc9vEhxu/+t
25Ok4JvRmOcCBxk4XOOnZ0mJ7/7L/cM2bVjW6J3XbwV2hg4msKtrDvk65Acy142Dk17LsuS0c+Qx
22tKm0ur7oHt0JfHbocTYyFEPv8NBls/Vc8y38nDmQeROa/TgVaBKFX/r/tHwueEI13crybZ7jYi
WKYauRaDRZix+OTFOYe3ZahzGp7J2hBcjsWBuEKGNxoG68Mp+m7qdEPv3UkxxAcQp1jW1AruSn0g
DrD6JLDBD1GudYJVLMxnWj7P8xXaYtB2wcRk5zRnn3gDX6001KY+qyb6y7he7S2mHyZ5BnCVclmD
OA1gRl5REa29kuhJv9FGoacwMmUIWLJxcM5Ijsw2yil06+EvunMSguFfCmlqet15HLK3INmcP+oi
Dh2/rwAzKl7OYBnkVxzqvfqUsM5xSaLhuRMhZvAUvqVLPd3cc1QtRnGbdcxkVZII9DqhBCcgrxUr
LEvl8BdA7hYizdsG3xHWdbSgqHVkdlhLZiXqj8aApbJ+LCrw3DJo/3E1+RKEQeR1Sptz9Z/+v6yd
KXholOS+1Dqh6Dco8HG4AYLFEDKDWqPvThF32G33Qribw5dpBDxZwpeLNGohPHm7cAcwAVxS/iBd
g1H6mxngjENYT1ZE7C+hNWg3MPgbJQJ+dT29p9RAu7Utv9SQvhC6YEZ+zjb2/kzp6ehmKWbfVg8k
/hc3icClpCGMGIqQ+FEugFWN0HdWeEQTaxVJyFuSY0MgkUPT/h07V+wxVFmmY5rsLdwFq/n1csNB
PeoKF3kz50K18IFJYp6veQE1F0utvGO2qIZtQ13yQm8wRsSfdv3rDYac3GbOwwAEnTfjU8CAxO43
vuDYhDlD+LeEIZG/cz9P2Ly6Chs1ZioIIvyjb7uoOypbdOk6hxZN0D/ae8dXevXJFo3cpi5tYIeJ
hKNJbuC0Ta5VgB8z58qlQBQPWjcBFzmyT3y14BQbJDAJfO0leyF473H1V8jDljZwu+Z9wET2zLJY
9E34hzK3XSnKJGa0e1DYHEbwcPM2L6lM7q/RQyTY35nFlS/HAGD1lTFFqNLivIo+UK7hI5BWbW2S
J1WX3Gq09LUCSnSm/n74tHsdKcS7RUdB+o26YwL6iwHUQQUPnjIxDZiqicUOH/RMTsewcM+Yiq65
i9r4od0vRR5woxVk/uJ0m9DGXQ23rt4ZKSlrpzG0+FqQz+8TJn3+Os6vwDtntFg+LY6/LN3s8u6M
0jTuIpJ9T2v2KosdNAN2GA3he0GDVoXPNc/ih9AnZRLG0XyChTZfLjqZQDqYT1DyH2JycaptM7tx
NgJXLGgWhCQEi+fkdO+1zpD0y76pi3QW2jioSqVLacZQSsHOerVRZ88RDd5zJbW+YocXnwwEcMgb
xfEW6T2HDNKTmXW5fTzc5GJ1dPLvegJhml0edoMgg0v1UYnVCost34xC0Fxkalv1ev0zYdOUEph8
DjrvKk7MxbiGvEob4zF4U9ObEnz/j0gbw6NByqnO6TR2Sjr5m2g+HHQzUco/Rdk0yT1M1sL76OBx
80X5P/U7ZyUS2JlGYDM9vzeaL12rcWL60ssALpU9lKraEVw9hn/63IKsNO58SmDNFv9cT1Y8vDce
nhzbxQh+1qrdJNOn4dK+BKbWKpGa+IM2WHZUiy3BgM5hWlw4r4ms5ExlAzdG9aaYxpJ3VgXS3NaJ
1ckwj1UiXONlErlT5f0gIcrMPmCzOCJgGIED7CX4uZAoxiHukLObWxj4UOZD7Zyu8FMuWj/QHDGv
dYDjeu9Q+1jbSJVJ+lrlfVFOovIgcJ3XPQ53tijOH8AkJ2KmX4fByPbuNp6jHEFCTayFGDUB8rWr
buznxoJhfgNcu0PFRiplbFyaDGxh0763VdtLcjiesH5mHJwy/QTV1va9cFK7SJDMCeMP8KrIJONn
r6+lVQqymlCj0FgCzmLn7MlQ/mSwI0rJPyiHAjRCEu5UPZI6LsXtVTUauihJHTy/4U2awhN8FLdr
TyYkVtcHwFAZXxUcmlASoBNgHoavDT3/TBvktE9324LaDkWjZsMcRQhacSXOUyXhF8Vi9Gb4VZ8u
VNh8En7Vw+SinAxzF5GxC/2I14UTwN5dK8mUnGA0ebCYvrZvjGcopJu7GkdP8fP1uZda7dpXNIwO
yn6R1pqslZ+VgvscXBCcgm5/0vCp7AcFn7I+22TJiB+GSDuih+C6W4E7GYlMg/tc+iGBA0tAZpbt
kZGGI11imjxhwEDkr3+uGgzG8hxbFeqxy+bHIx1i0J0q4IlYR1+WaDh+huuqxPh4y1b//+pj9VFu
MnVcIZ8cuec5h5DQRPIRfqaUuqTk86No/atFY1CiGgIj6+UvJPPNnU3rysJiZhpo2d7YNh5luuJi
RXqTErmDgbTwgurEeOxP7BTC0JC15wqJMC7vo0Fi6dCCgPWKDy6+cnTevgAAUPy3RwYjjEv4tbXf
d9hEkye5s1f/fdzwFYvSIkMY5ofCcKIWGSBjIuvKEB0qBW31DwbmAFwEpFiLWI7sjxnmHTM5CmCk
XgvUQAO0tpx+sKw2oe4MOn9PGOkH+VzooZ92flr5ABYBXguGNCwahb3uzZn+4uNPpoxezQQcmsxv
1HhSjyUzjze1Joqc4MVKYm6hrYhIUZMaBn1q3pYDpkkoYar7v64IOj7Xgw6H153W0IwYexFC9Jhd
7VwARr8sa0+zkHmLbnWtHt9ki0UI+ZIhrAwaJ/zWDKjW+3rmjCUImCdQ/Dq8zrQ0ZFaFI206Mxqm
pcddVzL3AAsEz8Ic6hYcVhs32oFJ5tQCSxjkaMFRu3nZajWys0/fUonoKccsrL0fb4PU4EAybo9M
Yi49RWh9j7enk80GSX4LwAWI8YHES5qflWLu/8WbFnc9jbq58X3uuojBoPjUTQie/uCRm/DEgDpA
oftaN/c6jKcmb6gAARcsxbcY012lTidqj1zHHEWr3cXMJuwdjUanOMLqIXxVa0NkDupRhTnzyWMN
jm3oAuDHUoWv6dYHAQd5fP2Iz68omuf2wroQWvrNCTY/NdbT39GrPm+mGNsq+0d7xPXfBtEsHISx
tLriXe/zWcBuo9vlZii7OsvOjBChvGglAWe489suV4da1vlWws2MjC/FO+R6YG/u2hsVgVMAzLm0
d7zGQlW28XCWubxQP1Bf7qKduNFGpAc7n+GnEsaBFy9qK9pVyVcHpEmmMdN4UQG0DapmKPHIWHGF
QG75ja02wfP099Zpecx8pIK6UcPlgnUknIrBfyW3e0y7ZorC4rB4fQjcYc+o/iL/WSj8CUpshn3T
6TnxOHPwWmT+uRoWnd+NRhQvKLLuzOL3QZoaqCXjn54bkTJOeKcATY6ZWFdVjw63+c3H7zoyC1zN
WIzIHRDb3jNgMvjW2RTiQ01jTnjr+ASvVTr6GIP4n5MHeVxKtwBvQhLfS5lMS4hp8QOxbuKQxTzT
PDFUxDwN8plB5YstIaVahtUgPQIfeIurF3tZAWw7l9JG2ywN7QLSQBBKWn+wZ1zkfCuwQiMROMWO
m4BfWVOkVFbPthuP3bri0bHUZVl58mpQUwYYgPrbr6dJP7BhYwQuVPEWEhP2RQHW1utwf32zELyn
e2bGnk77VE/B8AlA+Vb6f97NaUbEWbJDqhutM7NB6ZXA64jC5UenGRVp1vgFVi16JUtnQlDiSCzs
HI7deF6dfhMpSD/C/5h6d+PA23yQa+XZ4HWjiiboBXEdeg1OIzZz7V7Kpz3dn8UO2zFYO522sA6+
4xiepiCBkhqL+kxBGbIrsUH5D25YJdOFqajbC1EljbNtWLyzIifTukTCxBsJ/SSJJscvjnqq00e7
sCosKWjTrQkSaiRZo3GrgjaWB4U2/SmPz7mNY2mccirhuu9q9j370IThVWLNcnA5koDQ929Dn78c
RceBm0moQO6g3VrfFE7jBOhN+rBk3LSV3M1QHUgUFaBruBawB3Lrbnm4KmK470jTLlCYAUJ3QRb2
UZAkfsiSGEKn24hkhoKYhz0n1iKjnYVKHOmj13CCBge7R7DJJsseapAXrzveqv2PSFGNRmS44+R5
v/D5ESXh3HPsVU51AWihchg9dIQmatsMpBn6GK3t0d3nmEJuIPXagD+mczy38OdGg/0OT6cw0VRG
LDZRzpJ0ZXjipOP3kHB6aKPD7mgUqJ4gOGUEQd7YR5Rzc4zFBPcybNYcPRkSky+23eGcnUT+p3wl
88qWtK5Z9PrHSymTsB9OdY/kHTr7mSHh2W5TiGMtF1FAhupc7KhRlw1TLj5Z/IULZuN4+13x8MdL
ZGluEY4sNsGbu2LYYtTWS59cQCgqptS0iBnPTfTKHEeoxK96cS0HBktSaJWtJx+os8ORjZUu/Nyw
OQpJHpNfCzYID1uWizJ/FqrEL7NpPYzdmCPxsa0WxcUoEjzqV8C224APLSKD2q3pIN4OGhqKayqq
CVbsZ0IECZyroDnyhmTkGn6uwtS5n6YT9V+rpOONRYkUEznNu/0qkULmo2XWb0L6PHPEswXILjy2
P1F7qJOQQQKXEZhw1KJalSHcY9yU5y4ICuuoYVraJaeQHYB4Of+t2DkKzZ0x/bI6/kS29Upi/vqe
GciyPL8sM3H9alL6zduU5a2x0CijoNr0vg2fk0a+pFfHsmUzHGqNP0gQYVYdglXKeXbAw5ZK2ZSo
KmKdgs1+r095bqwiG2fKkafBwmWizReKGCDp6vEvCaNvk7kgEjLWZAC+0oRWXus1qbcxvnnySZm4
0bkD2BkTEmUO+Jk7gppzBO9yKUGxDPrItTGRuQvy3C1hFsKB3BgKwzT5mA5NiIFqVjaeSc2oGGXd
xLzophBu6Q0YubH3s+DkTnqokms7F6cwtexwWTlk52L7gMUmCd7eQIlZKVPd+1a/BVvmIckwlRQJ
horzFpTZAvCTkYy5IQbW1qMAcdIhfdG2Da6jxoOF7KqCntpuediPX/GehXUFNvceXMlpAxOeO7eI
qpcVX1/6peLiFBaPZ7EVDg5awGBGrT0Q6KJM5MlDxHDeIiYjec9lhh21jrvcDRi8zHudApfISuCf
33v0ncYlYV7VF2aE1FqsSl2cAyKxnESap20ESSB8DQbSeCImidRBBCRo1eRIQSAm6zsPo0ihxaXd
jU5p206K7NjE4DnPKY/OAZS3oR/Uw+foxYsfntxFqyp3G63hK5ZGtqETpw9+aW6TQ4KrBSVOwCnV
a4l/Bxqb49ErG4Qrxi4Xm3CX/lmyx9lEJYsheKT8fy9IqSZkpP7v+fg0e+EG1xtBTZLzIlF0VW7j
h+QdSNyam0jHIozhg5BZuR3X/F6Mf8lmmjkzgMyO9KkKnKjke2YlGxt9nKZTfLUrJZkXPD8w70F1
aPqdJk07WEWu0M/thqGM3VSKVKO79CZCUNb5I6XoatQ9CZsuSVxhyAE4TsKNX/hpWiA5GtZIOtVP
Hpy0I/DlFCBPZI4A85CrCeIMixbNXn19Vhqowb8dEwbEghldcDpT0yvYYNtofOIumhIeNN7ARAZr
hGKCIS66/Xnmodnr8qjGueTKH3UppZ1gU8cUNedGe04GJ9hZrhPy4tHjPd43Nk6T1hJ2ywLv0Vpm
KZUXIhUpp+7hQK3OuPaRqr6Ob5c5Xfslfh6aENXBjBqnM5nEWkB6wmZKspqeF444dgUPvBRV11kD
L1m7PdIN/08jqSpsGZP1mAe+EXW4s9s0BnRsCIOIjDy+hWFxVFLetr+yTOqjzLE8TnjPoZw7k3F0
TlXAE9MlnVSWUy2kULQWkhQeGJ9MwMo77/wyBCEmXq9eKN8rk+qSOWRt7emJVDwWriDplpl3JqH3
y5as9OX37hSAAeNp+BzN/V2s7Eucv98b6+ZlR3ujgIH2DpG0QW8Ki44MD+DkfgGRBpCcd+WGn9Di
hOnkPArUfXfQmtFMwg1miNIEy/IXKptj+u5JplAkwS3le3DoCMEoYNAzUL07kpAW+Hl3CmfqH0Sx
tBiTb2FNAN0ackhFOhY8R1IBnkKLhzmbMgVkGu6Iv4Vz8vboz2KYFZwxIqc0+q1SMS6SfcTZ7sBP
GRvkxKSxIsxH+qK0IdbNv/nFZM4HdLSPvqLQY7KjQNZ7Iy2p22lBf+Y9zH5Lf5Yym9pD9+gPgtzH
Fcfefu7GLihzqzUr7kHg2PKXAUqduY0I3+lY9gdxnAN/7VHkgACEErP35U8bXCuU/ZCEUniJ/cax
Qt4G/FiKNubJ0O4c4UaTfev20GnVu3i6zuJt4hFPRJuMPc9BxNq1qET8+fGU8gk2QcpnoLofWtvL
CxvZkBuVuVaFhnt2FJ2gjOsWWhCWgCEyThWCW+zJcGFTAoto39KBjWcn872SgEG1/1j3vswQsTi0
a89M/F4smKsZQzp3HbAFQ76A0BwmNmvpQ2Sy3l0rvt5k5KHXHqK9bI6xrGl0JSbtpQvyAUO16PJx
KtN95r6KY5XAUFEdwa6DuU/QqecyGRHicJy6ifyashfH8jKunUHpiW49IzkXStgQWfteFD0It8wa
X/TyfQTiGR/UPiY6SYhZGOYYkvOAXvROJiJO24vAIzZMCixfr3IkSGpNpHvE6XKyv1KsPj/vHv+c
AmZozYSi9s9ng+827+OXSuzhfcAiW13Y9c8hjCy2+e0FkT4O1CzPwDzssme8sTt0Bdz1E5P1Z4rb
IGxzAVXEU8kBF/74xgeWIYvRgSCjq7kRI2gcs+uBAijKU/aYr1QJ0pbRGm+LbDX0Mid3OgV3ZJd7
WYvoZ3uS2m7XQ2JDOPNCA2ohj51RT8GV6V1lFGOicZNa2+3qzRwnJPsVwG0sHSKBsdpnIugEvvlX
v961Y9mytV8UhJ0+1SdwpbF//uATeOSdsJHQqxsKxMKhIXwltwvPwL1iZvHQ8FvFeaZMZKFACwxX
Tj89s8hWuTiDN4Hub7FnVRJjdpw9hw8giaqeSLjd+uOwC//MXXCwqKgcLp4VsGaaJ1/0qsoZWLEp
IFOFlgLuOh529IP/Sxdf4QaSHpC3MNQTt0nGAnAYaOa73chjoYzCsnK6hLg0A702NvkTVLnrdxqu
YOt4RukQek+yoQcjiywYPQ8LM5tJyUx3yVfQEUxKsNB5if57VVtsbm2Uu45JeWKFV8yMX8DfjUxz
hvm+OAIYW98vg9SpjHK7Mao4l2wRW39mrM/9zU+7IsIGS/r6VJbd7i+s7P5eDajE6ByLhc5HKEA7
oLfpIz9L7P7fhu0oHNT7XENzyDVcFdvwpnteWLM9qCv7QpKgt9fk98bVyqYrarrmzOOeI3vdNIXP
igb37r6aVev++SKPVDLBkjabl7ZB0ja+zdWw7J7a3rSe0TyoyHdC4iwDAZ1X/976Gj8qGBMNtpCz
VF5YAHkVZtIY2UeT5JnJ1H833yNA74PxF05UwpcvwYt5rXQ5bHs03OT4GbARRH5VxevFvPic9t0Z
XEKO9XArJy1maHbwkJsAaFCq+wjyxQLw3dGxzlmbsjXQEj03+nR75pdE/xo/9YiRLS7pCmjR1g8G
zQB7Np1oCcDqnVV8bWnKVo0p+FRhiSQK3nQVzbS884B2nKnjjZCnRhj+mfgg+oQ+uggWgTDVmj13
P/+BPqm6PGvwQitJ0SHWugCcbnxivWzVGHwrUSUobZ3omPDiNzjhAihgihSHd7Gfl25e2J3ZFDat
We4Rn1SBYOdzjUMbH8TZZ9Oz1URtDrMSAtkksLpsRF+ox6DacCAcogwC6lAiFMV8dSmov8NHhKY4
HndF3iMnzLmkzCxnmIggcz7LtZKwAM3RqR4K/0U4z2BKRQh8AMfsc3h7AAPd28SzBdDohl6MMtFD
BEO+FAHBhwQzK6f+uwZhTTOd62Lbi4HjtBFgFOjS+MMcEuHlhVRC0/GCRBSIaVGr+3q8wV9eGCU3
p1P+qzEAlCYk36i0QwvK0v9WGhjO2mjsduajXyqBPv1EEkfwFwgjMHde827KzsXRIssbV/NPRhj0
k/w3pCSvFbscwLgDHqCguaLnwiBdy4H79BGr4wqJHsrsjGmY+nG82x1RmvYL75Kra9kAslEsMVWC
3krDESagPyVcSyo5AIyXMyLTKElffw6rFOllUdTb9fK8WcIkbyVm+SuGHy16f9uGWsnO5Dgtwvn6
TmLugYHyLn1KQnvx1IeOSKc6H+iRvkx35ZMSVQjRjIeLzBTMbflANa9dKQCMPso5zD+gJgvcUp0s
reU8XaZHAZQoVMy+WBKA1X+cV4dlDaRFJSQW9StrtsWtV5tAMhugZp4jxmrSz/ngAZKUHo6iZM/Y
82XZwQOApBBWFxO1Iig8Y10nLOBBxxBAPreFAM+AyWZeFEaVtRWo8eiQHytFzC0N5F61HAcfZhDH
fCVtaCmOIpYc5UkART8hpBNOiT/ZhzsmVygEJZ7yauOvaRzVghCmR1vFfD0x9zdgo4kH3AfgcuqD
wT0l65C8opjzirZKbXcGwkuo9VA3NxwFxJI1pQwSGZYV2JfkkXTa1MaG1OxaXD9FwIomlWFol75e
N5J9ddXEhlNYI7O/98SgXmI2f6ufwrCrNejCmhT9JEpUdw5H9JVBlfjn66anyYeHe6QSJPnKaiol
9QZ8CSEbhwz8FBCo3ACD0OHaei5N1oAM2c9GPRP8LvgTBHtNiKMTrGUaRp52lfKPxSYXtQuBsCvQ
3k8HzaIS94JMnWSOAdPP0ySmW0USY4lDrg92hdpTujyPPbJmem2bgHl/BeeYR761JlpknJ/4cxMn
wKbm95/hqVWJ7+CpXQrJcQxdWWYri8P0nYwHhWbtiZh7lzNIuCu1SbR0qwqKp3sIXJEZmdNW5feT
0YOBcq4ZQB0sYQmKAXGSIYny9MhPXBddbkMJ0XGBCC6ZvGCTMgY+nNkC4S8EsV6yEi7l8FCbfcyw
wglgqcMaVZdk+8jh1A2rvUkemb2W1dLE/Gn3dMLbrFzWMrh9xMJrykFSVLobOEVok7HvR916ZU5z
te8lh1DHuf0GGIDsyPVtLmGBSotJBeWEPk0Uxh794X/gJ8IX/rkwqq7zSYprKWFBtrjNV7ZDnpU6
auTp1wOklWvEsCqDsa2lFG+WGCFj8a1dUSHvsDMpG9NdoGKgBb8s1CpGE3oKxRav2IDrFSndjxjY
sEfi8ge17gYcYVhSoa7j5N8uMDIu+3UtZ6H5D+/r3S3opUGCsiLiAxuf/ibhMymwd6VqyIh6IsOK
Y0p2xi3snF/qEzABFDBgFCr/jdj+hKDvtrxNVuatP3Mx2tjP/DU28z/RWQsYBIjvQGWAZJHNWbt/
qTvyQy1HOD7SFw0yGw+cQF8XKdaVmF18aW9O1C8TQVqtfVgwD82pJq1EwxuZII4cmmdZUa1LA6ee
nRqNuLcBy5ZZEr7UFJm+ObjDgtVb/cy93Rm8UKH9BObhKeVMYHqN2VvsVieAiuZX/be/rC0qEX+9
5xHK4yTjOJ69Fc4Z282fIr5H8NratJ4mg1RGEsNBSA7w9QBq03Qau/g/R0Y08YFv/gYLIH5fM3BQ
mtLVPIAN17reBkQaWa4VdjLuVAvSof14GwltGwPDGt1W/Bj+PdbSlMukoTId4QypNKmF/287j8pt
/7Dp+6XMvfcJLLSIcOGK1UhDKJRRm+J9gqrvM+eOxTIymw939scjd2HNZqcf68IDoxT1TzIWj3je
kNiN4w/+5CInIkycdE9dCUa2BNW8MetK1tfzZJClmKkv5nMiLi70+C12xnw+63eL9+5ATXkCvIwI
d7nKA2iEmb1L8fit0hf5np/tczm/7SGnVHvpELApoeSaXzunC436oCPo7UAwXTTzY13S3rGAMXyD
T6BW8/bBvMAfmzlbJyCdey8hxDj7cP3kIMIgsurMyOnwMyYKN0kh+NWTlju9uWCJk0eKF+Zb7bbW
MLi1LU/arKYWTpmPuE2JtLmF1kWBL+5/1wwxNPG+7OWsJ3XCm1OAm4v4f1sAblU+mWYeNnAY8uAJ
gYv1jATMuxk8DRtNEpZwkDoiyg9k9mMduCiZfQCrKmFvU/gQhAl5bH9yoS3zv+rJfgD8Y0OV752E
Zxc50Llc09pDcz5OQjaG42X1BJk5B2hY20jIztII1qidOtMUY27r0DuFZkdCm52HzpSAB4LaG9ve
nRtX6nwRoY6BFUZbB6M5ySCIgM58xNbrTAQicYiQYPXlebg7X6miQo/exgYS5Gv88Mlaiu7bsmU5
/AWXlnA34b99aqp2c5dlkjBYQx1wiw5eqX6VvlTMr5b/1Ap+saLnbEwnbwFXk4oPoui3F2JDMZQ+
5cFEb/e6IAYdVAoVMtIYuOYO+K6Slue6tWHt6fGvtogBrnXxN/FRV/2LWOH00H7bR8JMDJnaV39l
aEqfkAaXq3A//sUKguCCnq6o5L70zCgaRbF5fk9vDkgit34b11XwMbudVGAEXAtMXzEvVwxwGwOa
jvwtOaitRRBoFvCsH7iGxJPmzZhp7TcGYs8Alhn8sNmkj+v1V6NqbRA+HxWbYY6FDhDpcbw+/YVV
lupm7JIlzrsdcXUAWuz/mXRPQXiisuv9+1QTx6q+Au5FYohfpDbfZixxjYKTYSw2RuvppDuFr0pp
Du6VLC7qzREW9wP/C/+xdfYK8+ysWGkqgEgziGnUXpah2G7SecRP9DjOwT419nrF2RMfFV9nnLaU
HAds97pc7JGoNMPR0hUoypup9MQHjY6u39dZxsgWTzfi3bX5ejAEzMSWOc/4jUWZtYP7Ux5Vg/DU
bPL18BujnT6b6FWgtmW+VqwgfPAOH1oaGsYIJrltbGEKz5j4Ipvykm2aW/Tg96J2d83KJ6BxX2L7
kH0R/27TwN78FrmOBe4tmeCymFp19NFlSWdm7nBAy7Bnfrbe5xktn/c6q5tKEVqEeT3f5AkHVnuI
OkNb5wCSTPTDCejeLL1HgpcjT0+AYUOMHPHnAyMOGfnWNwJG/gP3p5B2nqC4anaVP/AQI9ugjpQE
yXfgyJPM6n4G7CZbVkJaq1AOZ235jSf61bAaQQ9V5/y4Z0iZGvVrmk/8V7jLY0/QJScdvToc720B
JmRF+YBWxPaU128mDG/0fzO8UnRxNPeC/9cRX9aRAGtykdr+f2ZJU/Bsev50MOPefrT6Bv8xzkoY
+rdlq6eLOgm6UI2byMzPrWfKcxtqin1FHgxhd5HikU6o5UGSMYjGxJnL2KFgq1ZcofyhQ4uiSh83
KNxl8XmWMgzPsV3Kuy7E5NFy/BNa7XC5lHXe81zeASB2dv8y2EyhDucjXD8VdjYHavfMtoVLVbGR
jjrYmp0BmCSTlj/azzOR2179pDNJW0Qq7ianTE6MZ1pvfHqDvjWyEIyte+s2yDe0Ol4paQlcBJee
lTGN1Yp9CE0T65cqdJtL8Y+tIa7lRoiyNf84iqT5luguXYFaUrvfxYFhxBU8qfLGFYfc5OOeI7Vc
j2piFSzHzqQmGgCZzUbNm9J0dZvfNCYFcIplGd8ntJ0ZGy91jxhrBIq2Tk14up4klm7B5+gmiTSO
ZXjH+qGgs5YN675UxGUeXBciQ+LrM/pI4wxgTkv00WwDcB2q6Sh7DqaamXTCWGxZgNV4CN7M0hmI
nkLJ2L/iwM8rxf8Bbpvffy9EXMr0l2ok5jcAjgxwqNR+/lR3QVLIbsMlrVqYk/lDwfJV9Pa/MdbH
WJyv7GrRRDecm2GF/N6P++OymgX5z0SD09Xg9P+VCCvKxTkKx6BExaNDwcgN/mwSytt4AUxiR+9I
Nm7jKgqCsoSSiHqSdMff0x553Ba+JHD2XmoA66tBKMeyDlMJsv6Ez2jUZRx6zJrWA3+x87aSrLIH
e/xSRYCgoNoXIVImUrca3dwHwY8z+HYRsj6MffDFBxNoq2aY53CiYa0+SqlL4noUcxBBGOfOJWK0
QFAZs/ei+GS1LSvQB40lqMExDlcTgvrHbNqdSaX0KrsJny3pCk9XfaO09AyctDjq62tUs0cLDOu5
IbgtlkRX9TpDb/4ZphYONluuSE0w1A8uC593F7M/6RWYPkMM2DOzPjjW6ydYKj3uMiPOT9RuPRxf
drO9haiF5nKgM6LApBVBy/kHnD+GcnFPM6dtI9lz7dm47kj8IMXgpeJ9qvSoW8KvYDkdslJTr/sU
pf27qVcHYZomexxwvDrfTPAqcfhZyV39sWlmP+kbqqbcT1GqezOnJVK66g9A3wvcQ3k3IkjRc52s
mvbRdZSResJfMNRtCrLBxTiU8fpxuJ5M78KM9snMhZno7lbzi9evsowUto+MZLe0vC6Uy5NymCp0
lkhLOGgW2OcboTIv7XaDoF4xeucb9F5W98NONvuoJ1oiivha2W7gl2gsVA3V4p3m2jxAeyOHxgGV
mXDvIbVnnmAEFPA/YmSFYqSvnqAesmHPRRxeluu8FmSW4nGdZuxPdD9sYRQLuw1jh4bVDZBKMqdp
68wLgncMvho8Ym9cL2/w0oTxU0qFefLrH06/pmrlGYaHz3nPFnqEiAHzkkYOjSsqTwZoqlDKCRIi
DSNMVyJFJlhf0svfrF2mHFANgHNFxZuMGMvRa9VEWEZsm1FOjX23iMIxB3zqDWnA6bhO5UwsKOsd
KFXzotmCXh7dPc4BVR+Y/GVINm/LngYhGAjse0swxkSGigFIh6bZ2472S0AlFSywaSgl+/Wrdzqn
7OfDze5WUHwwGWmqj7WThiDrfrba1ukOXaTeR0am99DuolqSfxQPdHItepEO2SrirPxJb4o8x/+H
ewdaGLQPJg1ZcyGn9+BfBWeupS1rXBpT7/W1qaD3dU5MRWMvKDWBAc+MhWpoiSwULjjeBitXCxa3
2yswkWk0OtmaJClZVEUNRES3wlPwEZmnDFu/CremEhWm3rqTzgV/itE1/uS83XKHjaZcFZMs52Ha
Xe/l/yvh/d4S5+Nnsg4sJjDiwXY7fxgVXd2aqXMMBuVL+DUHK5na/JQQHTuGWAm1hRMgVeag2e7x
etLGJwYAd6FX9c8+I8NUJiyg4aBezNdDKlPRDtZY3pasr2gcc2O5cuJcbCLOvDPijK8SMxBdZLav
6e7Ltovc5LCn3SP0exn1x+IrLX0ojqX1KSQe4P4WQEJvXrCXlOXK6G46aA/cykLwIdVUs1wnAVYp
TsFbg2PyCQ+76VJfr+W1q6WQpk7dmmiQ5yI9qZlUcHCOQAiA6a6C4x7r4jARvkm+3QoqPCbIBiOs
qnDCTDU9P7OUS3GAZXpmZlyDWATEys6kZM0rBiW9LVod++raI5aqjRLx1fA9S3Au/LZvUGNmAGFe
3cGudSMY9gq3A37OqabZrUIA4qx9tfYYOZ/ymhkhXwlkzVkL23TG4PM+0XgDSBxLw9V6zfGr+ATL
DqUW3h4BAoPlgZ5nB2yuEw4oJthPaS//gXwdz6lih+SwdylvVb0cya7Wwmh2cRaX4F30M2TfjXln
CFivJO/Eap1zmkVQ4IF2zfYv9PZoZNT4/HPcM3w8jpFPRaP9TL2hR3uA4cwoZbXp82tsJbtZOW4K
BU/jTGVnAJt0cRO7INzCxEO41lGEpX4n3LEG3xqmdwUxnM8LZlI5+nvbQ8d0tJckN/LqVsa6gOrk
g0pbI7yiHA3YlUvCPIZsuSf99vDpZnzhmGafJ7/ZvNeQ2MNB/Ija41nspK3phXOaJGR+zGrcvPDc
oS5TDf6QqBKoZVlOzi5mr1BBSR1kyvxs3gKDfBiC7aV30bCPO4CRTwC+xBCYL/aDHv0W5MAYrq5L
3azsmRaf+07I/W98Cc+kkRLyIxlwPRJQ3lAM0l8/TvPnXDxsm3T/xXd9of/ov/kBVLgayf0NIh8t
EXNki+ZF0Hobh65Ra2FAMuZ/a3uvTIrFtTEcyKTRrtGPJeascpqEfi6wHktLT4YpL+9PNJwvffmO
rfU1IK2WCj7U2dE7Ud+I2vgCa9VU5YwXoX7SUDYBS1MYKWArdY1DfKvIReYnanvZxyWOGYE8iGkY
1IjrTTaoYO9Lg9lhdT3jLp7tyDYQdLllCCggJkMTSfk5T96AV8wAXEq9MOpWt4RSX+0NGetkEISY
4QJ09nL98SfwuZ9XC2C+Qu8MC6kRWXvPdTsfqpaTEPVhVmZB4t6c164yc6M3XMqmqNRroDjhjz1O
l4Te2CMaQ8rnGFJJi6ihfMZj6GXRyxd+oMPy32HBtEtDD6998C2TVjIvgR1p4hWV/QxFx4RhceP0
jwjfRAJ2X0UDoRNrxrdQJ886u1eDx1k+sFmC4d+ZnxlLtXTGGqpbwfafy/UXAbsF5t5Up4vFr/xD
uGec2uLOg8/D3c1PS7FAxAOkBwbAyctx4mcFNHXSGGHcGsCPGjFXA24x0LNyPKO8Y1PtDNBZp7bo
i8j0sOwETM2Hz6lrfLVUzw+F0wrD4XqTbtazk0PWEwnhrmICzR/nUL1nWjzjeEzBLrimh6soWe4P
qz6DZYhAPyhKlFM3f3EIITnWV3mRwH1nRW4H4NRCNr1D5ogo1ss55oTQOgVRny2IUA9YThLF1Rw7
8W7buwO/xJgiftebyrweYBbp1a/J2pGGwkK/qZr/BQJUsFC/ZHPK9voYUjk23MbPpVwwzkGOpJv3
bDv3YHFWgeLeUPRp6CCL/QxbMCcifULv1ShlAOjlgP2DKhPL2SsHMzwbrxv2QaWNRGV8d6lymHg0
hJYzPTSPvuWGpW1JruhBkhrNSeECmeqW2AYmGR745xkVwZu/X1mBu0/LAdUz2K0jTQgfa22RyKh2
ZvUpVsNb9D3DdnqZKMFf9BBcr1CKoydXnkVOu9Atj/MEqinCeEHJWvW6tsNPI0kZpFEH5Jyv2vt5
GS9ZKfoazfLmagHzzfd1nf6fd9vGDiQT670xmkGy9XTgbORFOs0ZYk4TBF4cIO9fXBxZ7EXOkDmh
MFVLkqaMN8+1+IA+mmYhzfJhQ2van2uhk8CuC5iTXgdKj50gdVlrIS62sTmC5jaPGTwalGdOXn/p
pxDXAjKjniQuX6K9/DYOK043Z0I+MbJVmb+R2UXec2DJNpKwRAul1rxCS3E+BYUnmaSzjDi/zLwA
kpfvKNkSYu0LXa0/KBPb9YzbXGVXR6KHcukhgOfowqTACnUz+o0Nx5FkjTFz/dVGTH7vvOZAJGH+
cVq5Gk1kaOrszn6CyMWZuIx4bw/J9cW2jVUVKX6dOT3v3/PJSIHJzz9PokI7tpFQmE/8BklJ1O/L
raNCfq7/ftCZ4VT/yOsEa/g8TSr0x/sHuqECidxWP749R5JrYBNdZdqAMZVo3xA6bUy19fBGJf2T
a8KPVnqREsbm1bYqfwf+RtZxwCLBC67SJhW7LEBfvS3oEhviN9PX4C9REzytKK7/Rz3VHIzWUC33
WJphb2R9AZLQwMmstL90SNyWadRKaa04DQAbAkl9K5tnWDmIeD1bckZWBPgLPjoZSqrdc+99X5Wp
iQ6y+zj4ypKFk7Sq0IWsVUj4VmLs+cWaTCDc5XRBRZNHLg91SvmB1OEDMl8nYVYl26nf+GvIQDiK
G/9VvFzy1qMH99F7qQa2c081pkrD1hDo8bnHo9/36WJItd7fqid7+FQPVXtj25RjeInt8rHanONa
qK/MvlIhUm46cuv6GCZ8nzb5i1o2QKzVEl3zg/zixW1hmW83xgXthPZ/aZd+LRuVgrF45Pqo+EX6
vpsms6pSzSNUvO8D9EB+U8n6hj7pxZL9oFyWYGUT9cHi5ZL5LS+siPIH8wHoFhv1emqKncy/a06G
GH70Y7ItdspEntbc+xbNETxTpdnM/SPYeowgmbB4+zG1iKjWTyeM2RybJBPcWD6midoUaCHdWhCM
nmdMC3xMhRfrB58Oo7k/2/GCAsgxVxT5JJhRzE6X+SnNeaO0QyuDM6ME/tgUvS8c4XvJsyjoygzb
byOaCkYlnmpcjGgQ/4wPXMDqEn/LPjoAj6/fEOL0+Zmc3Z+wBhXhdRyTlux8sXP0tPg/DZHLFG25
3XlIycQyX+ZWn04qfm5mle/pKvJBvGzOAbpJ/mVaj8RIQiUUHz76F07rOyZ63Xtrs157pPWxzbjw
85oEhEx7MVJMjGqXpwyvZRPd8YAVAt3BtI2PgUpTivssElwdDvvbE8gFJYm11KE6/m2XEnzq6vkQ
fHV8svUujrO+PHVpjHwy1YHOdr+2QE4zAzmrymeiL7rGcaZ5FyFKgNAm2rYY4nq4naJp8Bn8iQEy
GsRSiMscpTSUz/uY10MvGAvsqlBG5r0ElKCbdztd9AacHwyB52qMjj62OOES2+eRtlUjhNuV8Wfi
Zyf4z1EPQf6VMWIsEJ2974TSheEIXWT59g6juUjuz5FqDw7cpK5fdE/pVv6Y1KToqtiw0V44f98u
k/2hCZoDLOoMWpDi2z8/59GwSQeqishVh8n51AV71vgVIkYilIOJmqtKbulea1dm6Ezn5gVjt25q
tyzzB4T0ofXeqdss/YRuGR/uCACg6TPMeOqYpCDwSUyrAGZgn3PnjFnwUqUGv0bxhi+DKZTAp4of
rflGr7M86ErTDun8Zc5p4UgvWgLgPo7rujlpThPPwP6hkC35XrQkvgDxUVEl71jvaaelOmBYxTRI
zVZ1hNhgX9ErdzO3py2lojcd6UgnUMHO2Vh+Xt7GQNlURZLv/TFlip29br5dO4jBeSsAnjecOHl0
1+9epPvCWa1cpvOs4E+nCcoa0TEbj170nMJK5RHsOhmYnGWXupMl+ST5dhgvKIVZYgpHuRvwoV10
khvJvjqpTEKP/1jYvcywEX+mNvOtqGFAmHviDy5wJsJhvhprGRnSrWOpuLulXuYz/gfmUON3fvuu
mk/q9oVL4nU5BJPfE7Jy1rVeIFbJc65IODp7r1LjKUw8+KQ8YSHRLEu72YCITyzSXM0PUL5N7esQ
SMMgSbEY9UMfOmJEg0jdQY8HOWfnG10PYiJoGwWGToAntxVQrgTq89nd5nWoz+uSz+lA01ZlTsRv
AlMeVCU3wtrDETcpUMEj0WyzuHdEWFyTKl0RIH2iPmGAmH/WZutpROItTSaIJIXK6acFQ0T93Wu9
5F8lQauCmRcbsc/2SyguPkaiZwEERTcQzpkN5N+Q9VFyQRcckidboA+UnBgjdxT4FSF6sVfNYwdZ
MIUcjFuK29KF5CHQp+xXEziVxS8demh1q+WoKuqr0omefuroBX6zWTYghb0gQ/iZiezpUAtsov8z
JwLrcWHK7XJzg7V5z2rCLMlEhBt+VKMkBEtR6thflhQ9KSpDmvQUyWfJ8We7iFfRr5z13xNcUWin
do3oF8RZb1GWRHHEHY3N9vI0cTqgt7zC/CZGKJfUFMm/5OtuuWOezX82OgcegA6osrutvZwqdBys
A2/tBz/y0KIOtpokVO8Z0oCVo2M63lNzqCeAlIFD8n86jQi6BINvZi3vcY3lfjadx/TlSw95i5on
tnx7dtYP+d56QRZ9pBBCBCaHF9Aj1i35t7BQzEv4ZrehULGouVgGaPFzdNxWYKxdVikYeOKcj1YG
tlYjL32w0e1EHA26LqFLC+rw1nhdugx3HogvAxeiqFAbymDIg7GKlpj3oCWMQWqH19QMkqI2y7Ro
Ev5Y6WgVy72EU/f30/1nawAwa8/Jg3f6mhcdKg28Tu+Hv8R/Am9MW41vdn/z6/OHVSB7PTAnXeT5
WX5TWZLd43dVcq25qHJX96LQxunfb65sTQm2tZ7bZ0qiJX6erthjr79tQKF/shNMTrjQwloeqgjD
8qAOXonol78bN0LGiAa3c4NZXPUWVZdW+qOaX7HNdP0MWfAX/kwa2+VSNvx9TqUIDxeiF6crkTep
qgD0Ha9Rn9LOXyi1WEoK7u4i7EpDtmLZNLB9cCJuCVbgb/GB8or58rSCkYBny/BPnn2rZUGeTVT4
FISNmXDvhNLML36+j7w4s1/ULHYtGbZcJPBJLFkmxxVGF2jNxQTKjAGZdR3apkywyCIz+JxmiRqf
26VmvuWEWPXq+L6L9NyOGCIXUxIRE3ovBZlMaHWmylmV3QzAvP9A2ayqsZG7ETFbjsZqUV4e7jPg
im3hDk7+gMdiRZXDZirSEMYlifit+ZW3sBvnCT3vuKN3MHDB17QC1tuaceHz231vSgpm4Iscsxwk
FIjMAv5L436Bfp/OdI0P0eoOfTO5RJcnK3WTPInt3bvY9gL7cwekPXOVoTspBM0b/Xw9QPlbaA4P
dX8e0zC+CWLPA3OEViip1D+hPZK9Skf162dnDN9e2ClH72gY7/CbQzCfAEmx5Fqw+5VdfPixh6NM
Qp0C7+tr357ztt5Hdl7bL3s1Cg0/HRZhbhJnvKT+hou1/axM0ArqPcX2RRq9ICCIZm6J8IPvd0NE
1TOgv6dm5+guYR3TW5q30JV2uFaegH+7WvOchqyI2eU0bcVxvre/TOjsY+o3N9dsSiRnpfQRMnkK
AR9JaHd1EYrBwTmuaFxJ7KVVsuQXwo/st456oNG5FXnsFU2Z44sZ6owYHp7c+L4+f5k3et2Gw11i
wd30ZDBXnex0CQSEOp5xhUoRpRFtKTdPUQ4RZKL8CZ+7K6qrbBcz1Jps0O+FhOiUUPq1Nda3Wtzx
Gs99romHyXbLdUCIDWzW2ktciRpQhhtSiC4BcZVBnqjX77HiBEIVR7Ld/r4BGjqk8G49KIv6vLFr
IYXsHh4bRPRvbTU0C1mpga1UJcFfW1jOK+WmKOcNfq+iPlUuIPIYNIRf30sg9lmwilzWbUDs6VON
uFxnmGz1albmARsdrtNvLabCt6N4JtPiNd8xMSR9QjwIgSoC45txjQcYyBVIq0Zri7eMez4TIRX1
/mIWU2LJ7OHDwZE2EMyyUIvJKbO36SI15oFQ5tdV9TCwTmJzvbVKDTtML1iZFzstOjFmK5bXQUjS
MhG9TUuyl952h75LBWPe/rmjpeT77kuVR9vA/9dG9eWsk3bn4xVmFpl7BemFpMiXtPa7ygPKWOgi
EBN4F4MSfGpyMqidWyHu7kRUBkGhMebR9QfX5rSaKDa2cx7cWWZSEeYSlF9EvFHyM5jNbL/OSyDo
NLGxRkC7KxGp5iF9smMpePKywW8u6eDjZoIoAwuewL1NgGbzosvEaqANW9yEdZSp0Y81cQ77lVeR
GvYPv43Ia+Z1YlU1VS3Ea4ypG/isFph0FFbRIKJHNaLo+Wz4P86qafBVNVLKDGD5qQWIH+NnziwB
ZmqhVRTw6Et9dkBCADT1Qb2mARJ2MMHu+Veet67ACDhLiQNOvRgc7jqP3G37r/2iiC8wQ2aZFIh9
qnGGYo1O9usWrHPjdFz0gTHlWC2kG5Z4xgqkv1naqPovwMEWA1sJvWAnojONvFUrYVxMwnl3gAUW
ErTag6SSaJH+476vh1hGJCyxpxwzkBwQM4AcUqkNvAIeiIdH0ZMyq0k3fmjEz44mtj1/bJfd/4ng
NYk0PIsEjYfLYhbKe/hHAV3Uu80ZspfFctSFrUKyny+XWOlZy19HhrNepsE140lT7LQQKAOaqFjU
0wS++HhPHEeQfhmxXQJAFZMTKk8tCTg7Uk9Bwo3kuFbCUh9f0kaGg4cnjrhIQXMGdmv9AVF9Sgau
Jb7OVdUVE+W/WB5O7besgIuUPyqA/1tzkNEtagU0aFj1G2MWnNl6+7XC3Q383LXMaTqg9fg+8bdC
NQLcAf4DG4rk+1BCCZ9f+/V/YHBlKQIUMGvMa0qzZeXTce+QMgVHems7D4Oid7dIXtLL6JNVuRFH
H/nbfEWAkjzEtW8E8JKJW4UmQSvVmEozWy4iHsNNVUV7eC32xfnYB3+M1m1g7/XbiKkEDQC6DlJo
zgrbb5zgiDm4Tda+nWLvgVbhpFueRlQRTVGPk6FdMlQodwenfANhrJ7opmYdL1hYZHwb+KLGI0z8
SYFnVoVb+7fgBLI219M228uoxB2tinBe2mX3FpBo8jfFeQ/odi97hU99Rn65cwj0/htx5se73YRL
v/IqoQgdAgWvwjBQX9lyNap/DuWHk4KPNIy2VBXCF4zDu7vHRP83sgqVuJYIOES9DspZoDi1hGSD
fEY0sy5BVPqiTmbnTD7pn6Hiz3fT1S9sFHI7eBabzRwuMEQwztoloYKDhMiEz8peEnHAcmdJq1uK
/U6L1ABhL0MUtgZQWn3qb7KnavQolk5/UIRk4XuLrLC2FZc0ZC4V0kR6peAXvVFsnr95ZVEnDBHU
+ystHPceY4SieLMA3kLt3vczvE5vEYXs1M3MXeKR0kggmWRfPP/WGzOu7Q3IyVXHDm774bII0UgC
BNSCE2NjfcMk5U4OijT2WFIHXoDRgrkBaznJfhX9d3Ksercf4Eu3ZDACgwqSr+zV0lkneLHP4Tpr
ROj/faQAMjgrC29vECCcifiXByK71sVahFFEs17ja8LMeX3hKXbELeYwF35DOt5ym+efiuVjr+MH
5HstDBtAwd+judptV+T7L0Qn1KJihcz/uQXxzHB5hQuM7ObmqbdelBDepS1ABUHi9yutlIzWRmYR
D2KH++gpEh3ZsqfQ2ru5/wC0No4PTKlhJGsiY/9ZmbeZ7sJHFKBxoxjmgE0nI/uShtXcS1WmBKyq
J6PRt1HFxw4by+mzXN8DWAHptiR38Uaqs174ZJVf/d70c3iXfH3CWtEJW9PIqz6Cd+oRWgpAVTs/
ggim2wokwLDWAj96IQJzB+ClbUEyj3Aah4XsBih2dHsR5UpvVGcwPkvez+N8ztGli3//CDHxW398
dvwrc3Bf2WgUtQAcLkxFiH9+Bu1m0AUfJKGXuDc7/tQ97QybcVv8REmgnhlkYe8W4Nv1z8N9dXzS
4aVc02DJjTZ/zE7u2MWOsPUQiJZ2qg9sGxBPwxQp+tO72VcBjgSfdOis4V0gYj4Ko/+S48n5nM3/
BuKSnmZBuy5OchqKznzIrSOV1Cs+zlwdF9ymQl9cLfIkCcrXowjJe+dz6xp9lK+g7y5Oz5DV+koF
kju/fKkvHX5AHHsPnCir6R7g21/dlNdX70OMVz0lwBGzCJhSyR9dgqyPNUNwQDuyHKiccjYeOG9a
F/DoKOIDbWkoBKDEWTsfCBBBOtfi7lqhJpL0e+bp/l5iOpyyVoWMZifk1ws2rfZrj5VivgLzXPqq
C6WvoG8ulBECxmt72et3OnvoJEfIvgwL/FGnVWVYpmkPWsngRFBnp0UUJBImS81uYo/n3YLicRaD
1f5dbKPJ2a/P8Ah+6AT9fI51Lh1Q+hAN0trXPyCEJfs07x5Xb/KlncWrKpiaLGGICkWqmCPSPmYW
OxJZtigt4825A30VF/3bX5iXTZHNhIdCyJEGuI47FD2WqqBnvWK42QjlUaHn/t+uHn6/N1y3dkEi
oKw+4l25uSLlF+8hPEt1loA2hGtGWhV9DIlHzUKKkp8ZI3Q9MKH7sNPijipEnuOol2XChVokz4yw
n0BTiDQO3gBzdZZiZnOvRJut+o+AnvS2yokwztloKNvSmDxioSHUpPOOjbsklQkQjxA9xP2WgsQN
ZA5W2kXKWtPclN9NBvvJbmHEvK26pialrwbXeO7hpDl0SaZdP0Lrj7qGxHOAG0D5P6xmss8gLFPW
yupSNZohj5Yxqrf3VSBK0i2+yTeohYosSz7CnASC+72zedhim8ypTbw3W+8BwDhv5GPg790cf4AS
ScofHQbNSeIVlJbXST9emuY+WpVXdzGlQ0oq7sEWmFTGuzipzHflRAQh/VhZF0A6o6VzGJWURgUq
H7IJUKnNQAf1rBeLR5r5uy246lrcDIEJm5IDrP6DWxlgqlfC+qv3TZyB/IRS6/tHqNE38QaH5ZsW
6u4Z7I43QTF39c4Tjbd5I5/bHPhCrQ548tt2W+3UJfaljCzqx/gN9EyqDddOEzTiA7n3syp6adVj
1Lw5NtsEF5jEj/E7ytxJwAvWgwMDuC5ZH6j+3bcZyJ81AQQjOvIg0uXtkhB6Gz/9fi+U8NJK/iCu
goc+zcrFJgt+jM36+5Njq4vdEm3cncjs0H4ck4ueBAvaO637JWMSmgEUJ0vxj1HCZgcXw+PoihB/
oT7KUDjKNCPM9rLVUuIiSZBg6/6zfo+/PK5xhEBdl+gH/qfwk91gLkk76ybOyDkLHZ1xCiDcBcOY
+aOkDn/JRvkHDF19oaUJNPq6z0pE7umd1bO2bpPk6ww9vo/5en/svU3yarLATv99v/dkLfcHcjnN
gHgPJqfWVjeggPrIlNbSoK62H97YfT5WbObKG62hRQ9bZ74Vqf96d43YLaImcjgLmREmKWCsDLyt
xZuBpPLfcUkehangVaDl22xaKtxn0+WeFHTf/WgpyKEjHQV6p4cjfQqtQkq5ByBmDE4toYMKhMzy
W03WZWTuK6HN5aVjx96u1fbYjKhih7kokKITitFftuBsm6PC48CSkJ6uxlSig9TNCC5XmUzQ6ke9
FAr3pUomPtByRBHXpq9TzyRa410szaoJZdg3S6x2LM62THNieGnli7q5FWzJ2bd5Q8dVi0imvwIs
koTDjQmkfBBee3AVx1oIOPHY7QMCSwEwMUF4+ZQJJWvtov8VgwkPyClcGPSQeO3hk5oL8AOYEfqV
NT2BL7PyzSYohNPHDDMOY4E4y4U4dccMP5dZZeANMFR9qC+fKtS574Q+Sry8+cIvZS+dWKWoWYD6
qud7Kj/GhkoB/TGWx458lr6rvRy6GJivcql3YaIqIJaVaxxl/qJJEa1sufycCWbdfZf8JBG21zhI
SH2gWPKg4MYt+aS/N++4LvFbpnr9fzgAXpVCbwkbY1loHIqBe4C6Ic9N4ueOko119ut68kD6uWML
pl/+AxHlLfPHOEsCZ02d0j7jR+t2apqUCZUfdBTk0WbNekEDEUzbqt0Qw+QqVnC5MmalN8f527Go
FfXVObRiF+0KJyQtDV/woM9uapBSLum9Dcl/EFSk8PK2BEvON+0EuF1DW7F2eUt04a/9/aVmjAJ/
cZuHbnnBT37qAq+Aubaa08UVrYNl1UjwH6GiUsrgkXFlyx5U0rHQJ9RQ4CY4XR4B38B5mjf34y+j
4WaZ2h01pku3Z1vmuEoVIrJzLtO/dVkd/k6zgJA/yyOv8aoW697akPqDyDZ1V6KPG2E+tapW8QGW
QrpiUhKXYjVwBkX6OTZzD+q9UcyDzuFtMiLOHD7RvPNeheCiHx+M0ls19wy3xSnO+M6hYWvH31hk
lG5VLM3Ovd18VtR41D+hVkdtmd9Fwoie5+XhKBp3dEKht5U0QD/pFK0JwhAWQbLdebgBpheuvV2R
pf+3wlHtjq59ZZ7apmafbx+X1OFTlvPTuPvLT6XTRMtEUMYEGFIJT5+LmAlZHGjsldyexlPjgqS8
nmeNEO+U90cvYUdoB3uZSgpGfmgPkVUBgFU/zyg7udrz3YJtXlk2+LLtDUOUkwWR6BwE+J3Gd5ID
5cZi0ESblJpepinndrFci7kt9tZyCmvKQyEJmvJOKH8w5KB7Oh4OR828eVANMTZ+mdUAaNeGYBTn
WkDEWiy75L/rpzJCMSQEW+g/+39wQUQ/dAcgDcMe6/k7gMBVkGKoAHWjjdtNsOdyZDkYz4uu+iGw
45F9jtgo8veThjWVRQ+rEdYkJPEV6aJZbhcO+5GImRUBBMoDsWMRSstiCzPcDnUZhNf0XAioPIDV
Xw5q+jyudTpoqXOz4CTdGosraSVzmLB5YEcBOnjcVEGnyUSmaVCkfI36+BlKhR/oYNBuDZfOtg81
05XTTm/6AM1OoJYf7hV6ZrgpjXzos40aMFB5Z116JZ8wBks2mRWFWehUKZWpdigVvpPC1a/D5eYa
LLuHj7NgYM4yTdYJBi/Sd7B5hLk2QkBrOqYFJ12GTxyOd7aCG+8CcROctQcGy8JmEVrLBvcZJfte
7ij8YRlZHJCuAaq77lrK0eScU/VJQJeGLxL0ygqj25HVWFvMVkV3Qj+KcOzn4W6FjTHV5Mk2jD9s
PfKleT70qCUhGUWpSUd6Jzw4XMvBh6PKj3IASaY5BOjl20qc37xOK8KcH03xveceBZejQzY+HrOv
6BOJjvhQP8Ux5ga31P9kaPSUe5MJ+0JroE1dhK5GNUZo1jHmfHtbeOD7Y4EyhyIHEJhkbJY1UW/G
tRXWitLpoaeLulsM819M7h4CXoD1/xdQmW3IQDhRNMkkyCVD+gTTk1ZKD5Ypmrb6mQkv8z+iG6gb
spG/YsgJI+9QObEKU15EsMWYoJKQf6gwR72wP2WCIqx3Vdyyubv1CzWK7GfLQZuvO4eLW8tDxzh1
clC/pAkop9/9m9SW0bJxBXnWKwG0foqMJt7+fKUiHK8g/cGvuWiPTR606DumjNo2Sy64lVXGrRVz
3ChHx7nfYw0yog0aIxP3zT+4HN6/WwieHIeflwi5c1pXIKzLE7xjMgTG9nQztSkDEhqLw+fSoEyl
cb9/bxDr77cahKrEhwkGExgms198mzjFI+eM+eMdWOFNkGDQGLnIRdNVqZKy8eTyssC7s/CDOwcp
dHmNf+reHOhU9EFtl/oAn5u4KxmsX1CH8GiMAnVGmlQ6ckhr3QQRfpN8lCYiVT6v6TlPjm8zhnxa
TpJ472mtHI01avM2oruYmSsryflaL9M0zUBKuhlld/RgG9+eamNaU8NsnnEFj/nxQNuoX9Acg2/G
02slKMtMUZsoEdrex4ofmPLKrx2JfT++2maKOCH80m4/Hswus4GjqXj7k+XCveqBzFH3KTSpA/2r
IDZM3xKe+wwsMGSU9pULf39c7UilTGEyIqMQ6OQP1SzsQNGNyTgtM6YXHN0h7UaYkLATR1oVF/7y
8Zp0c0ii8aEUcePyGfP3CMuoAkMc9gwGIKkoa2xt4m10dx7BX190SGpmC5LHXmjcpbYcNaboxC3Z
bK3AyMst8V8tjof+mPRGc1XfqiH5d3bX8zJbmEIq1aSsX7DoxJQ0cPs2jTUdY+myjW4URf/Xz8fZ
2TZiGKCZIXiC+cFw55WpR3IK6veyKCj2+CEWvN4UQfXfMv6VK3WBYg1iYF7+IOLFuYVulgj5DszZ
6ryHA9RQMY6GtHj7Qpx0g7n7tMEYzHi4wQJyrmwksO39o+3c17ydWZ/D+26ynBceVPBYY70oszlw
GklhnSX34ToIKtPDkzzSZRBTdecXlaK2kCKLpJkFXQA7H5leKNv2qzjw5rVTN0BOZZcMNdF3ZOZ4
ASIcG7EOJ33HDbDSm4tmygqvlCvFmJE0gl2Yaz2aQGmBemeQLA7cw+Ky8FMzVGKIGOyurKf8ymDO
OW1Kcqvtf6IX1o7+DV5PoLS4vT8/l84UFugfo8O4JPc5LzlT8/sqk/EBu4aJLx7Na3ZOnfMjfMCO
0AjCAlmNxO8kgaZi8cgPjPL9DH/B0ndXrYb5TPktIwuXIiob07f5NzCaQU1ts/uUSkNLsB9ApypX
643llmT5F+sCPsojGCzVxQ1Qq573i+uLOfxUmGHDznotqYx7CbJR2XTdl6ZXQZx4mgYcxK8VgEUw
pNJki/2Fk4xqBXLdsyJ8sE+rDw8WL0GbsJTNlWK5sdR+mTh7em9yfhDQD3Xpbuah/L/TbkEcZGLc
NDXsyd+ZP7tNcwbPeXrOpCZ0ceIb07h3JOtThe0rmfnTpPcKiyQBvHCuPCjKvT3Bcjcmt2nBxdif
h8ajTQbtEXUB957tILwp4KzIt5vxyYKnct/Sx1A+ESHVIdsVPfF+x+rEJrufYm+FNA+ec6ys3bsa
aJ2P8GIkfPAxgvipya6am+eYVDzH0Kml2J+Xayf7qTyz0Yv+PgeedVL+5wE9Gry2M3ilNYQmTwMT
u+4wYkxjgDvCOv+qx0JRKmTMtLiaG9b3ljPPQYdg+qfoD2vmPT5Ysq+8Db8HqecR1XNSgv0dLi8a
vZImsFAeb7BQihV5CDwgdMGSMD2tqRhK0L1vlfaobQMhBku5Txl5Chuqd10ovhklfueSCU5nAY5D
8gSAPjXD7apgxUGp7aednhDqJkq13ZUcoAzDl1OT1QKPpOMF3Jel6mS49Nj23rLqFADJ7dQhxzcv
DTWXf0LKQuQLgQFMIyqxlVIvSjp+zKjRKip2mDsFxtXy1ckMHcRr0vjSBcwGYY0Re+W4xWSCW8km
4lMQfMD4ZUwMGWf/WXxNsA0++z5tWyEUVeeRY5cUfWFZH3ZQGNhKCbIeZJ65fx/4brEaLQQZFLYX
TrxboTOeXLTJUcsXf8eywDWAKiEfeDkC9AFeV7uxR6ylbAGFbgCZAUmueKJY1dFvUii8D2UYzNi+
Oquu6vBSIzUOb/e0zzkGhgj1rnoaUVxSjLVd43c9xWX+T4MhsoCl/27GcgFZpzlP8heLag9+mUdn
QRT41aCwjWgB4zdALruXraZM/MoXtirT6/yoWTcCGC8jrS1scamYdGK7zYy6JuLEdWUWA8moLLcp
Oo3Jlmvm9GxiaePDAsVPiw9l2De7GHduEXNyW5dId8vps+oX/XrlV/PRm6FfxgcH5oAEXhxlr/5q
MFWNaZW3PrIiXy8pBsJd7Hzyas0OIreelaHNI6ZNjCe+vxT/49qZoZsgIGxe+rUq0cLt38e4PTh7
L08alWp+ajL2EojLWzUNmDytaIWkOikaZXOp2AdZxwQ0oRcQPVsfDwiIDfxpitGkGEFshrtpH0X8
rUMm+bU1CfHU0WTcWbrTOYvYLSUyqdtRY8x4zwZjvrkpDBSNhO5iS2g6RN4LAPOWKxVm7dRcwnF7
/epWx+iRiqL2DrCj4F0Ffjz5e5ce+FnB7unD2Lg9Xv6vOqsfY9Qcz5xJKGQvMmi3tVf+7pE1CPOJ
Htx2h5AQJedGwF1iA/fS8r8CaDpme3B3SufXJG+izRMAe+eitUcCjCdPtKVHZ6ZlBt0zdD0pWPQ2
z3Zlnnvo7SrZzRNjxFLZ/fedQbzHTz5xjEtdKafLldBNW7Evmec3rhYGSDKHRihEnYB7ozOiRSD5
to7/T/5glrBAtZ9KtIZmGFegDzIuQ+a/2CDopG9QIPziSQMCsnEIJA4iSVRO/vIbYFDAw129zITT
6G9W2SKBF8T4Ofh51XYfIJizi3l5Ph6enB+NlLn04SOhboRGbpeClBkXL6XvTNVqY3xwif0RqtE7
p9YUmX7sdccDLx3eNXGsxhiQIgWPntwWwHgvObSlaz/sqEp5/iHe2DiUoOkUcqptr4zzQSD6XA02
mwIyOW+xJq9IIFnPkI/bEON8RpE8zkHVUZo9P1Y+jBqYjBGXzLQKQAmTzC7gZJWlAQqafub3gd7A
zwNddjjdQ0PUCcRBn4AW910YoJUlHAFI0dBsPbs2HktUeqgVNSn0AAedUpjw+L1dmDN9DigH2YNb
7EKOKjprhC5BAVB62Ou1zGsDFNFmu1o8wyKiYxmt5JU0aBPBEwgDgvugcVUiYfr4giVIhfiFebKt
Yqc33c+VH1GoBreK/E2T+VjsQycuKag6/OEmAAzR393RRFH+gWZ6zDxCHfzEFHO0Ly/J3wxmCvmi
e/nrni92Z9N9UewSJXgJqRSDgyZrbd7+sHa18KXCJChIcuJEYIMtT8YIIxUU3zw79asW2mbhDZAJ
DY5o3MCW4f/UaROlTr2ybKok/HgQlwQP7aSuI4aaEK7419obT8hdgK9ccjm7YoThB1SnEMqG1z4j
FKR0moM5YWUIK8JXwM32xrJuL0OTU42j97wfmOcgMiQs/6/3TozX0SCT9KRaMY2VuDSF7POqj6Il
MkmtJvNdocnY4R4Sf7x19g+mtMpnoxzV+fduZUOShSb+YsojoNBTKQ50dPhkhN9oxgaI1dCVuNbP
BbO9DkVowkj/t+aQOD/Hukgps9MsrG7/WrJhNG6/ufJT7Hdz5Jj8dsb5n4+z2kzBQth6EK38odM5
JlktKJkw59574oMSwCnkJHLzyqsZgd6oBb6A0XO1qQjkrWpOC+zl+LEFckyVwpvPEnj+1XWd4aWV
/dPcWU5BClRpohMh3z9AKtwq1j6RNTlt4m0HymuMenVhDZWwivPT+AvbdC7sA/XBU35BSnBjRECe
HTy6N1KqzOhDRVbsnR8dRcxWAWtaGuA8I17EicwOfynfha8g299DlmlOm2dXSdizU5W8h8PY8HlQ
7tdz9cjIo79/TiZYfHimVtY6/W4LJuFaAB+8Ai/2+Eb9Uf0uH9AnODb5hgs65sBGWsBt2/6jL1N1
UBEL2W9QqoSckdXznnvkglxMZoqM8UwXn7YA3XwLQFR7idMrinjAlwm+0Y6K09jbKuF5pap8M5Pv
JTGKH5hhjkg5jcwiWf/NHWqJpjuN5YoSEFDWcWbBAphFwJybnUE3HGpUIcRZPHNyIPrxrG163SWN
yFSXKeFlCWb/Z9+lZ5ExIpU8uEvJ00kSgO1qO9I4tfJskeQp50wxztDctd3+a7SX6Pk5453Ut5MF
zEvbBXA4pJl8tqEXti3nRnFREzv9c0jT3dNuGok7yw2oqRQSuqNjaHgh0e4UAH+oEzZnbf36wkie
iPI85USlMqLdGiq3IRdggdFNvLNhUhLEO83AkMPE6ZO+ZL50SUDnrOo5MpQzBeW61IPpJ6ybSqsj
fIvugPl8sWFKK9O8c2Z5uaZM1La39qHPHjCiJQ80VAiD+zY/FGRHopFsTL/Nj80TRPrbsM6uYeJm
w//vr3vqK0PKH5H9m+nLJMkR4c3GEeXskRM38nSmysqbpKmKyPQycBPIukFLXiu7KfOUsduAHwtl
J3Rs42292erCWWxfJH5s5hjcoODeMfI5qSdNR49LbxCXA39Qk+hJulkAonNyIAnqCOJdKgHC/oJQ
R/0VErQ6TaJ2nKMq02dRwXKEXbCzTSZBYhd2M3em2irGoHthW8bdFSNn8u8qZigUqd9CRvnPUAt0
qVULYaWQhbAwwck8LkvHKIZbiIYf0iwMC9wv6VISyZhZ6xp0ZrRCw6KOqICb5ChFdUc/fZkO5uGi
GrnTb3GX5d+aoFijwq2eErObp+RzDw5ORGB6aIt4e5tCuShTeVvQL7nUfHNCVWhN/vmcJolOh6sk
NCC3h5ScD90ihMsGc6bHucokfUuCsKMxhH2hv2ZP0BTxoYDYHsHJ3lHbNeohg1nCA9Z5oLGCdA17
qa/ezfuBB0kUkkBQ9xtLyFhQKqNB/3SAEDcwKmCMzpcyPsybhFlZKIfwYIdedG7pfr4fCUSzYf4t
LpqGVjkwzsPVpw6TCAPLKFxBI41TQWWs3iRxS/UpgFAfzmheEO3QLZ9Rqu0aYiiGtsx6NXZ0Y2Nk
7Xrkyr5/Ua64S+Sg16TBFvyzvVEh7T1Q+0zjLCIWvmmgZFBHHxW3zc5TfnwvQP1TYmveonS9mBgI
khtdf6tEXiseo0zX5gxnC1n1sbHZY21+vJjVQSHdOvWFi10g113z/u9+Bu+CI2gkblZLsfEn8+hY
tqu1JHJHBjadk398/IdichHffmmmL+xVpcSqwOUVgAY5AVIZxDkAG0OVFh2U9XwPV6ZR4LOSgEe4
OpDF/8oiurOlNBQLG2fk8DJiWokLuAGRemPm6HE36V/BbbLnFti5Nzo4zkIntro8TGKvNWVhLD3e
nbreiOCIIsl2U9w7G0qEvS6P0IcZOoXicAdxTMIdLI+hiMYq0GBTsnjjCzSd3aX4h+zmKsXfR6g9
Ph8kIYo5Us7bUFwK877r+ob5efAiSj/xuzt4nPkLYWd4pfpzR4zVgn5YD5woRLZrdpYfdiN/YG4L
vXO9ZhAttbSKbVlChgKPkRgiMs5yIG9volb+PwOAi+g9BfqsTGZC418f1C/kWVKr77cX5eCNvNtS
8VNnU47e69LeyHc3CYiPLqcczF2fsJFBQasCgId5AVYsWSUq11zMTLjdMH5Nu5klg5zIw1EWzudd
EIz1ssTOOOCyJH22NqDn5yLgWNHsBwUQqXeGmDxccSfVBhCk1zBMdn2Ri6rup/7sOwYQ2U3ipW/d
L90nbnz03d9X9iwwSaxrmgjSaVox7HC/cH4tmwIDvXh4Ehc3VkNJdqfIFUT9p/ZJdywy/oPIoukJ
SRYrX4Ppt7pbAqsv69FWMpDMGpYavozi/bRl+KRvgfH8M+tzNtY91Apjt0m6TrY0TJP6/AO3zy2B
huba9xYxGPd6SJ6EwPlo4MjgtXhopTtDbDjH0AtpG486+V0g0IxUa5YuwPtpbASBCUOOWQHuiSZU
aH6YkRTXEmlV/hMvfv6lE+1E4DOHZ4lPCEmeVI5q1gDSevmQkf7fr7mbj3ezzzlo67Ec+Dq993Tz
3bos/ZKHwNWVg0JpAM/xqTt8Vdj/ReIMf7/DIuO9IuAflg6JfUKtY8DsnDwYoxFv1mggHb7jLAj+
vv2XUzFd3d7muur9eMpH7qp9W66QxEaPEWA8gBgXcKy3o7fbqarEY6oJVq6x0GKqmMkzEXi4jQVG
DQH4BRjrq+excsyWd4Yih3fiyKQXGQURbgtXnbqLlbdc3Um+n44gw9CZD+uR9pKraeA88pve/5Tm
rwRSjW8B0lUevhh/TqjNaltWK4PjSf6gKUQ27bnXTXDktiT0O8LkKIRy/25iADnS8eUIwk2zHYkv
soWwppP0ekzMj9v3GRavBc32QJ2ILGxQOqkQaBSN8KHLyaanz9yD7zMNxSQ88UdCiLgd71PFEJsG
iJPVTkifb1QRInZxp9MULzietWImMisHI3sQqkQQVQEqXLTGvU5IlOsJPqU8VX2XUs4wpG/+iAPa
+5YQm3pKj4HzJzPp11uLyy9x561E7xCzeIsnDCN6RztgT3JIzh61vpT6IgyQMlcpS8U5sK9+5Q9I
GZo5fRsdkcCCSU5wQKTWS8C+PHGWNqadCAJZaHGYuG+WUqyWd3GG2I1XewKs1aV5GyEI8SlkYqz8
cWH6kstuuqgXdQR+1Lb7kWqgUBBkE3TbfotpQD3eFq0P3RULVBv3zyNDVp76ZY2vcrbr5YgTiFL1
8PJPy3aTlth2lcfrlpKILobUr8C/qkOH9QD7GqnBBsph+slfmpJXGROdxnpZpcdhqraY20os/p7Q
595gS8jGmJXTiixkQKERs7RI4/6qKxovlxGhPJ7TkNrUqyDl77Qg91DrxRpTuoPIqxFpQQiEcg2w
lVwA5Kp3D49iP4zFNfo6Ou18JWlZt2zQT/YyMPCGdtzz05teu0FlC6oIoS5Ac5Z7xdjc7CGBQpC2
HpTpsE3smJLqEGKy+axLTZ4OPwJlmj4yKnYPK65bZTpjANZccskQp6wlywFMYPwr3qRL0Jte1eJ9
ZX0lD2R7w+l6l3CcuI1Gt5uGEEJe4rqIK24OrpT7m6khfww4v04jlaqXyYCDBE0Ho7zLXtZoc/fx
OyEIT/a4olcUFLZScj7rFXCPMMgMcvPw/tgmuH/5yPfuz+U+l0+ngBZk00tGQ2gL+24jR0Vz6D9f
WuOCScfU2IFXBEW8XndeTbPem93s+0117+lNrgNXyeOWIlkvTLciihsfGzhD3SqDxq/j4I5KShVH
pt1CUxTsKPxwHAVaybdJzTvtR0zZrc0qGodbIsJCPdqefuTdVX3v1hniULn5ZwQ2CkngtC9GkRS9
4mq3+sGBZgCofr7wXnItBpxzlOlegmSb4+4HAmYopBfyt1mHeprYZpIFzLp5+VWwK+8aN8ADDKek
oWjuFv9JTT1D+WQN/AZEAEuu2BNtQNTjHZyw0X0tdDm6qk3/766B4LF3abTY8OrpWm3lZ6HI+LNa
AnHhi1tU5mDsThpJ3MLE1hVjIAOuBBRlGQsX7L7qmj1RrHPNPrBp/3ruJ17veuDQWu6pJrjZyygk
mdGOD+0FI4BlOfznZBNmx1K6FJxMIFWEOUpLbzkt8pBijl2p2kwbg09LIVJWZwp/KlBUSkVxoUpM
4AOkzs1XORxp8K//QFADSfgudQeo4OklvLGTeLDm1H9d8AXG2CNoxsA9s8X61RKd8fagdjw6e9Lb
KvuIpUFVgMwmAYDK7Z7Vk7AUuWiDtTvFFylYt7NOUwVXyR94C8tdGzdIFDB/nyaYTwBk2kDh3dn7
KSOrDL1qZHkaYiuH4shz2NqmGl9KKq4cGulC61VR3/YJLx+ihrpoK14WbCxSm4QXYHsm6FFHeO+U
yh9ChWRNkHZeYeJBM7txGUPJi6Hz4qaP+RzUbi5e5ilouVUE4AzhhxdamALBb1ENnjKaWiFa8ETY
qHdqqe4MikUtO92RJdVx6qFncEvExdmGi3lth2o6SMqXfZ8JFRP6LEhg1WQkcwW4v2UYdx+3Za6E
XWfVA0EkSQjxBYdQR3bAx4A/hJIEIK+e2sJ1DwtdCFeWu0s7PR5Yc2G/fHDxGhp/IQEFcwqwAvU7
MubBQ+j4K/bVqshXCK3WBaUHnkFFrjV5fdp2ILZj0L/FwjjJ81I3prd2f53zPjBxt+GwDU4R8snC
IyE7TTFGIlBWJcx+anNAtR9C6yox4cszwngpcwlrdp4N5QAhIbvEmvz0D11AjNEeAC6pSemHX1sX
bV4HfHK4PtqqYKBS96saWSJALgdPARWNqvj/6wztxogjiGzgf84holNABsCjflCSEJjneT+mh2gL
wrv0QXQCP219xAuKNYV4z1BGKIkOq4HUTN/sdUFOdhv3orPq/6Kp29Ap/z/FBiQYm0/pASCbdRMV
u6mMFj82grHv59NzEzO/TA96vEi30beJm/m871IvqsA/zbS5ErPsNqgGGGzJK1E3WWZCo7NvrIcf
kn/k5YUMET/zfTOafgS7HBagwZY4n6OQ4T7vHn4tq0o4UWTvNUNanNwpeBGvcRJ1NFcwyVAHHVaH
6NdlOreOkfyWYL4LMpmX8uQV9dK3JcKtqhSdRTRGqbdRA0C7HkCEY9M8Mnfr+BV8Hq6eyaXy5su9
Nxs5epaKNjmcNaqR6vLSPPxnwwOKxTSz+Nnmf3uAgn4+qwSk6fet4KmRMj2ylFQm+v9iRugrrk+x
O7GH2ySOmdE51w6XGt3SUdgyWxOXji5qe5ATJei8MYElGv85GhGl93Mn0xJ8eyDPpgWjN/12Nkyh
hLbNE13ZKCfGDQ+5/oN0s9QTJ07Ca2/lc0exhOdJQsFrQ9MSu3dsF3p7Vlr4wgyRNn8sOagBxZWr
AcAum5eB+xeold0mddteyoEqiNovLHnCDjMtdJW+L5dGIVZDBGz0tmeBkQNB5PfLOwLBUid2fgTa
0GCgrOqvTuQYJdzN7xApyfrtBItK+T17pHGVO6dIj3F6VDZcF2a1wYisLK6OV5Hk5eX/vGRadpf3
5DAzEfKKBUjNy5lpfBl7OGN22BF0+gvx9ZwPFk0ywDFkMMvScROA9bh4Lm2Ow+Mw8MGJfaLHSzLN
wn/FXRU1ps5rk1BS8/Jjd/Xbs3ilTcgaczeyzllKPYGKbMmDplA0VwaalhGTgvmhKxUvtr6AT00Z
gOARoii59mneWszUQi41/GSWP3EzUJv1M2nPSk9sc5NaahEXLAiuqwa5S3aDn8k/xG2v2BNd5wFk
tF65azA0li1JzumJiC/LZHwDC6GnAu5D2NJRfse+s5nXinzh2OxMM4rBcfSPWWY1KERqLuykxUUe
giqcKfSlN/T0cWIbeGkZBseeZ9542/Kw+EC8tFPeu920Rz3cYc9Cu9/2QtBEN4VClVAOHFKH2Ijb
RaprS+n/lwNitUTUSGqKdK5p4r53RX8iNSPYDxzAAozfdwtqbX0EcUEKiVhIebvzpzZHCKFWuDGP
EDTmASEvXVgnQbz/0irBXiCdZC34aqpykZSrMQsK0hxgIu+Gowa7NU5lthfI3d5anunIh1g0TwzS
ScR2qe2KIELA4oQzwGLzs3BoTm9JEsm3sRUXsMeroZlwk0SZw79B3qtc9bIiOhPYjI8u7bFyWBrz
Cx6G4gJtm//Ih7ADxpLWa8EnLesfzAvjK7jgPjbaD/6bmOdwX344QJCltXuSSWC+zTkI+hxvtuXP
hfXMZ0Nuf2baymvMb6drpt+5UhkwkfW7C6suHA8UgrTj6lz7y76+aS2IfS9iutLpfmZoDzx1TLcL
pB++GlO9KjxxZ6vqxW6M7gB2QlGQSWPK1GZF0FKMPDrImWxPkaztyAykviL0V4Lb3nZS3w/u07/X
fTfNl4/YyeiXjoJa7pnOKFaEF60mxJcamVhc0UTcgtC/3CAMOlV/U/+Jq7sEfipY0yaNOPdoisVl
yTMIoZCQ5pqL7cSEDHlLgdwgHeGiDNNf682sJD6e/+yJo4DyacnM/0wTMYzttnZQETGEpgzEqUdG
T9W9icRh14rwYDoNtf1Ph5SQNqi7szPZvuuMJU39AKriQvAhaP1ZUI+s8JRDQuqITJDsMMtD+kOq
9pwpWtxgB1zf1AjH5Uhl8Cgy3eLsGE3AJrKLWfxLkx6TZ8xasCwAQ2QLd0/u4rNEhKHE8hw7bHiw
O/zTOGyDFUuGt9AUmOLBN3Ox5qtf+MHxcl5FbH4SH2OT3XvSW/tgnGBdDgSuy1+jUHAEnYANZlGA
D404i/6rRceVyiTsOdeoIkWhwNSLTwbUOY0xCLnOtgA4QNomokpRCP73O59ubDwWdWvYO6Umlik2
S/2x/bsh4dx4Xg8Lt8FxpfMgMgPf1nv4Ziqh/Zz2LOjlaD27YiXTNESa9xojzeIExwpqXvw8vqgJ
and0DNDuVxH0U5pmsVskPIEC1Y+fcsGut5coIViVbwMKLk2j2lLOMkX1Jfj4b4RLkGWhHGkrnjSC
pXPrEXQnw77HsuchphOjuyXlO8kaGEVNR6vVLh82Q8OlkkcsytXNUf5MusZPthYPj8MQ34bAl1/l
5Q/prAVp8Vghy6iuZnY5UEqUqgJEZkg1jsVrFeUHWVz3powy6hJ1WBm0usLxzvKJvs5mSHJPqRQU
MZoXP7oS2s8/cEs8/kq/rQfEI8RE1rE3aL894CAgpZB7whxobAECHOf6GbBxvJAylSXR5qCl+HIO
rQQmF64pAOM/Y8lv7IMSXIewKB3zLGYa/PtXxVu426hXPjvAyJCTyL52h4UGTuBPQ52sRXOzGGZG
QsjzrA4tASRsjXRQ5Z26O9OckAC9jthYAcrXj38QUththJORbeC/2riwDnuGTMprCRpPebRO1qct
86FPspYgyd1PLH6NLiqjjhbW7FZu/grQpf4iD8q1dwcTj6e10WGaTqsm2yhjfq0NxxYcr3AAfrWL
PTEKOOPbfzRVKDd+2fa9a/ufWWpfQHfqRh0+GEr59gur6rTlRAsun0dEDt8Z9JUbiFgjkvsDhIXr
HYGl6uklBMBVjQbnL4Bt+0z/tDxMUDRxzuyPPx+UcriORrWZHWB8GDmH2aslB3qlm6x41PKIZicz
rFw+t0RFffB6/PVQt0RqvqukwAp4VLGwPjkBb3eAZK+aK52TDMPE4RZKJS3Rd6Oka+ZZla/lVTW6
zFEEfUqCxDII+89kajfOjJod7taFwvz9Vma/2uKKgSdAYdJT5gZHe+2MVDveH2jPwLssfx5E3N1k
E2ae/Kj9lAMhzxK3ReBAPq/SXN8N1s1RywHJI6XUXiIJcvcj1Dq9rUOVBkxp2DFGNhtKHp4KkvTq
wrornTeI3kRU7Qyv8bmb54cxzZpiA9A636BNL6rChTOHV9ZNNnuJy1lrmGUlH2SV9j8ZSvoTuQh1
ruX6psGhVC0xRWP4jUlgOTivIet7aHJP7QzPycL6+t00oqgrCOdzp1GzXC8tIPjT2JQQxZWmadwV
20KMvgpKAoT4tF4E0RmqUQQ2KM3pksqQ8VfLr+cy5D/GOrz0Mc7Yxw3aMoOSQSwB99ZUp+5IwifJ
zyLSrh40Pjtad0xCBCtludBWYDQDZhz60uBo7akBKCfKC1j751HsT3t1BYwLSd39hHHsbHbjREtD
Z22WRDb2q13DGeWi7Ie+o1nIq/HLJhQ3KCiLsZXS1x039a+tVYNW5OgZlus0KLc84xJObx9Wg9gx
ZEjHIbyrXMNBvtrkgUNmMU1OaV+QQ+7muDK3WSFO/TtCjAcrH6GO2xeFd7ycZgYd/d3yn9gkakY4
EwG9Z3mkK/smrQlNNrOzewlX07+AJRQ+d4/9eiB5bJDkGgKsuaVg8nFVWmRfRHm/vdqAw2UM9v/j
UX9Oy++RhxnKLqrcvFGcGOYypN31BWQRB6Jbvn6/dMEPk/JfQdbB9rcN5LuaNbAjpMDwYdrBSEa9
Zna7sYlS0BlcAuhAAhbmXOja6OiboVYxYFhGFSX2WEWGQkoAd4n0uknVqwzviJU4+5SyX87ba8Yw
fgQ20B2Ou8sOmA2YnV2xzhyU7AR/VsAlX93Sm9HmZs58g2tVQZ+EzzdhqNvjV7frWpxNNs8o58bV
YDLRp5eXSlxEBhj+1uvMe7IJxjsVfn3mkrGOR59YRS2q7jiGHoXAFL0e8zEwXumPuN8GYIKPVApU
+RuiwuEO0DWRTqjEtS3MAoTeL6CKfaZgVwYvy2fY32gh1a70q3p3sZbAjDvxB5Ab3q6THCgHlHjk
77qMR4mflXXYxviM4Z1kEk4YFulJa7HM0DTXTtIlaKg6DDaOT/EDZvPwh51J39txrmetSWruowJ2
DdIz2aJVvui4EgWTTtRzg6voBM3FeLU7IvsRrrwhfzkGEqMkRUY1oHXDgD6Uv2qsb6TgbWpmxhjn
CWv33RvA4uJuAZC/5e0ldJA1DTFMjRzd20id2pIfQxIqXNyo9w669I9znH7dQlxYeeLO/VFWy6eR
sxRDleolgMN0A8YZDlz4bBNdvuYWOz1JLa7k7Yl6FjP0tLznnA3shIcL+qIpw0lZhZqvcF5Kc3Dp
KYY47FOxhYNF/u9U8Dc5z8sH3+HHAOGPHAc4vRaV52HWyT0lRHB31ylQd+11i0MNb3z5z1xbPGhJ
buvuX3SsUOM6O/5MmyW9YUCbmQVBVpLLRmNSI51IUfUwBAS2qEwIIDgkcl4aLz/efPQp5UnfRU3n
1TM+ghRWCgcQmTvA00yKmOGdKGBYVMj63RlHvDOYedYRcb1N2Yly0vduum20Vem32KJtX6atDe24
YDsoU3gjb3NE5Ntr4mAb8fk9OSFhrT0oHIYQl2yYBVqDZUDC+NlIoxoLMC2QM8mZ6HvjKapSMZPU
bl1gBdO5pLVlMH5KuwE2RdORCQbp4NdekAo978BQ87IpbIlap0IHHl7HujbtU6M2iDZ4XnDruAAl
Iz3I+tgZf9ZrZSr6dWW6qNTQJILGLOgEfZFo13GFm4zF3H1eH5nqkJxi/oVSx5MURDyQxhZJSHEc
nlClvOJpd+oqRTykg/x0/XdSRduzls2s9CHd6IZemoO3VJXPx17Op4625q9wdm8/o+DUg+OQUwB5
TS23ZhOw/5lceWZhRAaBhNhxKVF/NJdVAd0cKdTspY4CDRHem4uX+tySFC1h0GhRiZjYeO1qqtKW
0yrJWKLotg5xb8Fz6rfDDxZPYk36VDNufd0l42aWb1NCC+B+wERWrxVZglY2OVyb8D5hiAJml6l6
2xXU7JSNHqsrHT/sDpA8JNhnGKUGinFAquZ98kZ97pOMTegaf/ewCHElcSyXMgEm9YazlqKki77x
L5G/W3uDoBI3t85+kotsF4BvG1TfMKRuYN/U4eZJwqSzWc23Cu8CvUyKtVouxc4mYmB7bPoLQyUS
woKgn16XQ0FdKDYu1tQCRTkl88S/Khft86qjwwWKV5mThbde7WJ6/Fyg4nqbjqhtbPj8e1U7hcHa
aUSCMWo26tDVdOB5TXsjyJHSpVGakcPSGbvQ1IrqG8msdvz2ve9s+8TG7iLumCRmhsl9M21oH8FX
Z9ET1I5Mba+SsuqhNl8k1lvSVFL2WK+QewuHy86TV/ZK1FQqE1lG/nMIxfbbaItI/g8GcjsvahPG
a6z2IN7kzjnnxqnbfkGL6Jd7Npfpa+4RNlYv5jEbK/A48mMQJvJ9IpX3YmRs64txXm0816hesCyT
BLxwGYvbJuIyviR00q1h3fDtJS0WcuyTGjid7rjS/ex1DuI7SJ/IkGDbwgWeAJhhB6QjBc515EFd
5bdCSc/c5Zwjnbdgynp63qJfV5jhP3ZYL5BH+nT2e/TDo7zVIw76jzDW5ReB0ebY/YWDKjWObtqw
2eZDlOnufhcbbBtnNZnh19sGd+YmLlFeTyIZqRGBoIzVC2TcaGf4aF+c6HQgaEcL8APNuB6Zk/97
s3BKhGAP+rwucxeFZp47wWieMpkT3vJBD8bFgQHCAxzPWCSlCuUPmZl9evloQDXXufmMI8wMCE9A
s83XQStZmHI+P9tEJFZGEPxUCe279l19RVK54YPNBpjDpHrz5IzfekkP76QeTd1rI+qE7AmZmrZo
m0gW1KUrjFhr9ArNdDnhviFlkZ6ZXOIuGqPkQKhIaTE6aLcs4smD0lSjF487NBQtDBYyHWdfNPX2
iFZIFPykVjNtcDw6n4oFeIPeDhRJRVGEUILnp2IOkDDnADkvM6HiP3ZHDgYqhW5cLbWqhDh8schm
FWLOB+HRWEyaDj9/ObUnrdf2zwzR2jmQtbL9KCUJWN5nQH/G22ephaZSk3sPyUKIiVgvCPSWoFWZ
DUoJ7cb2bIR0Xs0oTyZL0CY5RNGlldgr2e39ZMz42AudxyvYWhP+Hcrog8p9HOxjD4baumrGNCAi
dKPrs5nnwqUDsez8KqHKqOpGycZWChUbWOyYao3M+ota8kMLObOItm/5KHPuOuX1KGxAqfsDGskM
mTSGK6GrMwVx6FJaGeNMr5L/ZvfnKMuMU1JVmcfYUSUMSBDI0pike50QEnNL8eH1U8YdpzzKcBCP
31GAMz8rOAONqoGY2TrSRglraV08jpoLUpcbFN7I6MI7rgitvxvzyuYSCT+TApj49I8g+hz2Jica
Smr+8pez+t86p0ktaWth8yRDoEcUaDgvZWhKektQKvsK6ZeAZ9z0f9NElu5tlfdQ/GLtSda9X95S
kttlxo5MBL8mDBqUJZOZJWijkvBHi/KnOMp9b5zqbbjcFuy9Guxp1wuUkuwS3DOY+hVqZl/G+VUj
6C7bniVoQhQ1B9VVmO6BIOhjZ2joTysvyzLFU1/qY3bZPUtTNKNqGwjWODjJFP1pyrKidk6W+LW/
7Uh8j88csqHvnp//L6A5SW/hRYungazaGPvQZ5co1TTqVLXtqOVVEGDKLvgecPLbXK9bNsr2LSY7
5CE/utdpcz9buEE4D3edIpzReeC7gPB861aqFudFKqzlQ7e4+bpwg6me9l7/pLBPHYpK75H1nPeu
9SHGrfug3gqwOR6b/9nDlGBBynOEnkEwEni8BPRd94+kE+XWG89t/VurkqdUZWWVF/88+OEJxdj4
k2aW0Nku+sGGFmiEPm0We/Cgfw3lN7j0ZPF5yERgzCRayevEGs/bpVQHX3m4zdNmqjNiUn+8hwYq
1osvLWJiIY5h6EqZRXkLfLNYTffPepjicu6IDBw4M1RPUo68PwzOIN7D2yMnB1h5zTW5a+Hja8lF
193sFjK5gNzYbnwFjWU+I6Amq/NhqX095hW12ERWtQR1a40cW8aAg7Mbs8QpcYE+FjdpawinoK4t
VKv5HiuGeH07EEgtxgfgEdZG5gGxxxwR5zXMbiS8E9xvVVqSoFj3VKtWUVoY3gl51r4ecHmiQaGS
twzdu0FZ1xRFVuhO5EzueJkjX6vHWa8185nyc+Of1+FBWZiKq+zWoBT4vidmADWUjef49QQiUM3Y
0flZ1nVx5oh333k38bIjLon1Rf6hgbNFHsarwxTWuzNzk1GvaCCFYKQbKeXUg39pgJIHcx1RF/kz
elqn8eaMuZl/YUVLvKuFWLwLe/WMzbmY/1hgpdkeG9ICfeGkiA99uPsbt74dgFZoiZfiQbb3lKGL
p3VLGXO4UkY5A/rM+t6ehiash9DqayOlVw6zGOOUGG2F51KKxRvC7n/bZnwB2TGbsMetVdRVYQun
HELFgww1HGviSUHimO6NBXr+OBCVcgLzgWDK9lSWlJAp1g8L7ZnMAl0ikfd4Z/dHglSJo9Mjw+Qu
RG/9WRm5e1srT4L/rN4QLEvo8o9/2jnoSR0Hf1j4RBAkaQULfDD1o8S3Qvx0ntKPLPC3jdDK5OE0
C7ShoIUplVqnG2juAkfe2OfAxtGvJfOwFXyZ2RafGAq9s2wCtGO6lWcBS4vtLv12sza9rDPM3EJ7
SAC5zozrj8gZzrc0Cjzre0uGzLGMDbTyD3oJPswlM56g4nzK0ykXXazv/oBXiAk3yCaSTaViEKax
py4kcumM0PT+5cyubrOLeub8dzkNsZw64BZqFfzA9MYHTF3O0LuDw/jQ/pK2oJTkh6DaHBQwKCf1
9ETfG5lwX7xksuqzI2wcY9/W5I3K4T0ndiSu3M3H33a75lZAKCkccGLFfya4gChnrW+/tDQ0/2/W
zBAO5QoJoH647h3cCXWVDDd9cnVUJgXlKVXRrn8HhJ00Tn7Aick5WyHdzBvPz2aNVeJF68R5A92t
P1QrA63cVnJvctZdEfiqHbZLzzXMhsGkUoIKLWjlFBgp9sa5jkdzVUXdZaZ7Uj0dC/6s5nYf+AKi
qQkFhF8DDT7y+I6/9ClkFd5kxg87TqvJzpX81OGys+WTFXKYBbHUBWgSqA4l19XxvFLs7+qco3jW
RyCB3eetiUmHo9J6EhAZXtqXV8qDS8BZLIfZ3aG7crpTHV3Zwf/wNFi9ygUh/hYMDzThPREvptZH
45FxTnKYG6PkA4Y5ChG1khJs2JA3JocFG3Sw8hr39MQyo+1Umd8R2gdDfCZBByFkn5ltSZOq+A8M
iN1mCVjOXP1d8QSwTtd/Vbe1n5Zhnn3V8IONL9ZzZYJ+4Ul5OMklcRPc5Ih+J4OrOn3TTkatXgGw
rQko7aiZ+JEJanet0laSf3lkUWkpVry6+Bbg6gMHctGVa3Gqu7IGjBNNux1b1tWNGavCU1zBGgR0
7H3I/CgBwY+4tBLDID1s6mntgbi4ktD3LzO77MNQcoRmnD8iSQ8a9ki/ngDOh8AmL+DEdB2EJZ6R
O+DlkwJDF8hncj6Mq5ZDeIeHIp23RPiguq6ESoKb7pSznTgZ1GcR+FhlCsjTdX5LZIQY6UJt0WFb
lby8eu3ow4vbrhA0sh+8svQ7UGLBYeoMQdUGsYUPiW46X+oMthvNRrDniOtjoPFSMPRaoHrqxek+
c+mpeiL92Af/+ttZ7pPR7mvtmu47tXRIV7gnsx7qOgTWM6tE244VeKlt23Kz1bMRq/O3HhNFX42I
8nEKhteFJwia2XXZadlfS9v06Tj1/QunkGddcAPKD8St76L8AY8vckbSE0gidTfO4K9NwagiKm+j
J4lmSL3ls4KWXbSVitd2wFDsvyLEwfYe5x3I/6ZnlwUca8bGhDOusVWEXQTkUUeuiFwtwPFMIRJH
Ja8hnrtg0SaueRGk0+Nk2PX/D8zaBgaAWvunSaO39KgA+R0pHkRBFT3p2OTHLjIOz/KB5f5XjZXd
hZb1aUk/8FkbaYWj8hTSv7ef/CwnEgRWt6ggYQUmHNQzGmviSxz7lx5aU0u/SR++kxSdD6vXWZjJ
Gzfz8UCXZH/Osdq63ygTgzc9lmwjPo4zrAD1sdl5FC+QHwg0dY2rSduxwq4LpxjPIscOzh/UPlz4
O7F/cYvS/Ubv5k7v+Xlpz/aF8td56Nkcc2qIzWUjAuzAdUNyiMffe0DryZ5WgI5VK8vBg4FYB7XK
Rt4faqYKlLu5R1ycvm/4ZBF1cayn39GqDIee03Uy4ndctEcuJlMoiVuIpJVxnSrsn+/ascrP0n2P
XuqtdiaB79c+rUvLsJUBlFo6tAEB5cmdffH8+lzmeUDY92x9wKYsVxQOank8WZIGTA8qt/zVfspy
gVa5tz+6Bd6mPplF+NZo/LK4mXLTt8Dfp5kb73nguTHUkZ4eJML6y5knDFTEgbOSgyGB6Sww6yee
Rm/Q69FI6yJDm0vEyuPkpJzZnAiFDaba1mdLppWLdVjcfzDzv833gl0oNMxjmnCKx95KICSduvFo
Iw1xUan2dtysJSwCQ24Wzofe9YWbXlgGoAh0UIqu0TNC3PRkhfeSe+1HbdvCZMXYWbRbJXFKPaKR
racSglJFjF/4g/T2bRmmM/H8I1B7TyYBAX4eIBk9LbmVJoqWI0OCgZG5ySdauVAzTqKwqVNHRyUQ
2/R9Jf+3z0DQsi4Dab1H/TKq7NwG2YB7gixtKE1f/XV28ORATn7sISYXiZi9RKXIR54MXRLMpU8G
1iTtphBvOh0WL1Dgp4sYvve7AZppFIgJ1NZD8XIFmxob/1/9bKdCJgdI59ZzzUQUXn/blYQ17K8F
oxZWSTGJjSeeI//nW31/zeMsLQHVNmzEQUSUD0XFzBnbX5UtZRylrPHAKjj00fuu7xFL9KmQZYpO
G3gweDXowk4xUVmGy0SwSt7VhTO72YiXE7jSJ070uvmwWGZfGRb49aaaK0lbZtOTFyH32jjdDtG4
mUMXvwgLTePNSAMFzj6nFrUDvZodM/l5+InjwNfxOlBVgytmRhTy1ipdKHy7fgoE2NNXgscc0EFr
BdVUmN9vgpps4DsnGgDm76YMHQu1wqPVkSWPWbgOYJyv/tykLzzvh1AxqRw1CPMExs2qYpB0GbAI
fvSV4uW6Fqv+d4NXAPEO19TldHsVJAuh5jk5fW3TYigyBhsIDffZuZhkQg0T8n7RRzHQGlKJzygX
qp+eFXVZC4PKNMAr1s2hdkRzoSjaNTBHnh6Mspe8Zo9+m7e0WUcalbbHCACEUM4XJu5FJt6t96qw
jY5pSTr1onx9BX0AkDKKbJAWhk4BvCzg4arlSmnwxP+tqBCw298fCbbwwneYhdfYH8ZVlvKjv9N7
srqKIXSvcpDlCiW1gQzf5TUkOKqTz9XY08a0FcMI26ttMwcspdvWUf1bMlW/BgUYiSbinT28GNTg
NdOhp13ltseSQq+Wf6kY5CZbkqJ4CHnGifK1ODZNEm7ZAWKNbwiAts6Hghz1MthD8u0vNsQ8CZ0L
ETSuzb0JzLeFzc+KdNMnLOzejEEmfFgkXdXiuQJOhTmBhkaNPcFa3PztzpLXm+zqRFJQISryV/gw
0vplcXCDMIugg2rUh66/ib/xhX9VnfyMVIJeuwq/5hyXiGHQLg3qeBrbp4LT8Bw/Ybv1FMaZkNLn
Q5J7a4IrHiypwEegG2JspolxkhJRJbsiF1RJ5wTUCafdmJKtAcJgICyAIzvQHEHCmUYjDn+FEa4m
hLQ63tglJGJDbmwXvXMvozJKLTOAzJai26VQdzJqWfzey/vY4wX06TxB3m5AKqfq1M6ri+6/AP0r
hNX5DSdJ7vrrXX/wq/8Wxk8sda1i77NLUaRccpmaqU5xN10TqdeMyMsuuqecNlzRCJulxNpfIOrB
JGl2PZ3JQmc3Nkhs2mWvjmxaS3k4oawDbk9Y6bZZAbYnLdd9c85dqILr4MN1KbtQ9JdlkmOm99DX
mmQFNlOU95zXZE8daPQAT8Hgqwqlej9H5hMb361GxBbKCJM8tqXr6KxQ8NfNcrYciDod1d+GjMeB
v1qFuleu0rX4KHVtnF3ag9UKwdGX8WETeOKsGb34hFWr+p7LnhIsK4QUcfjiAh0yQ8SBUuQAXmv6
stLKfepJkpD4RCoAe8/64DmXKUbm6UgXzvYyVlXBSJNmgwzU114vEOhTTUItW8iIJ/yyn73E/iT5
LICB9nJgJ2azCFKE0y+Hp6S0UGfvjVOcRBm0iEpplkMfE/7n0x2VTEnGfdvG2twWPOIFnaTJuQCv
SgCx5mRjZwC+YJgAwAcVQBcz8/o9apRWHwRA6wG/QqDiuvaQHH+CJnJBj91g/RZF6YTUdZ75p1EW
e0dQR4K/iFBtdnx9mEmDIUZtY4cyxrAlRMedTOcHwbs53CekWGVPN7U3qcdrbg7MxFR0bbEhvgMV
hhuTF7UrOrqoDz0GXuNk/2dvavCxfhQMyDZYV8E78g9LGMvTlbd/q+wo7UddELN72l8Wr2zvbLpg
SnmYHla53sSPa6jq5IdDd4ige0j3UAb1lNOz1M0+pBLyuJ8Wa+PqmHEjy0bKd6ueEvVXil4UdkJB
OoAtO5w7GUZln0fUnqYrCRpLicdg8Zs7Z+e1R9Cs9g4ZvwxTrsFwQ+K0wTrdv1cQQOoTrgrW9ruN
dIZZf8L6m8oS2Cw2wRdHlErYre1l5rdBB2EnT0dhvQwmUkGFoKMltVBtfz+qDslMeJg6aSNM4hHl
0AmtZf2trqMMbDP8ve8NgcowIxzGsCyPxszK+ufLD6hft6K0Sd6IxP6BBUI1IQsQmhC/0hmB87mv
0WkQRJH4WV+01LpBKc756sdTJ8bw0Digm2IaKiqvTAD5Orfdod5eK7yD7WYRSc3UAq/492s2QLlx
NCpwbg8YBZEVj1WC20qDKu4bF2f4KX39KaNjEca5BhRONpl/TlwsTX8t43YyhApltNVPZ52iaRJp
lDOd8cKYLprkEe/FV/dJVLOLUpr35du/yqt9/UEnc9X1268WuSp7uYv5w84VZmQWy07pzVKkcGZL
syeqlDYO5IppGsMS3aAuIRqjalzeOv5xYsUdYEC26qyh+PYgJ6Z81HIWq9i/47NPZfYkPMtaBm0A
0pMG5bF/r1ohk/7goNWhiv57s0F1QL7yHR6xSSC5zkZBS275o9QXegV0lO7WtkmEh0utgxf+3Fgc
r0b3NcglqB6AYj3rqqoOJrK7UEY74KduiqRgQjN8JswQXDrCgyipjHDjQdeZu6jJovmkIum1gluH
StjHNOdHsdJagNXl8uYD5WYympB4b8ymKRiZJYq+SnKskkPnNEhtbSZGPNjJDgxLheXKhetajbed
AdAQZbHrly17krDeCJ6d6I7GV4ipLu9tYk4MfyxmqsVQKNuzdtmg0Ua0zoKUbe6mbe0HPITLliQy
0auvwXQYxPv1++3yFSnJJ304yuA0Ev3Da/R0H7PQZ0NsWAZITosbr23B3JQzmHUcZ2mU59J7PCzS
83YEfuKxc7f+lvdNPuO2veGjoGI6L7ukrI2al8FYCIMR6gxb2bvBmhDn2mlZCR1Oorr++BuQ/t4k
hRwsTvveoG17G3l2a0nfkCnyw7Cpn/cCUEh5UV0t+7KWJNVzNHGOw6trPkYfpUH5/wV5NZA11Ieb
XY3a9qiZ4mI3fUcY/i8ou+2kl8vTTxh419tJtqz82su610TVf4JOwmNdYHZQb3CcwUv3GqH5Z694
rUJVFS0m6j5jurklSHMA6KEx2n1e0s4LPnFwoUUFsCMNex8XjMaOGqr83QZOBbFOV82mgyUvv0l5
6hTbvc66LIcxhYLJbCClwxeqM7VJj+u5Agg3nbLNxd8OZ6t3CLL0Oxfqe+MsOadn5+8q4vusehL3
VbjxJ+TRvsT6YGQeljgwY4q0hGMOPQeazx/qe0IqCPOuSs13BpOah5sllCHF7BZpsTQ4nhs/cht6
Q0uNiG8bEBFTZd/vxIrdSrlpxxDgm78+IA2VFl1YeVB1WBLrSQ1RB2ZZNfyAwgNDrl0UCcreKDGo
PMLwiUxHf+dXhN/aF3kftPlsaO7Wjt8bt+dUv4tSVN92dijOTTNsxAadX57rtCi42+Ew+xlAxJsd
SVq7jRgEKfnWTgn4x46uAi2MYYsNit+EnXXUmmZcAVujJzCAO8sGE4wc7RxoeH/i1yXcxGldSHwB
itqo01bey9+77i9cVRKjrDlGax8lGs9tTB4B7yPhtnaGAX4L6+VXCqTrCqnSgmJTgznG9L/6rqLy
yKs66paKb5ERSc6DKlgLcOf6UOjCw/b2F8thS0JqcLMtUzTYPdIyS7E1cACVkX6WA9ChFsbX7esL
mDI5JvoNwEVtrIAH0SvxX2C8JLujBfS14dI4rQTwmu9LFe4o/3vsCc3nGWur/mWYbHxEP77S5Ax0
6T5DGxyRhXMtBpcSL/INUg2Al+BO7mZMDP03ufavPGDQ8s7NlIRwNPjtX3AiKpeah5vxjx0bR8Fc
NtQxg7Y06CDlQx+8FXfsZrA9PhdFE48iP3NhpOh0TlRikRp6IVINuhInZNusO/QYxPBxV2bxqo90
qc5F1Q0NZzQhCzUeH/hqMX82NjPefhR4vdk2xQfxM8HXB+W9OikcAhXCUZaH2iIj97BQuJeLEDq/
2+DkaHIgHWgJDquqO/w1p3yGIq3zU1OmKWUtmZPmuXgARImfyfsZ0h/fcBsyaApC8YzVMY9BFtso
O3yomO1vgvPIY6uIez4+d0Yzxctl3Al4nCgtnsLFkTQ5tf2u2/8+MosnyJNAvqtJBtwgHEouHUmL
zdCSpxdgcMbgU8SXzUUPDcKoT8N0KtGiUnrtAgZlFqsM5aaruUdK9wh2mNpJmCO2beMsIlc0ZCZd
aP++hJJkZyS1D08h8QzOXyFY+pQulLkxQwUbIfwT/zBdqSkJ3AKHeFabufbvtdMLsL7+ushUjoks
nG2m4bWxqYzLf6UmCIJQv+AuV+MSR58SceaoT/RIFD+sTiPDfCHQQffQxiXK4JHr93H369oW9NB7
Lxvw0UFi9kqM9rXOeuRzTKnMvrR+VLhSXNMPytQSCDeWuhukt3pS+dHcYfZXseNuHoXeDCmCNLd4
uBs+WRzvh4L0w5RoUsy2o6dEsSrKgt8jWIb4wf22QqhLGlXPDMODDam4TkyE62vJX3rHd/zCud+k
VVZ64kZwhnVMl95C6l+RQT+FAGVJ5sLWt8k3COY9hWzREwKzcwFQDruEca39UAXCni+9Rirv1AtR
Y+mEDszJa51GEPRYlfPGNTWkUUt/9CODcrpfrNGReBuLw1rzNUpNSdmcl/rkfmgPSfRfoHCdMgW5
YSN05+tKF7fnz10fY8/pzEgP4QmPiboKcuMiflZJLjUkpjYggSzCNi+2vZK4eg0GDznVpPmCVoVx
HRapPwiIwh2i2c/BV754ZsIelD3CGf8cksqKXVc7rUWUMKmToz/DPJN8tn35Pr1lX+8UDsD6hoeH
V0PLWPXStqvEsswPfRPjOiw848sLAXZX7YARY4mDbOPtUfZS5KgIoaHP5ilgZOrQv7YCFk9AnVnc
2BUzSDZYQoxxNbWxluVeKh63XsVpjaBAC7Rp24Fxzk5UD+8xJRQ4k7zvAtZr0JZ1z6X2m64bpTa0
tg30XcgvwSowLbDqnlR3Sb68VECjKxAOgPsO0y9iiqrVWHJgky6g8rQgjZFme5rxRTmE1Bd8rppu
O1fvy4pEu13mbjAliCItRT7k+DoOWOpCmi0wPBDrwSw8cf/CXMLh9tTyo+7P42WvQ/puxgR3w1z+
F81yboVixw3RaS/bBKbyDpMwnV4lnVphS/CyqkWyHKEzDEPRacNoIa/o26/GiPyjdLLV13x9sFj1
RQDS4iPUCgE9Q48QwlX3OVaQSHOgI0qegQ2P4qZfQOoyZ9LhyENWJO1HlwMtBT8bXKB8J1TGk+an
OI/rDwv/AKf8arsrByJ8hifwfR/qEV0RFAExS3eR3iKfgtbVH0sjzrQnZLXKpJx8nBeeKd/h312J
Rj/Luh2p2MZenPJ2GiQMOct/lz5b6srHrgMpIaix+s5NF4eFVhjWUVLyzLERE7OiaAITwYmufDU9
U3VevlFEn/p/f+ht0TYIpygzAViBmoeESm1MUPHScMEoIwkphqJmO3TVa3KUYHiItWhNTklSaylN
uX39/4QKm3rYmzcVEiC/DUhyXbt/K5QTZUTyFHcebMNrQ4TEmPKSOFSwe3NJkXug2ingxbGSuKBu
5aqZ3HHym4aJibjjBNsHQhTueOoeDm3uqsNDtxzlOTzK1HuXAWpLzbGj4N5g2mOLZf7W74iT3pwt
Q7pd1w5DZVMeu1CBzAfvFkCWHn8xg9NAedE9gnrRDpImTmts5DYhYYxlJHP7Qf4EcuTFqUmdVRF3
APrzOu+33UMtdewLiyN5zd5nmcAQpar+kEdFT3ZuFXbxlr8gUXqVpl+d4YDFHFWIAPII5Jghv3rE
MIk+Xy2KdMG0W49V0PEAWEd0vpEeEFo4zymzcS2b7xmCZRSJr8bTyNdlC/oeaSl92yKCO5n7RwGd
iX0uMJ9ooBkSbPuUo+mQ/58hop7D8x/But4MW74Yd6F10esjy909qC9Q/gI18eZ2SGFPLKC8wfH3
f77IHDurHO5FeRewCp/rehgcMEvfudPlrLPjduZ15xCjW+KUKANVZ880e32A9gcyDXsd8W/rGH/P
SJ+q4Vtzby+/sQ7ttIHMLVDdsqZwr+5oGfflKPElQ/y5nkEtlwFHMxmHgfTI5OAnjjqZR9iHoH5X
WDPLeaztA+MmemXFpqkdfZ67RouUOgHkNd13FnROF9byTQrrBYwwmjUlA9PMiEXQLCCcwVnnYh2b
XAB9z/UeHVjqjft2zptqgvcZdDtpkNiyJ/rc1MdeT3sCL6GBvB3mvmsOAgTFN0VtFjffWAEHlRys
ZvYVcmurCOxAaVzvjR7X7mMWeEx72M5dmhGyMg2VB/0147+3yQFc7qV8bSPDfXYEwzgmpKcOazfy
n5scwOBR4+qbz1tbGLmvySLuA+2oOI+QlaXjZtjchgfTUCnk5Hy8bGGopOvxD/FC2KbbnRK3nmkh
5ledKRyjcu8gDLe0YyeXctEYmDdzQeGPt2O38Z9JNZ22LwBTiOeO3BgcZXe40pGLkLJ97mHyLuX2
d0XqLz4E38etCDvoBaVJ62bZAhYsCKAOLcQ4NB0PLsOPMXDhCXc8SgV7xStOLnjy4G/6YUC/LLsB
YO+1IIk+PbZLGf7Pw4PXWRyR7naL0xaylg1uJN31lCwvfnDx9jCtOINRbH0HPWvRiArOdW2ORxKj
59AAazCSTAw9ZESdxGgbI0KA1v6zIu3jkXZ4sl5OfisG/y6HTAR3qHX4ViLejtua/qIbG1mHSOYb
adO5IQwQXM+Jdeoy3PN0KAWn93TLakvpUjWNEnnEjOTby7McHa/t2tD5c1SB8v4wjfkYu8LeTF2f
++YaBfWVoF5fgKQL1xZLuA7Dm6Wl3R/bxOTsAbYIor88eSwhIHKCS+k2VUugA0M8Q6I76X9L/Hby
Ogz7hBy4zrSV7izrw/GCWJB45o5XDZBnBFbB5fxfs9lOWSNb6pbq3/dnMzK19XyBMZqyJNOuvKxa
MheOqNfgUPk4XHB8Vr83kcFVsRRPMvtuJig+b0cRTiZPHCGZ2Og180wItKufr57ZyNL2+3erbC2L
/UhTIU0Ljou3vmrWqlAMsBFAcLHSUOuyxA/kHP+wznzWqpF9rHomJsLuxAv7KAzxRy1uu5fuDrLS
aNcmIP3jNAjHVh6gqNnH51rE9kV3B/cb2Wj6ShWit/MVjmLrQoitslgTwCjxIGXJExFAcx0FK6WG
2MPtxvDhftKgtx6h261ZVKuahe52r/JSeCLVKBie7Y3grSwC91L+NUnA6TVIAfXcA/aPQfuDC9JI
JOzspfcufEk60zNdc6mAt+GAScTUh5l0Qr8rRZG1hA/7f07UjffQJwzQJRH1R+JHUmGwbhF0m80S
nS4qKC1Vp3TeMKN/t6DEr4JEGE+6ku67K6aL8viUULZXhBy8qsmxI/A7eGCNsKy5b58pSqnKOGEq
EHVuxdsqVYD9FU3LYP2XPTXx1k9WRW1NcZ1dgzJSqnR1ydXNYm8l5FaWz1CEiPpHOI3KVDdNmx5S
EJnkiZsurYvUd983jEuAk2c0z78qXSQdvVM3HFZUMv/nBKIP/L7bxHzC/kHi378apl15F3qMNjgP
3RGxjx28aHMcIa67vnXuhKQXqv66QIkCFg8/p6+kyP0etigX2/YxoxaFq8hoW6j3LfrOiapvq78o
DdVaUv4kv82NSC7XNaVKQ1xk0P/Tju2pxoxyMlWsbVqZ17OcuLb0Pky+u8IY+EmXSnVysF1FiBd1
UyFHfXfys25yTBwFvE5s5nNGhwW0qZI3qFReVNKtTeiLH92fuiPARW+YOqbprrYlLxQ6GArCtE1C
a+9pSrKHtNZtKNT1fA4tKIcmiQgjhFwBvoGMB3wscBA4gL9fcHlVCz5wzPorXt3N02cD7KhkbPG9
jmFc/jyxXWOvz7niGJpbPAByR6WlwBP4OeSroEIaI7oWOgepLEb2uxaT69dt3uBx0mUvkVFSsc6x
VvlddNXZRsgKJJioMThwiZDhMEdoXvYJ2sZHEXyO6vAbvG5EmA/4TwC6lOpbXlw4cWqwa2CXCgAl
1VMssccNGAV6ny39Gq/bSeQSrCW5+NyxT/90f+2YsXnQHmiMy5N1U211QmrgXyG8QybETFFgdl8s
5jXiGGgiPdYHjjzooh3hyEZjU0u7lhrw4d2OwXJd2+vvz3Nlks0lxdJmDl0DZsuGUPuM+rqVpDhw
+puLoT1vvpBMGQVmNd3sUj7PMgHco0/jgrqWwXEL96UgG6oEb5qr62TMJSJOAa95ctCgNgnO+FsZ
MYovrnrSy3E+renm2TRhzsQJkf8SBWalMhjikgFImiyblCFkX84FpHWZcds01VJks/aaIxNWgONP
uEDBBkXoW89wHwjjtpbnA7jvaoaj/MJV77SJiVeszpuj5b9SsbwpP/+TtW3QIgB8gw5vqa3/uHj7
XNSL15p5J/pqLUf1g9NYVob9EHkcqzlmFSHqV6N1ZApNZzz03JK0v1EfechL4EJoNdZ2HPwKw0ou
sJocNJ66G6rxMW17hU3NCoekGSngaa4pZ2/BQ94cGKovoQabR4af8juCG5lVFOb6TyAiLZqH04z+
gvcwBqBf1583t+dX3PxsH7RTI719v8ChiWN34jeg8mnRRg1UL7jEcd8qmeimbiU89mB/UbfPqr+4
yV+S8Up5ilRRlnjcD1mOu9dPrqeV3eA9LW0SkB5ZIw/e64DWN7bzXquM2meJhJPPMsK/DBZESdFx
EQxivr9mf8mPWHg3deuet6g/7kUN9jxVlTkzTswaVDRn55oGM0WmfqbAsTTa6lSXVMPaHoTZ6uKU
r/HipkIlcdeB6dTjuNMr8yeL/a25C2ufy65xzW/8zpr3NEAv9O3rygg1hmmnuhOcRZLXr8AUlyjJ
9xapEJEC5IjhUOuFFUA6cWoF4Zz07sDpOcnJ52TELfOqn58afOgvUrls9arldtCv7tlhnLiSKbg2
Qy1MlkEqhvDLnzK+/p9993F8cu3bvBDRlbFZ7+9Aoii8PNIjiXMWQYq07zt5m1F71/aMtWQ5RBmC
Py9Q10v7pxRH/8pP4I3kp8hUtrkokW2a5rzu4y6huGYvl8nlvCg5c5i3jwlDQwKqEetv45PXxfV1
jfnnAY9er1j3uYfC62JK3VrN9SsS5mFFYqo3ScpmrjoJYoab1Wvl7ItJe4GtjV/Y2I7NQ7+Drtrj
wbPFf2qN2+FLof9ag+Zo/uh7zcNfB1G6XGZg22Nrq+vEYFKULFZzpe9UPb7E7UXI2a+7nJvr/R+X
Yp7N6iPJslX4QaDFqFowjmKdxd7gKRsBbKWGduh38IGWtxdre5Ytr0yWD8+PWudkv9I/Q6wclgFc
o7v8E7GsTQjaG61kXqcHPOtaIHuoSeG8vZhukbV7GCbcgh69XcN/WS/rj0F8Cmp6+uO6KZModUFP
TVRx2b1XzU0UVN7q37qP1j64/1JXmCjSf0JOD3RgQ32E4Cn4y8bHQCVScNmrBDuYfOMob//qBqOd
9nd6fWdwCjM+6H2w7p8zx4QH2QD9Hv1RLAe5ky5bQTypCpb5Px6mEX4myIsMCNdLrQoIBxhNSQCt
82t23+OMRa9fRQkmXKVisbntWjTMD+/9HAV8HGwzKgNhdkrJRPmXOnNvCVOh13VZkV7ApBFvZ/V0
YqIr/MFJ9DmRlcXYgSUeLrQkyIl8KgFn+awNRmITP3hUUvT1BJzhH4uEJhwE/EqVYEJTHSn9btyI
2NG4S4Sj1/Xom+I0BQmOYSh5JQoa7paUdzvX/eRsmriplDBE4UVLpMreNFMXZjA0rlFGu27ce58R
Capll7L9FIg5A85c9tMUjl3VqHpE2cCl6vkNiRv91ew+IQfMlj3jWJEoZp7NoF4aIy4kI+V2srPS
1xKhFxYmfxphLeRSXjaNVOlq2CaTW5WrPn4uGP5BiPTJ8ql4x3GT+J5QTXsBWOFIxs56f3fGeAbS
2+OyrSxuLNGRVc+iMkly0nRvtyOnQg6TlTFcVrgA7jmiQuVDcZcDamIl1bAPycFg9wkZt6x0ErhN
Ftd5hIy9V+hQ0Wys3+o5oxG0MnEa284dKyy1Qcpl4cd6cWMD9s1UkMW8BTmcywUEB/bq+KXO+apU
h4xGcBuAN/dO5+lsrABnLJ51CW+TlIYoNdetzKPRI9+cu2bzcVBLNCqageyclHeb0yQbl7p/RR5r
C9OxJxjfQi9rzMG5j+cJpTHWvLh4bi8ABvuEGkCSFOVRW2tFc7T3f2Eo1ta2ER9ofNWUpJ2raMHZ
BzDE1O3UDBSzbOBDuOj9WJcTl9jzgvYtDsY/13Ky1B81VIheszzdKPsNZg2yxM706hXUAeDQ4qZn
PJFFuIdbxg6ls4403O/25sPKJ2McVYf4rEUl7opPNfVFAvesZVQZOocPrN4IQ583Z3DbD7qem08D
V6m+qMmcM1mF1rkFXtn0YMjRoUmCCCJXeq9wVPaZrT/HT71uMjN45Kd+grWqqUYOhL26MQnjIx1J
BqBydqzQoYQxFtgYS6xPXbg/PeBi5JdE9Yuum30fWJr5vvJbeBHjUX5fXHphW4fJPhA7s8sh/yhA
W73zTRGxQPclMY/AxwuelNKALALlHJn7mfEe+GVUl2o1+/dclF4XCfZMnjK0WwHIABxzuYB/xNUe
Q+Wndb9eA0/UTyLkcFPCrKBVrJKJ+S2YWvN2PhSBooCj69pmNbQLnkRO6iU+hQepeALpYH6IdZIt
iVhFl0TVzEV8mY+mht9gzei2uTb4uFA9kBDIp10N82HkZdgpiaStZCW5kleMKX/LodM1WNsBQ9X+
6mV7dbD4DnXcux33L0kCAe8R0WlAXiT/P6sXIN1KP3SggTzWDHcxaQ2zXfEbxFUldPC7Y0+XJ364
Tu3Uf9rZDqdQy0PomV7qrNMmWAF9K4WopRIMXYqHl4LZ1/OADT7bQIEwK/C1P4dJ4/IgMm6awNL7
T0YOyUXT8tfORrPRvR1YhwzsOR0mrRFnlfwUkyHU/1t8DsFmxc/5HA7bC2Hp23NvMtS/2yxtPPu9
rNUq2SBmOaIyQXqMtXKE87gtr9wjMwZTrzEUBhjPB+fT6Lf+w8pcUCwnTiNk5wuM2c+APwfLi7et
mUdItPkkzVnH74Q2ZwNq8o+upjmj5R4W4P2Lr4iS9j1IKpaOr+4AvEEpJjRUkIUuNtSDZ5KqKz11
BQHMI7wfObua6VdjU0ITMj8L3RBP0iRtMnSBxA7Q/K7VkYB1qUaEaZAEDpg7JNdaIfmPZuY2KYDY
71T6lBbngCWWXsTefG3ndzF9MmdjUODmzU+j1tzRo60LLAoN5do9Wak1xVQonqn2KmbxhuH4sXx0
nJiUVwhiEJLP2DP2cX2uEUDxf4U5b8vwBTq3bwQmDNHJoGUTqEWS/14pgX/SrUUqBO2PHX6+EL94
HJjAm8lEs0XtMGf2Jw9Px9gxk8yBEIX5z0eRLHe4C4GZ/bAscsD8vUQ4taQ18Xo7zjTf2EejV0Jn
MQNtV1SWPDPcpuzM0Qsa7z6Ju/xmbMVTbPvbDjC+lIO7eDKOnnaeE1zkgm4N3csjTCGtO3jio3ik
GApGeP3GzEz37qWcS6LVTpmNo3ubuIK1Y9aDFdLoZMReRy2G1nSnR8IJPc7sIGsj/8ZoKNyeU0Wv
/CfueggS2Wb4ZLQaFRnitS9VzdxOJPvEYWIM7DOMgVkFulojsZwmzAKgBPc+v+5vWLlGt9YbRYbe
8pwhZRSw9Fm0dVjkon79L0gALRcyx3X+FRTtviKcNSvccPES1DteXf0aBKtoFj34zX/em6wLf0CJ
YNMmoyEQfzuhPffgNXsX4ao7fAlax21xMoWBcbug3FhTlthgqjyyTf/Xt78zbx5ZGm+1grsiBzQe
xVXPX14SgQ1kjEqhhB1QeVenihRTOuSPglJ7BOV3cj9LiXr4Bv8ZCSCvYg0c1i8DOMnbJG2fFHtK
dBN46rEUFY8BH9sVmR2SsujfwPqLmfW9cvnZs/eLBumZUbESUbfHWodpPKLkwXNyqtRymnc+Z++y
8o3yAwrCcCGWN5qFhF1qqva5fcJd/ogbvIl9dX1fo5/9RO6kpYcQAE+fcSQc0K76Z2TMrrYdsENJ
z4ho9wiCGtpnHeSdUQp3gZfp7X94qByotJ/8T0WYN7SFbB9pSWpj/I1gNDAhvXc8XorhAMC4KEZe
3IZoycPR9qhmXPJqOBCLX5EnRZWGm6hYoskPIwlR+iceH1V9p9bCPgGTAxUZ2tgHBa4fzkANJIZK
Hb3zxr8EZqFJ3QS6JJIKKD5At4NGL1GiQ5FScp7vV3l2CpjdERPPG5EzzG39oa6Llxt1U6ceDORD
sAFZYWNYKhOaScT4Yl7qRQOAUdqiOhTYWLKmhiRQV7GvZ8EWhRFT8rrAy2hRNKrJyYkw0PAc+sCt
OwWW77eDNXVN0Pg1Ul5puQXeDyen0WWDv8T9rba1eDHxlaSdYnhRnbjWi5R/IDeqY2ekNoFyiNh9
LLdC2lIjJFgs/xvfoGHfuNCag7r/PGa753BNWwtsYLFvW95ztx0i6dyavYP2ogqqO7hVAu/fvscJ
AUe4szBQ+ETtlVaKmTn0GlD+TXtmmdBjb9X8GqIxYcBKN6vmMW5+IHZChW+T/mG2LZWMLj3FrVmy
GGD7H4rdKcXnCBgyyJXGhlOb9U5K8nsV/Jj/uHRm+rTTa0K0WavlBI69pFrdOhwH0A3I8jx6kbGd
L91BDlBWTGk3//5JZUBP/N3rB/Jpq4fgtDoNdYwvxlooHaQyPm4npyGVYdP4tY1hXgQVM0jKnLRJ
Qv6XgM5YBH6sj6dLZg6x9MJFMh5YGMTB/Pe+qvB3Iqmra4OdQN+gulqkpfYQj3d47IAuVjIomRSD
2i2Lr9sMxTjdl5+1mRIsRS2CsgrirlAxNQS11W6fMSoe5xndhyLQrHvRz2L1z6aRxj8uxWhBsUc6
aIUX7svfHOTikQgiQndS1Tqc0MNzpTGIExt3lFnFDVa8JDyJNWxc0kTGLVt3iOyzZOGkV9OS31oS
LwSv1tgbVWgNN1rfz1oDL13Y+ZB+bCfdlcksS/dM8v8/iXxsVsRbH00tfu+o4MxdLk0q+rOz+65H
uKUh1hPnMIQwJ8ARDE2dLYg4oH5F+Y/EzbVq8d8pbwSrsmTg5BdAutQG9nkSED8rsNgCMTEj1aEq
w70Ne7QXL9HjN9NXnLVbpQlBb7RRTZmJpHa37fwSFgk74GC+8Fws7wi665EU3JZV/OtPVvqJfYtX
kmio3bA4uCqv4pbedY2YvglX1I4GWKQ4UCaSKa0UBNhdbtIWl5IRlEY9Ibbj3bj7ZrPpEgoiNvVW
0YJKaqLJFoIbLXc25TcuK36r9DdiT9r2/qcoxLvcVDcYRfGeak8la6NXo/jwbh/AF8xiM3shDo2Y
M8NqjkGbwZ6pzzR3ME722w1m3d4yc8D/XXjWcCiFWv/MGbAwGKNA8VzJEzefnP3PjcvXxoysPVtm
A5BSd4AJ5TvC1yBQg4bphr+LdMPL0GAguMLJnXzf2NsS2WoRY82V8VvNp9Oy6fdnSGPLP2aNi2Lz
XrnQh0fUXZEC7JUgnf4eYh0pksXALYiPVHQOC4eWFbaOdzKhS01ROlpNXh/jtVuyPR9anJV8Kxvs
T0oruXvITMmCEUWJ+TIPqwBmnAfWQuXUaSlBfIUFbLwvewwsbmOjpcsRIEJbqfKblYWcatQ+YDRU
KIXk2h6OM88B9qLN8dwkzx9PGNJfQkNb8SK42kc0xHFbv9/LkekfwkokkGf9taaakKqaBDD0rjeZ
aJ1Afn8/IDveO+stEwjD2XMvPRpcLszo+FNJY7sv7B2wuxGDmTTiBRdBxhshT0zsNcghiJapd+c3
6f8anBXYmCALu2soP0D9PjMR0hAjblC3SLSLiUMeH2JC4EqrSRsLkbvW2iim7E/wf/J85qBgb/qc
agYA8BQH//uYZtcsDlfv6xblcdQTId1OyQ0eKIwTUetUdHht8Io2AAj2r/kE3Hc0IK9E2cZs/Qt7
YM3hw9K/9WPhaXyR9aQnNFZvNAsYowWTTUS3SMKciRmtaRakMp0xgbk3cAxX3Dix1UOOuzuTvhkR
japzc2sAIBrOCz9M8L4stiSvFEL5R/eMiPQACZWVjXZqtBwFagPNILJunvuueKwADAS6KJV3pD8E
QIFiQ3xS/KOqdn7uEnYUBSZ/JadKlXPHtFGKb80WfYRfxH/Y8Lv3W23lJSghoe6UgPHxZby3uN2h
P0Zxx6+WfI997AOuA4dzQ2owbalP2CapkQwbXf8ioO++3GkO01xMa55MjoVQrTXqCDEnV4M52U2u
hHjpOslKa0tvFxXdXh+z6rjsmrI2T1DhXiYxmkwaHz2UbXpSwsGyt9JSE/P1RqVYJC8wvp7774z5
jEAy/Phb9RnDn8umEmZaLLXmtW70xIJXQSulxyH9WsmZgotAhVsZIr/04KG97akpHbCnAzaK61QU
FEWDQXr1WlYXtP2hBTce5zCF3oNXK5DahflQUu+LpvDO97/o8VLJMOvL8gb3230ccjdtvXA9W4JZ
etIrPUf/JT3jlC/QWFfx2cKus4XkV1RLEh2PtL0h4fDC6nNmMWw3lAgk09Usc3sa+HmpYNkUhkW3
I+GGwr+o5ksC1ctyC0hlBXiswA0PFPqMTFt32ZiPZWQgBqZ2vH8pZGgz997R1QljG1R+2OBCo3Oi
HLLnstvSMA7tM+ZwJdBq1rEidByrqt9pq20bpknXtshayYCxIqA6wI7IJnLyK+wbrkQO2znbVtln
paEyIyOUATZQENzQlv3VJZ3oUB5ksY142ILj/0mOt9Esl7iHNS8lSQ/425g3vX1eBQJeGZ12EZxN
rVb5LryTg+dFJ19fvNCNEWXMXwjo2XdEZ4e2Aj8AvxbFzwA+JCPaGxK8cJFD42U3eArLh2upGF23
I8JKgavcHYmgtjBWmXdd83a4yUQtQW2pcnei90qanU3GgIer9gtnri7Vz6Yb+03el2K9Iha0TeMm
MH/MK1/Jb3/Klg4x4BFWg8lBz0ILtfMdaBUcMY+ctRxnEI1OtT/26k+mdf9ORVylCoktqMdKA4uZ
eLrMlCO83i+WUM3xsFaNPYPIqw82RnK3Vs2MnCCtmz+2nDnlmV7OOF0X1bO9ebyrPchb7YYYmtRI
OpBeMiA7HscmlZj9LnluElT/ZTJCaM4FE8Kh1jppg4mTAG0opFMFfXiO7qTyW3/77l3v0LUK+U8O
9LId1SjJ1OTdL6Iy4PqlbPLJVzTxkqGcg2t6g/oE+IFMHOuRdumK1Vjgkac1iq+2aeUrwTDAnjAk
XvaIfiCk82AxuP0ou/+8lAhCiECPpJ7O9WhrPlgoHmu/AZ0CfzQzRGVa32wvaB2upVQxu7/UFeSr
PjchsQ0pFmqBWYxeBULwvL3WUcoGmb1miItjuIGZzxCHw5wEtAwECfeAutgM2wLVLnjOnAYIIHsz
Q49Pm2ZbYR2LbeTFcSlSu4K1oh+pVApbJwt2surf2kXc1cxSM17AkbltrYceXFYLwx81VxEJQcTs
HneIHs2NoLKmAjxFQm44jXX5jzEr4OeATpRyNAjMdyijA3BBoUSQJXk8X+qGmvr66fdZ2v8gghYi
JYrspxXT1Gm0DWSD29F80+1OPjR0KZA8mh+wwaLEivpr1ktBZ97x6cVyUKgnopLzmyR99U0/GoPT
atIOtWSMC5XS8IWTPKC9Fj/FATJEcg9GxQ4zsRiv4ZvkRm5NHK5fiByQ5s+dQroGTHSAE3qcDwnT
jCJyZtKoVsv4Y0MPZlU+WzWkIAWEaVyJZaRI64Dr1W9BJGtXx95r8Twd8aFzzzO9ZgcrX5nLq/SZ
zEWNRFJBLk44kYb7GYxojHF9vGtLJQH7/WkSLoH7QQmAjit6TN0IKVQljJvpFbXcL05njjo4StvK
C6N14xLl5or9Hgh0irGqsXv0m9wAsSHQdFYOJU78ZEUVnhREsmc0YdcXDiq1tQ30LV4RtM7lRTL3
62I9XU/n2m6zYLOo/WdOr6zJnv5BArGygTcFN+Cr33eJ7J4oVR3QVfmMab73/sri/D3CRgrLgk6f
M3h1g0WmsOBc917/haMc/3BgpzEqu9+8PeWoUQYS/lfm9Aln937P4dEypLDWh7S+NDVJTx0rTNCv
vWhLNTJQNAYOFhTn27zVeJQIpkS6PxRo1tPC/vMz0uoYRO7i/JCVWZIn6J1YS/eRgfIwHoL9ALKU
k5jhM1rwrhrcJojvNWWoeefyCqVj3QhdyC7Qm2LZFOfRHmJtpWoo93+koW/tquWVCCIa9gmeQtIu
bxW9crKIIlgJE3QcsdWiqVR8Xt+11s5COt0AOYnc0j+GiRuaGn/djLawZg6mwDxLE1zhaiJ7g0zD
AkOqd1qoOXoiTaN+B9S8rxcWKNdeD+XiTG14cAHJyj1Me3ymsMPGMIRyYOQQAG2aCm/PPhJThHUl
QtdembgO0KcqehIYLN2UjJ/EEI6/trk1c3L4CLEKTddZCEvXHkiyT7ZbbxjsmQMaWKBYwIizcVLh
dHO91uONDIqcTJhNuYDuuXtq6D0Z/tm6WzWlr+st3dXhBGTA+foLTcHHyA7pFRhRNg2JewJWfZjl
oFdyW37V3O2Xb/C82EVqB4AKSAuZ2ZJPqmjOLG2YvkSpl35KI57X2XcFmnLjJvsKnYDU1RxEFq5Y
QaNOxypWp9yiZJNAZaoE2HY58fLG29oO5YShZPNNqBuE3lUH/WLqiB8ZWGmy7HIgr0mnp91hTNRL
IbgNFN7GHsTSVOCBxX+5FQsHOuE645r5tySxo80jb9ymyQ2Q5BWDloSrH5W2E8flQT1Rd+KDzcwf
Dtq4zTAb5j+i3+JvPbizsIX85AI+H27Q4hgIU1667xHFTsg7Hz8RsSmQ9E5h5oNpE8PUi0XnSgVl
dLscy5YOry7F0Q0tYa34zMdhuEAAzyYgNjFSeMJBIUR1qt8pzzSCJ7pVp/TKTykVLM0N+OkOQgGS
XsvtXuBovJw7jty3LwbXNcORsEd7NoYhTVvN+cbH49XVHhTkcdH63sp/W4+jOjK9oIz4KmxWENXG
RzP4ORs2dlvRAVlj8yIVSJ/WShJaDe1xrVhZRpGOGmX0CHjIFI1ctLdoSq8nXS0ArxTwveYDQuHT
p38BUBKHuwYRZ97w2CWX34pGalnqtfKkXdX0+nEjaVG3bKF7wYAjVLcpKSAJsqGxb6axLdxrC4GX
Qr8XO34UzZwQujCc3Axe63hzypQpNfWh3nKOrDze1FGFG7j0aSdSAoHf++b72JoLb6BWLxnOchDM
Z83ZhjJVLcip6da3pbEepjvZ6VKF9aUzlnzugjEAQqZAUoBRzfcBmVehoAFsw/cR2TAS43gY5QyT
L+NYml1fjya2gYJDKpxRkdb+kgP5YjZA/SZ9u9bL1dgo3SXuQ6R335PjiYk4wDgxxXouRlGwWSxC
UQtAl1SRW8Gf+wi63mnojFK56jv0UBd88TKZULi6nDPCVvb8u096qX/Mz8rvkFaSwMcolBhXWN5K
B9O3xycaTSm9KIH07ES/XBE7ubNd8+W047JrGDSmxjQBkqnlm9gIq01zmjgOVEzqcxTNICr5rjUp
bI8hbQ/5ENCoZHzTuwUwJczHOWBNe94WrDriq0NqHhe/0y87KOYSX7QmMeAmft+CTCFnV8IshrtQ
uZdHIhzLWRUZv8bAcnRrz+QUn0VLaXEpNWFVfJk46W+cazI/8v2ucSTy40v63xo+nCDBGMxiHJJZ
gJLj9QlMM7X6uqCxAihEfIUPKTRGPGK3UFpTwjaLHSq1Nbez9/fnyprE1cUsLhfb6WuBZzLB/nTG
FHymNGMjn9u+7zKdDyxfHSYkqesib4iCAyegq6OcRloJr1U/SfHBhN8xDjwPU1cIFBVulcKGOofG
y/0EWoOZahkTaEw7eEABJGrdsCDN9/l533dDzZb4IDw8GcuGqoMi4VYVB36RtHTpg21M117BbngY
IBmG/QPliiDPGtZB2ShwPRwEl28Mrc6vdJhf9mk+B4TNORgdp1ncDO5IqOBFppBMTB7+2CYVFtWg
PDDFLySVFGz8dPJz+NrMiKeeQN/1CzBdZVNOFmU82mV+I3X7PXf6EYHfClvs5ExN1PC51KMjHHTQ
MOV7wET1dUPrzFjtTSY6XqPEA+xchiznrQC3oWU6FXlSCVCnUc+TgtvBjcChZlo9lUkUlceLmgIl
5CrrcOa+Ob39QJGdf6fOgMsY5YM7H52UVg/+8OGDGnWirMrUd8mZFaO55c2/G1DlxOvsiFh7EMle
WoW+9QNY1HHFFI+G6uIsgHs1awUWmsRb7K51CFvnZNX+uvNcBd9D9LxAXO0W3lDZWxmG0jpJWEPQ
0wQXnVd5ga/Ng0RhjhsebyRn6KbsH4t9hh4QVNAYZ/ra115F1pSmo1EvPZb0DUz0MklWVRNaeDEl
ZkpsptKSUHykTkk+unO7gCg8NKRFVU9YLE+CWFnG7sMAO3fy5xf10W1R8vtR5Bqoju6ZrPfFy4HF
z9B8St121Rk1nCOI6Luszb2k4Geg+OsenL1cd5mkOlUb+NW4aI9VJvyHBM2qmm6ynnsGWQDgOIaC
IlnKnOQLL2TtOHmgWz5OZ7F/Lc6JWuMURwcqp43l8VOPQzMT+dgYBqFxE/FA2uKfr6IBSVc2q7YJ
+fYudt7sp2yqOHxFYQKyhdLjnQiginyWdFrWqvHLZtPTWpDnO1TDj5ofYh4L4EwOcPKnznh0QtsM
is1dT5vofRtphTt8En/WjTYmYbyaqUSFZUuuAirj32iheGmEVnSY884qg/0Unzeutb82gLbz7Gj+
X3U+PQXl02GK9OR+N2FTA/srIl8j3AGgLIXvYck3QVqFUTSg339QLRVfp6s6Yz3scSnUef9/1s2I
w+iNVixjaDZT+Pv1k7vgLx6tDBV8DmWYCJmJuNGlVZ/m8iA3AGooyyx1y31E8Cnn/WoFNV/jSa63
ZtpSJAwoINsy6zB0HghBisyXEqbtbS6Pg+kDFiPQiXCa1uq3HeqKQfOtH/wPHcX1Ab6lCoJIyiIr
/EAqrGq0F+jxpsiwe25tEcld0d+v9cAuRl7l+WI4anWdCllOtQqAq4d7hqzSuMVWdYAibNQL0X+b
PF2E40+YvATwvS92TcGzdyDOqYFSCnScd4vWL6E/dnJoP499Vup7UdaGlMgs6C1bTm+2J+FwuT3a
RWMHOPkStu/wPNycj0txUuAlBhFPFaWcKLvqtTtjGaiyj7/TvXFL6YiZj9vgXn9EZaK0S/QPpP/M
Nfpox38+fEo//edmh2v3DKxw6QKngmNpSdLRkbi84/crvVa3CJAhKqonwOcpFvzhVrIeZ9cnIEhp
WDYUZwwH/8wV+K7taGEXK9u3+2CVXlSCmXzieENfXTgu9QomXuUUaMuohucIHcITSct8Kl5rtVug
WGqfjq1oQvZghPEmjfM4ZVDg0CKIZAMrji6DiTQPVK1oNrB6WFslE/tvQDlLy/ff5m+BO6h5HhQJ
GXKNgt8u9fYe4JSSATk4kOWVcPPu6BUAFmAAuabPnY9aexw2thZ9zYKOZUQyjVvSMCS+l87j/ftJ
J0JKcT2F/KMmOvO5w73APPflb2h5ZqHj8lUFSM724w22TOh7OekccPxzFdfF3hWFjwsIZHcjCJUU
rw6APfG1KDHwommILuvAKb97wZfQWd+yA82T0phzAXFzyRipnSaqeJRZgl+GvK3YB5VB9/n8t5c3
EjwBmP/BdCsg3YcPBO0H4Ct7iLUUpkw8g8V+eC70LGKNOPdzTaF0mFgm1E0apB5EDagFqEpmDUMR
pvlgb5webmdQ/nwY1DsCmGOPDG8V2tPrmbiNkBLkHbYNdy/sSQYDo1gp+ZvsSkjqonfAqYf3t3KH
8cvA7QXMBw41IvMVHvk5BoB2Ltm6Qq588xvXhXUc+r5E7uLxpyY4Q42cBvNAYHfE/cvXnv/rcv6r
1EWeCaK4eTom4jO/o8Yz74c6zU16mh5qaOqw/Y8P2FvA7ott7MKccNyTem3Tojqan60pekEUecxZ
5oNFFnAJ7szdUhoTUDYRr9LbN/bnoOMBcd9HQPZCg0wr3Z5RUmVG5RJA7dEQfepfQAWD8a49q6fe
wVMy25eacsSq8aFzkQ1uOPTPb4LcAUWtdRllAfQw0PLiriKST5O8TUijxBjDuf4Z4UBNDM/qoKFC
tm+TiTnp3CzM65wv7mJmcvnOQxWfPIISHspG+J0m5D3B1c4PyUtknncm/xVkfbJ9AXbjNKX/prwy
o0App0tcshJ0Gk50aMBziLmQjIMaVygLgJEsSPld0+AkoSC8cgL86MmMBNFxvKOxSGwrjy7RrqKH
TkXmfuclwO7HLAieFKkf0QhOC6YtH5cg99gvrRJ2jlvR/4Qycygs3nRTpjwJsRYMvAspKfmlGxMh
4J5iNqrVCsUh1gtt9mIKsrY0RAsZfJOgXMyp5vRW819mSXP2//12i2bkNcfn0YFwN+10QgZaHMk0
KldXleDHSkYQEepS4opzvKO213+D1I65xlbQVthgrCsNgy5Vmu8gMpmFDMCRNU0aXxWPuVWz/OKU
c7ozGO+qQTIJRbKvA6nOQhpBtjGdK36yJJjihWGN5kynlTuMrhhQZJFWzCtlKiZstH5yB/Cxi5T/
E1H7chALxOV5iuJ66EB95XqqvvlxzOkSYHrMoW0eVYNwLdJ0IOxHumM6/qykIyzdcYSKc4CjOZJZ
mjUqoq8JdXCIw1nTyLcUh0ZLw5YKNKwtbOrBTJqfDqLxS2whnWR9cFq52+5MNugPpnIa4CQbWrcf
lBkKfPc74iGPE8e2IE4gijTOIQZhPNhmdxfx38lumS+wvbBR/eiCen65Rv302AHuc4d8P04YibIr
i/wzURIQIYdgG3p+OQD7k/darkPrfXpY2AclybhyKVDsDpTwlkp4Mvsaee5mO0Z9WQoY4CA4d5pj
n7no8p3X2lbQAWSzi9Km3I5mdKuNPg0rLENrg4gur8q3WP8DT+o34M9hG+MGDtOwqLAjMkxdKKVM
pxH59cHCW/oddxaWCT8zYBAG68R/UWPrqGjzxsr6SRPr/I4lnPv1IPzr+wfiZQPc6mKJs/6Y+wxA
5O1M3Wfp+1zQKSuD2Pz/dkTqI8uX+svG2LqDMgAtlqy4qk8guydAWdq6jFclVFtk4JgxBo4O8LIE
XDXJEv2QYa88VynzrCvBqVisD5lDoPV7EF/w+rVz8gK0toU4aOiZ1J6e1svnPD2srnZedew/Rovk
pfngLfXNYfnG9TuF5EstCsImSMdXK6Ey+VgkIj/a2kUGQ2ZFLvCA1MKDZ5eAQy/2dga9PN80ws2V
KRmOpnEtwUXrs3h50V6SZfoFq9UkXbGOWaDKfEcxTarewrsgNwTVoXVaanuZsTqhksVKSJ8BRX1j
54TC2YfoEyUd1BTO1PH59ppkFsGRrJMRIHfvPy2VssYOzo2bjRVcgLjNgvx4oHG6sMC3WLJZ8wPN
XFLmSCjfV1Xo6hKmPzHcbg6t/I7lOnHTGKLOPjVnxqaz30hdYTYEWiuJcTYSO0CftNYrdOAyQcVI
en71lfwQCMYdvkKrcu2yXn6DHAxuALYnjb3midNE++WqYx3EXCWlPoxT1SUozyUromJwYqy/1URQ
oTYrxjn+NDI/KCMXrOiOIWWzzSIKOD3h2Ke2lDnsZr9IaLHOZq7n8j4BMTGK9c3nJNtRjcl0Uw5W
LEj+LdUWc4UYDty1juqB/FCKH9gu5/UcF4S3Z/Z4NQLeyyruORvp0HUyNeSY7aLaRzvN19P/T6Yv
m92zop86doBwt5C7h7f0+sgkYr/yLLB4+hOO2U+BV8v6DtWYCPRTKl2oxNO0N730+eUkIXxP0Hcp
W7GNDBQIeX12p3zY+8DJAxQiilcBnyYKaFWhx+7+VilXHiKOT0a3/kLDinWhFvd2Tp3D954r8SUM
xH3Wb5Y6FCXUh8y7ewglwdRchjJpF1hbjPod+jJIT5p4ZY7QlXxNggsEJuKkBUBzAGAacziG2pj5
Y3T7bozs+drlYtK3jH/uQ9U3SRvjNYOGdXRFYwGGx+0c3/F0cxfiLJqWamrl3qa/LzKmq2EmMNTc
rpf7w4mQ97K6FEuMEyPuEoCTXQc01w7PN1DxzVwobZBxJRWcOVFJp8G7Hp9gvBH0EPKODk0Kvg2C
BDotYsruQZ05OEWucLKCRK7xMM8SlQ/Q14HtZaXLqczbaB9f6oyA1QGFvu8Yn/S4v+uaq6AyR/os
RkIQHVOseYbR34NdB1W2yqvq2Etc7uDrBh7H83P2RPJ/NqIDmMMarSorQFisKkpyf1Bv1lZMdA8E
ETfT+scSmnNjxGcPGKBLE10pZ/RQE6FICRY6SxC07BZrrn1BHpd6GBpLGAqB02B80oXCdsmas7iH
Yj1fHniJUQjt1iqz/AoP/qR4kyqeroK+afun7v7z6porXzxzwybtfnWHssqXCInCv2i6hd2RVwk7
VZOvfWVYlsfZ4AZMLSp3lBihE7ynFvTXjIs0272MAY5BWRFdSsPWnEIlt2gp4uT4ofgIUr+Ol7Hu
10B5VjTpigVHdJtFhO4tKl9RV6SWCVR1QJzqbFdrrC8FodU6QPi8IjoFNRBGBDoSws6K0cV6RHMn
9vfx7gVITOzK4zEASA4j82pLUd0Fp3bp6OeOpa38Dd9pQR9HUuVv4Md5qflp0qyHq4l2N/9BAvHq
x0/3la0M4Elg6pCXBYHv69pFnmfelb9Eto3AXTomoD5/fZ4HjI7lTtnfU68qSd1XYJZHc1tWtSX4
ZPbixwZSAjkNzXtkHo/nvJRYaXgni6OjtIolqA+skEf3Yu4pYuCahXaCiwXGQGhuMqe5Hv3w8OKi
ElFQ5sYy8r89rAqOR06VFFoMS1ITsN0Cg8oKbP5t/2Xp8qNOM8wPc/qiMIjiVEpaqjH2EjUAv0XK
QUNSiGFUphaZvIss6N91QigB4ocKOJPXPXQm0eO+GzMfe9iXR0GWYJbq8/2GddOwwo+TugxZKEo7
eJ+eZsPZXkOF3UXeOVmFhjUfwtvvAFvTywbFJVlC1X7gJ5CPFLNwy7TawD4ONprZmG+Dt9txB5if
JiETNDswL8Wyhlo2MciSfwqFsIA1xJD9ZF0ynLYmP4KmsMjMFHD8SJRLMbEC0UMh5P9+R4Us6GHR
Y0zsm/yFYSmlu7oF5HfgjkpDwpgA7kfaIWZc9InOs/i9uPMsrR9HoUXkjtHHgcUROlFV+9XP8EEK
94KpBP4ZaEBYzcelARrHnNx7Ykd9Am5CadqPG3b5c9nUBFvVRiQxu+aakOjsETutcy0Sql/Ko+NJ
L/Kzudep43Kj/VDllFgmG5wPfSTOklADwMrOzN8VRpM8pyi84CoL3TbuPQEI5Gk1ichQNGYvjeuC
Pkyrug6gu4mRmmlRj6z700HaPV03gMug0BJybT19Q6VduEmhFkoQwhuiaeZWqX5M1vbZ6GFtunTy
Ey4qz1P7qWsurRoXt93/NeMWj5lxxRcTs/08jQJHJdNV0vlHI6blX1ZL793VkaLXGvPayXdaVdvt
ZnYQF2tK8T68AlpJcIEg4uAd38Ky1vXBNWtyAuBcOPJCLzJgZCJGoRxVeWon30beARxdtWNzzu6f
KDkodHqVGteCEToeJ5Od4wod4doavv/VNZfS6BuJKdHCGGCdoI2PgEs6cTLsEdBgbdhzT8IyXQIj
+jtT31Z5nxbq5cdviYEDt/B57w9/uW4T7jiZtllxNoVq5was01YpHrgaorsjg0rLJjyAZrhweS1B
TvCDW/ha4OGe02ii0xqe7rycfUB2kgV5QL+2CWHyLyhp4HQBd1fXnt8t9lKWGDlkQ2Oc71rL3GJt
0QKew5B5TSO5tbSpP+2jOr63+khiMEG2KrLSpzjf5hOURLfBXCQSX39JD/yalD5x6F0GRcy78ocE
R4JbsS+LSrtsOXcH5qzP0PLRo7KukzMQqQAERVmvQBbKQVV4+D2+LgvR3mDd9GYc4lVZX4lA0T9c
GGohYOn+eQ07xreKXgIbBKT91rj7hU1MewDdhTDkpbo7CMrwTWCDaq/O00xX8+bj5sxpUAuiFo00
sGzEL6+sc6QSqWcspoqQjJwmJbWZ1yXzSLehah/zH/pjrNaRmM75m9Ni55jIQoLcdDosmBim6Jlj
m6Zj/ccCroh4QPjWFmVsBCvG01AHl0xZYYiXZT2tO/P63Msj+ZAdybS52mxlSpYgCFHHjtj66BmR
43RLwlMIV/4FgicGXGXWzAcli/8rWZxD140DMgRYwCPk5CQlqmfkXTilgf1UTIkF5bV1/ZxRccI+
lxEVpTEWhPNM7hVHH8ONYxrvQRm1YvYvxK3Y4zIp/K/u11e0VXEZc/+DhuVKQ5VP1MOXKSKSQ6dT
JS5PEaYIiUHc6RMt0fRBzJSDCvoHY1t/UBQo9sqKtOOuz9D7LnUKODzLK/+/ApXSdfFjpDHnReiL
cG2HPH9twD2RobhUGOAJoFsEW2hEcKTSGVhNR+ODVFKQ25DCPtZ2cxP9Jc+/4w9J8rFibIKy3Eco
5z2YRjX6yYc8eXtPcAQSS219djouUPBOuQCSIGZOugDR4grAE/uymcfMN0kzChMxZzagrYJhzzSb
uUz7ujLOrynKHLjBLA95JaCwlgAJcwpWvPNgZLZBAxpRXBZrTzRX7wiCAzsoTttCDM9LR1iyHm9g
pF12Ln4pXOgkghyJcXSZ8Svi2ZL6Jwwb5IuRN5Y75UMfpDtKlr9GRILvsLKX7Q6XUBrjI06dsub5
HVabL5+jSBSwe5LJqGPx1kadHNL7CZqCuZG3D8FkesRsE3cQ+8SzPp2kym+lcx7JwZwJmwT+V6+B
/nVHIIwfKey9xZMhw7um4vFSyBDB/LhFuxGT5AZgnyOktEoPc8BvxlqBL3En731NLVkz+o/KFDsP
K7tSpIH5r1pQMZ6/zrh4h4DmA1f4F+hRzL+gCj5Uess1wP6Pfu40t0mUNeTurz4tUQCvooTUlMwI
xXEmAXTylGff6egyL/CknTBsKIUSu3c9EfWm90oEL9m1xyuxNwneTX2qwnLmzg6hmfm7FGRIvCQH
tkqs5tKDGSTk78Na+mbf1CuBrQ7l+3XRVfeTiXkTPWMX2vO5a4frlj4eSRFciBnpX/tO8riEeodG
o3hTnOJ6iehhbM4sI7acMPN1hj/tdujUqWsFxsUzMvzdA2/3Bhi+BU5n9V7FepORyB5keF5Cyv29
iKJNGMEhUuviWagY8g7pd/NbnG9dqe9DrsPC0AR+iygy7tz+DYlfCQxD1jUbdvlmtqZAFmeVrWTZ
UVTQkolEDhgPGdMBZKkxotpohNLUlKxmmzVKMhVnozCqaUX+4U9wuGbQB+FWBxGxUXTDgE7NGWAb
s8O0s4aTNKoPtBsZhUQ095vgdZTSgii5rGQJaTs3Io1aCvCxq/fXfc24Evm28NPl33HizHEzOXMM
Lxlpd+B5kvxR+JLowV+Esmjnul/Tb+vkKEPf8f519fk6IE3GF/JcQS7/1pLOs1BbzysIuQRccL/v
3o1SDCkAyBJZSLxGav7v7C0M863cERkbWLxdoOhCWcjEFGFg6OHMU+bdfhYxrDBQeRIE6NOHocul
FvFwCTzZa+KKN6dt4weEMECEkKVP4klrKSmaPTIAp95ufc2dol1xABXRCPa4Yz879xb12wePwysS
aUFqagDBPlakvqOoAMru7cXwC5jvqRxktnriZnfF2AzrIeW9N4UOeAzZLiY03sawYQ2eVpNmfJ0Q
BfAYAYSxlvJjwqI2xrjPlOvAp/r+5TzoQqgLRw4bb3cGPh//tKf8HOHiHL7qdWObh68KMD8NOi8X
qsevZYvgb+1fqKkX0M4+4T12+RTk/JZop8x4Q9Lf5K9D7/KKThtS9iMgKB+pefEmGBe8OrHC9FTs
Xqf92G24ls7YWfhPBAsHpdvit5ubpaMzttRCOOcbweeo7S6XFGChfeNOQKaquQV/oekxPbHBPlm9
1wl5gXHOwMR64jvw6Ph2HS/9eBWEMVx5jjPRTrHG3zNbqsfkg/B5SZ4FhUAkx6pmEMK3vo/83X0s
ylbzdZskAxmTQxSallgjnnC1Hmx2XTCWDV/ByDyPJLELTP37OqYsSy3lArJQCkIgFvXv9SJbDvNA
psjQ728IMaAdfqGtVz4YCrnQJGLE7Ur9rnvRWFtd1/FfaPJ1eoJOVVBy7ZD6Toi5uxsx8nb7rlCv
7JS7vj7K7MIRJflDbso3Sj+9ts+Nmztt+AUna2Y2azvD5KV00g8kJU8d0lP/mPdznOP6mpW+TTb2
ELZ2905eY8j1fYnf5KM7ulJUD1iXLFq0xe3hx2GzCDyBgYOilEWbLxPowxgxpAH9nLiTVOskhhKD
DtLgkNmUhcRjGwhheVIbJ8rNqA36RhH11n9RLP0pFOs6JyroWn6bc1u8MkVeXDIrErPbmIt2zlmR
vhCfGpmhpy6mHq6JmPMRXCVi1FItJkOWx6kRjjh/EAX0XR+D8VeHxjWcHqQSTvcoI5+FFgHpGBVY
yquj+75OOB8uPS0M+o0Al38QFJplfFhQ91zWJFJTBnq12MFxzMZC81ehz78YsfP/noobISqiaxEE
ViJS6tD8rKlAD4tbfuLmQZx3mzQXQljfc7cwnD2Y/kCviaD2RYKgHGCzULNajnO51bkb/IvDrfsx
JWKRilE7Ohg9atZGNvwVufk19og5xeLXuaNNjE4tcnhqnfnh6Ym4noR014+N5VncO7Pq8PJ5cIKy
+bc35EY3KO8pdbDMqK9FBEySpCh6JZTROP5LDUVtjGv/738WLELx1ZGHro5qj6XK2vk53XOxsBvO
WrHI6htCS9Xu+JQMWb1+4KKJ+mp9MTobMHgCuwiHAC1qYC3id3f1D34h7Ugo2e1zgHR+D0QzeO/I
t4MqH7UfX7ueclwmurOYKtu762aCfMYwIA2PZSYzo5STga3rxdmt9TPemVlG06FbfyZL3pYhqxFX
fZed/wknS+Czhfk6ghcHpeyGP7BCEGpD57z/0+eCIMJT98viTB5A+uQxAyz5Ga9LBPV0s5xzRrsm
DmgzsbC3lZK6SFdBEWKoo1MAYM6g+UTwVPCgKmZC8thcsThuhAj8MNtJquPwBhsLzccW88duiYMp
FzL83Jvm2lVtl6tziEvzkD2XyGf1PePW16YdPkqyx+KkJdHmq4l0TZDUTPCbqRDfCpRJ2ohdk/jN
pqHQuqveieV1oWUSQ2MPRwpfbCox7dDWwytHEora8Lo3XZySLdaoox9wc59RD/EIBqltEO/xFbHr
fDwBPfu8rDafidAjdl9j7OLBtf+9fMiIzj2yXRFLYZOfa/CCma57ZaIAMpyQ59xQ0p3m8OPguC8T
sGKWrCxB7xEcOVUQ9bscQyPAeAH5W/QnATRc+3/looQEkdX780nf9klC07j3un2VsnM7drK9SygL
xpp0i1qF8QTg2xJaNjK+mIIFvkvXHJ8NjizdmRC3xWK7RunSvtqPkpIkLPI6HWXbISej6fqLNGYM
kmvFJkvWkC4L4S/f81P2E8delw6XIZ6GeAXvuM0WplWNiQnXJINcDf56ovLdDjCxZKMNcJVfu4b7
U7R6aZFsJ+2ZDE3823BosOpIHYkDnjmrOb26abQoMkATF/bPMOVAKHRuv+3H7m9oMoTNaub9zkdv
lpaR/Z4JqnN+EApuwanDfWuLKM42aO4jDwHPY9ldOT5lt1QgxAkkDzv6Mv09holqUcEwxudJLAgN
z8POWZrsAKy0d1xau1vsLNirJ5JN3ijs2UG2ydksTXuzcrqE/5und9VszgxJCFbXDDd3VOB1NcpF
KMs4ZbqwRUS8Rppa422Q0Jhb4RICLxxWUr/tcuQqmxaGbs8J5m9+HAaDrxfwG1TkGN5cQZf7pIaq
DSX8KviOycvrgl4IYrUicIFRIFKiaZDKcxfMdvtIXsJZKYlPCCrHEVX90Lf/F8itBb8y4jtimVnV
9ye10EdPVjROtl5m6rCzs0gqOnn7fkJW0YolP2ZW5Fzy/TFn9uVG6nCwwVg+mSUPbMU75AsMU8b8
2MdxLygZY+bm58d1Oan2Cu2PObW7pHqZjNxgWWTdNOx/jwIvqRXoOnBZ8uw0G2+kPD+11yYc7e8f
s80H9/i5qtwMbL1ZQeooZUzFda2PoZImVIRmPSG2LSpAMEoLJGPD1yl79pbw4RLni+Soi7gC2jkr
iEZkmYiF9lnr0AK0Kfw7yJOz/4ioCFEQ9TxdZpJKWLOn4PJQqYWPWP6soZXPepGfz8YfxrcgTZ5+
o/LpENB13lIqHnO1FmeMXrM8fiXELQVOjOFAY7Ebdae2g6/m6aIu8qIebMkw0xGdzPQuRCnTIBwr
nVthHo+qyqjaEAiHoURvF4UmwEJlA1VKzNyCViXEZD0pm5ayTx+rib5J3VHstswqLDVc1mjaBLUB
RLSwbvVbndiTPluh/LrIqEUmBL/Glh2g1r44aocqD4yMlW/AsslvkogWGKKYQevQOmOZvKbc7DFI
lKh2FDCC/0I7mYmPeTZPnQ8M6XoajjjBLyjrpbVx+CaXbFWk+5l82+A1PAmi5ufWdjWMKvxL2wm0
2z+9Vj30QxpzVWo9HkrqiPOWJWB/3wfiKzCaX0l+/uk3hksEOWP2fKstpsWpm4PJQumn/uXL4HGj
I8KKAUMAG4qRo48Qj+xle9LuUXd9QWEZ9GfGMrQHtvSPtPKM0q1mFPGD2WCp+wApPvbHF/r4nLKx
0CDnSFS368pVrPZtb/1QXb7I2fFvbdvElDhTZ/k+H6O0+Y7oSD8VwB5/3vccfLK/UGhNNiCkDthi
ntFc1UiW/tAgkwKyi5rSi2zK804GM3yatmo+zK1XFrvIyndHTJxJUatt/0hMtW7374mZK8ufciQj
Y57dHN9KccBwk3DJk3TPNfI3ZeRSJpuziWDIBJigvq5tyOOiZo4IxXJGOrgzdyCKuaFH3QPEEEau
PDzUHjy/otnpphWMRtcLvBJOnrpUMVrYFlBlmauPWeKdufyRFfTGWntL3E05N+Qy8bjp20R7hn+o
04Pn3hRQbD4YJX636zc6JLiZS7HkxkpnkigJA5eLop8tWXtBHa+4U8C4AhdHzpjHdT5DjA6mSRbv
qVxZZRYsXQnOL0aURwnYg59us+d9rWmc6aIb6uYGsS+Hor3ttJMhlS8erZaiLfHigeNedBP1VGv8
IGBHkK7uGieifih8dMZf40UtKzmT54M1SXoLn4131z5AjqrYA4XPSVsqnCqdudC+3k3HroyaxNUh
/D6eCZhdmPwLNLoPCJbNw27FYBp0XIBnjdybpVr+Us0S1KlMKf4wqg9Fb98GOZY4gAzr3GXGmIn7
WtFYmeULhsSwamgg2MGupdZ6S1IVTjogjhs6+E+lLfuROK/tm2/I3sKmaYTxVU3tY1IQdhNkcvKC
AzEIqW0Gqeyp926LROxh1AYSXSrZRV1QrqVJoIdH9AGfFFBN63PJvuQAVtAqDX0929z5FWcKfDa+
oNxiHHmmGFzjSvMe32NsNlr68ZDKSGUp9zm9okFK1P3PU+KqbYtKEuIB5reS2hDPgJFC5VmImYpZ
J5ti+ib+EZZduvEuOHEgwQnlmvSc7KHYhSusNdN3W8xZd+4jB/rleRln4T739ecWRyOXrtIQXkPP
iW8SV0RILbrTGTyvK3yUgjO1lmuem5uHPL55eGquyhbXPKqY++ff8CqmEE01rq067DwZBc9hNZBn
aHfE93N2gtdX//nW7oyMeW8OaJ8LM/vmAzG7YjauNeWztHiKsKmaJ5AL1f9cgOPvSXJ3ktW6ngZJ
0wATT9DfGxr0nvgBl+/0GTz8oVAE1d+I80OzcVS6bUjTrjhWy5EfpQQ4+53K0h0rGvVNRPr/yRVm
cAAS/PQ7UyrPd6AudIVcCecvpsID5DOrFDrGWIrqnk+7bbSW6ENmgyl2xks8/336rsC6XCAh2Hcx
5vy3106y1VC3T1I0pHNecdXRX7eQNprrgk3CNoJp6JaIgbTt3oOjOmum236n2bNa9YHyNCSYr3Db
eYjIMf2zvs2pcmiUecUQDg5ZzFFJFOhXIZ9glhym/C8CnhTUsm9GDycskxNS5BT/f6zIEvCWLXri
9tYRZKWyxsaofq7OVAph0rXO9kvGNcGNw4uPEHqjMsEqmnB+szYu+iCiiKlw8YzdC+WW6Qua0jzK
XMa959luDVcVvTVwEU1nWSD2bFTD3qzQxXXl5+6l+s00YWWMO8liixN5wN0yKdz6ihCQLnYIUbOk
/Xc8HCz2vJU0/Ym0jXzaMcG1NPiFjE7Fq1eOyxxGKnwhUE57H3AKmHV9VNYfOCjfM0FxCvWGr7ef
oZeEpoh4bPIpvyVgUcDSPYbyS0lTAmjqNI/BiWT2E268LaufUJ/zGjdGC2ycYqC9ntTSAxrRmCnv
nlAR72K1EV6la98KNfJMBR+0VGsD+dUXRQIKZGOqT7qZFmQIXA5PyzO20VHU4ddzbU67DSJYC/+S
8o8GGrhlaKH8w7If1pT02JL/t9cS6R9FYzhjZKW6iRdendZyqh7TvwA0/GXo8bzPxci2DeG8OgGl
DZAw4ggTymrPICDk/EWVbubrCyn/vScGOB4oSmpWQAWBr6fLJNtoV4IgcH+xWFSW01qSfec0PwH9
xxKO/G3tp2tQH5VcCTNDLwD0uaHr6eoQQncjQj/vaU/F3Z1fQ4AWX5KNijmfAnfoazcMdoRyOVF/
LQoQBNKCyrXFcxsUhe8hlOyVj1NNN46x/mefTM6NeWMS+m+Ucyv20cLKC/s6TcNq8mrrwS6nYdoo
bQeXmxaUr2dGa7mTGqYW+RNBCtgKtm+PTZvwcVtmR7KL+gK3XdePnj8RMQZYLq5KpIVefuH6fAJ3
P43L34BWY25PL2aYNJErqqi8yWZuvovf4QhhLHK9E7v0ET272ydnEdARrzwKwkGZ/ebfcQ5IfbGw
8DyRxthHoLWoEkIaZKk4d/P1STPBsNLFrSLjNpDqrvPX50RllbEXFIhyO/NTNvvkb9HeyNNBppvM
ETHWNOKC/qv5WJUCMkE96bODGiEW6Q8a0pOy0JZN0PZpMm6AN08mTanabWijSUjYsKQztrEmCuha
W1ZZHTzfS9UWa4zdj0QPcwnz2pKF19nNPPMHyHlTmYDofUlcHeuFCocUrNJ7kA98aajXDh/bNBxo
OpHswG9wozzfvyczEGPqEMBp+xNxDqmX3KTbgZSrbMZJINqHFXoxECQ0i51Z/iJWPmd4HBJMpior
Mk6jE7iIMSpVhFOi3YQMx3eT1nOdrALhyeSDj6s6l5puWpKn3RQp4qYKREjJikqsiuU66d9uxfLR
z9ucke3RiLGSz7K0WN9CGivFKtaiBQ4ujKQJZcjPtxmXSsS9hu4Nbzr/sCEdrUM82uTAS/g97yMj
ZpesYHdaOq8KiyZEFlXTiDh5ndZr/7jXtRYct4jt5g2x3qiE5X823PEX3bWGoKcJvWq4yBZk9mAc
P9Xcwr1hiYOcQ1uJu2fCkJwVleHSV8UNx2eONppjwohnMhwq/cI4e08PP17qrtt876D+3rNRbtMT
4vRGM8h7PwBA0iNSMh4P5cal2oBui5IyBCjqu6bjcWONgKnG4MzQhZ5CKOWb5W6kB6lIjZJCv58r
xQAzmlIY1HZAXkWacXKl1kur0C/D9X8ZFT3jBqPLsnAeU1bjT9EHVl7vgv7cjpZRTQlZKt0r2NjL
YfRXh5hzVMGYoTt9Ehlj5Ck7Zjo2ke9d0s091UTpnICy6HpePmTsz4bkAnaF7sleEeQNkmXVMepa
XPzPnE5vWRTSXCswNrQmwNXf4EJY85vZlCvuMEe1dMFxupwqKHH4HsvqvUKcfX0100nBuiIZzJwe
66KzsjCd64uANK2eIRx6nNU4ZxyPBkzG7X3Tg1rJD8N6sCORffqhZ+Y9sCwYSNSVVcdzPgGpnCw0
TgWYt/n3Ugbbkyurik+lSAXqelwk5jhCSPA44qpqGDlw5JC6lbkGzNn+kvJrv4q0P6pDFDmkSBS+
cXKT4LKVQcrxluf5EgbeEfecjWtIqCvDgbnFizvxw3s890pH9IUct5Q2LJLWfUUjiNfDQHwVquUi
F7RuTDJT0ADZU2muwxnqsOMhaC86ItjKfVRR8XntFDV9ZrmOBuOVUQbRzv/MWGcDJmdjMoFnf62C
lTpuCSiwcMT7VdhT6Am2TndRCZszdVzoNGj9Ni6KMke1GXCTZk3ERZNEBghPWSMtbxiMKvRZAsiP
kV/XsTB0ryqI/5Wm2zehvwRBUIb0z3LxLW3m1rAz8a3wEpd6NlFcJplAZ2FfrKkZr657Tfkllqul
xImbE//kkH21aOD5ps/2QpFCIl0EHb74SgYydE8Y6BquzWHIqo3DTLRuS0esJA23PJbCz6S1ko9a
7ywcAMbB9OdunAKsTxBq7sIrZWrPfStu/cYyRXdce/xVTDvG3ETg7/pRdrcBhg3FZbbVLWmq0uYn
iKnDQOBW+G57G+CUPk2Q1A6mPKTUGHF3Yl1t/kWLdNDbhF5UQLX5BPEe4eO3yATh5GsmHuKpflNr
CdZWMqUuIodZ2I7Je6ZIMt63q9ULET/HfD1KNXDmtdY4fa3HuT+mvEwM+Eh3sxQ/5WmCIEuHSV6u
2kACDPV8Wp/yp2qAkfZCw9r9PgZzhyeWyIrBGrf1KzU4wbzUpzdzgrMuSxXXdix8/T2pUHPTJ6Gs
Bt8VOkiwDlqwdbaZUbwKAiWtP1LgrZsEX4GyDcMdWIexS1gmCzX5mGoxVLql8wSElyR1S6n6G7kZ
imo8d5Ae43h0AJJYr1dzbNvqizRWEaGdw+lcmHd/jPqhtn5YDcZPp3+Pl117X+MbSKqvfwIfbFnD
WruHzoLaLN2Ooqvi2d4W2tLLwvbynUXGjuRaYh851RBbJP9M86R+CH0HplRYWUs+KpN+aNthyXtf
l8s/tZVLfeZ7uGgl7XdVTeTJdW7B4AT93s8ct0mXTJmNdZJ21ZgI0Pqx75SJZI+EkDupdEhTIpQI
b2GfYujq+WSH0S8FoZGdHKIMCP0h7ZNczeohHS6kKUPzlhvNtglJptql80pVecJFSUwQZ9eC5A+N
qkcHp5Al2N/nCbFTs2k/w1y1HavyN/SkTic/5qhuu2NAcdYk6faS2IxfEhZ85hrHSBwcpZbF3H5m
HUo/n0vK6L1w67SOoFmSSDKHjF1tmC0EuwOqUmIy6XGZEUzIZMJ7CQrxcK8JkX+f65jd2b5i0muF
pX4Afmf8enj0dyttO9h9bHon/b0sK+UFoFFv3STex5QHNGm/B6ln8SnlxuafD9W2XVFg8BOZndnY
ANmskZ4DhON8KtrHv63Cm8ZYX0DyrYL/MUEFcg5tGs2e3DwJVarOt0U6j5AUjiIJyMLX98NWamP/
+hHV2J5JygKUDM+pyUjUoNoXhCD5uB1KY8lJZN6jJEgwog+5MelEDvvnTtqPxUPY18onMgDYuRfk
MLbudfDSE0SpVRPFbn4Or88sZoDuU3hopDG9br44wHrWGAd5g7G0ksjJhsTlGlhm+pVrwNOmWYvb
uwCrSDpvRtKb6MhkumRLOe1HH1NNQwSe4MhEAgVsd9NgDFiERct3vPZ+wBubOQ9Y/zquY0Nf6L5L
Uc0hI2H49PkcsiA6bcjBmajE/eywEQoBmrTxAlEXOmaM/a7QM2Qov68PM7QGguunaEKhpn/wLP1f
f/hr11mnwm2Bs0qL2OF5y/1IDE4ptmuYwRGocsiONAaaDfnYEGmD7/PFXAjjxeMYeF8jznsXuSFw
S2Ii43z1ltY1otnrYv22Zqz3FVQ65pKU6K/3hCFabiJg3TV9bCKwewTrqoMFkojn0xNOGFlqY1af
/s3GV64s1y6g66cOGaJsCDqHjnPK+OFNAI2mcsl8Zb7+gw/jqzALeLzlzbN7mAy6qsnmMyOHUEZG
3pK3vu0ZIGTqPE5xIIISD+jkolJEzrmT1qX0j0XcqlN3s10EjSA/6pt55VsPSGh3iDEBtMgBkT+R
eo4t6UBbMBZP8/yeLWOY96TvlmwOmT++p4THPgY2tlMwrOLh5t3ZQDBZAqqiOezRhOoBn4EzEjoc
nrx6PUKVxynBBC0gSQf87veZLfB3xaqhTGgnsC9zlwURgeT7U7NUfiA0wTYdWN3Tk58XmmWXNGg+
jFIyTXu4/HY/xD7kaEgYxjIZgeWDIosqdVk1OlwrFZjOpRMe3H0zjnaGoGbMBmwnxgTwgzBA4GcZ
EpdoBIJsj51Tuv81erG2xP/9Oe8IYb60Elh1SPJ1HPIKKZc7INLGZsY4LqCEcSD8gst8+b/lLfJa
JHcgac/92HMGFfI8ym6qEL0Goz3wZgI3r4LNW1uzUvqzTAnTHNKWeHmwSxHXR+2PcHMIp475+Ilp
4TDFkAlqRPt1UwmBLHwEOgn0N+O96HwxSnEY6PKgF9PMb+FTi/bslrHAgD2XJPErzajXVWG6BqiV
MLJaN9CU6EJqcTiLXibl9hAJJusn2b7nGUJ/tZCaJ8YmfC73qUd2PkcfkLFaxlHJ93yN4Sq4KvXG
VwpKJXdOquO8G3uKR9Xbiv17kBsuub+KMMxAO6eQYADiNsrtrgwL+33G2sI4aQegvk6rUjazOydB
5U1wC3E7XXnMKKMhbjNwmBn6mhWWSgVshTBd4dP5D9jysBh4YysO7rE5y2aX4XBqTtt6Nvz6I5do
mcFePSeheI6mUGK98iN8IB2iIi0CHlhfb0U0XGuaafdXu7qpJ6AeGKEP0phqyEgh+iKPMNEZx1Md
BKIoSzxYll6vt7aLQPxg6dM1NKKQgI+NHfbh9DfsHnMvSP/IsaYD+6q9J0y8I/EXVuh+FEHqUXLh
LCYQFq6hsuDeZvRYZyNtgnhQMSy2xwuBA2ATrtoLst+C3VBr7Au4nq1LH90+8cuA1Km5+yIAKjwd
bysfuIyIVPqRc9icazs+XUGQRdh9f43E/8GVXm4hqcgJcanXCKVfkG+rR8y7VQbYQB6ZKh7yMRs/
2uY8WyKZAj/SRKKIpx+V/gkCvlXjHpvVL9UhQkbKP0R1r0yGkdBoVNaos6CXmbrxgERjwbrKair2
ObbaT6ZZKLlVM+WxjlWOWefKdyKku3vAwFGdOHvzLQuCI24afA3ltOYAu+RNWyTfsyXNrZkW0mcG
CpFSa9Q7xQ9oab45OvVkhGM0kNH+ksFzSPOqEs+anVGXrLkLQgAKxr72MhDaLlhAYMi5XvZ/tCOj
9r+Q8V4Sj/WnzrdddT2Ao9URFZNDdp9FMy6HF5hNN3oahMNwWNwszU8jbRzyI/ctCuZC5uaHWqJh
yR5RhPZsB9cMa6nTU1WbGa5aOccAC/hxHcNylfB6k8TtLKBK93EAzkfawcfRz8BXVpooErKO4rvU
+w2IG8Ljjt245b4EdNFmQri0MoF4+bsqhDurU/IPgsUWMjCvjZxwAxZO08VQwRB9w+PP+FDqE179
4/jBaNUQAtfV5JNybMxOJIdU0/mSwn2gaDO7CAZL2PunQxXyEKXH+gTzxF+0f0ehUQefVVqfDysk
dqs0K7xV0BW4MelMsKFg3nrCaiC4Q1L19FxSoW+0oNQtYuf4XGyk5uPfkRzNr+v2KCVUYRZ91w0/
ph1AIfyUMhzmuEMccMvRn6FZ0H4v2Ud7Zw5XS/M1974oQPqF5EK3TGJES210/BV2Kr1GbMwvxDqD
ffZmZy3X/pcDQQBD2/5wlw+NacrJ80gXso33TjnrTpT+wPM6J3sVZg8xQlrQv+cTKTp5TOne1/GL
MLrdnxn71lfjgwwf4m3n2dskTgP0vZ4RX01IIg9S8ddy1th+NTkabJIjEzSoWZCWO/OcZoEoV9RO
svYRIPqTePyQ1xig2k3cDBb1ZkfPdrCG+tiNbN3H8i+wD1VO12iUFQktp76gfaZW//spPrszzCjZ
XS3AdEvDEvDx92ires1WTgJIINU92PDPj71jfvAwxXDTM6tEnjGDalh2zfFZzXqite0YIQ2vfQpV
oxBnC/dzO+noGK+wU4tdr5mUPPdHYcmO8NJ66Mx9VpZzxU2uyCogkP+uRoHJYRDd+USuP7uIvs4/
WxqjSInaV/agMutaFMJdAxFIm+oZnjBo50qPW0TlWW14DaHKaloWd0JrMsS4uNrxi1mOCOz8uISx
tJ3gz7fWUqQ+MzuFar89RcQLJG5xWQ7852s+lmpSxTq0IT87OlMLTA1KtR42kHObMgpDJzAPTFbc
ftqLIyarTjTejBdtvHaVXVk/dMNBLyEuyiHhEWzljqCuul/Y/imOmO9lRo8KX9lKZRkDMcKbLB7O
nxlPji+J83NQf7vpz2jJfPWfb6y7NliELxIpAlFiWk5iLDbKutJv4xUOX0FPlDQtGXHaHVxSDn43
VLaHkDSiKSscvOvQjt7PfSTVg0GcgYIjYdRJdjnHW4SgSN5cNcqaUqZqBRKsZL53ChWmDS733A5a
1nEz/Oahs0pVMp7kWO44L2/0mdWhgb36Z4rU+S07gjZeCZR7bY6xKiAtLQi5ut5uwo1/ZdepfNpd
4ZN9V3oa6SLf0gwy81NtTqF12bBWyfgapI5EbmIzgullIdLbzeF2TQS7pKFHDGPWIsw5IGaqzZOt
NieWJm9lbegugtPyxGEFKYJ+9Ml4dzpgSTMiIVjnqSLf8RH/00S4y/nkbijNOQ84vh7wHuZw5bif
vLYB/zNfX3IvNEVXeG3xd6IdZ2ACwyIvZM7/T0qDdaWxSuHAUKMCTna4VD8flw3UwjadqmKZNHgy
lyFueAi8yltFnrIfPebH0H5zmLz8awzOqAhyxKMHuC1ELTnlg0bUdUF8A20dzRenTj+qit1cFs/L
VfS+e8YfZUwUlVyjo0sBRhOvYL3SZtQyXf2h5dnPMIuTShSxx96hOP9cv63rjnVq8TeCAoR9FdGr
ZUOco5paEZJzAhxTXKubtEQvLWZsDnUyt+Ccbq2PXHsp3dVrRj92iM1qZXumA377adGgIY+MP476
pJaXvEQ64Uei/x0b32n/5iOnQzn5cIfA8O+fTEd5BPmuZvaNNFrf6ln+v35RE7o9pAoWhkBSTh2/
vhrh+r5KA95oiJ6cc1KQZpU7Nu03ySo8N9Q8KkaepZbvN3r+74QvzZqEi5NcoWKNt6+7AkFDN8my
34ZkNDNCMLnmO9hBXETEI/t4RjemHpIsaE1bQpVQyfMDyR/F8TlebhYJ7r6mBTsh6W+8NIIXxxYZ
HMEeUdgaFaP3O0PGAnZ5ae79mWG/LdYG8gQTqou5TW4Wt+xngynqcjYcW49san15vPnM892/iPR+
rPFR9us5z8Weeo8JoeYX0b9lDcFjapgcZ7KyFX4XaQTFyPjo+y5ctF5WRVVGYS39tUcrl+hIt+tb
LU6AAmtBWLQiyDX9ViW0iAFNI+3+xlwZryMrxzu8xjrt7H4py2OufCSF3vjoI2a7ZUhh9yNgfyoD
yj29XcDo2+QlHzq+r+Lhw0w738AcBj2oKCexqkCYNCB+DSXc2AdC3ZbnJGrmXLlgud74WsBYapSa
GwMn2YuuYnO/RTlGJ81D6ArvVWhbjuZWWADFtUdd95eKNwal4+PhJgZu2c7WwRl/QEXhQbhTbvQJ
HPsCcqwFlGPogMw9XkeF0d0qK37U5v8pn1YaMYW3vE6GmGELk2Kf/5sG+IosiKtZzVBuIKQfyVjh
hWTtWksDA6rn3pEQt/xVFr8Ez5I6Vr69Av6q+L4BjBpZKf6bLI8TGtLAqRD3VEgynTJruZKoQ/ZV
JxvR5drMbPyr+Y7+pgJGAcVjq5mWIsvp8l3u4zJWl8LMK0NC2HbTleQb3ts34ejOTExR7KAdewPg
QdgqvvvrOCotzKiltFJKKAEIa0lc+jmZLjxtnch7ivy2s0UWfJaDDHAHIrJaJ+XqplvMzFo/sPA2
hTTxcHF/S2jhKnDFB/WZzn5FkTQ/uF0Uac7xzekZyfT1PgLRO+BPSCA41STGylCbm6PEO18TDWbz
F71k0stwS26ye7bM2VIU/WnPhHDM3uVxAv6DdVBopoDWuD9BMqTDWkqnd+eJ6k7OBgZYz6eFMhq8
2OAl65eSbdK6tdDpiBXAa1Fla2MxF0ofz0Oke1L3sFOOp0nKO4Bij3LrmXri6gw/8cjN2XAdghYZ
jSY8PrysItjMhPuCilMsprjwyrUG2q97q1avjEvFi/se/NJrHP0si0zrzOmYGr2RDVa2xgzSvKf5
7oUuxjzEeKcTIdGll418tpNH97i232dt4nTWO/H1rMXIPxmy9pYECwvhT0QqxyaFEtX7p92ynk8d
19p2ZfXeahuOMA9aDcZxnOfgWyU9g9zoRIgqFN4rE8Afs6e4zLCR5Mcu5wdFwJ9zQnYzhFF9ixye
BwmG9fvJAeyfHHyFeygFgF84tX6H3+7G6KKffaJ4tOVfDPTqD1NyY8j3iQonkjJWIqhMmB3feXXS
qKnmSU4CLAw8pWRy2VAg9VMrnVMAU7eyP4gQRgL3E9uWTTR0dVMGDerAJkqvqV5JuyC1kVIF/l+o
mqcyWKLoOK/Lj+7D2poF+mHYg+pyBfP2ZUVuNbEFtXOQ5p1jgeWu4w8eR/twHlYfQ4aFXCzEpR45
SSsfYERKxV6bbY85RYDjaNQCuWqKR8DMoI83y4v5x4Bq4i/hQh4DIu7WAg83pdqvMfpyX4arT12G
VCFFGxVqgdFa1RosC8HsUyQI0pUb3+833QbWQVkmGUnUUGWDCUaFQRntjNR05BYkB4GaaqHxj46Z
A2OIsUvR+DRKCVcTdPzyOC+iWnIlIIscmvM3Xbr3WiSDnxfi3nGEq2lmiiN7Y9gcO4rB+36WL2gM
svCEHrf9Pzit9cb6WklyUHdi/1nhUYyHihFJov5u6AY1v4BdrWxc0Kt/uVPMlYLrh2fAF+V9E6VB
IPC9YkY4J2iicCHqRpvMZ6sUyqR6XCcuX+4+5oIe/Nkhdv7g1csBjv/VmyCVzqVcgLGy13s20GrF
HTLmXd0zc+ikoY8zgpfJZtmycIASI+j+KF+KYYlQBTW74AI0P/F0iNyD53UFRByhf8iCnysGJNoS
uJ9PXk2nnLiyL76n2pnYxcGtMAdfCSwZiiv8SUf52+xA26TLRhTrlXuVGzr7Mm2Echz9A7C0j9Pk
niL9YDwfSlI1gzU6DE2G/yFweTVAWsVyo5WhrwhUCvqDyRwdo3K6IS2MI4c04l0RvHKmSWWija8X
tbIoGvtWTXmunELerhS/qSLLblQGmPcNRQrX5ZcOF/j4E+/tJ7CI+ywNzrMyT8CRkmDy0OYDH1oK
oUXpcPRcsqwOMujAnHmLIdBbP/NmpZL4x3tT4g9ff8BrbHvDZ3EI86Whrw86ao8G4AvFonnoQXWx
GJQgixpa38OoFBizU0D6BGFxFqD8Pkmoa5Rl8LaBNeKMoG8wqnvF7FET8dqIn17AJW4oIk/xkOi+
MPIxxD0PYeshU1RR0J6zLZh+B5CbDsiB1IKuMUnXt7IzWzAVOVoIPXs1keYdGjsbJf3Zq0c92tym
X2WIQnhRnx9AymrNbjWiN7Bfury7Sc2zQ0EctYcxI1BkJyp0dsMPeLnzBt9CYXn1U8Y60dDmEUoW
TjNMK7oAXFLDfOlvmtyfJ7zKIRqjpw9T6EGvZB5rOyoeQdb06qXtaqumJ+Xdjc9mQOvKoZKaGGNu
sLk4x0SQWzRUvA+dSXvF+QwOJiTY1SuyzaacQzOGo50nYHcwnVM0BdtUePMtHJfpJYzrhLhnBOwo
e3bGZiL62me1q+ViiO9pCkCM/bm0mzTTdZ5+kyp2QYV2H/0PAyJiiuULihltQn7wSFuOVcZB7iNg
HzeUOPnHA0puHqR3vRRj1x4vDDEfevktUmq6sR+74pOg5R/o0q6DvGdiAP8hHaYtK/Aiou23Z2TH
nKKghue0Fjig1Kzhlq8J3lXJk14DMBHHTHfKty6zJI8cTBUOn3M3QhpJrYTACTldUAKToYFW6DAt
Ho54IW+hgEr6yrZD13dK9OERWSP8o4Ii/9pRu+0eRfeqfFgPfRptOuSMyiu7nBCixTo9u43flDZZ
MuhQakkYYoH0pGDzKG/RFKS715+suekXrBtD5XqjUTrOkEcW4oTv9TLJKel0pXkfAYWxrKoX/olh
dkbL8nje+mGG1BOddVT7D9Y84m7DvB0PLW4sDQr3obiIqTLHplbtQSfmcS/tQhp/y6BGl7somqX6
76rfo5znBGieI3zt2eUD374FcHuefcyy3A/JpBtagetcMUvPD+ZshOtEIx+QQ4L4LeQSxV8INyMs
Tab+HG+CWd/+3VR9ImBB1g+1RRz7FF4w9nO+RCcjPvsDkAZR2qGTMC3bl38Nhlh4OcCBt5OZPLe3
TYLYkuWnxStrN0S3r1/rr3QZmNPU4sT5W8TapIAnBsDElYpmRA03QrMjreG7esnkbhHQjsqefuJv
GffayPugvAi1pR3Asi0PNuwwvrrUXSTCMZHhQm7HKz76Jc9uXB+1IEH2+1qoerSuiGWTCBerAi5Z
xIzkEnKxnFd7n/Waawn/bve2ZtnuPL7lFQ9k1f2pGVp+cl6zvORW318po3A5dGJn2v71TT1TU3qj
836e3OtnsTQMMAwjHMFGS6PZ5Cp5lQ7TJ2SAm/CZy3QAr2jLL5e6CfJMsP/lha03Vvb8Xkfj+9Aa
yVwugxdb8sVbBc2wxbm6Q0d4/2YsNUgcMOB1PzFk48E3C0prSPRjUGMeVKJXLJhTDmM6vOcbi5OH
KjMYjzLuQ8vR2AQ9xL3xMPYPCrt00ng23p0o70tbgo/Gv8ecGn5sr0XP7EcN4Yk+y0H6TsURs0ET
9PjEvoag4pbVrWAg2vw9hP5O/6+L4o7DmujJAB9O4AxM5rZboHlBWKzfG/6upWB+4+JZyFtBobgo
ClqNtpyko9Fui3I4siQXUcKJA0d+7h/MGYSLFf+FknhSe8YDsUiLIExWkhaBw2mRQNOkbk3brsd3
WtM/6vv+JFW5Zt4JS7xz22LtHZPtbcHYTXCd6kEgj4B/Gs5Er7+5WYsklPafGbeR5wFRkgkvWAGj
2x9tNKqVGTv9dTlQWuPyTOL2MOC/Me3+PC2cgCJYfuKEztpGQW9EDhryrfBBwJFNrBmBYnWzFY3+
Yb/3asXhABthNH5GDbZzV4KFDMQMvSiNUbLfdQcWX/FvjaM8T8LRy2eGblGT2ghIvFmXczUr1Tb2
AsBZQHFQJRDPf3FV1yBumG4LHX/iogPZLYGgeN6sppClhuAQyWzVlDoMH7aZ8Z/Xf4qrgl0Y2G9k
WgYLVIjb2TUFnwvBADTl0CXouC72VbgHKFHosipCFCwSEPyCXfqsz08mAINXUuIGU4EQdTrOMU8M
oOieTA5HDYSxNwTIjFojbUjtgCR2Gwv8G9wCkEMDudgwm4Wnym05G+zvaH2Yr0vLARXASRuJ5Da7
OdZ2IbevNIAnx+rZ0D5WclcnhDR1kOoYYXQd/ZA2c/Su5PHfuyVTnGBcw0np8n25Z8zLgetA9ESP
cP6xUEL/klzt+bWZ4oxSbJVuNhDWNPo20/sVCpdlvGTo165CiEodD+beQwIGYIvFmw6JxgD1d4Rh
YDGUQdTHhiOvhbElYasRRmk5jYR1LMmjOnYDQ13QSLzJuOpQI5AwCaPiXYIC3nixuml+bx9ILB9F
7l0UVvar3cSVChsJOUEr0tgKlUKRelvU2al54wsBTNcphJ8P5kq+Yfokn6Lk2+lOHuhD8rv2/0rN
v8mPQz+m+KjJNBhdf7VXv/omnrrohfLLOkHbBfGh474buJB7afnWJiMlqq9OBrD63ttcRk2XAVUM
mwaWl7xRu37FhqWjjcS0LoPD9jBQutL3mlaBnqOL0/FcARAyjqJnpXgH74GOwnffAxDU81fYaqXO
BKfD/GvE2lyoEVnDf1zk9cQ/K2d3tmSKZ7vhYIN2GjYU6MguqIKlPvoq6co/NZABrUaFZE8O2tqo
Dj3slMLSWE5D+K3Iqat6qbzbIWU+4kqj7BWk7vD/vhjg8zvmHElyAJAy4yV+Rb+1Gv0uWLcNPyqm
uQXlxfUvERZQDoaIJV/3DEH4chEAAm9x4IZ6OvlHQCWyZn/ZpyKSp299FaK22qFlwSjvyndtrWu8
JSRILLVt/ksDjRH7XIcdbBES9w57TK97PALeug1hPgyCvWRe/rmt7xzO6ahMEAOwLLWBuUrDv4P4
qisxvh0ArYHE3qhoCIifjuhhr9AQnEUkcENeSFfOBKjZnpp1beYAT0XHl3xzcCaYhp5MBn1TJW8V
8xcI3VUeb3CBXZ/x6rXpebcfanf4PVLy/B70lAtjebUtOLGuQcErN597vLtayOXUxMlzewLTyVAV
MLhazr8+0RK2PA1NAHck8BDQX3HPYk8uyHD0FhBu0NMEQUKFOqRDFHeYwqShuA9YVmR9kFx/2tBt
iwn/KEUsePWIwsqqKnzzzysCscJxA20Jpl5NewUSTQOQ+HCbvEJm0YnqNWAiVDTiK4DxxXuJwlm2
Xxlm6ocpWusNe49H6odEwKYl9TAsoeLuCnhKfSwsKVMYNRpC6eivwB7Z6vB4Lgid0OqzEx+7LrK5
iVjNV63vwG2lHx+7Ithv5gb3MVPirhl0GCppY5GiJaij4uO6M3y33NuZWNkBEbKOrOupO6jx02cI
UI8tVyjeCkFGL4ADPXFTq2tnxFTIs6VkDgGNLPV77yVvoJn5BHqIUcnJx7AIH+HcKFGD6ZA62DlC
AO3MQgmLdMjR4PHj5CA75CzpSZaBuionPYSlhD47Jt54XGuCuO/R4JLNufCEP/tqt8XCYD1RrAcQ
NO631IsMl4+agXz58nWkVEBuO3MP03qx8XMZgAP7wbxAM/oLojGmn5Z214fFJZ07pmB8w6VwIjww
j5Xs6DuR7LcK9dOrI4rNgNAibCLh1WX1dYgifxIelDndJFrEiduTWiHfgpVit0/gHax2utfPpyKr
bDqbbHMpjojk8/pdlMmiWQtP9WtxBovjAeHrmxxpfCp7OIkd128dkt2waXa+TTTLSZEPk+XBHdFB
ewKuD1CZhgpKRDOXPG0Lg7mD5Yg+x/inWgXkeG24ipCu2iv4hPdJIWnnTLnQcZaaqukQAwEjYwD0
c6K+9A2lK/MzxDoTM5Et0i3L4u0DBjNBOjEuIq0DW9gOzHaGo26Si/FSX4P2znfQ2BIbtcURKffd
ei7sZa9Ppebl0T4HOcGVapIb7vQuC1kgcfmfMzyaXpZ8T8RE9AqHqKWPDXCCoR7zqnq/dGp9+G8C
bj4CScEFsVrhGuU02NXQ91MOUYje3c4TgUidY2EzOQiiIYaFT/tfQZBHdFT4Q2wN4OB5blRiDBIy
XdNYuXTGjfsI+HbAlHjp6UkFZjVO6PcKtG00xRnTkG8lJ1VCyscYGvtMiS8wFmgKxjBjPdEndvk6
AojfCVHK5VXBGhBjS3dnO9rN7XzD5O658NDL0TiHdpyK3E8ggGSDBNxuk3w99a+2elYj61Pe6Tqi
BYm/QXLAHrzo+3OOlT53Ri0MqgKHECJHhdP9Dck4h1jpaL3fA3BkpvkWG6vWnUpnBrJtdd5+brsu
bNaMN8Gop9AylkavLzFCv/itMVC2QHZBNqsu/Tr4ve91JZIA1EJ+SqkC6EMM2tBTkmlDyQjdcuxj
phd+s/AbOfEpc1uKpJg6Qi7RBP1dDGoinBugdjHyHdVsnr8bx9RFCi7YoL3XdHJ8+H3zc+v1SCIo
BfkEV1dlku3E1V1uCC/EKdJwLd/MPvW4ep4gP7wx4hR7I3F1hx7M1S7IA8x3ox0EvG2YRDpDRT1K
HJmTMu3irc27xIXg+V0jbTbkpNQwkO1s2n763S97A4OoWE/zkhMDR9AZm2tE1R6+F/0SVSmeMGWb
4pf6g1Z2dRggSshfc93BZqYxIMBCrxYgtBK2O9uRhguP6LI0aQv9u8J40hc+PhgVZUIwx9Ywu55q
s20NSOcFE2VQjzrtGlXSvKeOSuxXS5LyoaPtCBhfK1Kj/EaEDrVms/9UK5X78OUuuXFRkbaKnih5
Ztr0z6DluCXyjSaVXLg71I2SQUMtzFwqAm2ZBlyo5tdFAqqVe5YUcCKB/zplOtN0zmKcjB3WYnAW
LNhPcgaebdOemEiHR5V/E5JkzxB5NioTDW+Ltno1ps1KpcnNlFrrWYeIgmdtfSCI4JcI0nz+QEhz
z+w7IeTHPKER6/2J8iU0M4wuXeVnPFTjSeb/0G5QmbHcUwPOqLU5LXqlZx7Kx8MwBcjYTk6UL0CG
sRJvHvkxII99Hk3MtcDmW82G11kXYSoMgftDHVhUysjwrNZGAlqQGsZfwZr9GqbcVtbwF9y3qrmR
17NvgpyyBtRDXtU+Cz7DkmPmyWfm6DJ4jebbXboAIj8MJkK4a4+ATY7YZyMh33Dy5j0tsy4YrU1T
AziKcV16CPr1mHOF1wKJdUya9D311coNgyDcjmV6O9UgFKvMi02EvFydIaFR68kJOfKRvXFn7p7J
QKda80Pg1f3vnwxljQ1WGOa9jAuduPA28e+PLe/0cAMUyRfesVNkeqA2fMDP50yINikPfOIvkjf6
cJH7U4IOPL0cZ1i8klwCEZHVeqvC9CNClWExIT5Gcj7K7t8VA16ittLFxCgq1WIadTCuXQDb3br/
WgPXjqchWSZmySR4rsjv/ygsZKpBsAlUBJEuNO3GvNaSXscEhyReH0MizEVPQanvBQrzOkpcvndl
kfSrI5uovanKEvrcI0jwZkuRzvXRlcNe5ybeHhRwa7Rvv/X1puQvZSi6wIY2f0CVALitiWk7Y/3N
2SNg7jYgI81UwTwVmcV3cnjlkxvd4FsSnfV/xOPYmlKiBQ2hZjoglT+VPvIpkwhh7PDucUiWmTCQ
ABB4ysqTBde7QS62cUadjZKj34cjDkY9H9t/HS0sEtCQIElhNrxiH4pcDsoJ95asspEwkjwIcON3
NLAn3AhOKd9YiB4wts2X+M4vA5em0soTR74a4F12H10/IOxJVyPrTg8JIQEuAZylbNn8DU9gk8KD
7V4iHDzZTFv34YgqnELRNS7id4mPGqJTAI5L/AjVd8NT7H5tQSpL+lyxEAgnEOldRjSwzUZkUbNL
kOi/LTv7WTN4u0qTaoPEgWgIBJVQb9nBNQTa9vyp0tEefVw4b/VqfDZoS8fyWxYeIYsRhpdUD8yl
CGBzF3jx4pUV3WwUFsUJGD18jyBz6+33n4ntc85pKyVfBQAtzrByzzL/eBRxUFsmm5wjhsKR51tB
SnVthjfo+KBalEwKSU4u3Cbx20FrK9/ctWwf8pVlwQ7eVp+UtZErB+QwK9XstSCm664qNKPtJxXG
re89Ea/7bkQQYAHbHWUwVdmxMPV7SG+MijOgHgRk0RmcL7nyz7AuYLY731LUfwLwjArOjdmFuIYx
LdZoEoEBAhZuxZPU4YqoBqQj1IFvuRa2cB6fmQSmxHtgFzCWjRPFZ0qbfyKDfIn7oYnAPjqPj50I
c6Xv/SjSpCGdVl5/MQu9NjASGC/oe3TqItBBGw9dVhVuD34OPPJteJe62AmpMKOVUc8mstLVOEJ5
yAt+SjRwNYUgeAmnnUjkAYHqtL+QdXIy9Q7zGYaGS09BUP90++GGcnSaZNUQ+fapZP82Cl/UUAlJ
CPRIeWId0xY5NzqETVFWaqZsUtcsqA375Ioo+tNz1bp+rLGQMPR18eR/K+Gr3pwoXFDrcWgEk5wg
XMR1kFORpVhkqKCQF0xfskp0KrQ64WrMLPS47QI04Hz7aurle3Q+YlAKEAY+A8VmP2gkeB8xW7j0
EY3ePcYYnuGeFAA1MMSbnGIMKIrGz/rrBdzoRR3M3AgmobLztqrZG3v5p3zYnhAbd8Li8j4kKSnp
6iv2VVfT0/6pX1g4zNX26Hkd5Jke3bnpjtyDEzxmsbsltf0V/nv4cAAtDDInG1hfnmXy/efb7UUK
LL+Wj49IU1dmbhWqp/T4v549E2gplVFmpXxB9ZifJqDm7FilUYBmBKaEh29D62KKafTIvLSRktiN
epwjrXRw9bCQTJqikBt4XJ2ppPLNe26BqYAy97ZonlN7F9gF2Yc/mtQaJcpOc8ZWKtTt6iaaCb/N
jCoiHGiG81eprhEftwN+qHp/rANRJ4DCWBTrY76xvm0Z/3Qm8pnXxcFMs0aEqdOAiZB1Cx56CQid
FLXBKAUYIM4w8uGcAIWQ/f2sjRBtzQ/P/DdmeVJe4HakEX7bD1rwYqDsGRIMn0KBHZ1SYQ+5cVYj
zBQsnR1fEFrLap7Pu4BRtCLtyIyXTzyYqgBzJJ1ZdcFgzNtKcv9oDZSXrXdtsu+j9ln17zdb55Tu
hGRf3rZaFHvBxeB6HFeq0ESAEuvDsU5xYoculWWNYajrdEt38oVFC/bU0JRe3HZcY2ALqJhsHaOE
tIPm7UXkD2CKDcrOf3Zd4kOkIgtOJgAYkhpK8wSbzx0DN7N2h50mp9buHq3dDFykkSXjvdWsV6kc
qDl5wwhzpO+jcB6f4NVQyd4ClLEfWQMUpv9Y+PhDhZxeW7wMma0U6DZu5Qhnp0SRrPej38XbGS6v
R5DNuAEK62zQ4fo77nCRZFd8/eOjH0HA0n4x4U8TKhME/kKsZ2nyYjHNR+seTYggzTyJCluX2iWK
HFyC24cTP+TsKY06PSUyyDtxyy7ffPzCSS4us4XI4IG/PsgYxCKZJ2eCnrLjoaiTqSLTetjUGatL
d0k/bDZQrRi2kQe2ZZ2TbrHgAqmalJk45/Ra5oV0UTwXSanQf6PXB5Apj17ihj4IpzF6oUHDmn4H
yCXneI7N+0bOmE+Jze72yOIiYjzHZVfIishebNqnK5heNMolP2JP4AlaNjdh4l7e2WwfM7l4Crf6
ZtA1h3JYG7x7Y/BN1nA6jLVuCteCCaxaeZy3vvjPPwyguCF8kvEF6Of6uYBr3Y+FY6cy9MFirjSi
K7VQ0y2qJGSnvDuWVIMzIqRpPBoHv2Zr5IhAD8SMsJKmHrcG0xfWv4dpV6omMufL3m5JmHBwdD1C
vMctN0iADVcx83kHY/dgPC8Bfq/WATFbZgq5mo2u/5JUW1EHMG8hIVCaj2KcTUXPKf1xLuAZfqLe
vEy0tyW+wWOyeANwoHJKFaspvoAmjfV6bnWTAn+goj6/686dCtNyGxiT9B0d0QDcIbBmdHWqU+NJ
PdwfFS8s00Xr1JHHOikeqWodG9NzrEnT+8Tbwg1wOCbPYp11y3AojMh3eoeSEz+mdCKa2OWHR0o/
TnY0wrEJ51Dbv9Pjp/A9J8avXhW0UFcwGn9mHaEOnxlX3dPpC++o7/qles69GjNMY3SubkjoMms0
lk/krOqV8+dHEitJwuchXt1u4b6rmihYQ5U+2YimuRUGaNM6NuB6EU+1sACbvelIPWCpyjLY+9vU
zFEZiZ+wT7rB/ceS4Gx8pNjTQOvZjqfsP5nP4/wEf4D6mzbCmkJED2MaeBxrKQJRlfaxHjicnfdf
oyRMYQlqO4neaTadDakQFryeXitbWHWt/eXlbuTY6dq4lDVwHw1uMSAti/XUTdg2td+lzg7xLhfx
uJZKqYcbK0UQbzyK5gymzOBos9YGoWWhB/fx96/O5jrs4qI539IbQON7t0w9CZQde/qF+rHlL0GT
rZNSiJY/IFAzdac9czCh17fYhcNPmk8Oa8I3he8hWqSMowVbcI3huBnyAgvOZxykJsYCTaEZBzpO
goPg7yipme8TvaiaK7lWVPQYQvEHfSjuGLrAPGRBLaI76QO2YmkcpKO5OoMq6LQwcKsHGAnTSRtO
Kn50iJA3ArmKmS0D0EIFbu+fZyuHGavn0xre7NYr+EajmqWpUDhX2getU2fLKNghqhGY51PYyZ4+
mjAa5NOUCl4kmxALeNsm33BFmdfnBlPMmMw1t0/IzhlqupOeP7mMghPovUqRhoP5F/wDaXQ2HmjF
Sz39v62Jy7w2jFiUqmexaTGPylLLDOmqRga8NDDKt6f+ojJ/K2QG0rf+3jD2mx7SxK0kbCeccVu/
04Q88PoxVh5UQ0xyATcYhatJRepmSGm99m5GZz9bwz8OhllV3FNdhwEQMU9Y5MAMFxfLXCTPIiOR
uNkMxvZ8kx8LMWC2Q/Shc+h9peCTSoZjXHV3l+KRM2BKakF9q9TqNoejtTi40ZlJ70w+pMmxSWwS
YaBXtk+9ad6upRVckBZ5nnk/j7ms3KY6Kw+SJS90C4+I5NNzUR8O3QzdWrIxke4pI7GHp21r8H1d
muxRJlbskvBzQ3Q0dbQhXRQlLLhp8vYyAHk/p/HDD466QLaStDNy5RM/vJM7I8l2QA3JsHSAxr6O
zI//+8W/jzGQu+uDtv+sG4tL2E5DmKQwlbMpvrwyNfus2prRlqVsLQuazV3RJPIy8W54iL3Q2zED
tYU5kPHfIEiGRq1p8YHA1CAaawtOqu5ovhs0bigACrJSnoZCDN8Lx6WZJerPYxE/Z0sMRNmWwjYM
HcKGYl1VHdxOW7JQmkMpfE/6vWIFESW8joYqqc8+S3lrPPkaQ+8RXal6lzQxhHcxcUZ7kHeSajI9
+ks2iZCKAvhjU6q8LuFkDMMLHkQ6zBkoFzL92OUSXzOA/7vsepf7KrNvWJKXqdOXOuI8jU1PzB4S
z6WHDtzZHXtblErHuBhfKqFDdJPDw3xNyDMd62Ney9ecVCCnWCBszmS838TOhTCdxs0DrtgR/w9y
8YfFztQZxOGR+7qDorQcyX0HfGmpsNxpFN2cYXVxnaCt5knreV+YzS8H4+Ph2kl4smEWlAejNUO/
8T+XI8GZGF7x0ziNWUuj9vOm1xG/DPhz6wbrKFt/lXNPnxh4sB6ipi8dv6YynjJoANPxSwpmrSK4
MARPN2EQZvrFoUkLmZPo6bQ/1i7hmnB7tR3v6eAuVeshpBevOXd/rQ3FV7E6TTqbsaG5I5pFFgYg
iMy/GmOZgmRjSUf0dKBmam8i2wkMM5nACm6WMkqSCWFgUURJH5WrVxSrqOcmizwqACwJ+jHGg6NT
2pKcMqBJDgJPudTWyBogdJN/dCx7jgA8UK4CNeQCHOL4FrA5kvLO+ROD/mjHoZaD9eJ+yfqkhbb2
FiVi0dqYqDv3LFQxo5P9cXjJFZFE0RC6QJqA6j0toDufTYs6Z+PivmEJ+2zgJ+96/rn7P7+vhEjH
8t3C+mAxViAySmwNkJUkNWj3pPc9Y1a2OidVKGa/KMCEl174zPE2oJXDS1mQ7ERvrI585ix7YiVn
Pb+XA4yDAZN9dryVVUZI6ShJgH/6LQmir5AoPakVeIj/rZ+0BkIJhuT8PW1y5cISKs2H36gpEbDR
aof/ui/J6DO4yL6GvgJENi8TF9ZkmK3glWppIMkQmhR1bfQjQ0Jl/b3lL7p9ZCx40wPmCFEvLH+K
V8VVINAvGEFHsncHwvDxQqi+c67DH88sYjwp2AHYwso7HAoSYBjnyYjZHxUFfy6dT6zOqLS1SeQJ
rn6aX/DkJegEmM+ZnrL9wNy0gRzZeigs1a579tGxEAPbtx+EY2eN9sed8dBSY7GPFqwtazfvQD9P
Xzc5PpQtrWaAlhc934yaKIKvg8D1XbjA4eKll6UolTlN4HsPamh1C6C1TrVLsxic1lbrIe82/Q6+
3MOA6snlS630RmwmMt5oVLYSBSsxFwD5VdLwyanan8Mmt2QaEkVFcBX5XhDwpAq3TDVOFkAEFiaT
s/jcakejrOVRobvKjEmTnOVYs3WYRuvoDJO+rYJRexS0MFDRymG7RiKyp7IUc0CAEZh2rcPPKizb
cf8lFeDzvND03Z7kRJ1mpBAe7iiAIIq5Oqpmhr0mYMPknk9tq7Oseek1Uwq/7SB88vN4F5orkZue
Y6uegOXqev4orJtqJgg/5gZNIArdy818yrCLn0UbrNuli4JMHOjdsq3iCOYcFxd9yP2guU9c5KiP
xa8ogdOwqspCNSb7kbzUnCxEjMnWVkjxur6Jnag1ei1UtuLoKuMXPDRzwqUCg4ixnmD7r6MMI7cl
5AdVOm4xdle6MhkIsG4RkuYaHg7e+JdP5fsCvf53wENpobSob8fyQgRXhZdBCyQ8L83WWXli7Kx3
hyR7g3x5JX4FeFiqEVCi15mjNGsOiafHPwBPopEts6dRg2JFU1YzDaCepxvCW+RlNNceByUXkmW5
dbzrReVJcfo6MnpX7p646TywEmpBdobLDtUE1mWmJAnnC3N1vFLwi2w5ZCq3sWPH1vkFEb6ILnBl
Abvm/SQvGEk+DrnFYsYnEnfsCI6Zqz5S3LO7C09i1dV33XB7RmvtH0vhW1tb7hgqLVdVnGB3Oz4u
5XW+65HBXmYKW5AIqIb9PPwPwU8oC+OHb/RJKP/Xc8LCxODCnFucS50wT2ggG1YaqnxGqU0VjAl/
c9wWXLNYG6Pt2C65fayXOeGP+Sg3rvxc5fdIuFXi+OYe55ZhJ2PUIKEqgt5jq19Bim5KHk8xPlhz
EpVI+alNjFuL8N3zq5NIIMFrAQ0vKcTeH4QlmGXTnvcPaXhxWsZ2uDORRyqP/9N/oSU/ZRsyH7+7
Cz4XOtNCAGVvlg+1xIJ7Wa6iYsTBjDLcIy6sdr5Rn9MXWS47655K6uHw8IzwD3elh3NSd+OAHyAG
sHTo/S82etpeNF2v8v8XaKEsTMi0GSH2kCkUkUKuVmQw9/maciglEHWoaCFrMiUBQpkFdbTHn0ib
h1k2xlaET6/EYgFI/Vst+njzYQX4XNcthL2831PC3uqAd+rUckcpQ0f2dbc8SMQrvApY41LcgJeG
xcSMg+lp1FUt3t/9zSa0wzCyTIGRSUo9W9V106Ef2Panzulp8I7Hw/3zO/2BmKVCOeIfh0k5MQoQ
edw1QzRW/yFcvnG/kYm5z+HG0a3bGgrXwwPreTY5Pjh6q+8cs6tvZSjMKRxOgFjR8+P6ZElmU3cT
MGavYkrC5olSnUc+EG9gFCnuHAVNpT8CQaaSV9QJjNKMGv38a9MLjw69YqptNpmSIPySTy/juWrc
mHhdIBUs6t8s00RAMBZakHz/LWWzbzF5wjtu7ZKdfPERgyN+kApKKbEm2VKOeMkVetFFQc/rjdQp
mcFSAc+qnmSBluZ2B4lQszraFoNV+0v6gNGf1fnU6YxeuD7/WGwKI/sOhFvlIiI6dvzmu6dJQZUb
DcqqfgcevF8z/RBRCZRQO1i9G3sM6Gk+0R5nyTtiQB+qFmr3GfmgBxJFFH+5vPfbMLsunuyJjEVh
orYLS/sXkYGNISUOvDM0lYi4vY1FhC+FC6A1423/3u4W/AowJw84Hpj0mbcBx4hiNUpp+TywGLOS
/TRDISXmDetBk7Hy1OlU8aAa7p6aaxNueJfrJBC9dr5nQBTFU3nmO3qFequqhb8gouDDnn27MHnS
WxTRVEz5kcJOln4qcy+ufsUYfkyPCdY86LsjmeFlh0ZHUnrc+jChCiU4L5KsrN0Na2z5MzdUAHq9
SzPGRFlkwYX3kr2lfCnVzozfc4awLrOQtoDEC4cuKpXIWuAfWVYOSZl6hHv6WbGx7+bIGbn5n3dx
EirR1f9Q7gOC8rTIfDmsb6Uv5Ny8B1qj4fRiB2OdlGEam8UcITN3DjEdFq025NcykJPLGCMSaGJr
tdgYNlmeNFBfmk10on7yyyhq1vyY/CYsh9J48To9k6jujqJWC4pu82++IuJOF5IIMStNBVTFLj55
B4GwfaMi54ansbsKpHFZOq3Cg/R4JmuPsOeEmaL4lvbBTXOUyY1K1Xm9R37kWxAT3aFKuwfv+SqX
5Dm4GdjxIi8LmEk9aeOekN7b9PVRCBr/M7Dr8CVLCLSvmvv000crps9AjAJfHczIZrOM9oRE/tUA
/JCgUQnBZlz7reUeSfbGTFaXAZWs4fhJyFltzWD7/pyWbi/OcT0NbgJsV4YaVFxgjfo7GQrb3niH
xSwNBIoNRzm0pHErhW8TytjVcgN4vToTfZ4fyTrluXpbM0FF6oJxl5nxRrkIAjWgzb6yOXMYIt1R
dKJvNBlogh3JoGIPfmm1JJkv1WufVbxGHkzqIU5FEZxTFdj9dcF0cnaJgAXhCnOLYopOhymrAWoV
gw4oL7PMRyWHvrRBU1orU9dYekygx0qg336FgohadttT5uEkdxk0fjYZjvkrlFPLip6UxOPiSeex
zmasKnE807liXQSN8ZdKBemyDB96S2x9r8EyV9OuhS2ZuMjsEus5UyfxLTENx8uN4adEY06XJZ7s
O4GnszNnCQFIE+sFBRb8oGl9LvzgNwVCJsE8xST6UAuqSPV3uYU9a9WO0wwLFBnET5QMww3+Ikc2
zbhnsuEsensSXnJ/kFrK8IUaj5n/dpC4FGWBfslOfxEAmuojOFO0miNkcmES6jAsYjdUFYOahIeV
TtbQg4bV5y1aeQ06TOcbr2kRGYwjFFXMP63QV72hnx/WxqYnDn4E3YzB6f0C1bXm4EmMA/SqaaX9
BhR1QOkcPYPAj/6IyYGpjiDvQgyjFGl9CcyBpZyl1rRIjuHXQApVEOqEltUc8Oa8FDX2dHMHwGhI
t199ShCTvZ3p0HhkTloFRnH2h6jBo342s0T4uF2hfeNutgMZAbbbKPqmI+h9d5ZeadLEgXY6jLzh
sYZnwtt37TTib8eyT8ZTHjQd7+KYLym/Akkv9a0E0jDxMepv/JikqQ/6YOW+YqO2eqg8hzulS9AV
kia2MScQ2BYxkZYSSlBNfGVEds0AiDMviKAfU7P/xUd6XepchtJy4GfcnrNxR9PpxhVYsvcZvNVL
umzJy14lBZJJgnpmg/HiWTKdZiXOb3p9a4EZce11xo7kzfigEelcxdG8UUUqFxNmtnUalfdvNCzD
tkPmG1i2OH4m22RL/xWUwhe1YBA3ISUoJIWfwKiDK9IhyC3UiRnSwqpDCYirRN4TO6XZDpnCaj8E
c5TTzDv0T9j0Uwqn1QixEYqCQK+rvijE0lasSLg1tnolkd3WSHVfrZQPse7H7AWx0lUM3sS37fPY
w0JAzioO7EgKvUuIa+AiWrCnSBM9Hcnsq1uBTKLi3u5DQdqYamazzgq+Mp5p0gFgkexm4l62hVPD
KOlEXY5ewfvLGthGauTZLi0lSf0fAZTkSc+iV7CtRupqcDiki0ZrQbF6bN7E1rOCJvQxtPvVmN3W
A+F51TG2lR93YWKgK5JOwnOW9cFtacZD5riRl3lQ42gAKdtB3ZF5OC0jrj1ECcbjT8Il4syB+jq+
qQM6Gfkv41ThevCZEEZLNIKKjuuN/X/BDFajomGvL4pSai1Oc0LZLQdJsjzDiF0zmONlrjrIpUFB
w/j6isZ2V+HLAjLoVAerPxR9AWvpm4Ph+x6bKRJvFN3IW3xwwxzFBybo+B2wG/drNKgL2NIkbQlm
ZYeMHFRm5uSXWMNcL6RGYNWyUwV438YM71qyFETvQ5g9D+zxiICUoR6B5mmsxlSBkfvuKjebpi7+
R+fvQN4eVDdn3ZutPScbMBvDZA2xt9ZS3pbeWxD+x9YpmPqG9eUSew6RvywkJXu+h+4ihTlobiDI
C89RYGs5F8wR2GMitlAFoIbCzYhS2t5TpXdjykgTo9ap8ZPGgL353Xgtn4l1mYSlcsdqB0imS9IL
4zmZRST/IUlkTYVLMjqLpX+mgInb/VxoBHQ4hlrUHm+wISOVv0PVW0K41RkpnFMrDyS3949WFnhj
zBDd1Je0+TxnmXnDRk75LYr2NAYxnRi+57jrDowRofnF88U8zzAUALpCnUkEd3GlsPwYriWI5ZMP
pI4zN2lKdq8GJJfCr4E3YYwTvPGUdINw6tMIw8rn0b+pxkgWe02bBZcYIly1sXDujf88sIfwpkvL
jLBkUABBdXa9VE1fzQUF+AmzXjODD2XKsmR5uWE7S7uxAPpPfoJGzzfbOfmNu33Fe53OCQGym0N4
qKg87WX/xTnIrOKGy4KifkxSiR4VUAqYlOMuKsJj1YaXskXnvEkAcNm6cfxleZcjM/G5Sr4HJj0D
VG0Hs/eCILf3UmY80nIs39s2YmKM+zuzwtt/c7IwgZFAMQHSo3hB1otU+flBOdbpPFG3m4QCmmKF
TcXhoHzjigIwkJovw+5ffMp2spCsMGd4eASfd68AStuVmSzJL6gvAEBOrI+9FYqmXTzEY/K+tZ2A
PXnTNXuGPXHsNUNNpC+rmdgAIdiaaz7NVM5frvJzcknXELGYJ3RsfgDr/7ROJb3Yo4uEvRAp/urS
v/LxQBysIsN1Rw95I/vKlVc7eElaOGvEMNyrYMjnjGSxZ3sEfFaZ+/wylkOXzpfsOPWWzgFvEf8k
AxMXhmbCeL8dsLVp+QrN7vZjjdqVdmmVZFAKvrj8X7FOI/N7DnEXhGmEN63vXU/+F+x2kA54y9AP
M2rPgWMY+Nf5/1IZAzMe+JngNpbOZhrrdiXB4Q4tGGlSzVoe8eMIVpuYe3JDx7lxZG+CupdntSPe
a0zxMX/7Mr7arvN1aT6EJds1gE2CY5i6mrgxc3cDU0kZcOt4NQUbn1dg0rK/f9S1mbWRpc0jhh3C
59dZiBV7geKbabJ/o+JtLERdnOdAR9sVY23g4AfkQgt+0VcMKs4Jwb+ii1I2TGsMFkFXUEzyJfAg
Vw0meRO2Foi1krrCTrLjbj5tQkVAmSZs3R/YA1pId8Rdeaggw/ylXV3vYU16dwg+ot64ehG093Vr
ZP9Es0Cum9cOp9xka5rbjuP3ZEMxEDJ+AMKfJ8qWpOi0NhOwTxOzhil8hvl4i2SJE77Zp2fSGeH7
44+ReMJErrxc9jbBeYFsSLpVx43asEnyrcK5xLI82Ylh/V985Q3EBGHuVYzKzWEs/NAbr4nx0JJu
j0KnrEcwAf4a85WKydwrbP3R6oTWPaCoxEX9v/K0B6MmOSXys8Cn3wlEzDoHYDQrowFnwm5GQ78B
3wxlYyBbsd14O1OH/i9vF+wwGsf4yzawHCQbYQVq0q52tj9fBSJiSmQ3lxDbI9ab9ir54/M1GcZN
Nj/lgCqrPihOBp36eLHxXcxxnzgNzmbnE0/EPG6kKEBjvPRw2130duNRlKspzdRnfa4geqUo4XYj
kgGcbo1ngldHdnnQVOIcHE/IbTQ3JX8J3gdy70M34wVH2FFqb05Ir6ST65/2Lpmuu3h71Ikk/gx0
Ob6w84IEn898uvycvPxSAMEYv68O0jEJijPQ67jZwCnTqXCqpV1CpwurXoQ5bJn1PnsOJWJA5/YR
oos+eEEuGy4wzgYovMGawKRKdlrLIIiq067QDBTTby6qPFeVOdxYJntK9/MebNgQw3WuT7GBERbr
P/+KL0KNjPp6zMYy236XSzhkSvK2FpktE+wI4q4b6YviwBqA9EL1aWb6KZLBBFrnZESV3txvTiN8
G0nkkwU+Je0W/6uazk0jMsJX3GkgUm5HfKtV0Vg0THs5V+AI7Dh7QamdgCtLK7kK4Ouc2celtSDX
ybBCOdZPXeddQSyrfGQ50YYwXnoZnecwNHRfY3vs6tRVWEXMosJVUSWOThmTwhYQ700ujYO4auuT
Cs3YMQuPI/IGF/wWQ6QCCo4uUWPwbEiC2Nez+8NTp6vJQ/77zyHMNCzNsG8P6R4AHoeUZMv9V1Vo
X+zUI2uf7lcT8TUYeue2h1TzgoyvheQF0CKo7T/mOejWDQ6mVuWDpW3EuUiKCSiaNbZ6UvazBqGw
TfpgPDQnfiSlghuz2FCE1uBcGYF5Ci+LuwrgAsYK7U/Vf/hNmFfroDC7oETU+dyrT7wfsiC4oiUg
tczC0077dnAdnzocngNW3i6836o8CgfaJNz6LF4+xmScsz27nUIAbsEOyOAkzt7DthWe6h3kjB3s
ZDkxE3OM4wXZoAtDdW5z/FnmII0brSyZZ12mCBLNgWXRVNKSGmurucA8Yxtsvd0W6UbGF/+cp5+7
uiT5Q2C34Tw/nY7P9OFS9T0/7HFhOlAMj0UgJGHvSuWkXbogvmOlrVo5pp77P9mIbMHgSdg2QaOH
VC4Quq/9BtVzPBmUtH43pZyJep1M3sDZlJ8ur1lGKlNGz32uykQRlRh3GgBkFn2/ikdrwAT/MrE+
BK2qp/KXf0OR4jDYPOOL/b6bydBgkfsxeI3aNSmh3i/cxU80jSX/BZRoGF2FAZnUTkfx/xi03wZC
CuAS8xo0neMDG6TvVxoUlYuRFVaG0yj6EL86wK+XNfOVjKk+914deI5JOxtZkCgzelHWMd7qlAT3
bqK+pLLfC/AOKfOKrFa9+8cZa5kTE7V2kaWnD+nAeHieFQ2HLvZ0I3xLCRZzrJHNKxsu8KOfQIk3
e2L3aH+KElVTFiw56Pnu9p1MsHLVpu55RQA4GrajwLELcjjZNKnNcjki2+MptvXV629JceP5P3ds
opR1WnQqNBo29/0dgabF2ymt05obSOP+CCBQszfxvVK478U+BL0Rp4ykWrZd/W1flxc27mIRhfq0
YoN5DbN1k/HM2OWq267TpjYxd/3ejTnFyKGTOA/1UJJk1A/IxSkfgrr3x8XEwywnyKHb1z5qebNU
Gran0ZvLnqWzcnff+1XwrGRmI/bls2JmgS9LQjBdKoR4mGPgnes4p+wS6aqvmODQLqxfnJMxGeiq
7yjQhLgPxt9meLd1iEcZ1oVCf+IBpWKLbD/Nw5WB0jLt8c4LvR+hZn3tiaKxFzQQRS0Aj3iriKLt
PA5LGhgBcBk2ivDoe1TP/kzgMV2IXytinMQNeIUZWZkJO/7inrOtoeFqmlwFg3kZWirM/BoUlnHk
dJprtujmoxq7jSBUKQyRBYf0S0+7GKVOb6Im1bH2ndCBMCz2MxWaw4J5oKi1OhSmC/KTz2iWTxgk
BdQNfpCR8iFNpdmMeItKkIF/vDpcdwiPJ91qlY9EiVQe+eiexcWjx6kt2zpOigQdQzrQ7gz+voGc
uURxn94UnpeLwlD3fIDBNkrF4ypY8hYRFnXrgqGxkhJKvyvUz0Is415TTbrRN79MqU3/wMtsmLEq
wBbe3LDZSbHb8CVUCZJIu1vH+UtpkI/HdCoJit72GAgSTEu/r2SV/knTtUQZda224m6Ol8T5HiLA
V0i6/ivT6S++2xG5tKa7n90u/TMG2yjkgm7kV9W+9Xq9LpHq8NFkiRdLJFiF7O/hwUd4nKRuAMWn
QIQPIPLfgMyanbMB5nrkWpp29kZb7VOjIGSy427yeT2KEAM/h7bJqI/fi2mpxzoFQriz1Xr9cHCg
kfJFy4yJByE87SQZv1G+pxkcXmW/g8OTW0Lrc0Jraxt8SuI1AAQhKWx3zcUVK7qoS2uZawcGcgK9
pVe7pqHa2bgRAq/27z6Antu4rWxEULJR86IHzWT8TGDCsS4VpuF+sMqkv7HLOtSuaR1nN5hwu09q
7vq00BCCI/V6szQjw+UXs9dEj2SD6RIu9AUWYWgzKLMkKULs4sdnT5llQIxye9kiOyCf9Bu5P9ev
3Xbeb9grJcxPYmhMRuiYuEDjW19f3D4CD6z4h2s6TWxCYcgYZ2Chpt8tHHDCiLmTh9EQv9MI/01p
3UIbq4Z7Ibe+Seot5iaHLQukGIcnTVK6V2Vm/1DThEkaAw+RpoSOBeKWR4fYmT+qBkxR4Yk7Pc7P
/5yMwzirqHQdpRbaHuMVdkoB0UX3lMByU6oVQ+i7LcmwhNSTxkGBeiE4PVx/34qJzYtl/19cVvb6
Nc4ORtoHADhtrIfvRXH9e/PjO4/8sgYvvF3wOBS3Vszr+g6su9hSAfPlNI9MFMwYavv1ZBSF9zHW
QQIpqigDljqmOnmte8ZqxTOulV9u1EyrZTlSBPR16exxzu5ZY9SDNiv7WSLXBolcOIolWrVkz/3b
vGIIi/X7siD5A/yJHeHs8gnVj65t7iNyk8w6++sSxe9NeKC61xiwrqe65/7sKDyw3U5Uxes2ZLiB
Sf3tvOT1FBI88+gGznjbQkftoFrtbccAyxodRslMQbfZSj8o9R1Vk/XL17LJahQp8/Q1Ju6jwUQS
M6ZUbpsE6nJH+cP79tmIUx/Mar1MKdtPj0VbijD87cW3FMYiorye/sMpxUBKXacHYviO9N9hmOn2
j/Gwb62FfO1bqvKgUdUCyBYVFrvO04cyWYUZEfCPEFzdW/GkwGKYNyy8uvD2HqXWf1nz8L9yBwBH
GjKCfgikbukUJ7AGJR7sqQpYEcaukbBhNeZ1P4dKfpP42c7sJb7afo0r5IQ08w1t84ZVcBjnXBJP
TLL6aqjj9D3kw2VZKDTSdFvmnYtl4PXVD/EXkQC1hUrjCUyZiJ7RWMnTXMVBADr/r+21tGALV52S
10kF4veGyHDvwhalydTER+vTZaQebejBk+0MxzR+AXUGWDdO7wN+LTNF+rLWpzk240C6VpFECKy5
exttINq8/pKZCwFRgsQ3oGF8OOsrzcoEg7fgZLXQIRXuggeOIuC4+lkk4qmshWmZbhYk4AtAdDSb
EK7N34SuK83k+vAYQdbEUITcX4ZzT64gXUI4bIpTRhODn6V/wOjxI16qTWBcuu8BWXXVjuERJtup
VCDUcDwyIpcpauHL+LORmyKFUNapni57lc7xF/Gyg3588PTEcEb/ZoX9UfwzD20/0G7M5H5AfvYi
IrDQTqBgwJPEx0KCRT8ceibr3AThCzJznygK3CncrkxaYggzWpeyKmPT3hIZPG7pX3FUGgA0rNhS
hQCu/IyRUIZYgJGOy2QcE10DsZ2ukDfwWsvPYUYncIEzD4db4/zYezK88Kt6ceqiMbEHURiIxkCX
U1+iCTre2sw1geq8dr5/NKGZBNuabMq8FACXgAVP/o9EM7dOzHh1TUllDD/uY++gXWPigY11LDuH
MqkLeuL6U3AWjfPh1bw4AbbQDupPMTO/NJWIo/CcmMXa1NUgUZ+5wBXuD/nxn2AghA0uvA/mW+JN
lh3l/GBbJ4yWb/A066/GZtXkSzOvD4AKJMiklMMTHAFjZ+Vpkx+n24aekG9IIGS9m7ThzMicRNjo
rlakSriMjf1GdRCsL1U0aEwNTdJfRcNJrE2O+SApCxC4M0Vuk3ecOV4lYIHfMXErAPTv5BLN13oD
VcmHI7ZjsZf8J2rtShxnIrCag2BC9Xi+OgAzYx7F1Q+JPv+XKgyWo4GrkQfS/Tc8+ElaEo9nMs0A
HUH07Fgfal27RtuZESpB4Pm7AOC8gkgC+OrbvziHChb+LvUfd9W8EIVJjWEIZDP3912DXdvmltVM
05wsc20bG9h6iTmxOQ2eIiO3DLPn0XxGtwHIhg7RqFSeiKfU8Zx3psOpBo5bbbf7R88DQozGYf9l
Ub5cUBIV2Rar7T8xM6pfpqrOb3On8M1ELWVmbFDa3ewjUvZhw7IF5tnwPfC133ZPNOcSTgkZuUjg
972R0hWdDdEUYukL+xPgOnvBurqn6U7hbYph1OU7eOFUX9H8aqT0SRoHdcQmU+7Ma3jWVdDYyxBA
ub/MePTMVHamc0btAvIDBFqFomODa6pmIjy1GWgn0RPjG8CdyOK7EeNXfgH+5ZdhYisWhks+bkkG
ZlV8aPZXtHoN5B7RURkYSTmwSt1vHTNBhfwkdn1qfvFWwxvp3wsgWdPYwx5dGIG6w2+KHo3RN+TD
4qItRyZr50fce1CW2zB+nl8Rj2bnKbn8yJRRGHyD2YdrdASaiGxvrpGFQlQCkdTsVSX/lRBr0m1l
/tgEC8CS2cA6sj9qoQvXMpLOqY9w1owHRFvxqBEq6ynjR/e4T1Ma/E+M6VsfB9Q56atg07Fn6dNL
CyVEauVqc0940s3JZ2fqqis31S/eIbcMJgkL09h6u8j/iOnYwVkzzfCdXlJ8eGUjaEiA5zwXe1mm
gXSigS2UZtjfRViFhdtbjAapIbPyouMSbmBn9hMA0b20DVL0UWybLqDwem2wQa3QvCiABJ7XRfsh
stWlQZw2Yb+Hq8JmpDv0dyXHpMUTDDbjWcQhP2WE7lYLOepT/7P8rnEFr9NPJBA4g+1o88nH61Df
D/M3wZCx/85UbCYsUCTExDhgQ0w8Tc2/vMAaGojFwfEphojXYlE7qjhdKrUndn8PQ/6CWVoBUMZx
8wV4d/mhVK/BQg5ws1OpNjDkNLohtIwJG5iCO70MHl8oaUXX3JJA8mz0vsfeGvavX7AZz5gYeuDn
8DT5TDDzb0FJcpAZrdW/bsvCvdsH3Hz1oimGakZwEfWkDh37+MOc68JMjuJVZSN5gVHc0QNT1esw
yGKwug9uAiVI+lBdbUoJtl9UdmM5DxfFHH9MgaK/Tw8z/KOfR1zK8QD4FDPMb7IyZkq+alC/GIRq
M51LCUAm1UzjlZYno1MFxVxXCriqpMSZqPnLkLNaM2P9uUDDMh0w5yHXAEMRSjUlOBXxZ8vkZIc3
AM4E08eyU1Oz9hjhrrPz7aS2Qy2o017oRS8AJP3BnAXDZhhcsUTtZWr+ovPbw6oPrd8Qit7iqcp8
5cma6BPB4QqfQ6itLxesVp8AYtUdqleYYeh13MPVD3auZD8wiFV6OEDLi7kvjsdTcp0zLlW9LKQ6
yl09dhpbtqvTukKSACcic0az8Mg5CfJ3PV6RHrJEsl1YNHTcyk/6kELuIXs6C3GTGNiLtzHccWSU
fbyy5wEzv67zXWaq+7AbxdPnLOMFoQHZw7AEVQGfRzSyezuT3c+68K5FI0r+CQov2XHwrpu7g7y+
dcL9WL2oXbCDpSQlZO0CZIgI7QtWu81IvYAjBHzLUvth+pRqN5pLpimchVuQFZvDaVLogQ0HI9s9
EH51kKzxRlQPewYhpb2IOSjPYdMmw8tNgBMq0FhGa6/xZAljupRzuVXbhFImgO4WcEZa6NyoRupZ
tLwEat0rA8Zp2FXXmCLJh9q3TdVzH8Q6C54jJLk1Fl90ozaaXO3uYiRdu2Tf+QLxGXBhKwCDe9EJ
ww6TZGccQpaPLlGVsy/6lM+pIiIpm6sGbnY5BmvXNqnneim4UHEhnAxhL8ZQt7HY6ZtgeIA6Gbnn
OaH9LDtPR1aHx376rZXzUXeaTb4mwDblG88wAmZg8j+znFqWY6DPokcdgD2bwnYMCfS/tYj9TooN
EGeO8NtO1XjiwB626zUJfHJN/XKrWLGEl5HJi0T46g6XB/TvPxJ4irhsyrYYzuVBtNfErhUv4Coq
VI3uXt3xuoj0c1iVmdBF7jhj+GqoXov7ue+SHJbi7/pFIJGM6FrVncwFICf0O5bwDWwwtmVc5Hvx
7ySQw1nEjaCgFAujLtqa3wGnkganwnDnDcJ4R7OPNAZ7V8o9PesDzcrG/9X+deKDjE1te7nhAOjD
xIkJ5aJOZuK0tPPy99G8C4E8vU+qHE53Bi9Jzm41OasyB0D8LxAg45/kY8VvKq+12v3TfHn89XlX
kbI1xuXkEzM6tC6C9aWcevdvRrIUQVRNHVMpCm27c2Una9Qlwzh4gMscTkJR/liIOCS9tPQrq6E2
ORE4H7IsFi6X4EIggSzRIESxTXwfrWmnYUV6RxO/GUAc9y1RQFTyFWfQ+Y5cS7RrypW4OoW4eTsK
21Qtx2Y3IOtAmkIae9V2QV/lW5GZXPhCrRStD4MN8FUPBB0sgF7ideVi1cJUgazHcyuvbF8fFvON
sB3LNwcm/dZkkhFyjmo+CElVNxjmDbAFRMuxIsX/N5LIzY4sutIqwMetNQR+2pS9BmhFXvi7xIN5
81hQb17cce7LYONkcR1DIiDgUiZLs1knGvBQJxq2eFTTHMCBQVueUpsidVd8tO+B+faCqogIFUEj
2tU4XP93wQbV3k5aASqqi7+GW98XobhJo+EdbHbVo2TmUd4s5sH+sUPROFOtye6Lbiuo6MNQ67gM
ASCN19/xBfOfziLQ1CDKHB7J/+gOdpo9NREabQ2BtgFSfQNm9ubh7Ssi81p13vnnnpr1vNQ3qcL0
JLhXyCAqI7nS3R3aElGEkO+gbtUpgpZleU558zxLt0qWBqC2QaxES2v2m00PAVN0X/lrWJmrQQCw
o9Dvp6ShpGw9iURXQ8pRQs1fvG3lruPmN6L3Q9ptPezh/t4zu8GwLjkDzBLNMzOhudPDgoqnvgAq
4ZRttk/uyOAsYh/9XBVcHTaPahwy7yF9MkHaqbJVAzojsjbtAYNSOXvxEOuu1XflurjizIfLq+OE
oBTnHdlpiioEWPQDKMHLVtvoGbBETFURgr1BQnnagD4iT+/p05UpEL7p0j33LQuqNHt+nIwETy+a
dBkbnPdCyZx57UdZ9RYKVmPt2LODGFdKAFX50SsVck8b5205HO7cU8YPdccDQR6cpU+LoSLd6pbq
E9IPw3Hmv4NWi4BNUcTtMilivb+7otqrU3xQDFA9aKB/wOg9A+zHoSltpMsQ9jxQvakRZKW++FrV
CgS8UG/zMzrWUEb3JQj9Mf5Nql9GqYY1kJ+Y8975KfM4M2rG1U7VHlyC7D+gHuJlq3iiHD5hPWkC
2A5vvWcWd44fqJyMZreSrsxmynhtlh5GP1oqyFy9JeJfL71HiLrZn0jJaXJhpiYzLwOuziAAHDvo
XNGaF+ECRje9zMBXr7VYvGVJbTP07BovjqKpOgwoErld8pWIBy2aiNQwB/DdqjZ2sP0HkXzmf+92
+AiACorHlLY2VhR32aJPerx02dN6IhsL1QJVdYibkKvZmNXcdeX+qZzDAqkLyRsno8Wrcuexj3MC
zlrzG1ndonzG4QfZr6KHMvvZojqWeofO+pph5ArAmemPf6X5k3Tif3OPSyQt2e3qhzetXnWHHsXU
icFWKy0o5eH2ilSQFS7bY0ABsLzCGg5Df7fsC9vt7saUTaBXzhBeySqYEMqB8Fo8W5v9VNUfGyjw
CeJEQQPjrYav8urosE8VoyDuKwPVQ4ZFZvNhmh+PfPB5JZi6B+UUapLwJSso1MCQptM89rPYUJ1B
olvEXd76Gw4aPvBced+GD/GcsIBBw4Hk056kZBdiW0TOEOwcG1FpoQfXIZWXv37Uhxl6RNyczvJn
X5l159eAKSp4gag9dzjnJcezxJVhmENvpee4j+yIW/j2IQo1FL4r/57eaNb/T+5edu+M8hDqhOKI
ZjKrTEBq2BYSa8v0kt37bhAwZXdXV+PtNNzrvwZ4GO15TDlMIuqhp0yO4V8cHNUFePVHs4HMywr6
tarenTQUBjwTKII6/f1I+BRt52VP0XaeJPa31eCcG2hNcOhh5qOD4u6gzzGtw3as6Yt/masB1RWH
DRfnqDuo+V20r0Urcny1RNcZQ+aBjZo2YHQa+X5K1o3LGmNkBgvEzQKQGrnBD75jsf6NtlmLwdSY
ZXlLFrpVnydQqVAU4ZWFioWCcMkzGgFQJrFpQfCBHiVSFrOnFRCyjvhM8INy8x+0BsR7r6hGH+t6
vt6eREM2KvPcTHZrMvHMRbgavSlwe5ArveukV697GsHNMNrjyMi72oGYfKLbzaWOU6n7ODyHRmoN
AuIdHUUu/PUNsml2y/r+jKxdeMsiZIn2nmY1tZvINLyqSvFLsb2/eYSXo75jzUmSr88DEzfQUdoe
ALx8bQ1+h7ZQRrr3Q9TzEP4zXm91VABYnH+ekHL9Gd715fphP32wNTkI6xh5lOiMKaY0HfthfcVX
iILPjbSzqbGg7mkG4JcchzdwzF8ZJGTFXj216ujsD63qpYlcYDb4z3RlCW8KaAjP6/1r+V/mEY19
iJTKPdwtYspN8chcz5ZUk7ZqJNcrdNbuggWMVX6ujNVI0G0wUGJEeO/5vAzywVh4qdbR4G9CZ+TW
6EAVnHZM7E4oxu79f/IIeskdbJiKwgyvpdGhhEyZ447f11782D14MLZQQ015bJq6Tzj7Y3iVab+x
v4cPsMPWMQ7mUcLoEcZgR08cOtFJvKxs28yVkYcrMvrRzB856O1vGK9gflHqKqSmlH/EyOGhbiX1
94WUGQ0RgC9KT1b/IuD286ai9kJOy7EQQbOplOgBauDtZrYonSiya13lXj1/uJxHQ3la/PQ/kfLZ
QxztV1CGxm0HGtCqJBCpZYcnU0wE7iHq7nBqE/kYuu5TLsEoTjlRZxym6gEC06CfD2NFNDNNbBxP
uWfBag1NI3S7WpTcxsY6YJ9UDlkuj9PoH+Ca6d8eB6w3szX9XncWMmFo93FIxfnFnfwciu+zNK72
UfmUGk3idInaKRNcc8FbcEJ/P591oZngGTkodQaiAI9blUSa6nBgdiJYu4sr/vdJCc6otSlNuWHW
YDh5fpH/gDGtu7tLdeoFFXxrkFuuJ5MBWXfb7/AzkzUDJeLjOG0eJV9JbWSmjvZWDuiJIwXh3e6b
ntaweyLXDSXgMKuyVksxjjmNDRUDfSp1boO7YY6N/sx9qu8OYP9ShXK/DGq9qIPwK+gjhSstvKOS
NDyrB8zPgnvTQdcm35q9pMfixmLY1eZpdZtbykPayKo7As509QSNiHGA4h8V9xXietL/clWsG2OR
/ZGFxjon6/USXRAW3O57s9GlOxLwFfAZXLAlq5wdhjQUD7SYp9VY13+MlT9t6vdbt9tl8oYCbX88
1yUNEWScI/r0Zz8l8ddsONpgCm1ia9Ds/nE2LtBUzYf7UHPlqoJVLPHdXIBE613GT9a6Ar9GM6Ce
BUOIpb5dLRdsoGIC5vVemS9fatgWXhFgG1zcros9Y5xWghKHnGnipA+K8ESguf6OEROyCmQKOK4Z
SrGPBZaUfALyjI5cD16/Gw3ET6GxWl7BaW+TNA3qgmAQhOhf/PCx4zE89X0HQOGHR3hTbanAKac/
1CAZg5QK9QKDNnCmvA/NWsa37rq51kqUcGMWTkuxirax0sddu8c7mhXz5Dp1KwP8yaDzRt7Prueh
ZNvCLSYxQNe87MfmtbfhpuBtNwz66sjh/O/eGwub7DYPZzLstGjMGUcytTRfPWhgqW8ExxRBvMXa
W5JAZtM1sVzdRk1pfCrHmgvfvChKZ5VUAEJPLS5nK1zrdpIVJCcJyjxy13S9+KqO4DxsMIcAEF+P
pZMWvVKkc2DPawwnHb5YMMNh4NX5pMxTWKEbFZuKBVGndgvWGM+x0IgvatsW5KyjyDzO6dvB1OJU
AfpT1XKna4tZE1agGPWSWrZXA3SR9++1ur1e139DinDgOOMAkOqwFT/3Ls/umf5/cwmm+eijlazz
csTxv91yj1ZCGETfBnwMHxQ0lGbUGIhG5cNCl3idWQ3reJQZ0XPP30dSO1oSwlaomZzISjT3dj9z
c6Nn0a81vR+FML/32omHsM67JD1z69tIQ1haKIh2LE57nbmAqw/y4pkVTsWB2UO99aKLEWzY2hhV
tgFhLBM5iSPztAzW3azuTB9o7NLAZ6FOCR4LTmZhwiIeHbybE8+z71urzhrTHaKK4nPDQVqGHxO5
QVU9R9Fdv+ON/3zxgIJ3d7zfe48auLhAn4okm7izBSURHUxyFDczBjXa1ldZ02WHmTyW8l9B29m9
PliWNShTs00kDcltRyLCr+dkpvsZZWsOnyiDIvyiPczIwiom/l6QZze0nXg5rUW3m8mkYKOgq9lJ
67nRIc3JprFMIec51ULludg7+aUawAnDWWM3bSNUjcyoQv8fE6Eu2B3Vss0OC8UO1vCECJhcut68
pVFr0gGWCDXKR416VcpsNMZJkMU7ail0V0a7na++UZzMNQqHsq6TwS2TkQjUn/L/I+/7jDVsRh/v
1Q44S7LsFeSh7bxKqVinH+GbUaNfV1BZOIO+nM8brmfz1kcKp4xkeUAeU5iM9ydL+oag981uTENw
Af5s5Hlvfyb9JW4wCLN4xgDeWyC6BgF3pQzROgmLsAtVywHxWhfudz2WguyYpNCHml6saUqQeQ4o
Sub+qHua6koNK/5egByfvka0dGgQDyIqOCOm252bSMEgTnHbl+E9fI//RXxIH5goxCQxd5nOtXaO
xCocKU5aVd+mp0k3fAQqKOlfR7bysswUjvwwRq/sgXKahENqtz2fV/rgyTSH63KwzVCfXxKYtSY/
BxfZAAbZK8dW5X1df5I/2MHHcB16Uy1zKKSfnE4cKPb2GP7X8naUSBHw1pwjK/37ZJjKSX/khFZd
/d/rG9mImLaNajGE8i2G7DzoShdXBGdNU84YiZVvzTRW/qGnGy9uqLFrbis3eFGHsu6DVqYqm19u
AaZuCBNLM0RvpzmQkP4IcqTvK6/OCEQU4teXRVCppGEmfkFt2VJC4Up2uwP9B8+xh6xKoPSC9hmQ
bHxkEIHacx3uczISTnUorFvpzBgMqIdgwN/wm56SnNLZ5dmlVQZevg/jXMjYKf1HnEqgGmogZyIz
ahJJJne/JDWOd4fzt41/k3U5NFprv8SJeQw7TUHjx8rzOXKGPsmx1eNFfE6GfUg819v2jN1iMJn5
w87ClbielLTIQczUTtEBK08UmiQD++YJyfbNuWB6n0iDkilhYfOsFnLMvNRgPBZs+fDr3prZHe9G
tEOoCslCxL7no69qO9J0tz1PDL4bOmGQb6OBaz/23ueLNZByOOSNuY6s1Y1l0xVEAIHGfKp1MQY2
9w8Ooem0w9z1MmDvBN6RjlbZn5BO9EDrdTTGCdKSfiH871fA2gDOcXzxz9bfot+zG6PxCVTLXDWi
17fXyYXJu1t8jLyWAtpIR69mSFW8l6ZRpwbraDJnuB5o13b5B6QcI5RNnFuuEUHSuHtgwZ8nykRH
tGbmN4Q50Dn+uIuQfVhyxhrSs0/7sFFhZNFunZR9g/N6xQKqSSVM3vU8CZXk+lE8B5buw7f47Isg
I3sZjPlaUfrZ1w8fZKxn3wZLt8FJtRxkWPlbNUFgDOoh13/11ba/ulIDuLHDfNaSIQFMz+hX2lQy
8d0mYeMHMmbVA9DAr2Pf7Xrjma+Fnoth2Ur3XMuUqYsY+0zDZmFNvHRbXJm1W5DXGOOdN1KCiGg8
w/4FVwtBr6ij4hb46DG/emuE0Mn076z2z16EbEnaMOqsW2fCz33aZntGJQu+HfMcC+4Md6ONcgD/
KFxrAB3fcgbh4oteA5YghlhawY5upkzm5rf1Vf9ux9sOhC9r5DZZ5y5DOgPBieA5g4A2BxcDLDLK
REbLY5d/k9Y08gRdNbo4ndGBMibLXZhfqq6AwrnN7OJt/3f1fuLtnBBNtFXbmNJ8HNcvYVtrIQhE
1KRO5MWwycbIEuVpBAQBtXE/Ts3094CWc1xOzkTdJN9rNAIaETWUGcXDRHAIvcqG9iyQp351nIrq
iNVheGqBgFiKPe9E5laZlY0IaIpMAnK6m82DG+AicszhBkkXt7nMs3vca4LLH93STk1Zsthi0Sc/
eQ5uz0HbZpaDko2+xe95PxU7Cgo1bSh9f+9NDaAuTfLLoP+hJHaJMjTh8ENDOtlPNsLqUKAzqyfk
8JYbr0lY7nFmF8XN5i+IGHqpOH7aK4rSk0aSWDIru6ZBSaztqPXsO6sFsJI5JsJPO3KK2val5pGF
Mk3GluvdbOTcRLvTSvynzI4dYaiZKQ0Yomjtn2bUqcIZ14z0joQ2B0k/Zx1dZU96CWPJoMBh2jKK
vYXWlRnj93XCvmgK1s5Jce+xdhnmKQ1VV+JgSJnv1wMZM0fEXoaHnmkXfLvySZ9V3e+o89SbMMMR
j0XDq5Jru6i8ND3K5W9w/86/pAAovSMorjMa6RMfFMvetkMOVnJ1uUS7RtL2Jv/lxWx+z1ttAA7c
bRPsoMPfO+VLzWDu4/VvXSfMENRuRqoji6pZ5Y5WEgwHjZlfwbV2Ox6UxrEUOQopCCe/l3yt3pFp
HyhPhOqScL9oavURiP4PyUjNcTreoWkw/ScH3vtr0dE9Y6dSWtpM0cIG+Q1dbKKMs7YxcReQtX/J
eCEMmZ2ZTlfvW46QZ/6ueh5rAW+npK+9ai3IqFY8WPBestbW/6xzQ1TeyRijBO9/0DiHGmtRCDmY
ynFxplash76FXd3YGJvZ4JvzgSiMJ88sN+nTl66LRZ9+q81IXLfamYUckfkeNfXxnmpMKSr1sNqO
GqquM3F6g/W4hzc2Bnn+PI3BMn0D1vqoQpZvI9s6noQDXrUX/nIH3j56KgVgc3RZ8WzL9MXeiCHB
iyWzQm7XUSEsLJ5d9wl2QZYnlrKbUDMHIl1e4iaFEu8jY0kdSdER38ZwgTybOD9lv6/ajop9prk5
CRtXSPk+INNkNSK+VIXnKUQuN9XV2a09tccuzQrDcTb8lGmaFbCxTU8H8ComzRC7dbtgKoLgMKhI
jBmfDGCa00zJD5Dj6Vcm/gy7gg+nQLN+FFpFyFnmjOb7bllSnBzdA/K2/LVT0FEg4I0L4b1PO9Sb
gGQeVjJn6Yy2OgV39BP9BmXi/Gj5xXmsErOIjScCMet59fe+kXSyhIQp17dIQXtytFw37qBCAefP
musqRZcdkizCZQwvzx/LyXGvKsjyIMurHGMsystDS6uV+kVLeaI8ytxm3cRAVrE7dRJK8c2waOFY
R+lM9ElMXQyXoIYfn11+VKHUzqK0jvbLKyfZghqcucRQ8dBUxtrDtgN7nsB15IBJqItCVV2NjbMA
P79u174pGS6fIIcw3oF2WB7WBEp+PWXxB1dI+zpV/lI18sk/moTdrICOOGfcYGRKXxOIgn06PXHs
QlNcR9/D30ykVmcCgCTtS2ZX4ElOgYH63zLDMKmX2DZY/hXLh6eCZEsIOIOsGpxZD00GVKgIIWI1
xNl8dcFZbj8/lJkRRM5wjpAGV7p5QDn67XaHfpwlKwNLogFyJUyL+ONvMNpxBjr4i95Lyr054H6V
uZ3bLWJyradPEV6u0u0Cigmm7xx1252N+HuTRTSdlOl4YOY7IC/dHg07TS40k4r+7iyvCw9FtpxZ
czWkTqdZTjc7FEcSVmNupkQvf6kXNjhDswbd93c7f+5HsBKQX81DnD2y57EvSp5SwVDC8SakQWnL
wrnIWJ/6yh4f/wWnvtucnQD/OsIW8FHBadLeXFzgQFHgilc4K2wvM9dUPWrcU/ctCkknCZIQF/Mq
TWNW3+yYg/9OZePBJFpe8lngkiaYCmLw8z2P75Rv8gTs4RSoIX+R0pSMlEFBhFPeS0/WaN2OsX4v
1Q7z29GNMfTxlmN/1Vd05iR7JI3mLLNHsF+3lO54af+EM4Ja96t+sfgtKp12C75BR4WX7VgtLgsL
yuiI+7IoP4p7qKi71un6QvxFJtvbUdj4acXQRZOkM4w/aY7/kpqxLsJ8uNywsKgWw+NJkQdoeOKK
Syr+qXU2G/MyvTWwXxvTysQ/x4H80jtoFsCsxBA8nTKaMP/pgBh1q7pUC0D03+vakETY49ZpGI0q
hVkN3acfHfeB1swuDiAVbO9/s7iUZfuIcJj84BOdd9aoYJB8B0S5IohpAOSB6SHzXMvnLKNw33U9
8x0119qoOMq2buFaUai6Lr9MR8KvTyf7cFf9/2y41mAIs2ttlW08PwdgM1JufjMiQpjO3Hti39O+
vWnJWbwrSISZmOmbLQiLyz+Rw3jLWrE0WblA5crE8Bs4eaA94uxUFuxVx91Zbeor6XZ0xqC223Jl
/OsLIEfly7RtAX290BrpFC8x0qmcmFX6PZs7DVYzs6cXHsOJ2xVnorqiXey6GcqIqnF9VRMexAdU
HoK/2IflG1r7SPY6NtlKqYm0Rh8J1TmjMFOQA02r4te4EdXApexgVi2Q6Shy7N+8HiP0KdXW+MZo
+Z6aJTDre0HeX7ruJzAr3EnUHJSprgZmMCjXb+JIcyYTszucTJwp7EYDHL3H3FaLd0gxdBHQ+NEL
hKFvbn1s83S9EADG72Rc5AYVvxpL37hLPQFI/LKxdtLZ9E1Wa212K1/SOz89Dc5aHC48gjuFmPGc
V6UlqptDQY2wM01Gzye2BZ2f5eAM+eJU6etKSjN9QQiM2PyQP0xYgYAbzyOoXi9zZ2MLCliWusJw
X2gKqqNVsZjtmQK3AraDdEa7Ny1fonVmNso1YPV5tS9TDcwvhvt4RyTF2doc7KensbRCy0SmQu+N
GcSoi4buV2uXnep0KxmHYDp20JqlqEcQCwasT6pvnuVSeRtesUslCde8r9K5NfS8O7ECOEUuSiiI
LAOJfAKBTNcbCeqke/QQZEpcaqEmlJe06xxzyB/+T/O3K5N9CDy0rFW7MhVjIeK7Xo36q0ljc9op
sb5cFVQnkJnrU7Osb3VyoXNPJhto5+r7NksihcR24B0DxkSY8ATpmRrvhGYPfBeGdLfoGvvctRFu
7az4E8Yuo7Fm3fqpGfPG3jQmxz5lA/Fa9IwK7P8octk/dQts4wqhBVWdjOWHsF0Hb8Omvaw8meTU
tNRf7Mrh4HY4ezsGOxdYDHZo85dFCONBvcxPRsOkPcRePix0JI9AoWGZF2REEBuyeiRe/aavw1/z
5nBHVjPjL4kIt7JZvO+01ZdN29gHiWT4yJgkns+rutqQa5SiGBAge/PPNwR1pgnO4V86bay3MvUc
PlZihJ4yn47+421Xvc+tAMtAZg0QyHliwECZ/DcTiAQQoePd8wRh0xtTWl3eu3N2aS3VMMx85SyL
4RdaS5cL+zzDaKMvrpKPi+fkCVavyf6mXkSJLG9Js3c8+XSkSlaJcASEHAU6Y2MRkM4clOeFGJmd
qmEBb/VWumjSxpXsX1x8jFQmDQmQetk+nmsMLGrlbGo0VhMT0QtZnz1tT2fUdIISDebSmnmCK2ti
7hFIgzEjp6jOeeDgSuWOmvETRAtGBYzV12v8C7Gmxz8ZTmP1fxLVZmADQ1xhGDoU/+n2Tgpx+u8N
cLwnRLwPyAJ3+QrSeFwecFrydiow5L/SAAHUcP/ns3ueCzqwyVLB4/nwcSvMN3zDhZCihH6Ybj+7
SAABjOXeLYVr0FJ2XraPoWQrP1+86jwRAO/MauA1nfjBuNBDk6CkPUPWWYFeIJ4tJUSKzcdLXfdB
b8E/UTXwU1KEsB1K8fEl5XSXcBXQdoxLo6X9P+6d12TokuxyljEYGDoTmfOZiK6G0C+RPBt7CBai
wlgSy0fLYzv5t/ua6InHLfEMocidM3ICPJk3kdjPHS3tu8Lfm8Qvpv4tY0i2EyJkVpMRrILwS+jr
+DyqFM8NHzTv7ylnHQmA+XIbGZS325C578GiwNHKQQlyEMeEaFYJIdXeEPPbo0UzF5f4ELZHRlrm
0WduwAGYt63qTRdRRrtWAWKWyO6yvAWOyEO0HVI5rVlx2fRaEENmuMUtjJ0DXHHv72E7IBQunjKa
paYFeNsLhXDzgdC8/nnvg+YO1p1H7JLsJBCQNB+kldQWvkD2EK68Ffni1u3TOcZn2k5xfpNB6nqt
5EVyYZCFf2IE9V3LEzEvt+5idN0n/Dl5AmIT1oJxg3GYptRyUEWkuad98OCA+5CQbGPCBnyUomIw
dg1zCyUUqePsZ5LXOCaaEwGynLE3+CloPIKS0Pseq574HFsC+87GRV291MZ63R8sMdqmRh8o7zGf
QBYMQtrMXrFckTJ1zUBtH7c10NxqpeP1Ncakmxxp7MYoE33mk1/xS0YkdK0LjGAlUmvCPHnm/zJ3
5FQ8zSzxdpe96xNp0ZS7kFREjFlvqrsbaREqBEZL7yJrUIPI8fj0zg+0pnNUvITXdm9q8Ndmdq9b
hdY5e6RiUc5bk31QWAxPAh28l+OqFqxr91HKA8YxBNZllUg1BHrp+5D9vnbCwIp6tGdD/st3QURG
C3MOX+vNRGNJPc5vF6ZVfcdC16D/w3+qPShqXAslyKDyO28lco9S0P1TFaA36FuFZtS6gLcFSiV1
wIr3L9DpgswTjby3HpRCEQKhCYIc3nbxsBEFQxDfxpKnrhr0kzsArawYO+GwniE9nsFWiY0roGv2
U20t0rm/k96QxO/5yZ7Mzr8obVtpkvnZfTp+oFpkQ3aOyF2b0l+wpmz0TC2/Ltbc5f53c5ISwVXB
uTUSwiBaXpAMapNy1L71O7O57oLUfBylHXonyOcKxED4m4xzVo2vK80omnD+x5WC3DeanyifrSIp
3KNfdMeweoBL8lad03P+kUWZDU5z3BQ4K4Ah5QNQOUQVcEKRx1cMvocZaZExnoOiLjr4nQk7MPgz
ZoVW4fnJWvLoWWkF2OERS/7lAjzVm98ZP++5zNLx1teaW8ZF4WwA6cLmmg4yiOtlgpz4zPF8RUxf
oRexYPNVClkvwh9WPBr3CjrBa1Mwil0R9ban3ST0qMJ60qHrgQKUA/lIPNVnkPz6owK0EGFrdRjd
HdFurMRAjxNitnczh+gYai58i0JbtvGoetpE9wMhUpDmVHD7rh7ofO/gwM3YMZSsACFFg6N/mI8N
S5RlH+Hspj+tO62BNwtOgf34IzlJdSebMpaNSDvvMC/YSuFSRL1DOqi3OX8bXGSVTTS+7SviuJLZ
6vzNqcB+afWZ68i7EruHFOSSP/K1d8ymiLWdgb0A3mqt4y9TBoNgAagZKphtMT6ZHdgkjIVpfDUU
xfqCaz+OsbpQ6gry20Gw++02W4amGNLeiN6i8dEg4KbxZ8DFElwaafIsVdhQGtcitDItK+CtMgBq
leGzNZFNhFCZhT4PdyKNOtEhuBiCySiY5HC8g2OAxoZiN4a9c8d6iF65O45lKfhdbKph42iSAeOv
EdZMEGth1+XdC02PbpJ34M2u2PeWu2VgFdaKfdRk4F0gZySCt1H1PSYBhqrgrC8K7/tlS0STwEVQ
31GieflxaHbeO/UvqwJ1en+tjQbsK1ejk6uQNu589DGNtS9McrsBgMCvpvsOqacfhuTjwy1Z9Bei
L1bUELpMl40jajrW61smx1nTdmzAAmHYzjLlySCZwyLbbb2x+89htRBGZP0q9z3zKDKAEIXNZHez
tHrqN7XhvK23Etai0XtqqbwDpUI0gs6JIwzKqb3TZh9ZZknzcHC4dn00zgAFEYnYPAKbnzlLJc33
czW+mQAnjOVajIGbBCUKePBPCD50j/+j2dVDwjtfn8TUHnk3qfhdtOZDosiLn9ITHIH5hpK4ir+X
HgwSTK9PXxWd2wKyZHbElcM1b6AzwF4B/PiuHylF54h+Pa5/k3HaNXxmHLzcRwGY6GIeQxQGVys1
OKTJ/P6yKXsjKiqCsYscdBgl6lHH8GkzaW+fAMAz9jr3UEsvKbnGWxkcy4zAwfsAMNU/Ti26yik2
CzRxJJuDZUH7y5QTdczRffP98QxmOe2gqfVNSOIPnXSM0/vLgkLlcVembpglW6vxZHoIDzN6Nrg7
nIwZxkXcz09UAxkFdkGcvOVh2bVKMNeGU14uKwoDXpRD5c+MW2wsVtCp2RK0HEamHMKW/X/DuNIG
9qf9WNdcMzfAJ+mh7Of5NREiqiaFoXT/W5ZXCP9UJrwg27vg4YxmwzF2N1bICi85z8W3S1MiYIj7
z/qR+Rz+CMH+4L7zZjZXKGzNm96oYwXifkBtNSKUNXdzlMcw2Qxo8XgIAUCIHohdxYJUy5Ed8z43
Iw+nxiQ7QjOjrNx7YaD8HnImBwfSAn/Hc8OyrJnhU06cY1TaY9yVF1OtpZLSWPO9ypDEe68YKYlT
PvGTWvQ6/VBS2jVEjutGTPvURhqulzTPRZrfJijAhyi3UD2J7i8nqq7/gFk/qD+0X3b2HyjX9FTM
tTat05KF0bi1tr+fgy6w5CD53NShqDQhZaQf69GbKZSWklJOBn/QIBf9gmwqzAQj86vi60xO/nuv
3y3EWPDWpihY06JjVWtMmsQkwyIgwm8dPBGiRrZ5wLZj1NXYYhyN2b2nbsoKoZBM2cyiDy5cHqf/
KMbvYyTEqwe2We9qDKa4bmoGdhCmE8kmiQWXV7LYcfJIpEAnpK/J0iTQk2WK7zZCHT2hPzEkV1+C
ex5h+4nMz6B9AVBx6KQxQYXh7x4mTR15NvvANRFf0qxvYUIcAn1Gz5Z11HuxrnzNpE8/TbSTd+G1
kVmekQ/piK54EczvnqVeOwts5oVj42+fqUkStRxS06It4Bpb74PhEJtSZZThK07QK6DIVKEITSqj
LpqR7MzDO7aAgHH00VTcVKcDAT5N6c62S3i8OoPB7TsvU3X+GuSf2IquqEpkUWDGnLa/B5eCyITr
Xtom/P31sTXVulsRt88Ni2sTWIQlg3hSRmcA/u+hmXyyUGyZIE/5KS2s30dzLLJoBJpkoz2i+JGf
mNhh+VwEuSpnFLRrh+JxgQOeqnSz60B/v7b8a6iW+891xeX/pHk+db7iYfuIrw/1EFo33JzwUbDF
4O3Qj1A/G4KJpUWSydMrCNON2dn8MAMPR62t+b86hsk3x9MReYnMrptUyhMZPO7tL1Q/wo4ydc/J
DdWtPo+8x5vG3OfQT4X1K092ivu5wxWlJ4hU4jSGeV2ejYDCnBCLO4puvyUWc6R6Pl3FgWk4JHNu
eJ6slYjU8DcExTnxbn3qmg20Dbe9HAQY9ghH/oNRlvKIn5g6SaziS/8SLbzZ6PkrT9bW43+D2bv1
PvAnPsWZ5zAjI+eAar5jarUPOAfJoGkg+LRe9vmRcYlescemWE3G2bR83rywrz5KGmc8CdGA1dac
cN5JZytxRwYH2/x/RXt1jYT3vdlU7FnOj6n4a0phjkqAgYeDwJO5fVRAOWolS+UgDGGt3Pte8Y3y
h16KAgf4/rsCNF94k8lvuxJ0mtoE8rSIQcnAhznm20SXWP3hfru0Pa8KxBJ13w9XtQYaC5LUcIsX
nNDaiQBINMYfxAuuaGsGvUNyN0TR5k0XUOKWqVBvxvx1UIK8YzxLKhzCGgo4Osscbytz+SGOyh6j
yZ/vaRVVowQceVB50jobFJPXLSKXGkicHJgFViHOaDEveTSF4R/K8/SrP9YENiFmQUXCITe3w+YM
6ZDYK10J2Z7gDlXdCOymZdY+twZ6wMjBgoKt5w6iDqRxQSnB1dyOGp/VfQBQWRnov940xieNxDCG
Qum9X+gqgwydEYlfPTOE/0y7yZyzvDMfWHt1rPAQb60SwtpGWoZMAQ19XWYs20AjeQtf7XKLpWRc
xOlf7psFpByEUkNDr0URVavNAXJYyPCjwqjPaa7HESAJ28BP5c4XHdjUfpRfgyN08WmQgwgDUBTT
6MppnR1mZsDqRdzjMqiu/XDiCkbSbgzQgGD+V3m4sCy6/6yldAnpX+UoxqJ7L4jvwzr3k3nQ/N9O
9d04dkfoB1GGI1jYrbtWj+jgGeinbTBMZYqLXFWp8PAFRfznBt3fNjtRMrZf0fTR+dji6Fchc8Z5
K/PBB8eLM/s0AmzfWPxv1dDNMvafFJG4QUPc8TOIpbHz1qmoxmn9ZbRhMloiWCGzdMUVQ4DqKt0j
VsIonEzGo2egLSNfF6+UC+Q0eheMwU7NLaoC2x4/keHQU/Ogf61qfVrz4e+10rrRpyO6TRNUJfrN
NcSW03yFhf0QyBuYZMOwbm5WCA6ox3qBYhE6ylfHyo+jmbf8TZY7OwsB++Nsb9+q6TqM+XxAotGe
sw/jWlwCF89Iby0mxZDXtpymgenwYhxMnq2EUkgYRyJ+88TDOh20xx2g4Sus+vr72tP+Fyln9jto
iDFUay1wUhYfAU447fzK/IN2evPztu2uWrxpbtlgiWt7CDoRH43LcZfBkZTOZkkpBo+afxMoAlEz
OJxXh4zujRMre7hHZj8pLVssxbkcTTtDVpmAkNO7k+jDyr6vNEM0nRJspUG5rgTgcCFxEBiLV98e
1Lw/jjH8laX97++dJgK/xRICJkoLooxeG0gje4oi7jnN7S4wRVCSdc0BU275esOkeQvg/4ZWmEv4
Su9ttzUcb+On42skhepzPaARKbI3izwrog20rYbr0HYkG76hHVV+iMssw1YFzWadh6k2XA+ouKHu
KazsCCRUulv9jWGkr5sGEPWsHX6TcxqJInfoHbdo5lMScFV3lWlM3hK89+vZgLX6j99e/1oE0TtB
F1rP7QQmBTSr/cZiRSXLHN0kHBIJSzN9T3P8pghbflOjKiIz8z3YDuM4s04hENLz17qkmDNxOGqt
n1zMSYCCy9O9o5HwSgiRxbVAEOSM9WqHpFxbHlUsLA/357ZvNyxnPGhC3OvVr9bnpaz3K0UzmCPR
H6lr2N9hvKJLNKIc0vzD70IPmYY6pt2qCZfqLzj6cs73IDDiP5Y55T9bEhq7tkuQNR1l6ziN/ZPm
UIX25v8vXZmlCYD+PZEWVWXmG7+BcpSxcTq6bVOkqx64ycfrlxEB2tqdEheNMVD6oTa5hTqR1HkP
XQzLyp+iIN0WI3t8WZ0BzimHfZrIn2+LW9C7Y9SU5mF7k0dfFVszhk3KVKbWswiqnKnnDsKj10CV
yEicA362yj7iPw8pVqwtHaGpjrOkbMiE2oaCds3etWhwInyZmR30l+lRoHEPS6HX3LnWdAKJvrWt
yiUK9dtMvcsNDAe+iLmmNJqB+5XeuiCULFvOnqHmwMd+v8+9U5D8TtzztowRW/j+ovjxgMbtPS4+
p5Hm65CR3Nkhl3MEmrXsmodO6HLrs/fhAPLNmsUoXmepbP1na8SYJz0kuRu2ieNKhyxCU/I8JLfI
fhWYfjj2NFli1mVjRQ+QAoMTXRa0+/NjWLndlsCW9MQZ4/3q8H/SHJtMjN9hObuw3yqdfqTVeBv2
O9Io+l9JApRItrKnQZ/FX7bB3GhyF684RnqotTJzDJHTIBE48qv11HHI4uq95bjkvQJp6vjL5wBN
TGPUnwyQf67hgJXGmnP/FjowElq108pNaI1GcBFNqwPvq2kmzYKzRFZahPXcgcYALI/a6HxJw2Wr
3lfFpZxtDk5gDGFw5LWo39v76+QOESJgwO1VbR1jpK8WXimhxFinumwR57PxxaMXCuFgb7LykdDw
PbjT2XKNLsgqj8UZKSPEYnY9emciq+k2jwrAOUcdbGhmbIapqf0yDP5kJxGJoirhB8dwQoanl57D
kb99FZKHu3ZgJf1Vvx+ddOglRd7OMzlix5qvnI0D1fZ7UD5nCQmSzoBFOgznehlg7fABag1IUbgl
/QqibvBekmeiuckX+2UXd5SlYZmew12sNzLqxnKLtiFCQ/YA5ZYdAGi8vcWOem9lbsVws2c0wjtZ
Y0CZdlPRcQYrmINrieUZd/G7J/U8A/n9EuAVWKtVKu9Ck1MLECtAM7ewQVuKoSQ8rVGpWuaUN0bU
yP+5WcotW+uxqhJX5v/yCh2KRYtPUsPJkcoWN05OtnTckyitUTBB2Z07rwLsWeFAKMrV/4NmIp8Q
v3Lw7mvtFQAqnHjrLqLOzj8CrVoAgLcHbJxYLDtmYf1jQWxfTpp5K2hIJmjyEF5NouTVWxwvzYe5
sbIa3/t6QuCKhZNApxmYOT8BWfJdHkFTC+IKhmL63GY/Qp+3hOhfdic/7/XIh0pd2FQ2XcqJKErz
/6n+78+cLWgo6W3cK9xWzo2axrbpnWpWV86eK05xh2mIjKozCPfYobkB4tl2Y46PKu9o0LXWMtXh
IzFBN4dK8GzJtbSGOlla21XD3RdMfk2S3oeeb0n4Vk5s6PTJ32llUq7psm/FMdmnKzwh5tiZXKXe
nOKbU6v/Wb5VIjeqGjuCUCMsZOwwowwBVPbFgBvos0R9r3OU9mjatN7upJLEnzlQxn1yZpSbsmk2
LHJBG7ENbMtDkxPGTD1cbvU4u7ghpDBnBFpeQQK/k9XWwD6HCWgRy37/5RCkaRWz1+oh75Zte35k
xYks5NDJXpWlMjzpf2VHzwvnZbsb3QnNcg6UiLUTK/i/JoShbU58DO2AX36LxXd3J/tsFLLhMe9c
DHkYUoNXmxPBBfz22RsP/7dxI9cCKBB0atxnUaHMSpvw6rGkwsA579iE3z1GFf3wlyqAnUqb2H59
hkJDbo7OHxufXOmunCY55Hcmnq+QjKNVNTlels0qVfsQJwH5r0HryekpX3Q91dyeAyCRHvoXB/s4
Q7tDr9EzgYq5FQlb/Aap9ddnIzUL1yeEgF8JnJyYe6mpKZBLmss57C2gyefe+WwRTneXHVpdAfbT
xKZykInohoEhIaYmAkYjhGwMHh8OblyewaQBLox4eLx1bWYiLZHjLXTgPFNn2FgxFcNk1i+cEYRn
nHnWulznhLZGfINLYNH60kypzo25Hq4exovNex4U1UJTDclJvFE4u5tmc1CAITtXJ9FiLXThj72b
YWtFf9Agdti3rFHKL3hhV9mZHZIIO9LkAaoWDy/OxbfrwIClxjUSze4eyygVyRJ9IJjzJNO/W9E+
SAM9CrHTs+5RJI2xKEisoPLQbyqI9QViKSr1r0k20Gy7q5fJWUOh30k0Hc3AAPRkM8zekml1+EaE
O3hIy8sgOg6TmmWc5GWStveurA9XF4xbEA73LF4nSZAEU6cA737VWzbKyZwE1PRJjFHMY3gYz0gy
k0mf42aXP0zH2hO1DxEy/KNy4BhEdTKr4MC3aVRabzYMDKRhIB8Gj4IUa+OP+BBb2FPXHiasECD9
8wpK+z1LRVncnHbq0UhV1+ppyooMWJpQxUOJbfIJiGa2SQ/5tUYblcFH0+OFsNZ1MEmrmVUalUU9
s5p1Mo9yyETbXM1DBT4A5hV/AuaNLXNN9BocvOB+eygpHd6IMsi9doK9LtrYReUUtu2fAjPZgWjW
QMJZ1HE0bSg3210S0mq6ooIGTH6EiHQFLgWDIgVL+X15skbMcOqpwYTuY6KAOLkgf4JxkcQajkja
kg5yAmPuwhhyx2xxjtOdjY3eXrpvq9AQAMXNhr+YK8H0xh6/30KQ3NfacQrYa/tcgJldk8+8ee5k
ibpOeoTPW1D39ayerZhGMxZ664+4h3nzPe8O3U8Fa4rEFul1Z7sjOFw3nytiRNjGUysQJ4rUpZQR
y8eBoH+pTBEuLb+X5QvU7FQ7LneZMoKRlh6/7q1qHIxaB6RyheHakG3oOlVcpN82tKrNIPf3aYkf
+HPpL6TTFbqO/x+J94tlQ/yB0y8sIlG4KO46nDKn/yH7xfx1xyI4gtzYNAlxe/JFoRADRCjeeeJl
fddaM4jbGic9wCeFfOEywOm/GwfPV7iTRUEaNmgkaKmqP36GV/Try3eUQdm7UP85uHMKKMdTxhdb
l2wJn+KzXCC0+dmOy6LT2mXMk1ahp8ntrBMn18+VsrqcL+YYazfXlewwW5TAJ3sDL9T0natWYRcU
Ed7xEldnQ7FfDIMcelkjg79v7I6MRU5M6Z0FRIWcPZnrUzErRLmxcfFAaoiyoYsv03qDiXRi2YsO
Pm1lEEF07/m+ThgFdOC/RtfpW/LHjgQdXfrgXiGcNoYlEyB1ekpKC60q1E+Kvv8nz0xL1jh1qM0K
WG4zdmJxWpKa3N/HJQi/seKvxz9Z/fCIkv4Sw3glrM9H9YOkqbQjao2bicxgziURIMkD3DeKlPx9
nP6mRSYNukg2AW/GYCrmNOKBjM1Q06I3BbSG6lEcaxlMExtIk4aZD5xhKjoV23jfI/gbccC3Pi56
8u7q7/FXvLA4wVve26Ju4dLQaU1oEjTmnqaHxhEjyFWKnB9GsGI0zRD/PPqOMxj73D+yjMK/xq3K
zKZhyrhmjOWxpPGIHB8SNNd82NtJzO9vxPbxOoI6Umna2notQ2HetNNVAytP/q2R+7KwmVQyTM/h
LalCfwdPqiEqw2WQEU7DDUj4mg/qnSIJ+JWq3gzjQYkGwnNu2towbLzaOtnJPsD/NjNNHF3W2INY
m3aEKaXTnxX1yURhNfZkPc8mQBjAma7yrey5pcAH4K7o7lyE+NQPG9NC9afMsv0wa/qL0gmPz/d6
b4T18EoNHhoP1Pkf6LgiloC2osp8lXJtwZhOr+mkBah+vTcJkTMSNiMwgYRJ0YsLWLT6mc63nscF
3dP625vv3XVBA0DddOAGzw350XUSjhMDQ+/g8pUx0Um4z0pPq+f3HIhujfS7HY4peGjoBaQImMIs
IjzCnhtqWCW25iUEWQXFUSGMPC29AO806mg7I5m9Bc0didtqDtJLtJn6I/LyNtiItXfWi5OBD7/s
IYfW5z9OLVudzl8SQqbJrdMx1UWGO1tAr3py9T1mfIalWo3kp519thLXDNhp33nfmb3v7dISmDmc
o8V7Hx47DjCE1HPkMttfAO0ZRDneedR9swnvymc418pusMwiny93L0pL5scARp5ipUysm3Gjd0bv
ieJW3hLz1Gw+jbOvNEmp8S0GNfcJVtwGpjXugcpGj0n3GiQieowG8gyCyH1mtnGeYVwTJ/mMBqPN
gJJ0Mn5DSilX6SXACE7+p0vRzBivs1i4ngECOb3Vr777kJEwuq+ETuS3TPehehtH1zTVNMPLFbjz
PgvAsv8QSxaaRFt99HqwWNK1qDxmG62llHg2QSnH20YNuBmtnkOYH1h92RbK5f4sZP/NodnW49Zv
/0mrAsPtEFpojK9KF0xCwLshlai4FnVyDXbbTEKLNzzoNyiiBFcZo5XOrtdKYjxogUZXyyJr9kvU
v8yHom6OgHFK4inOLtxZ1nTqL1PsiAAjW9E7UckLwdhmywwHC5iLweJn1yiGgJzbb11FVrrVm4nt
og2cmKUs+xaDWIbZWOzYiN8ZFN+qQ5BoQ7dZgBx9Cqu31ziAGU+TRWDlxM5tFncBl9wRa90v2GWP
pgWO7ZS1/oX00LQjkZyp7AqRiPe9XADHmQVS5eLaqlCH4ZTrQi3jFin0a/TwSWminM77PXSrxVIj
Boy0zT7+sA8ThPWOhPRySKsO35MOFsqWj1Cvu7Bt7dBOYwulMw1Blg9gMa2xWSoSLHkloBCMxFuD
Wiz6unRJQGcXPRpHYMuC3cMsgf8w3vrMYMABj9YQ3rAc5kkNVZ3fz5HcLcABofSU/LsxJpSWVRFC
tMFqjdOaI6XDSMPMug92VGRyE7a8HZkx02/WNqI5uHnvnm+TPKUqhEIDFsGLjAZNezJj9BBNiV4K
ufzfvG3iq8EzowBnNeGpI3dweEqx/qFYoiOuJNYfCbbba+1hM63IMGpLQ5q871HZoRfMZQ9g3WHd
i0cWmQPqGFx/HTdcXZ/UzarUV4xQDh/XGxAOzk/Ne18XEBflsAoac/eA4izxGC9vN3X7rBBfM1Hm
CWeNUt3X/TEPzPgWksr7+8DxxtSf+nC/MOd/CfF4v4RNoRHWJ2YSDioli+Vjd3f5Kvuy5sk5iO1v
N6s2wehAxmjbzd/stNYZ4wcSJS9Ao7Hxp/5jYSo+yjbp+vgzficAtH/F+6bfwUmm7ajivvCiSfhb
Z6f5nwzGMkF2/LD/8WrMQnVHYiMcAudwnb/9tDAi5gsAobvP4ZYwBMCRqRQ7o88kb2sKuFG2+NmC
rnAbnelCI84lCISDEkfT5+qjhfs1gOL600waB35g67KQTSexIQTTt+4k0TVyJ4UKj2C2Bb70/5ib
eiAkadrDt/38/0M/WrUtHZreERd0cj4Cm8Yht130tHtA781+/X136mLgkx745omaC2mItEOBA2CM
Iv9vEoAcBMhVkc4tUO75FYQ+aKJRmMvV4oMWPguxdFLeV8PpfSJFD8O1d6jjDt9DgwS+VAZweTun
JLuZOPE3PBMwkKEfOHnHZ2cfl1E1EsX1eC6djG+K9Eg5igF7QisvfWf+FN/5KGQUR5L5WQAa7C3P
pEic7QbIfrxJFUjzaPqW3TIvUUM7EMpDdmyjIwrKiHPXDx30AiHU9FeokUQkul8cvceopm+SG1xD
is6Wf6UPogWun1lpJQ1Td+mbpwzbf2RxVPke6nCVw+SObrA1fYfgXULGj5Gj+obn9gBiXumSDFQC
CXQJHwVk9IKSJydkoeWBKjeDre7VR9+F16RG87NThX9964zQ9L5iVZCGgqZj5triiCrzah0RxG57
zVkAVsUYTCcBTJXXzEZyWN9fDdZBGK6SN3zz8ZwZMlqSz/V3Fj4eFxNDRG/E1B31O8dnsDS0GJ8q
b9u5bxTQuLsUe0U6pnGWrhRXf9yXtHxG6LMtYfDVYvrTdPQNQfgJbVgRcrsprkVDB25bCZgBoqeZ
wBChdbzMn8adGK3eP66DFQn5GLtykyyDIjPc/r7DZiu4e5DE8ilSIzL83Mao0lHcvLNqHNcfNHcQ
wxfZa2WgGPXMrC378gjieKWAIXecmeq6G/0IZNhg/K2SbdgkF58vbabsByMXHH9qJEB7jAE/xMuY
pXf4UNXKAsJpIz6HP8ZrZHukF6z6bTf0IVmhKxZ8JxNDRjy2q5Dn/xzWPiVIZqS7HKU8WEW5iOvd
ee6ymGpIOKh5/0fSIeAFWsaA8KyBkU+qcC/ZB99c13ArjKqW0Xyb2T7cWvN3eIvSOvQrWHV33TOX
rHNtHTvUAZhgd6bX7r9T3/9pdd20rtksEJvdpQ74/OGI7xACkCPaLOepSTQ9QAXgZvcuc0Rw08Fi
p1TY5QL64U3LA+sz0N8eatFoMmbzv8p++mqG8OPDAWc1/fYCn3Syyai0o9R3EmoyAmJ/r7sXLiAs
q5AwpuWHSFVAlCHzZE1ux6HzviyUVLOtWzrA2qiNOJfRbxV6npi6mhh21uiHJtg7qojuA0E4i92m
SnX/Fpu5sxxFzswgDyWeSXksHRlVG3lTT0K0Tq24rCMN0mwsAVJIlmhT/7FK15FD6RuGCT7JqVO7
+93aIFx/lfabjUDEAE/s3oFf1uHfn7FYlLPFR6lZUaqYJu0VcXLrBj1iIxfvOtqtZE/WggGPch2b
/0FWhLc3s3v/igjEhoYjAU6RjlZHjq8P7m0Jpb7uGIloF4X2AbcDe1BM1iCAD8MS2I0NDLRuZeiG
WsZphaaqiW9NNtm44IdQcJqyQc8A0fWIbHnawvCRp7q7Tk4gR/VLu7jhLoKqvXPGCL2wUrnQ4CjZ
H/lOO+5J79pCYKoBQNZIzVmla/kxKAmjiwyX1cx8PKT7HE19RDYii0O2ASbVaDHhW0Ejxvlekj1a
5n5/yxQ6Db8XgtNv4n/3Vhbe4Gq88lY4LWZCqqXD/VyhMsWIvRHMPk1Mzga2VKaX+Su2AfOrstBb
niZtod84y2V2moAvS40gAO/WSFC8EzGGAAlLW1Oxeyn4TdBXdSkNhyCHnPQ75PV9WEqE/fS5Z30I
sDdp0VB1cs9A2z9y/0N0HAitA/JKqI1LRCmdYa7ue8Q0789bSN5W6igWtWCjCSdskcs+0WO/DFQH
dfmz8B5S/NqFY1/sX/RMO+V//H7Ne57YXmHFhK/FmRI8RIwgUUzop43BVYwQnJBDSsV832ZDxYHi
CSPilPOeM7nddBM0XVo2XyYrj5MA7mIbRv9hRUt+gRTvL/T6QYS4OjULMuHkQsblMf7sbME5XmXk
1oc8GPOzC3KG/9Q5FZ6BrrbifcuvVdGzsst1Jp1KB9QHmsE7eg/pMkwgJ0rCEZC45vIu9yWOTon7
y9OKD8EzRmgChhPAvEZGfo9MPaSFzk/biq4NnU9uCjVVBESa0wC0aG4N+yYIgf5lIRgy2GRNimE6
1u4/29/wWRUwI7BoOy1uIN41XkAAsRKKeSi7cUzkRKPmV5r+el75IEIWZ22SWLVg9VghJ+kEcjKc
qTQcP36EKqXVLIk4lVP0QDch0dAY+TKjS5lYUxKC+Wvk91FkxxJqcYPxNDs9C1NO0rZ4L6rh2X8V
cOVf8XKTtFyX54PknwMSaZOpApkegsuzrcrnv9HAk9Lz/eZa5OsR2mlfjSCZGPS/yhEc9N3Zx3aQ
jXXAJ0G58g/8+brcMptgntJr3BPST8gEZ0+uvM94k59/cICZDIT5+3DPgcHwxJN7OlxhKxf3yDaV
5JipgI2SQMcvMerP2mTBnb+9kKC5M9mC0roxl5WIoO5pqBNG0Vv2uLlwCmudn2DL5bWUTx6zcu40
l6B0eStvC635xyXdk2hlyCr5SrtZsVw6ykdARmYvQ5lhM7zBCaf9s/rVjMn8lWrIrtIYVlKcM3wa
DZ+BMFJSB+D2nnHOnF8ybTjeywU4OWplfNJDPP+Lmvubs7USqMYrmOQWFLERplFd3jByLLEqpu1o
m503wYsuWKJCspV9LaqqABYt07cZHfK5o00nT7Cm3nteYPHLhLqv0xNucpZgCM06gblHpIeupMr5
Xg3McyAJvyFVCnIdNSS4gCgwH+HxGrLIn7OkDheo9d5BuLslSgJLMoLqoAYMUPbwcOzB4hCw7yo7
yQ0m8ixnktUtrjJ32GpGcHW7D6dhiwN2N5PPcCFy3+w90Ccd1b5HIHrqv8J5iy7S/3ANxDi0360p
5O3CuVj8+nWm8omzwGIornfH7/0R6yrMjsY9XMAyygzw+r7GuSXBdXc2nlQjAwIQqEPI6cjWGCFm
O+ae3wuS5nrkL07+jtFtkRNrCjKmgGeAjX0N4+RleTYAMI4HOsT17nPuH3EuYJF8BKBLxqkC+wE6
bYVr7e4jyDiZDBSrRb+bYaFhi1n9vJs74MUjWOSjomNNOeVVWuTaKayuaDhm5lg0FPxAl1xeYn4v
IHtU9yB3vlYwaVQPukVthMkE7mN2274M/H3aS4rva69foYs1p+vxlrnTDc+9h5+B3yjmC3bChZje
KJsTNGdUXaCnFDhZNkV78FysuXUQAQlAvOWHfEgfQ5+d+G3HzCN/7y10SI0oFhU/jIe7mgSS8MGH
yWSbVKba8/iGckidNy9+SmZpHTgPGZA3Owm0DOz+tD2Amt9G3K+sGAB4fDgukhMDGf9ThVFiv0Eq
sSK/jnW8Kt21qp25i8l8Zgs786A3uoYhKlHJOyskhlhMn3Daugqoqtqz3jy39g2+Vo/lyqsmCxdT
5HLEJLc3ZNtSf7fgu1SqCPv51ghT1a4NKOjJZnw7wvaz00RgtS7AmFpo6eOjkP4oQIzJrr5bHqYc
Fu9zLpjMl46S7rCySZqNb+NehdiLPUSae5zDN+EKXF+PCLwaFz94KuZKiY0Nw3HcBFF3dBbYCvkm
rxi3L73BaQT3JSTGPuqr8NN7ayec13cimu4B8pZ6y+hdvNfzeKd/OvNVWzJ4f2mcIV78QJveTmIJ
sUb+7om9i2IQvTv2nMYUYRCHZrU8FZyov1NkRJS0cbqvq959gL3S0GB06q02BvS9ywctxfnChZsK
E5Lk7f1jgKBsDmRjFDkwYBqnlL5iQqylX5Qxs4wvaudeASM+z17aPHlVz5GWwtKeCExLhy1wPhAN
vwQC+ucjAGyQYFsz/qqdOwjabmB8mjsntBRtN8P/pUJoYC4myrN1y337P6BW9Jq1Iks0vGbOq23t
EIqlAOy8w1yy8k4vC69sjauzuPu7RESjZcgtOWC6Gw+5YoD/EglzCNJT6E6QTzJqvP5CX1yq/bee
0o6G0zU/KmAOdqX/+SYwQLra+4l32Krv85BxY1bfk7x17rxP03IksbEGndknhcsoSky8ClRBHwMi
FTR4t97fRg2TV0CTXCHz9dsAvSo78lO3GJ9mUa0+6l+13pOI5aepCXY3E8QS92XdhwJSr5LCgoVk
+DWYP9qqQHTLV4/unLifgyGN4WGKKept4Uaz65rsqnxPZtt9cjXQLWaytTIZcNib3OIwJFi2DIXx
qmcDn2G/92Lk4PMK+3PBWIKdQA/GgvUQR+w6AzfxtrX0cQOCAhrj4o5QmzJe44ijEquO1/VaGRbJ
xQstgRsEknZfwzNmirGY/GG9MeYK6KJkKmkUHATxge1NZPQLN6uMZvwsaicaIiXY7YY/MLh/UpE1
qzMQK26mSoi58sTcCRyIVPk9Do7G1u/NcbVyT3Xa+0BXARPPOG/Qe8MmhA2VpleBFYVaNgGF7hsj
sSkncRw+lvm0PquSYe9WQGiUOlfW63Kb+JSOr6/VynqNknm6qrFFZzZni2X9atkTDi8AVLtZ6czv
XPBRJ+VTdIurB3nX/9vQJomlDA7cdukYIS5twato+sbu9o7BJtmjcA17XKGg5Lm2tlvDm90M0ng9
+dr5PUo22tnWL0jAC/Wogl7rSWXWc/hJ6w6ufKJlk5CDwin0ezeSf+Sv1SfpEb3hI4yTHGoOHw/5
k6CVIfFyvtpX05oeZS1pqVp3Mx1+S4VbJa40iaqZWqZATMWunY7HWNcDeo/dNJkeNmhORYl9oiK7
S8rtKqXpavupFJA9KVi9yAiGOYE5gUI/exggLw//qehs87yYAutJPRYDcrh2KU2bnI2XmlaOnhn6
F9rZr6An8DTUBXeLlF5h9r3/9dU0+4ZTIQCxZd7+bMSHC5Od3aqvm9wvEzTszS/Jh96w+c7q0LrD
HCsfupXjWFPQxZvGdnJMh9y2CGGEuCrOIENx9z0d2iWTNvGu8gora4bzC4q3bpYdx6VskOrhl+Fu
T5MOpirYoYMc4Cp43jXE2MT3MrUASu19flAK5/Igq1Kfn5RqR1uYpgdEnV4eVSY5fmzFEz6E2ORI
bXa3sBTETE0/VbvBin05wvwboxkosJ1xY3Qhjtyhm5z0nw9Mq6/2/E/pLs1ohhb3i9FKJT112ujC
umIH3pVM0x3JI7bhwrCz3jxwaLwtxp2Hcn49Tb73UCi4SbyOS1MyEtd2hQE6CNfFTbl5+Ohwxu7f
0mIRFSc7oCit6jQb3GO9j/nNYf/eQtvzHfYUXw8BjF4oBCsEiwpK+VDYhsUky5DdY8Y9afTCAVK0
o7RWLNliuOheowLsB7ICEOVP53q/4YChV6MkmBa4OtqrxKM5QycgGacmofpC54aaNk16O/KP7yFR
0x2A6q0dEIWOQH2hIZdl3rtdvkEOBE9/TxquEHCGo3QOjOX5U+3nwKuqkbIcfgtsVZVyaJsgcWCB
PG6p6z6gmcCQdUrYo1y3Tihzv6brwstl4dbBpqact8ah8AsvM3cB7EgqEw0O2HoryN0STQfTkBHi
S/XcZa1hcA5jNhBwtUqQ9w12XDB0CKBXbGDAL9TFvZTw8QTTDQ084ZpTeiH4NDvG5lX2Sx90Iytz
zjl5qGHLXJR7gMMkyUgHHDIKW/5pwsmQpkR3Y7hfqriPs69HattgLOj1gRMwPM/O9CfFheXRB7P3
ycSCv/q7DQf1YuQLkwsr7OaRJKEwgJojfcWxmMLsVVYbnJVxNKDJBOZ0VyPiZ5sHqjKJ+P1+F4Ae
721dR77XcbuFuOuiET45/5bepDkiBPQCxeQAyZK8DgaLhZRnqXF/zWS5X58i15fWTIIcXaOyD02X
uKe2D44b2cMXHpXaNLVQ/B6IsPK1cdWeO7QdE8sbCUOzzJ1msQKNydbCxIF2KlQqLIBf9CwVCpPT
dBCa4vKjblvPMQT4wyGdyzySzaUya+8lmBAwBWn8F1R5ETPRQNQ9oVhwYXrkIfS64LdW2vzyn4iW
qOkaBnfsC/Yq8wY1CaHeDvORv0qm9EcXW8R1+pjS4uZb/jdCG4bkYsqtFU5x0EF3nD8n475tYNN/
WjiEBapJgtkZN+sM8bHtPpc0bN8MaCoh0j2PDUEPn+FPBhmvYuNSExlhZ28XkSy6a4a9/i8TMPbk
XQOYOZ+V7P0W85HHX0gYyatHOh7Ct+ekxpSNzX0sC1DwhESP81nwp2wsiufqJCR/WjKhZ+gZUwrP
ATliU1tmnp91QJpALlP6e/QwsvftJQAqovTzoNjTTcs1vAEk+nlIQcXzu90aPA3U0akkC7uXEVV2
+PLEDGUjOyZbPKurOacHEpZnnAOmQxxw2VVkWZrRjHfHrcX1mHie0uJKjVVpB5XswivdRc0RyvBN
WJGvscXZxZbxEwsOBWKK7U8NUG4KYAgGy5+t89Q7TObbdw60/DKHAHJAPceLrRI3TeIns3Oin6gX
QMYzGLSOegdfI118fjzTFqKR1WNZTq0LAC1lP/c/hNXRpy/BVy+xepTaWGLv+DqlI7tlQ4xpIGkL
XpfgHbYcrKQl1wH25x2aRQTH3jf3Az31Rxn+0BeckYtJScGOuzPRmbMmA/aiZy+dBJ5bpyFnv4RI
svwP1DSwlOPltXJktfV/rtZn2r/mAq/39q4kkLn8Lu79VHBygzBOOtaD/fwf4wsLTpgUmh5M3SP4
Kh5tlZrVbUFGZla5MuSQrSpnMJ0kgRSiup+7O5z6E60L14g9bR3grps/EVJphwHxPUKyCEl/oQJX
0Js/4fXcJpJS3oLR+gbxwsrNnCShqQYxTWJES9LmSQf8cf89IPviV3eVU6WQxz/lNV+VO5aZV9tC
MYl2wbriJ5bI/Um/nyFEtzPq4rHqfuQiKA5yiGHXmA+L+erqbXDbjuL1dNdPLOKaeljF5WMpdhx1
/mG6N3WPqjXW7wwI1djo67Yqh7LxBEkFeiePxVmKBdVvOEpR62t9Mw6VVowtTBhWGq5jeuzh/8ZY
H5ZXg+ejJ5YWnyIqqrDtleUMhMq8x3armPO4b1jaTLWeuJXQMngxfuzJVhA9lNS6lCvRS6TyvptT
C+a4zJfT8Ri3T+q3sFe7iP0xSysUADCIYAhf9SMEbiisEwtwi0iER/NTuHAooxPU8zQ3myOBECIw
TOd6+GYY0VQ9X8NYbIpzR113cxoSMvEGgoSsveOS3Ik03dTIZtSczECA1oyc+NmSjzzrzE2mqSFE
2a7KLaLBT4w/FKcj2hJt+b0soZsvNIBiCk5qKFe5sCooxulF8qstQMZBi8wKbsw51b28EEIXosAn
hZPGpUSL/X6Bg6AU/BPFVddELb2GT7GrUGtnc8QdPf4nlfcO7prIXpJYmWirPD3KkFmvYArWvZX1
uzANJ1R5BjwcY662DLkSvK4KuEcY6SfKCBg6MYHqHetcgAfKtupNAujbPE76Gy/tx1k9cKS9h4l5
9tVgeGgqRRoGvkw1+PxCCVmpb/JNF9pzj3Z9bSo0bCOP3WNRtm/i4upsYwMkm4X21iIwyqyQg2Bg
ENwkoWHNVZ8fXJBIeVQUyAeksC4czUlIgJboMlBP+LCDTRBG6WiLReb7Lyflf4THJ1trJCVCcvzc
I06A9dF2+v2bRC/zNZfWgDn5kjXrdAGyM7U108W4MFsk3WaaeD7JEcRVfkFXwHvbANeSPgzZGyv0
ffIQnFSpEnswY7oFRL2jISd9O2I6hL86oMaQPrvNfLPWiTTWz9Zz9RPe7cRmcWXR8dZetbpCJ/i1
OBvIN9YCnrhJOi4lv5zHfOH1RoQ4xN/9c6B1pZCHiDONaSBtARfv73fj4RGe/HfNXJPv/20MYh8Z
TUv2RYfcK0zRsDIWwBBKuEsdMsgM4i4Obn6oTzCzm11cir+Vq7op4nkLMy6EfDnxH2rMkpT2OybS
MDUGpTf6yMcno3nfx/tP46KIkBKzmdqtKlXZBVEuZ/NfprHSK52/zivZMdBi220UHABmYFbRhhPy
YBkGsjpqgO7JEY12Ugt2dblZelJlfw2xUEHND1HoMCq57Srmf6w2hAufQmvC/RBC0DGUcgtKHsri
/QNCL12E9KIu13HJp+8sRlA0J/WkmFh2hhRcyILMSQ3MNHwbEwdVnN2cyovK/GjSqu7Xk74DPa9B
+9Rdlt2TDXZcwQfwj7JozovBLDArAW7VzVmafbDSuLt5NVToEt+YNwvc0ehXDFkefjZk+dIhSpwA
qV6Onr9WYXfqd2AKCYVyZ5yiN8oT3Q+rpPjbtgpccU6qYSb0mVLF0JLYRQuMLcQqGGh1NvVnCMKs
p3q64B0vUOG5TrfuILG8lXL2uJ1sjECqQTUeDb1xMRoVdocsHKOEo2B7GGiV+v8TudVR5VsBpOEE
zwnhmUXTN+GQb67G40Ar0oNs9I2dOgyICOZdse+KRuiXvR5afscz0ASooTQfAqFZuC/9qcn4JaSL
fMqJFq93v5YhXEtulGrvGlhKO9hcp4zbARl88IumhFHeqhSds7RP3cqYT3vA8aNED+dlvKjS+Ope
Gb5WXZ5njjPBEYNOegBaIJDUr6xaLEdUcbyKnrfX5cApmKq8hHDr95f2DQ5rtAp/BRw96AMZIdRO
tGy400b0L9tQtyrqKnxnhh4h+vlVacHQs/HTvJ390m47+ZoHaPtmk+hJgmgwyaSKTC2uHDVGTIMD
llTKzYlTUzxBayKlReCdqvdcwPvC2sjw9V4W6BbcMIUjpRmaxDwXbDMfUNcTEatxkbeluie5Lg2K
fMPECh91WjZucWiET+qM/yQJgBIcGy5rpsY+b4e/rb1L8Hr3k/pxF9VXOM2iHtWxQnAD17RTIW2o
+IbqHI/K5sLuiICLMJ6tRxY6K+Amdsfz7SWjJ2RLpswgjoQIDZM8spCY8G1jg6Y5+CrWZOtTyGr6
JHT9VZtLgPHalmOn/xY+aFhhec2cEYRmGTdHzdf3k5fgejoLzvG1+dmUSAfH+OKDcply60YtZy05
s9Xjtf9U8JHYGTMN1F3mDG3yM8tGfCYqfR4bErCBmxneAzbRb2HtxTcpyJ30ixr1vYCmF7TvZuot
EqHK4b39a18RbLCxFeQhEk4tCkjvjpUaixByc7qBevWzdR/8PU+NBy0YqocDoj6yESBejb2pJUVL
sUCj5pDZzuva3rHpAq/EWiPNxaBZDkbykJDRVahkiMegTbWDN9Opfagig/PSFdtUncj7Qyk2NekO
qFjc310G2oxXU6vyf8OFsvtBWuWK3MSyuP86+fQf8DAjIYwZfNwMtyLgV27KTPFK7e0DYvtG34Lb
sEUlDBwXhocrTrNhQ7RcgjeRHWfLAbSeh6OxPnCBcdlCC4nDCZUAqj8Y3XZXzUvxqLKPQbagXgj8
oPaihJh6m+a26iw2v5RqewGgQKeOi2zE2/3BpVWOA7pMIMkmHGySzfcrocAwt0f2voIM9ENbup3z
otHoA5D9fULyWoD+fgLpXjpCvYAAjwx9I/l/sDOb7VCpiSfnx8tCOzejVjlKQmobqnC7X1UcxCEE
ysjsMsDI4G8UQiDWzV6nLAsW+vC/KoajGzi28KwuWDNPCX/qzwdRfn8INkKbJz8w3K+PFjYGtqeu
qtotOmXcOy0tt82HYTighbxZ52b4TK8fszsC1rP6CP4RH7Rs2lT1RFbquHWjlxFIqO0O+nOynlbu
UxNEC1Sn2Iiw+DL8IHz23KKJ2ExMjbiebNtp7oTHY7AjMBJHYJwWNd0mM6crO9AZ0aFXNXfdS1pf
XVniwK7NVCGF8UFB1vc+TEKIkmDkdhE2VKZCsIQGsGoVUmIoCaAw734HJWVkvNXwBVPc+cV/M5iN
shm8dTtV/Nz44vqqRLfaGUueBnwO/y9Sbd43Nz9btVfYqTFDsBqq9HHllM2+n4LkGG5rjJ04Q9Gq
GYPQdhKGV552wQJQfoOPu52J9y4uNGmmQGti5kgVmiAkLGSw/TJKTTxUQ+7Sg4yFVoYi32NEG2a7
ObrM9UsPDEckyCOFB036kFrlKUrB0fiLyTKZ21swUxjRrz/GVk5WwNoN2duBW4dy98Dt3ptCXc7d
r8i4Yenm7dqCRvsI8tLkI+ccCH9Hps2AAmGvHa/NYAOKxZ6+G2CoZkRWvTPTCOlmij2QURj2B5k+
xMH4WMphmR/T/bnRXrdBOhXXWcg2ZqH0DYNANdT73ElMAgX4JFqHIcgZwGh/YU7S2UhMgLC0PZ/g
GC2DwUjm4vlKmMbYQMgc9XWSHSZXY3Rgz6Diwe8cAmK1RS4BUJS4Hl4nSaMdoTbPiAFxs+f1fjmM
k5aupbE90RE0j0dNSuREDBl/GnLydRunqVMEko193kWWdBlKcrT5PKzYWjRAiM6CRcJnC27PLTHm
UttKoI8uUafKPNstJ27J09z8X1va8BUfd7tvQkcY0onUF1FsgLv3d/bOyn090QAMlEcjdBK5k+/a
g/KNDZ4elm9dVTkNR28fO0GnFG9YJ+FlfDxOEEMAw5UVtPre28gf9vqYAM17zTZcLQdRvl/vpqCK
b4PEHWC9cKkc1nAY9Yage9Cx05GURYDAWzcamnQaPNRruBovxaw18UHloLgHIVSPVUNolcTpfPIq
eDeLtxSjOEr0mVTSnxFkEU4dALvKvRcCvZhTqG8bCU5yOxPZTbjyK8BtPgv6qW0+bxquHEgEtIFN
NUPG3/gcyoy6KqfSpLLbU2I9PWGLZr93BPRSJM9eHjCezmBoF4fee5TY4VWfqZ7hh/uLgI8A4PPp
E5wLz0a2w+Gr7GOF3L2OYa/O4H+m3CCyfLr2ZRu3YV/521hTAzFLOYOeZDq/AFZybF2T6ezetEy8
wpkA1WBXn9hUEoFOm8SctdTUjS9en3ouS/CH6uheIzBTnHxCELbHbB+2nHnS8OL9kHVKjUzsTayK
TUNmRrD6Se0RyuiHquAas6BpwV4r2oLyk75OQXxosqACPzqSJBXkZILf4/kocpHg+0J9S38nOKpf
tqcO+0i5Sup7zKnPMTcJnku6O6jbj8ouOzWZ1AF9AdS3tinLPlVcqmLIQ4AdmE2DNHpJ9zVXFOJv
lPHWQ7pbfudZwN1o6tXrfgcOzhqLJu9GyZ/lrxS2WX2yv7v35HrVBx1n0BGI/uwai5ONBThJttNn
xYqsW21IE3IWn0fQZD6fy/a45ZYRbDyjcLnvrhg7oq2JO3GzkvVUxTtRPZxS0hrueQtPlNiK2Qdr
LUUWAV75sqa+pBwAWeVLcDcVqqXwpvJEYHD5H1cjuJJ+PTOdZes5UOjP3e+OM5pKah1XzA0t2CCb
1/n4SoKot+rBq+XERrCpFMe307TLi6PEDjd0raf2hTSgcBLpVrj0KnixRCehuVSbtDWuoHzm9wfB
e47G2HZIok/e0oxI+qyIQODFUWia8Dw7qUmAJbMyu+cPD/Wa25DYKdVlh9v8LR5wFfvZG4Lc7x5K
Hf3smu32DWoMKcxaqXXbzSHltkusXIqkq7NRjEuEhGJZdC0MFN4no0K0lFX9PF4D9Ju2tg9hD94J
GJV4czz40DVTx+DbqngfKkPymFrXJT1lMK03pnXKyQn8aefqt8/dq0uYkZQqNZiv5JSHlqhfLKuH
uoR8HQ7594D/nBOna4B68XctK7mF3p+C1w1M0mMh3MZMj8roVKXNmObYck9fAZWItXxpoYWHjNa2
E0hGTXE9ycMV+TCBVIIA7tBpF35+NxaIBfVz+AAL8oa2wORHGznYw6OT2WO5ssw5LkpbdUcE1E4m
VA4gw+wE4ateHSIClBwMxOJj0sYN27Ci9QiQIyjoVrvl4oyj9OTGzsLBIL91P6Z41g1Ct+/MCWZl
BAxGHAEzTkJokTofrOheyI4mifAPG4T4t745cLzvGenkLauE937eS+KmKMH+noAwmj+CKcLSAWkq
7jYAuFoTbnQOIa5BOb9rdnF3SdwFTRVMMTE5ReTEheZliPyzK8BKkzkfWwd5u30nfRzrdjdAntWp
v5z51H2dgeNhtvS1O2YHNIRAXRpbinzVbWtLV6frwSkmgk7sOsjIlDaRYGE3aSWdfMkmmBbmDy83
kqFaIJPnP4F3P7iFVx6S1riJxvIBppNJMMFbhDm1jEyIdkKR2kWqe9YNJkZA37EdLsanGjqh2Ywy
ThVvxfAIg9qgHqdYRZIuvyaTyFBtLYLmlat3PxkNfW1Fc0WQnFI61Xe3KBqUTgFsWMxBPimoTh/r
mFlsQyXIMralpJJLD5z3Px8G9+tG1H5nrmsuJIBqcNVm6uWxRoyRzLo9hmDtt3mIIonPhExbJv5B
5Z4gKm6P00JGhYFsHkqFS5xPV0rQxdA75M4c/aQvYDzw0gyqgCe0RCIWVKHAvmxMyIARhBc5qzN8
5cqblhqqxxdUr3OSC72lVte/SNezFJRdBPc8ekCarWxL9eJIRffoWvik4jMjRLE9SFOpxwUat4DV
Z0X4UlZoLjhmZ889kW3nQfYZerMn5KUxgIho7EdVtNRJk9A4uBKBP6Zx7DigssTSJZOYDf8Mkx3I
glO8JQd4ceGgyhiEdfxSTbXsP1sug7O/2OtNwj+pf1V3Xjag3g+rFpq5KiR3qmSpKOx9LT0iEwcA
Qilmje2X8oG1/deVYXtJ9xVEgrRZv9snx7juSarD+bZljfwoB0qzxqfWmQW25TjqbZx7/ztTpVuT
l0CbcMHdMiqT84tU5yyGtim663aJSLipoQaC26p3vcxKyQ0/+/cxWNEQQsYhIzHJbw8EgxfXkgco
eKK4WQyRyekujGK0N51jOLmOXqYi7zspj16H/AGOG6Nu1JKwtj1+bla1chOe82V7jMMw9EdNsmms
9TmWGWJOTLppNuU0JpgTX/6AqCseVndYhgrJoXKlPDdmpf51sUKYhak8kEH2POcFGqy54wH81NeV
oyA+WXHd3Ugqu73hH5IuUVJV9sCJBhuVQTRH2fnf42jvcwIaHve2hREbcjR9guMs3fvs+XXKOJ8i
HpvhGkrvLFeUq8Z66bKqE04bOFoHV51tbmhw39/fv1zLTHtWztwzo+pNR1uuBXNWiUNSvArLbo+m
N2ZQ3NH5viFYWBQkThzienD0qXIjERf2VGQXhrCSBJZLF6o4NiWpxVUE26JeJXOUL9PnKXhsnp8f
VjRxQ84Vi4cMjv5negCTUn0tYaD2NCKTLoVsQLkDcSeZ9cGdkWfflf0SUoHXaln3gv6kc6pBkwJl
iehGY40t31nkqrbTKs+0Wdf52h3jPJOlHt0dW4aw4aWK095dHimo/Q8LUze89lymhLxPF+G+2n+8
un+/iZmH8bUrNnruwr/LfXLNVNf7xkwI8f/lvdjPMGD/ygWcQYlcA71h02UkQ2D9SDxXT/54+dOw
sd0BYBDHLwtlAfg5zpP3I3Mhw05ekrS8gdF0mArti5RLzfGN0lZIkvLOLhwKcnVFhJA6lOB0cxzM
MbBn9lhrjfDSZxRhbnZOB8VZN4d2An6nsIM3h7qqzZbDI7GYa4/Mdwdz4YXqkDH0AEpLABenEBf+
e5zyyPkboLRnodNDkRHOV31ygbcrOEzT78t9FRzvhjFdjVVuRiRIWYAyKotOMLmIaSLvklR7Xki0
43mLg5z+e8i8CvPbOxrJVjPW0ncgrAAzy75mIe0fasA6gwOex55xzf/kjxBoKpSZbRE0Gn9dGsGr
0LODtdBnxBVcsM6oxvAUSesTt9ad4BlPQobgfOY36Rv56aI9JYRwrTQtamhrAy3VN6Nug98N3Co9
2Y0z8YNGLuc6dBDcobQVGw/7aTQMhCsFziVwFDhwepXXWakBuQV7y/g/RZP6IuYtC7IVDOGSWrO3
eFmut5swT3Y3Fv9nYuCNGd6A7q4p+5U7GLMLM7bV3xK81LnV2PJUD6sOrUlFlYLslMXUowv21Gqz
kjjO2GNKvbkeSRB+kO5A3FU5Z2iujbZ7yqvHlpmemFXJSuEJsJaivhrirWskyW/e80dIlN7KHWMv
FE5ZOim42Ld5YNDLGuTGrdpEw49Brvh7vcG199zW9IfA1Lk2dgKxVrCikt2r0BNQDXa9Lt/R71kX
8kAWnnXAI1NWTqBdX0fUVzEBRn+47w333Bbdf1LUlYWS5b+FUaK+RHoMP8NeXjw90wUeaMnZpeM3
jmzduKvpWVvRdqvHgIb+kYGcAjc6QGyVUPMEDrNaBvVTTiLlIYrU++amJgWO/fvZU+73f0qSFBfk
5Km0yXEZ9TU3+5cVdXP8oH8u7N4dO8UgrjsxMk+T3/sxIBYS3hQijhy/VbmTqOyASbOY/ctqxjNR
X1lla2vF7WXEasLLDOm17ngspNrplEWvkeReiFmLp40bGCEGLggpb364dYOvLC2/L/Q+4JghQgSH
3jQ7s+JKybHAcyENRWk/oz2j7JzP9l3wygRL1UCjoXo1eybbfY5mT72MlZIjg3oG/mZc26AsRZ8M
CYgHDFS9aVDAEN7YqhNV1/bK9h3PdwBU/dMsCEltOcflHGlJrTQoRHsPo4oYAezhEL3nbFobi8Qw
ip7ZoQwOzzzwKlcP/Crec6Bd0Hu2onZra5PxBAuKtxTCi9NcQ92UW0w5nG/MQM7Hw26yx/tTnKWz
RaMTgUXW++Lyk4u5mX1V0ayotkNyS+zcY0apVBfNx0ruUmNEdfiGUgHu8jvegb1g5lMDCz8rPaeD
U667GffgrTxOz9kOrfu4DQ3gWXGCIXt66JID1zw93yQ87/bNeGhZA26+mKnQjjirnQ8OGoXsmxC6
09Ot6TmiSdIEuLWOIlXhFtJ50zxqBkIAaZSo3gSb54ZTbyZo8Izb8JWrupuyuAq7w9TbIDEVmkJP
blWLeWQY9pJqO8VmwzA1uUwzhyAlt6/dCi1BznWKXSjGB7K1nlJRtB7hICe8gS1tTsW22Te6y3f3
syhm+TstUZDX8ghNtZ3CuQ/APYEKhyEcfKX9dfbgjelrovm0Ekzcad+e0eX2u++TjmyVqj01lLD+
HW1icDF4fvOY6jQJDeFzsilzKDq6dQLYDFPUCYyM5loBeTjmSBeO2CgRkpWhT8pRKwJFEBfoD3aZ
GNwin1vRh4WKj8Ubs29b6HR7xtWEy4lrznku3vjgG2o8jCTiAxDye2pAOzBd4k/pb+9Q089NfUMi
tDcKvv+sbHt3b6hzrAlEak1wxem95SARkqaTaOEOmYUe/3nPB+BPgCjmT0wC8AAO5PbyGWndCd3P
T0mCyES9H4OGcYm0PzWw0SqDXuaZG1B8wtYVFVgxp6Uhd0HlUWZ1oo9lQzq15DJy45RvCdTAC3O7
rgIS/Kxgf1Jz9LJHNdilg8O5Q4fFIOb/gttN376+Mm7YsJz18R18gqAKPgkvrSMb5n8lRsQYoZVT
RIM/7c26+UpGyqJiAM+BFpkMI2VPCteuQzD4JLQwXr+O2RYDshKQL5t8UEpTF45vQL6QJS4pxF6D
JPytvisvw9Dtf9iVu4wuAiW7YQ8+BVhmnff6KqWsOtlvpd9DqjdWLXehtCcu3m01UcOf2z/3Nlgd
FMP6/vrhc6s23//LVbmqOY/zrBl45DbEPPWudD0PKBVKeSuC2xuRbJGhUexF1rhX8uNIG2w8uUPT
DadYO8AEIagaXqZ6ccjf5aJVJ4Wms9q6GjGmLIypKqwe7aigxboDdH8TAn7R7kWaHE9M2u3RErg7
E4/jr3fYOzTbjv25yE2q28L0JY9hkw62ANQr9aULcCWTEbVwSSFi43s1yPqXhiE3QKIGa1R92r5b
vfaxeWC2tVkaRJRkBKN6is7Zt81kDiGivfTCewhUrCFNHYw0wV8pQHy+90AvxH6Q6yOndT/cTZZW
Ie7mNxzKo5BGoh4zLvHYO87oIlBGVu56rQH3XHJ5z8w0Fyf9ihZjBMZFt1tCoy2dZYAxdt6mLAz2
EbWgaLKGja9n/QsKeyVE7zDuqGhh6ti2XAmQz+0LqOphmAFyuwMGxF/yiANpAJ6pSKVa97dUkJkS
cobEsV7IPx5sSuzpi6OwN/G8YdPBNzWYNbQmoh1LHo0hRznILUuLsawS9PTCMQwtTHiuP+9CLEl6
cvi32mdqMdIaB1CnyPUSCHmZ9Ph9JXaqgpJYeHFiu3g0bpL/xX7lPK55olSZMlesroxbvsbV2OlU
b+z8+e4q78d1pdMfR8ZuBzWeb9mCwfQ1UtLQgZv7M9Q8xumcrO0t/lW05BVEoW1+6HTrJvu+nSRe
eqbLiL8aoQsFi5VSSnMFcQFPlq2PjehfQ298xX7WmRqtcTIOpTh9Y+mIsS3Yd4zda/zRKUuNzrDi
eKDD4v5EeTI1lqBWXXhdsXsFMXDX5AxDS4IF6KzK2Y8vmvJZgEJhhpD7mHrR43jziM50GfgvbWaL
WcuyRMuED/i4ffYKo9pk79AGcTUeq07ZDfPfIFSw4uCmiP34vX6F0Wk8R4jD+5J+L2MCYE46JvwG
tsUZojd90He1AZTpmj0yNuA5CMFY7GGj7/GWN3oGecW7vBfMAN9dG1bQfSfmxRl+xv21Ewn9p9W+
pTRWzex1c8yPwwRIB542RoGX9Q/Rs7cZFKUflYDnhOpc3qzClmm5liiTPGSJpdw0TqWL09DiLpXi
BFH3jrWWf6dRxuhiMI+5dP+8cYm0sdVcz6zj31IEQPdpf53KQf2bCK6Kh56qv5blKKk9VSGBuQij
OeNjkQQG8lowhQucUmFj+RADgUx9kvvUC1t8DTuTWKl9lkqJ0I+KlxgmH2jtw5h06jJ3FsBUcMgu
SHoOyBRvQGrgBnLkDCFQo88yJVx3pcNpZ92I91pXBNTgXYqcGtP5/OG4o4DeVhB0ifFDm6D7kEaq
fm2kIEreobmPfhFD6prkZ4sT5MdGC6Y480uxjeP3poFLGGIwjQhKsgmPhyxs6ZjiP27BJXIacRYr
c/pqfNm9iydolw6ilqyq1YjULkwA3uROfc7QFODWojEAwCu3I9lp7Xp2SMHSfA8Ie2dr3PhWmWd+
dGf5NOSzKRRK4/Iw49fPOXfQfx4SCiNmgocCD2SnPr7pJg5ASU/1YW+8JE+aCKapyrM7Y4d4+v4d
LLolwlbyxXtC+dZ02HYhi7hvqf9NZm80xuvAg//Y1aTQgzMY4GruKd/qXo0OFnHO01v0CjOJjkEy
d5ql9tusc25xrbmuvBhSkwOwf7bfLoUXcvHWy1/BMxQBZ/wLBF2SmchZmwNQW1nuLUbJZHcNZ1NF
05ZnTBw1DbRdpWh6sf7VrYJacoMO7IwjuQDjYwX7c+wVEL/OxsQawM8bJQUsKP4i6hzjfWH3tUiX
RBrd87yVWMp+WGPBpaH6LXJ1tHVF7f+h5ZB6XjTENZDhQU/t5If1vTv2g1f+myC231MtoGYdL84E
L/IQsACSGuPSaYeTk6je+2ms5BXm/H4RMn5N0sA3fcX+MkU3dUEBvPTaAhpzk8BWHfXwEJi4Cx6j
IL4pSWJapMjr5ngUy0lwAD/uOp9N9tbx84g68IStgc616Lx90Xu6rAngxNiNJ1fBoYsv0Aq0Ugmf
+gx9mq/DqfNw1VmVpPInoSUVH5Ip9SMQWKsFlC+BEvi9sBvxj7aGtJcyALe6aRcH/nWrNgNX30hA
5fwJefX5cjwEtpGkTv6DIIQiO09NENigVg0wF3sfLl+1JTSsm1gWxa4rYSL4swZuARxHcciJMhHp
umTz2mQmQbBHtGq1LhnhkKgmVlLmvtogBtULsRlT6DdsJNJm/ytjzP+Xdt4lvXaCGTqS2fiC+WLJ
FnqLeiySJls12dykg9P/T761QuzMkm+36vIsHzDQF0FIO/tCuVYnQgiL3I9MClBJ7OcOawtY53Gi
QhKJy8t4Vj9b4b0ML/2cYBn56bdBNynR8AZK8MH4EmPnKGyQzQYshXdAEIzBtB6Op9m9Z98VB/Kv
QeWPqMzc98geD6//a/haE9UAeFlM57jHxw0s6NdR0/TngWQfyikR97gwfnxrv/bBuUk8LcQetOMG
YNWz2R9bSOVNSKumqzjvU8jNQUS4q/arGoE5yXU2DaNRiI881Mv23cyZkf65LWDLNBebKdHqGPri
hk2UnyhNbDpYQ2yqvSyCBayFS6ND33XSw7Vt71vfxZHRmFEZFt/f8z2VMUbw8ZVPc/S5YaZHSeYo
wmXAPpMK54S+B5HtxblygGQ766YuxjMZl4qVCPdcV0z8s8cn5/IugB1jcSoEIXcs7NZW5AujSFit
bPFzb2EwzhcyWvyImhS3czE83s/nV/G1kphjMX1lRN/cnA6oZrT23aqNbDjn9DlzJppu62Pj/NJw
dDbQOj+SezJEZaA1p+/uzRcbamI6C5d/OkhkKqyluLgxJNWqeJ35pRABMw6yaBpn+Z6HJ5wTCk1H
XwlSAx49qfAaeh7zFHzj7NRNUdzRrmU7SB0NvvexTIo6RdpL9B2lY9Ei3SDkOHVeHBrb3DA6HueC
Cf9gDJ24UZm2H9k2Nvm/e2ByzRj2dnoXhaIy1eqBPPpEttY6wgi4SQYX34FuA7hDDlE1DiQPsPtE
yKwK6lJRzBu4f4/zyyO/daNnnZLZljuW3rIlZJGAskhhIUNuqIHcopKrTtt7peWEBebHUiBawHxO
KWJ1Qe8BWYJ4meCOI6FyK13AVbbfOWsik4MIQJhii5kJ0UbWMELpu6NLWJd1XXZ0rb6TZSf7ZQyS
QAN28bm8ItnDzQqxH385FYjHBYpHzq/t2MInvaFgH8A3chnDgddfpTmYlXp6lx+xDsslwD1/s8DY
ne+TE4n9lESrfSL8ECMu5sGQbdQ0wRSjb+lKIDaD6YlXNSRbEIMq7JTZf5vVnsaao4DDg9hWkZwq
oND52K3v1iBeappshJKGSBHX7lwwoSBUYohQwNAaWSrDHfAeGp1NNu3sbwHxR8RC+ClY8P1vgAEx
sFwY9FcbRn3bWDb5JjhfCdS/69XwCRXp4OUJwWlgnCpN5p+i611E7Ei72Mj+Ntwd2QumlCbXSn50
DbLLYxh2ryWLWA4qp0FQWsKgpbIEx/WPhfaPYHjTerccXS4E+5lITRSdsC4jKyy9jzNDVlyEAS0S
JM2ljxd3yhq0d1e1yEeba0lWPlJCH5k6zJeuSB2lVBLobbSx4XngchlbkBBy65O377KQhFRt7a56
j3LjE9ghlhyMnFW7Z3MYryIfPDMO7yFPfjTBUqIXCPgo5ObiG7+m6YK6a6FcSTLEYMKdgz+eQRNH
XU6bwkSIlXbEsKbqKNjzh6hO+8YL26JuQEWqqcUUnNff7aHM/QqnSaY9ZFPGeumGtwJFQd5kkFZ7
ygpIBIZ/mbhoPnXZOn9ewk32H5j1aparu+ukYHSgvn+RLSnF3YVHtsvioDaHc8fDsm+ChtldcoAZ
2zpELh1ZfBDCmgPra9HHRj22rLhXUM48TzfgY16C0ryRz4Nb8KpF/SSMfF/tZigIq26D0ObEXwWm
WXRwncV15VJT9G8S16gaF0/6tDiBbAoaYAeTSBXvuI/x5RB9u0DeuYusfh1LV4rT4VxuebicSMTL
5JwBH+44KYXp4629XBK+ZdOm3BSkcMAtyhcdWkOvIK9bPKh7QtGWbnGqnj3oURHM2OXpA8ks6rXc
qMHADeYV8E/TQK4LcuwQAEF0VEz3odjBf3fAbqLyvPDDXMNeNzyK41Q3Fx3zq9DlwETOVWwY2KhE
qi8R3DrTjoc/ShmuFG5br/Kh4hubEz7Xmf1ocvPPYowSdPtuBHsy/7FMbzNxihCAOOo5puD8wF15
QgcbvGFrCNYc5g3pGao+OWTwPe2XZVVmbdoDJtB9aSvPc1kqu6br6awePcGTqHqyl31IApe3Tf53
6D1HAwZWUVFRpN81pbjkOxJg1/mmHvIBWSlspIyo1/sn+MV3IeJFUPLK2nF5MFvqW+TW2+1Wcctw
Ix+UFWgZFKi/imfEgRRD7cUQxFEh+oETlkekee7yYzsRanPtE+VzQSTimbF2uwva7y3scM5j5rQK
7GEtcqJRWeqycM2bSw7XgCD3L5TQ+ZFE3oIAmxAy3KpqYgHi2YmwsWDBh/1pzVNEYxyf/Lt0nbwr
NKFyhDe+e6kR0Q6U2Q6Toxp+Py00XpIFGKEqQ1IQTsKFdony5SiH2p1jxDvfuUAkFeWSDkiDPxXR
QnzN4s4lHOJHQ9qn7hkENU/CvxZ326/Oj02IF3r5hhnRRKUAKwdFUTdcG/RCR15P0eI2IViNWsD9
y8mqBqCNyBNBvOO6sHoFyfD/3VSpIrUiVt26C/yiBZYj6uTNB9LSTTw+iNGxS87gP15MJbM5tkNT
OXMyUn4ji20mQ5j4hBJLPWS0yXzudwYVE4Z04o/wtKiFSzT2DCIJN3CeFelO3lIUBsJblpJXI7vY
2tiSaNmdJ5rYlEKsRfhfJ5nxzFQyqyFVKgdOmBsS8Jxzc6KiZvMwrNSHhsjBKjCGj1+ZC1WM+CBd
JH2vxVNGblWKP6XDOffeWFMO5MvUKxA7qLl4pA7bQcDWwPY/mTBT4nmAOgpITZ2cYG1wZIjX7d7n
fRIMDx7VXwfO43t4UVgLDFLWR6z9Cj3VE15MwyRbeg4LXFSnhwgORrsE7CaPCk5MD1H/xbWxFi6Q
tCXgOWsHNEPB0MZ6DdDzu/WRPdaNfTA3ZFJcG1svdY+s6r63cCQ2iBFxAe8KKVt4+FzCveobQIyO
lVQeVBYKltMCQ8NOH4TOo9Sq6Z8KA6UV0vYWigyMqQAAkUrXBWLYJb0aawS9672pYNpxcsvuBnZh
6Xhzj56aoaUBLQIvQskHLn/W2fpY4W3/AqKY3ue1OZcbktr92hZIifMX+H+t8yDohjJ68eZ1IlDJ
X9wwn+oV0d4RinfpF49jz5JvLDyMpIxLR6xmMpcRmKgAbTh0Y6fMxH7zNuBHiQIZ+Omx49RX/PNr
u7Uw8EhgOmQrn/N8hmQCziyL+UQFRVHEG5Y7VZvV/iHxW0oyeTfECfhMlt7ezOUIXTbmtCOL5g7e
oDnz8hCP+yyJbSrEWTwGSDrsQMU1Mw3qcKpfyIJ52Uw2FyZdWFao5iUi2MEQAxcwNiQsAfPWYl+S
24l501JEibYbezDTjgMziZ0yvwG0RhvbDAJ1GO+W3UWnRp5vQNvmiiyrF46I8hPsq32SYo6/sfNc
MOTE4Hvhg+GRH5sd+8xANtMh0FFU10Vg8HE+J2F/wFBJkKeZJQvsyVW4iXDQ8cyY+QnzlKFkfqJG
cjZ/L5cLZ34KX2N9zbTB7i93ZXx9h6YvTFv0BtJQlqAMf9Zhll2OqlMQBD4e8vQ8UtG7P0Cuihdo
ALQaFCaO0n/1Kfo/RjmzeTsqi8NnEWtB4sXk4A9odsiTrAhY/hObop+phSPfiJIndQE/mp5V5ln2
Vd11W3CAk3T+lRQ2boeo0UAYflwJsHxIwnaSVUqy75BTG5Y67b/IPFVPiU/tEiWEjZaSQeg/jMkW
5rota3HM25KR/ZAB3U4s8+4sCvw5ErhGd+RVhT9djZ1yP66JBnv8tqIiYs7vgSJFjT735uktuXJT
lQym2l+aIQb0sjnGT+QvPvRc2T3JCm6LFGx9VeCSiHvQbmdVkKuJTYc/ABdU+kf4I6SSYXf7vqAG
rJZBa8HCqt2SB26niOEL15CUZa+FXEwyyEUPlJQTrSmaiNPAP+Mlxa/+Dy3lPyNccMaofVp7dqOi
OTFnw7Dv3RW9AxOtAfCGe9XfOBagqurqeNYajN+3+ygXld8156HIjpGZTHzCyTqpuE2Afx7eNr2L
kF2ly52QWEpQyKWJ7G9V23dhdwy5++WkRaWeRNcTnG5JuDTWGtWOOJ2xUZqavd9xP906TF2d0Pg9
dg21iuB5FRvxZXpgtHNmV3SOHPOEU2KA0ku4zVQOkSIz41NQsEU0yqMf4Z6Nt+tu3Ff7NqmmFBxC
BcKHn4o62W8z/zXAWXAy7yU85p9eR1W03YGnpiwT1LKgn4rFDLAkmQn+opwmcuKxPW9vvBB21RBu
U3aCTAOjpgI6B4fHIgit/oxbTJguOWRmnN7u2zTM63vXnRNvh3fo+7aGR4Tz2v2gku1Sqb1nuv3E
UMDqga6jBaw++F6tDdwsY+9nk2GHeDvvZo6p7QCLZC2evG/xz2liFQ4W8hfMQCKQkAa5cXxjWacB
fKa3HzAqGx6y2A3QYr6aze9e8+HcuRg/4Cw55m/ttb11v0taIzvmV1il8FRL44aof+OEk3dCU0yL
W0oiOaXfB1R/u/7BQq4GO2Ss+y2rIftHULDMpLdBufe5jjSP54LW9d7XjdmM35DgMhbulolJTz6e
yucM/e9L5agOqU93U51Per4y6WQjfQTVhcfuUSJ1j7L1RSzngL+6OQU4FqIFD7etPNyMqjyFeedl
O24AEsz5YFU9FqnP1Uxf8UK7500wtzyMCY82IITSjVDlK0RgRD+obgozLOgzZ9UKM2P6p4MWHznN
lLnI7ohtnW1+yFHH8S1/9gMnxEa8I21gKopq7CSMDzDb0PcLh2RvtUQXDF76xgJyiT2HrHZM9j6W
biD7vfzqACfgyWRwJ5hrHAOJ7QEz5mC1eZyQK7QyOOoEeo1fI9DfO6qXZ3zulpaTL2A/4/ENFW5E
Tu97h1EpSf/TsRf7syi879IZ3aVfZhhDvQREUe5hdoth13s4VXv5M2Tan0Hw3moHIU2eaDi18t7+
TckolqS4CkLmuCNREP3XV5YX8D4p3helGyy6szNwikkKQOV7rxVDetRKF91cdCTxfeSu4aq7pZwZ
bbIX1qqUP216R+yyiT30po8Mx+AjgomgWTzGWrGRWaxtlsMeCPYpK4zitNUEc+7c8gHd+N84dLlJ
DMhmg08Br5XtjrAjFjyj1joD3VrKFHokVpdql54z+q6BLh6RwKL1oOJjkO+HOFoh/5kHX8azCxiR
E/RQyZa9aFwRka04KSmF3wYNP4JcWlN4CJkWhQ4aAQspdVuVZLOWLeJ8exnfG3Vbfbj6p+XfhV8o
dzAhByhfjpqocrx1+Pp1by1Tsb2loWppyP7H+E0EhmdzvudFzuyg/DMe/hT8GSjfzHKof0XxAdLS
iVf+sU1z6CsCI+FhUYjlwjmxuIme0EOHHlYk+SaO0xjUZbuv80acC7VCz+38BLWluIGjVlmP+b09
wfqVKCMM+zpGCshyJUR8Kc7as141RoclyMcyA7iRzileK780ElSWOI1dIF+tJzBljqLAXzid3XiO
cfh7/+WvufQeZ3sXmp7YKh1yZcqe6isLWyIqG8XKcJFAWdlngQnmg22F164CsAT9IBj8Y6dzsqSR
zszJqBANrZacW3UZbjq5GE/9VLuNZ18bGQPeH7NkLHAwLgUN2aWMDt6pLaP4BkdYScT3eEaNqOte
30MRnFXAoWeVJJrzMWVOUaYWYtrVyIaCVj/zxu4PYOBaegb1QjMGWGcq9slVLDmePzas/zo1a5II
9mB6naVpVjYU6FZPFBjXTHnDXMQKHypdiql6d2Rzo0Y1GovBaBTPBCI6HLMQE1IPPaL+2p4+LoS9
AA2YYm2EtVpKAknQDOyjDONdSjDDsdTEAATo9ShXU8A/Kbogl0Xsi3ez5Mue2IZGdtlvkFn+M5v7
sYe+OWiYPA5319O+ZavcXqOTujHCWERdESIXSDuKb/TuAur1BpwfQ/O3uZyldv5FCQtFBEDCKxFy
c9JhIoc0AspfIDL7gilQIKO0CN7jZDTBIh4Nckw23tGVUYX+w1Ea5mVFeSV2aLh2aByxrooHYYfb
Qo+ArafPTT2OSuAum5AgKfCLGeOGkjZezuTgCLumrVzbHghEmO3aEAVdGvgyoHO/FHdctDM26Pl+
C+USkZqL/d6BuHJLWUxXwaTRocTjL5CHcSaIkTaZJJt5JC8u2lEOQtnPyQS36SR49ACrsWRFC3hS
3LZl2LIQ/n/RUYCbSZcFOB5n4xs4ExVaxZt4hXtDCLCymni7ZQgPeVKt8YkfciM63VrD/kuRKlWp
QkUQ2iJ28yISsKgLtnsvB5EQIai3/ryP4j6X3Vn+YLz+91ac7zowAE7/FcQFFseI+jBPq4YZgztk
u+NBOQy8R2abGWZ5huYg9Fbavi+gddD8x6gbbwzw+yDdSKScV713EtSnFj8iKYK36yD/NDi6gMjC
8Bm5tgQOM4yDRzelUIda4/kfwdeNPBQzEbTyxRDNZIwkI9bt+J0+UjlQbG8N0t7+e64ovPzSsQMQ
QqNpxrN3EBJ255SNLoZRBpESmvTkLt6+Z3LpijefWqogPeR/bQfhiCXK5WNKsLzsIA7+vqMPppXs
j7V55F9yyLd7XaZJr3jHAPc09oDMXBAQ1rbMkSS2B+th16XD18babrmLBX5kEu6DhMWSu8lSJ1xB
bh+oH+9Z9m60QmM6K6b9hw4Li4lKaR5KrfWX9AQdocysgMkPLeFYME5QboTFh+/dGd5x8Xuzwqbb
b2O9rGJShfAKZazAD+pcga/Flf/sMzk1dSMViQ8nOD4CY2p3+EZ9ra5y9PKFC6ToXmvpAVY97S92
qBa+vTmln7zt1aAess/ufY8igAmFVrb2eVFrLjdNhQLgrlyX5ob5On0y7D59I14jhG8thSvnHq+2
E8jLcljEfqOoSUJvhI4UIYV2ATgDEE4rvQzH0vYtFeS15XGMMl+trxJ48tSZQTVUwFuZxI2IlQY5
dzADtAAyvlZBxTp7rgw8sAuyh7tVHk+pXPoddguE9WBF0ABTpxWpWXt0u4Hp3EhacIitZcVpo1J8
HRtHJZ0ZOvUKb1Pw+oPy9XELoqQEkdQREVvuxEHiSha+m8AThMnO4LV3rSk4hISC+/+Awigj7MFn
+gtuzqOVx1KmLy/A65HnXkwXkxkVfUdDPbv6dGTSQRu6L40PuCwI1NipmPipM13OL1CQCbM4Fmox
RaAa/lj3SUK0h3kwwvBQToJv7axUY1UN4lmw0p9fjwsPfgXGotLP44KFrx7N3p4yLuzkpRlTuahg
QyMLNWLZXS05cUke9qbRo9FPaEF63w94OsrEM/J6RIesDgHgYYF0vPvbJxhz3iTqZZai+Y0gH8FE
z7YZ4RnVJUTE4wQI2XdUVI1gfwMuh+1jJduX0UHwDqpsoCe+vy/Bm05tLfvIyIXlyFLlA2C/2XVe
vY6hpC/jbqtIx31wphvuJedoFX3hxOuTFt8GGR9E2yotZaihpLdVLTFIiyCvUM+U+JCqduYPNWlK
zKW+DFUZxGuMS402z2nMN2UoHfoYRWNxDYsCUjdVe5AHQRo3yXpEhqUbzUJypGDV7J6GhpDCOt8A
ZYu3Ou3eBattoKRfdEBD+nHjD3h7LKjJI6tqtCFVC+WLLssvinVP4A1SnyITGXyrl1ICST2c8Mtk
rNN7TqOeiyNtm3hHgTpqouqwkpin7H5dZJAq/a9HmOakmhRgODASlcBlM6cKow5DmG4CbbUPZDEe
BFJmXBjrJHlPixoSUx2RXFWhygRj2N/EHHTDW85T+Fm8YP23eKMSwL0Ulu9CPGSD6eO5SJPqqzsv
ee9hcrbi9YfucK1zDmwphG0jQ/WXzhzwSv45nDmc1TOBJzuTj3YSmSbFaUNH8lmJ/TVBKd5xdXHb
OFGpOPgED3lurnFJrZfW4a+XEDOpNh3qEME/7X3KRA3clFO7oF7rs6TQ+eB4z3DqQgQDqZJ9Bcnu
TtdYe3J1Yol7sPIUHd2427BKgKpjqMyc4Rl5HU6HNQBQsn6Zp2MzQNh3i1Lb6CyRptUwNMs8/wES
aMW+1A47fXHmmJ55lIs+P2JDCW/OMp9b7K22Nz2kuRCQ/zUj/G6s04fTzt8rJBTTmQxKDPL1m6BK
NYjNkqwSWi3WfjmgMYv1cyhoCyOduJ1PsKYdyR2KtolmRaadz0cGjGlAmAa7kkqupMEGPBH1eaMw
o19ynFwb9bQyv3Kf0zYGhEa/o1jGTjyfWK7PZkzQ3MSb0Kk9aJrwSiRusDdKuQCYiOaC0LoFnSSU
4YbpymMSMmHy2TW8laLL75Smx0yiVLByLO6/ooB7Mfu/BiaJz61vZtrTUUPhe28z0+FUoiL0sXgW
qabxoozLfOlEsbpWJkfVcihMOQEjSpunBaVJuaAKNgtyFXCa8TiZCBVAMw5a4szgfwvuFlR5K1eV
FQ5jwe6QqJNgRkbhksY5v1S1cg2+s/JvbIduCPz0eQZME7wJzw7uHfhLDyNoWk6LSUmDGkUUO9rc
kJcmnpF9KQJz5Uxz2jwXHYFrFe0arqVhJ5UlX1gI4Uvw2y5Bprdt1F4n4EguUUzVFMArAh1dCE+A
r8eY8WZT/E0jacg7KyazGc9IdZlRC1KywscKIqWRa1HTju5loF9JGlVvF5hN2n/eKQzCnsbAYKJN
3A1JBj0442RmY05Fa2xsKyZm/qkyQPnu7jBwpH5bH0RgqjTq14PPNrTX6aOTUct/hDE9DUvRbNGs
uObwErt1Sw7SuUZqG/rekr3ZEMFvN7j49Y5EbnDCD66Aa6E8RcNSw9BCeefMvUASa+weH/pDMbYG
k8GUc6MVHspTiMYPcoiJKp4um4cfRlSxz6etJH4dBh0ns6lJR7IIqayj9+sCwovLI0Igk6a2su2N
lee07tzxMaW1wr268G8yEDQ2EstSf66cuemP2QyLoJsY13yaFVYulV8StyuZ+bxCiJdC1AT9aHjv
0U6r9EiMwNH7JUuk21v3YgzWnQu51AkKcucgD7ZzOm+OcYpsViGji4Pkr7u0zeB3VkQmyVPWHMOu
b4CdnAD31WFplMa8vvnKRCev8ta1lSUNaWpk/Dg4G1SzWzqhDDC2ZVZN05uNcHcq2PYQlwvOeKGx
Q4JJzHQIId+jjPf410OBg5TqKB2rK0aHTUxE096JSDGjwxdE18f0TABQqEYcYGsXDtUGTJTAKRiA
ztPttmhFxZdz588EgwtnGAQntdCYV4AM3rOkgkMS1zzFyU9Nj4BKPrt5oh61NlNSvVz3KgTP36gK
vjyYqSDjm5mIa3eV8rStp2EXxDSjVDsQjs/WB8Js2rym88jfJgePAnTk271e8CmadBL9jZ0VfWwB
LtOy34EOPyBFUu6i6eBF5rM/pl2qzngHY+C1g6r/OSBo8+uDzPXa5IxfARTJF8CpWFKZed/wqxLy
H8pXbtXbXSAFwXztiNt3AbrMeLU7JSGBF5naaGPjOQhXdsKsCxnrbo0ouLwY0hcGRAkagqjQjOwf
YyAEsZbgaqR0F9vOGiB7T+LvZkHimOAU/zBY5H81q0vrXWOJ7MtVLWrF22cpmBS7tjNePkp9XX2c
bp4WcaUBkbUnSa/Bdrpyxa3IXqh1kf/s0hUL40sxZVVXbqvRQ9rH5rkb10nrozQNtkzQLHHL97ub
2sM9IERyY8j59GjQGLsFn6P0DaPZv44yPem2yvB89tcmO5UK8V+r/CTVc8XlfOyqnGE4apiXUkGU
yuiKuL17wzJwUEf3iO70tm72sbroKO4961AizzjxV5HN5jS9/2iK1oc+GuD3rOpNDFFCT1VOR8tu
KAES3GxoqlZ1CZqQNJNbI1q2647qToOPsf4Iy2T104z8nouf7xf4y1necQqKEo54xNd6jyPV6Sz6
j/wGoiw0hREzqnOB1wvtuw4fQ8hwkfRudDOTOvNDnCZP05auPwYqQ+4GXt5BDk3A7P1Rr4bK1xz8
4e0Oo9+bsPKVVtYZCROhg0fB+m0ClOC9UI8ycXEU4w7maGciYq/lwdwnjQWL7Nmr3VJPDsCoaeuu
YKAUS6NTOiiGTmhP0/SRV1ZTdZMqA6UYlm+aK9ltjmVp99Ye6LJXcHRHg+l1O4cjC6afGDSQ0WtT
Btt3wbj+e9BfA4CJXZ+tMIO9NtAUSRze0vJ0Fr2ZC8nz7rtZ/EylDCJ8CJqeH8RB+4k4wAA2GCfL
yT1h1dcKKdzla7z4ghRx8iw5+sq4TrB4N4OabVLxxwDCt+bKiJpojOHaE8aAfGKsjI+tT8yEOWeX
YT0Hfy153qL8EpUf9RzR+DRAZotVYs5qN0BpBcb3rlL8kfv6StiQDxvdE6aD/cfdTXpeIxpxGZ2s
OSMXInVKkFBDDJ4xQofl0fICFdHptVgHxJ+E+LZfc99W8xtGqR7Hkzh4QwAEs4Mbc6sdULMmsKyR
MYw/ygA9G7boWhX1cTF43kEoWHFLDRc/aTWaoTFhY6R2slpjNYl1TV8gMKSM3/wvBWugbzcsr9JH
JIluAE2JVtTjOwnMBQv1n2GtlAEoXQCqqJSteXm6vAS6NNRf4GWBOxbm9KiagJshtduEXf2UUMA5
L3fPNeML3zu83+EGxn5UI0cQQzFLbn9Xo+pusPYXtGZ+qBvwmbIfXKzrfFjIR2D7v0vTot2XJKvm
4AE0saNzhIa9sHSgeS/oMdMUM/GtfiL53OGr9gNN8INLcyYljsM9qLXnsYFrhMfeoQAogVeWKKWq
8aLKlnI+boE5utMgB/r1BoX3zHhdSLHhaj+trB4fB5zFlEf7PLC1vEPK5WcTqEPN+4dVGl7KgXrQ
uMnnUsUXeNiKae9BB2FSCynmrk7Uk47uDWKaDDvZu1NV7cERnKzDacYVZ4IUzBWwh8YuZSEfDE/N
oYKgAqHKauL70avq09nYAWqTfy1Bkdw8MxaspeVtEDm947/hL3YuDR2XkEukturB1Mr8ZJmUHZu4
ZTPRPaUQD+gcnoGXsPpFP/mBSLY7eLG6SHmfCmwe7CQxXSocc1w+3fRQrBPfAh+pkuPJFPGHvf3p
s4WcrzLVkevL6xHthEKnx1/m3DEW2/AzIawTgakDIZqjYoCLUoUcdtV4HkVoKDz39kh5WcUPNmUz
BLCg8ZBrzSAZbGzLFeKAyqBXnmvsDeiIOUdgfGTe5sDNw7rMhBW4fpt6kACunsKxdMwSNQ3bPNuR
hiiZIiaFPSVoFVWWhEsKlemRTNx3cQXArwB4wMIvDonRm7rUpoVx244++3NgTtdZ9VMFNo1KXOzP
xjx7bUkAhd8LI2J16vBMy9dnHx4i5sCM8b1zgB1uXrEFD8CJuRBfsADcM5lrqnuH6BCvoFoXVrIC
uyzPUF4jYQctb2+WT1H9TnLO1WhaH3jFVwxFWF1zaIY1WM+D1dGoratXueU0Y69rvNQQrbMB5bgC
RAEyepEsV6iisD6KKpEcy1hblBcqGA7mVgfUre6wPbq80hJRwKj053y2+9QQ1SeWAN3Koyz2eHYN
2Vp96TI4J3UZkUC7e26pLTefWIaHhvsAONDFE2WkUEP2JKnzYPh84y1nEceOaMy9y+sW48Bsx/9O
bTWYzTcEToCkwIuIsD9AEJWGiYAZtBIhdF8b701IECFuyIgdxg3M3c0Yf2QhYWhRvncPl2gi3J9f
eG+BMwReFkknHuZZEDh7I6KrnhMj2i0EgOIhVliDLgzzpCLGHZxea8+N/NyP5rqp2OoSVczMg9bc
WEt8+v7WCAUoxOQ361P/wgaiv+SV7uZsgHXwiamY/PCNUsctdcipiQcF4hHuv7LNiQRWT2bjdLKc
butAp8GpDnapqRHHpoYbRCl9lgPUFz6phPEZVjVKRq8e49zNuukyR+Gu6SfXk4CpGWaAx/ERIfLI
EeGJCbvSI1qoB5eF1Q7I1ix+K6deH5dDpvRtvydB6UEctcyLgDJpbxlbxzs4n4Go7Lx67oB4m60O
4Kcd25FgvayFs5869p0Xx1SbI6igJ/kGnpU1hTUJ3HNIQ6ZJdDQe+JbunPdmBH6FAAHryAoVphAf
Pu8TaCcEx+kIvJtodD3Kfanq5V8QpGuUScpxCJjE7eZm83GPTu2RFQ7m3yOL4i3WfbWc16RqRF6T
wtywqfd5vuASy33QQCrWtXIbLkoaZVbnGsVv5ygW4JRNDl1re98H2lLFOxBTKaffxRLEr3sk6yJF
/+UEoMw1Cx2zQeCvqlzI+XHfdGXikFjKuET0u+/WzI1cxYLBXI45lzuGETq2rmzsL5utt9NxwvyS
GNiB1qKX6BphATh+scs94iztrdVHBolgbE8JomoJZnFzmsOXpF1lkciZIdlz8MzLa1Q0EPUmYT6Q
IxpPykxPMhmiBCtJmq6PulvHLDXORsrO1Zl8EfJIYuE1Q1SqKUsxoWwCyCIMZmM5k60etpBdLXbD
hOp9HPP8ngS1zL/oi9dsDIFQoKWlGouNfLftSK+YUXdmzkWNh+JWgMNOU3K1S9ulUDknCg4h3a5d
o2uS4T39/V9aCHaaQxiz1FeQS4vbl/OcWrrvJlA2Iag9AbJRdgMlOzY2Zmp3CVKyweQQgkSTXtpw
pWVgYWQ1O65VzWZKYi2fFfrRUkQxqH2g3KKAleTgM2gH9h+TycRVlHdb9kblAAHkh2jA6BqF6ZO6
akLIPTGGvllvxhOJ3jy2BT48gpJ/JVSx/mC5coeHUoGIX1guRUWJqRPOKYXEN1D5QvUUUhM+zFao
KPyj9FRs8PtPzFJXWxxnC/hCo1BmtLTRN2rBKbG8aUrH1atDkHsfGhhKZu5/WFF1OGOXn1KULjLm
KbBFDNMGuGIp1qNdEGUO6heZmEQnbA1u/d2I+Kog8os9qUduJPvjrAOzPne5weYffF5nNbopF9vY
i77Dn3kN7vj/m2nRwMaYtoDXKK9irsynwuiKSxHzojtXyY85AfKCUmbgtDngHKmUjD1E5/Jy/xNS
2WJuvKe57fPiDXBae2VjYxfQeJbzT60a7JURYMFr0LytYB6u7/zqtmJQyjpY+0nJUhZ+Z+QTf0W4
5ccIWlxoZuwpNwiQVlE0xx18rCyo7Yn/LIUyJHYtrbevfP7RPqjR8mE4vUr3+5+BuyVYkX5k2Zbb
Jz6B3FRQHOY1dBQl/Gh4d7Om5D9PL1QCyoOhNYgk9W59t9Ivcc2OyVbjJyhVZ1ulmRojr43/R6XL
ZIGpWLWmff8S1O0zfDpS8/tisDDx+nsrK+hAq9J3ECzcnfoPAGKG2+x8ly778zZJTrgqY/AjdrD9
QcLFKyvz/Hv/DwCFj2EO20UpJP2B8CRrubwXXQxTialDk4A2+sKcFPnSdXF2J/LpK7Xd6Is6Z+El
xaavIXqnRLDR0ibySt1B+UD+ytdMkY/vTQP7uWDQW33M0kjl1JGgFTfealh/TJClUcu9LTUFiq/S
YcdZzsYYwiigfWu0YUSqeNIEbD0cKM1GQGC71qSiqry3NUEWHJbqGMUb4khDVC/6c8Rvy1PjyPUO
TCvkmBlpI93S4YCnpP1F1Yoi0EcQK5eSOEPmYBXR9LBmoFKxDRl3uNY7FZHTdrTdcsOs8UyTWhok
NsNcy4Ez7xgcR4q5b/JVjEvFerImNE4DrkD3PORtmJi8MddxKlfoBldLIfRCLstxf+Ng3QNebRcj
7JbyAwuuimdIXRPc/uu+7h0lBuPvHVtF3vP3SfepZwD9nm+APn+/zdihthgdgbujUcNiodPo0Suv
0Ly049+QGbLOuPpfo2s33y2Nl7ewAzGuKZvirOQZx20nSkRozbbJPNMTzMocyyyZwZgNor0ZVPCq
oPqA1jP6dnGAZhHeoC8PkUe2v8WGxt+r3Yo59kwlvy7kJS5o5wYOsfFAgtNlfmLWn0MLYHx1INgH
PZ6m7sa/K+EOwGELhcrXNpyZ+lbmPfN0YnM25qOmGhJXQEbmS73tjwMn2Gw6GKbEHE4Z3KS30mzo
VRCDGmEsX6qbFHw3KIc/EJyoVgMb/MVA1qbdo9XBqiZpr+tXCrwULkwM5cz94oamrNnuRporYMMH
9q8AzfBndfiNvMjFZKy/WHjUVNdg0AUenorInbEWop0XpWpgI/fZ17PZlxA/H/1+rJPFrd1Diy8Y
zZerA2uiF4aGNs7wpTEvDu51GaCWG2iNyfA5k8flGqE4IXq+KCMBNE6eoalQXXhL4DsFQL5oOZYt
EUZ8n2yJ2xotHAyhQxPceDUPDGlW/Vh0TB0oGYqrb5FdUmQYeCpfbtuCHV74C5s0COLk6jIXv3n2
0+fI/BQLXY9ha6vWkgQLskp6caqFwFO8sBK3X4u9lKZrVfar66TDV0pK4qkls41uXh6jPTxM/lBS
CRCHrGq4KD48mq2l4XZ198ekr+jEDpP/XqDfN/b7tuhaEX4WNy+Krwz64yFEHZgLlXGh2neSa7yL
GCU1EeFDYCcGCvn+edKni0ICwA4u1tUmXX2HttmAsb27KtLAnvvfDEpnklOAW8fpe/B2vl274RaK
H+DjK1dT2iKVZgdfmjcApjTHt889Qmm/5mM+KBr11AWBm38EAAsUHwsgrhJJpAQ1tZ+umX/LMzZN
MECwGucHdbtVnGsU3IrqZHNpclhDQR2pc/B+/fmxGb2NvpU3w0JkwPafi/8fqL4FQVzpEkcsYPHs
awCGEblDA9lpHzI6CusObKA/s5/6l/jtw9CqKANlYjFHKMviJmdTpnmfD/Z2snzXRifZ5lzMs1r+
tvWlN+t2p/+Ef5sSH/yXOK3QO31pgOwjeensXNbInHuHCZtyOXX3VTIID1quEiYx7hV0L2iVgaHt
vaVUD8Lf4TduPMr0KbC8ZZfIgiLAu8Kicqxc6g3WqJhU5u0c+Wy+3WyhxFELmGqJM4p5Mhbwz7X5
PU2KD89UitV/6HNgivc75XkceTxk4+M38/F3tD+2FlOiS16t85ksx6i8wp+Ax8LPY+dxCk3V3aGT
sOQY5az/UKquo+1xKJJ33DGW5m1kv5tkaatnvbeuoC3qr1Ph5PsZGSHFxwSY+aKSDAgi+X/uaacW
6q2Cs74FoJSgCF4pb28ECflgouPe8gyhFqKv3LieoqtXIDuJxmj8gWb5fUuQTisoRBs76C5KhxkM
RxDzB68j/ad34B48Ht+J6zx5PDJizJVC/w+qyzYiBN62AQvVSC9S/4hig1MDesB1aJleWVNFAM0q
PlXIRBjRycDhaAZrQRqutsWN6OgXZBeHHAH8pLpV36VcbKhkaRd4w4TN7CY4Wflbh3EbLZE9PvdE
9c+arF5+R15eiGSo7W3iYrJTGZ8zpBbUDLamZaQHoFo0Y49EyGl1suBByja+B7zYtTlWYhuHy6k+
jjdWEXYhfMNWB2yUmkYRj4ysH525xtn+vGUzF682pfsqPP/HRrIbfcbBoRGaveeSJaYs3GgtJ5W1
t3y3aUIfgdrz6mZfThtM+xRVWNuZXYlX4zccrkePLN+3B7pDhC+bDywhWH3s8liO+m8+XF7JF74v
UzTubU9kfrLfLkAqCQj9qtbomB5eR6sGEEMYS3OtyFQTSRAJXH+F/MKckV+v21yegwSmzhB/SGt3
+TBCtoMbzXWF6L57XslLVDISNRKs72IOLidI/irLaU8odlRcaLj3JPR9PLM8ZDRFDap+qj8WYXWj
HZ0yane4TrNrOV2xh3W8lhy2HNmFoHOwmARivAczD8UJH/DsnfME17En9Z8OAQeGhZhLl3YHNxXL
B4R2HgV0HyOVujLI9DTx7ztii4PAWqYa5zHwsaY4sZvPAJ+v2SjHZDQ+N7hp3BHN/gQHxbcjKobE
bkr4LrSJoltHZ1Orw5lA3dvRQnsIN99ls5NyWqBsJAOS0UPdE0WOMLaKPgzUYKuMLvW2vkAcPCmg
qsvyvBdF2nXXoK4Tng4C3zKr4JnrP/VwDx6+bDAXhAb1g7+eqwTGLO7pFXWJCayokDRihapQ5c4B
eVUPDgroRDxJcYswY5tTLAgc/moM/1I/D4Hxv2Xw/P1WZlcn1q6/KtTMTMZpj1QnqKLzPBLGQ/GU
jK8XWX23wnkiuA0RElaPjzecVK/RWPNCPZKtB4y5fw977oJB7dDxT9VOoJmXLtoDBj1x7FrbVK54
10wEsSO5KbhW3RsXVn2aji9MoDr4ajmq02Wvgb1ADOIruvLl0Baz4j54rrv0U/V92UufN/XJyJCn
Zitq3lKHUn5kBcdXZsKBAFAiWLVgEiXfttM1W5h4tjeoeAhq0/nsgz4YG3y7+1WX4ySThoRZ00Af
8IqLIYEU1GML816Ljt+1Tx5Z5TdRgTOJryCsHBO7eb7wMbHVWwFo4ECZvWeJ6KnXVCj49Ut3zlB2
41PNDaxU+5JTknDt+Pk30ekVIVTzchH1XGW3p1cw+KjxHEGtw0PRh+r68d+gmHQ7viGYg/OevAdq
Wsk+HtatoeEqkO9J7A/i15Gwg8AT6qkiRY6GBCaPKGLk7vVLO7F8ylClWYcwPKWHV3+91jBiirzC
gJeT5qSDDCMajzuPVHWRrySANuKQrvzQU0wBN3aGOvBMxYPjpfxf5gJI9u6gH149Aqu6MkJb8piA
xidUf4F9bDexqVbeiDcyjnbjj7n2oTOG5xLQLemg9gY4XlYYGLRowoEmEgKEH9jN5w8MdZ8l0Dl6
HmmYAY9Rn+CE33JhnCayPdyt3OzC1PvbHIPxfmCUlG4xiZb8OeosQJl5h1RBBVCZ04pF1sDDS+F7
5MitdLCupn9nzw34rdVGwKxW4o9mr0dH4RPwBAEWsxz+kWPgvlVDunJ6KwKPE7wuSnVjbd9ApIUU
oUdpn5dYSqe3bVWRM2/OXynfKA3QK6n8tRH3dcJuDdqCX8+Ms+jgua6koDK+dBmqiVcv9BjTI7zw
ydETxk1i08Hg5NDTus4O4EIuF1wjMiXons+f3cWRIHO1PN5uXmVKf9OpnHoFOT8kvQv2CXBXzVV3
xr8qH6L71UiRIw+kFPGnHVXQeRMW0cEjm1AcAH07g0WSgeV9MQXluCeEAXMaE4ZKO9EWGguhODXN
cJCeHsXLLXaU7NJMk5YCe40j5p5FR2Qsq84H6pa7MGZ5DshimrvMqQQWGMYUNcJEhOBzpluS34Bi
2MlqUI1/P1SfgLHX8HHtcU+UqTplkBl9fnXlO0R7FkBWIXNLnFRgta7x3v+/PfWaZswCsMeGP7A1
VmdF5EesqBZpLn3HQHbrbnxQzyVYxsddLfg5V5tICW2kres4GRPJ09zB8+4SqdIjZtBR+1yM7X/e
z4ynb7fjyhAg/MvGzruy+fNemYJEbW7qtDOmXHowEbUo4IQiGHQHCHC/MpHANXAjpXdHkJjGyAvD
DhY4q+IHx2qL3pyli+/k3aGfh8MAr0q+tXroTdhOQhvki+F9TW6NemrlcAS4rjr1jHGIFRW0C2Ov
oni+2w/5MNUeXbMCwpPUr8ExQ/MagT9PgAnLMDdqHSWgw2d/xyeRFsa2Y84MkA9iP9kRdRvdW6gb
MoaR1EHH3JoxZ01L0r2a6CCCpOm4cXkecaFOpPOC0d8weFf1SsrY97RvjHkm85CGm9IEs38noU5d
01YEOUY/e3RCUW/bNHyYFIOqgw713hjg9KotpoVyHUInf26CUCf+VFHyIjApxVm2EEsOMyDFXmRL
zK3sf3t6QxYOEK+6aTxDXr9wn4xxAWAOG3eWHeLC5pTPTmUJyT2LZ8cUL1WKJLx3xctKYeGxtzOu
g+2WOy5QzjHKlTxkcjqc+jgyMRrsgUT9PVO3a1sD3tKr7Knf59PGyg77rj7kPgkqc3gVLNlFxY4w
gnSeFWDLNxWkWannbUqySmV+iT9nfm/lA2m/SI3teLzxN4B5PEphOFQ2Fx1rNylbHbvM0Oo32lzV
pkJVgFJiFlDhKhP9OkdDrVn0rSylDeyVr8XBzAQFwkAICJT357WawjQTdBD2yZTJLbRs0JiBnnyQ
AQJN+VvLUbcDlJdfwELbMBth48JoUjRFO4qoHL4Ggr3RYkqvpgFgoHf+bo1k4izYu+l+TO8vAA5C
/pj39wK4IPRPZkH7Pk8zKV/iGWx4fpZbLsQp0u3QAGx5XNQtLWX3FmJaGs32h1ovHovBSnW1KeuC
szJsr1YSY+RMihh0szpNHsI4wO3d2edeVTf7vtlu6g3NHWT67UFwpBX8+yOMlbP4+hSQQwEsJq9h
v2SIjnPsslEU5WEifXvraqujWiq++2uQ17qjzAeRK28mJCCdfX43+YD+dd4ItOsvqrrPT8zbH51y
bzVeAk5kU88kj0nhpRBN9VnRfI3FoOellM+s1yiYKEZ53mRR9PJ1lUtj8EfzVudQnxtOp8v8lSCv
4NIn+KWDGeUuFm15Mq0X04IBy+/Szm0bgxN8A/mSQRuQNJJ1of2LXYW/NTJTvclhNCWlQA6Et0p0
qbq8+PmGs/tI+aevEz9iX+FL7Ep8wahHGWA2jcuDlgy6vXeBxDWd/4lTp4ae/CwqF8tydXfu9OeO
XYquXNM+GwtCcQk/h5JAIPckPd2RrA6N+eZ7yvJ39MvcJ1CCVA6JHqXV8bJqDCWnVrL6SC2C4clN
b5tXXxcfAXfWoWRpm+VWNL+ZIMn3Ek21zWy7+uMmB3XGzxSo57ml9UqMFLF/4qQJ399dGLAfCJpl
1NmBWTezjjbIFr6iwMg/orj6LPFoFddYgHIXqtx6c13ge2/kQs7wrKwPzxjB6sDMg0pwt75MuuI5
t+hAQKtGgUgQKDhLR1lsCnwc7irY86SIh0X2UtMX/tX/uv0JQTxDJOKs2hICPcYnl8d28+xLE0kr
hDrHe3mI6rZ6uTtHBAzNjEL8iBqG0D1O/4hucOPqOCreqoCBGtZf9nNPKzfPkAaKK2c3x5SSSEZg
f4t12b1X28G5ysbfmzISXkdzPTeaGSdyM3zAKj16FWXr75IRZAiWJNZDYwpaS1/epv7ZUKoU+SUu
Azw3Cngpj5Y5M4qv9qxG6sRTxB3eZWbq23LF9+zWa06FaI/4HmtlATYjrPPsx7k7gEdKYsqxrfSV
2IW/iW2HayDKcC8raTY0fpVhzYST50wErJL4jPac8wiqU8tgwFtwFi3/WUAYw/16LPFPKcBK82pc
OWrs4TnUu9gD03rOOO+QvC28bNH8OFllynI4YCw4QIMGK/Br/L7smAn0pArEhzmTLFB7mv91QhUS
p9i85+PjCta7bV8OvH59AjIV9T6phJp6ikjhVcZZjWuK2fI139xvLkpOhIhqSPiSgybRNb1Ej7ZG
H79XGA0qOOVHTb+KIU0LZegB7UcmZALecNXSbOnZVn38Vh111EhIRqtt/G1BWVyKaOQQsNVkKKEH
RMis+XqcD0rBKlL2xKIHqjtcD8AWW8MCPo2yrYUADpsldhwiFyFUthriAX+/ENn7kgpt4/sDaKar
BePimecoPYUd0hqZISDEG3/qPrL8LRDDoDoYs+Un+pCALwF40ZMimsI+j9+6MBxMeicd4mwwbbCE
Kp3ZKmfcTqDfrIdIr7dH/GULdrBv7CrIzraygRuyc3Jk1WugFEvxkuYf837hlIhdXctPpfBIeUEt
+61mEZOVaUEEC/yMCaWZKFqV4DcXDzeWO3pcQ8XE0mrjo7FNnY5rcyqVtH0NYnCwv57R0rC6Dgek
/PGmWKvMX/k9xzkrzrWdWgYGC4SMzqO4JzGzKa9W5MKGFNa9i6HZH5cdIf7FNumgxHWndHDIPGI4
cxpLlStxrhfpGJCDwbH79imTime0JtTx0U65FTBDT7sAS/0GyK+Ow7zjsiIhV2aVRDVgwtkgELzZ
PmZjZzK7m4V8NeQkf6ODYTHPZRV1KVNri5TRIdyoS07o5UH09WVRvberqh25tWSNXqxnUdt1FASd
FBaMZBsqspPwoiTCR20dYdfeqWK1seqaqxbozTXjSQoZVUh7hJCF1toWH2nZK8Mob2jaWvxvEXSX
HU7163qSFnuO9mQ26BPkK8E+BMx0/qMIY4KJ+WaXfwoRFYgtaJKT4e485ZGJdsYJNwZyqcN77JxB
DclIJsOsfegZakBncZ/lCS80tOSwYGMxmqpFXAXZeB1ujw+OXhK8vT78wB6sThLzX4MvNc2DDJwn
ftPxzq7l/xWDgfMCc1ThC4BZJWvMmef7EYbwYGc2UD7jNYoKAAykx2n7Jrg9EQOtHqpIgCSlzEDC
iu7NBokULoJ15ReYVsMeBRDdeKb8xBt1GrOu+TWBbOUC+ifF4OIOhEGDSvBYQAYd9LThE1PTI/MG
Sf5zQUskY+PBKHETQ5e/6au+YYDTIFoONKAhG+VCLDLjif1n9qvAsxnAQAd3RN0GuIibda2aB6Um
by0FDK1FTplvPM+SNLyRa4b74XwBO1cQqz9r9oF8k6EMm10b67g09BXt8qOP1pmrXbAUql61uQxq
AsBrSTicJWS3TxVtQ/QHKkL7K00hQBnHbDLht3QsDfSi4miAeRUoQaFX0cbBhBUrnwnDG48ky1V+
U2be5cCB5PQwdDydJLLN5e1NSRN48lRWfz+VybYxPCCvVJm5ALt7LzIxirbT3NiWmP73b3FlfTQU
J57nsNN80IhDt0BmVbt3nZaAYgUxe2LVm279R4ToxP8iK0d6d6FMRwdZiF6CkIeDMkTCCos7aYTn
pt33pat8p3iq7Pk8rRxzRgP2CsKtNWf68J8jJnBCx54owKPcFPnxrspG29p+463zHSxAQjZXYVos
Wa0a55krioeyfvKyhp/ZCegGzIfqpSzZBS2CSmOC0D4e9XuLsXU8ESVbfnuzm9vkLAG5lvTXyQxV
3h5Mn19uHwkuupbHiVGORPT+H9/N3fS1d8K7opVaIm7YMp6gB4b6MMSPk4qzb7yoP4e2Q+GI1S5p
kl64B8pnAp6FPiDo051vduJ5Y8ShlwRVFtbGru78g0xOAYodMUxjRbWc+moS5Wm35+aW1qAkY7zJ
K+4ZSD0Cn2y9h8jo55NOIoVIIZmMZLrycpim0Mwc2VdYCub8zZEa7ceG7c365Pq+hwlYUKdYCXni
HJ9JtD4No2o+WkYVGYGzte2ZN/CbasDNgu5JpG2qNarugYxFVytwJbWDgqZlVF400TyMz9x8wsNv
nl5bx2pXruATYPiOD3hXDd6pY7K8C3NET65bdn/Y8aP++Q0A1XHfaRTYEBJQUpmUyyaisi5Q/Gc0
eAYljPX2gE28W6xqJS2aq8oOVsEMWZ/Q7wmfjMPLt8gP2nFL6KqlE2fZ9nxaLIn8371AlWhlEWT2
sFI8oH/V7CS6B5CN4Qok83XPc6vFpWOGO4s8VGUOOhlBuckw0vYi+z05yvEl8BclkIOlBZkKuzRo
ZdGYK5xq5IGDY8S5tTYJNoCqFOIRZtROkSaUwCs+Yelx80lq9+E+M71vTUbWGc7NgfMKS7v45twN
wmNTEge5cRcOErjOcJBvIzPApr/s4hwE6Fz1rk8t7g0ue1Bjn1LYs/4qeCoSoYxv1U9u9CzypIVY
R7KI6mKUydLUdyk5TTP+AXDWUzyUSJ/5UzOVtvWArnEbsjFmszSqIVG9Go2fdDHvOYMn5hAm6AOH
m1aux0ebwae0+FylAw3CFLIW3OfG6Aum+H/imjSO7ZL+QOANL3Uri1P4q5WloUE3sYz6vVsZZVN9
DXNnb65aLAArq1FDQFykfceCcK9FfHGhl7ei4hqBU0TXh1Zu964xRkWp891eWn4lmC03FIakkm+C
KaebMLINdoLzU0l/PaRv8KKTq6Tkf/F522BFI1BPCOUll8HQ7zkzDIcm26qHkK1LscoXx8GNSQ7G
nNdXgjOndvQfWQ92rDDbdKD3hIBmscvmdJl46cMghtZDo9mGqXc1XtWUblkcEK+5ADSbuCKWOyH8
7ZQKQ/nZK8bwyYhDOgGEOqzqe3yJiVC0kqrl9fAVRPr7MXyJGfwny+nMsVFrFJ+etPuXG8d34WG1
AeYRgotaZQuvFqBObQ2Mw0+k2lOa80oLHJP3jpZI/WCg+5ubVDHSyR57TbCZPaz48STgAvqlgsAw
eC31JH1pbbJ+rxmAnS3o9to2+jmwBf0qRlEeK2i+Q/yPSy9zdSzkCHox1ZltF0TBvl5kIC0gBwKW
aAPsaq3llDlXl91HYI5tPkUTF2JQzGXqE8B7QhunI/Z4yO14TLLmNIujPumLamjcOQEq2y11YKWJ
HcfXbx7LzN7yaZ3ANpxdyrm1jM7L89Z3N0qNnB0F83HA2yeBCZGEIR/BSVoN89APnBhE/NOH9Jh9
pa3pFOY9wszIZMSX0er9qAh1n1DXoLJuD1tzmFI5jTtwq6H4DtF5SUeHHxauW0kLr4okbGt/9yHO
vyud8iZRmqOyboJviLS5ZIfHprABh836//rg2bHU+KpS6XJck1zerCfSy8dnH+tUinajDdEUV8lj
VoxsEJPqput7Q/M0Uy/FuEdVCuW6cLblAhPXm60BDbOuZUolIBvMobG+0b4dQYEr6wtqMA8pOmJZ
l4/TVCfL9t5lUVFsMam3hnW8iTwnWEShCaXjv3qaSMFJhUAeHh1GJrW7YfF2SDUPKX8n8aUiWM/J
DxRoh9FuACE3WwvHbeyk0no7oekeRxh3Xt+baxKzl/T9WEXXBW78UParxwYYCblcSfY59fUv+qu/
mXt5dCZM3vaPpAQ+tQbBxGzJh5CM0lUhF67cRlgcwzeGXeq0eq9TMH9zKmfnjqzlrjw+aXNqresE
ng4Ry7erB3hq6qmgfgXzIEEU9xqZV+X/pp618sJ+96Vw8FAtsDzlGPkBSzcp7tIQxo8KSUdJzarV
qJV9h6dmNm7LYyLCMaJQSxpYJ2YUrWV4m85I61nWnVSO87YIDqHJnJIb2dwHLs1DS4TRjP7u2RCZ
p2bLxPr0Nvw4whoV15P4dYy6XgDOl62Vj56UnVRygGWQH48f6MHfV4aUyxENr35u+vBUhj15IHOv
1Vxuh6CoSsbQxywm+zM3bk2WPMHh6T6G6MvrBuw24mG0RL6tcAADOkT1VsqVQDFLAclMFm1TEB7V
K4iT5vQdaLOHE1JVG8MfV7NI+naWaKNgcsOE/jFI7mfOcEABaxO2IZPSWCxJtJRQ1Cg3ZTT0k2VG
tVgqdossUo4apusUIBZJsh9Z79AXMs+0Kltvqwne0wyOerpYAhtNrbKG9IDqcVBpJWH3hbJwc5o4
JzYoX57+d75DFgqHzinxIYer0egV8CF8FuiG/nhoQNio/truLHoSjO5OIHS9csgNYVekZEgWlmki
kom6qSq5by5LN2Ja0ikatcww6SvJuz9ATE5bgirUF3pXVlRwSooTLlXR4hkryd2xNKQqA20Nyi9z
mqWxMIk4fcW7PmBTmuSwH4QgbaSdsz6zYA7mrNxLOfQoiHxc9upn3muneGXuAFZZH5f86TFkvaFX
ognWE8vBH8Xz2/9Hnm+kBpF+/xlfeV7ZP3pcTFX0Syi3aaPToaipKS5Cb2xlVW7+WdcNxBoJpsKI
ea84GtyYBSeYGToi9h0udDOj5Hr2GLNwn/r0JaLyx+gLQ7V9T4uM+AFWbsLLbz6VjaACbj9x+ZvZ
HaOM5BolrP0hUs08rZwF3q65BzxeLWdENgJWzWKr+12OXdZfFHbK2Iq3UWSc37rD7VOpFi5HaOD5
1EG0U9qkvO2QnkEKMvWfUplHjEPPtKAM/KOEZFNbSdOYQG8JmdKm4RTgdRPAh7sfQ7XOOKR3TBPm
eFqDfmFD3FfgWD2QgMVPJRQmtRe7/JbRkTNQkhJa5KBUKWhtOvSRN+kUJhl9DAI5rpLQZlDOvoL6
HbbVUkCGaJHHHAsHpIhVQg0pox1knlm4qVQudgZKP3g16o+r+ul+R15qsRXI3rNuMQD0ZWfyhVNM
aEmp5j9qaj9NiuRBiiY1oxwAA9VD3WCdKIYLec9FxbRJWF9n1YrjBNYgEHLccTWeRpXkKCr7VUEJ
1l4pCdXq7NLuTvYVDlS39vPrjgCMF+wrMYg6XNHx9dgNRts3fY/Q33i2OwzHzfmfMS5/vz9E4Pqt
QbQfsU6zmsSToT8cmWF0K2VsgK1L4EMGTAHJjZMy/ck7ONilhSXlqUhhQS7A6Yu6/OCkentvWpxp
CJx/yXYTmkpso+c2bMwNJ404UIZGPVg0nA1gAwxtxq6Fu4Ca9/sv+VGg46BF47RXSj0KlPrUqz0s
ziMC5HaUaHukiG957gYp1N7vp5zXDD/JlHDobxSxlTIV4OtEVE0Xq2p368GXc58fLczhLhZLTckU
7kqjFKko9+bVSLvU4537pEjxMVpfh0ydsP/kkm6+TfM4qw17aSjPWEiV+Xm92yDXp+xkkFPkU3aG
8ZYo5jrIxtnN6XKnsVpDeEwConqb+3c121SA1ChnJqqhMQFwbFsZufmmJ6obI1Npx3XopbNzPKb2
s4S4u+cuc1nAqreRoRv+zBXGVLnt1lUjYQ/Z7uPF0STtSWmtm1h6XCr3nuCEGU2l8jnmhzrEscNI
aMayfD4QSxZT4n6lwkaUCo92NXcWhzDqabbPG6I1jxXTuwN41f/HaWjD9SMc/NuE8Xf5qIbaRZCm
dcoouTbCmIRsWBQcAnZ2Ry5LJjRLqQo0oHEIWHAEl69jyyqLCFa84lAAX4rDfnWRndT+A/sYiuAT
BkRWU5M1jL3pggmvWqEl7A+A7CUlaPGeX5j3vWsC6BiCODHbh8+kzMj0jXvoetQSKxhN1y1jAq3h
fzH/cp3+Tb0/P2f9uSc29RwoMVmWn7ihaSiGrwGny3JBFRzJrmVZk+0MNY3q2RmQqT6DeqqlV72U
AnteRK2r4sq48RewqrDfNiNgw/DpW1JBpyGPKx6sN0RuK8i1sGMAznrpFlJP7F9zh/jMsWmTGIst
gsR+GqY7Sgk0Q4IBaE4sM4U6vbHo9d+wZ7Lr2CKCZQ8l3koo+VklZ7hUG1rTDmHQb3PQ3rCvpCrW
K2/AZdlfhgGoAFDYkLgQoBB9SriS2UAFQ79hvWqZSNzR1sWKYNK/LC6E4Xkvuh4kGvLaRXPt0KPo
kOhH2O+H1tuR9V5LkYeHoKWU79GatciH/swZVnn4SS74LDnd9cDe8xKspIvP78YBGvcQC7PjHAhV
jpHBYVyiNf8PxXp2Y8/SfATOeltjsxrA64k/2k6R7Aef5U4N2JdEz7/+ainzFXqwtqkycDGdLUbc
yLIY2pqVVL4uLVPVL/ylFOjljNn83gSlxQy9yscAZPAhmRoa7ztlTIS2o95Qkf3kBACorY+q88a7
lX/4h1c1ySTl1VlSYTKvn2sXOvcp3+RxYVo3UdLYNbzyMq50DRZs9fSC5UO0V18nN/r+WIwxDp3s
Etehqyy1+OIgs7JKdTZn8yUSc9/utoXDEbo+GHkW0IclRNEX20N/dR+6P1LYbShlzZJFc42a/w/1
gY6LTsxJN3CdKjPGiahTORug0fRxE9sNUeDiG8KoolrxaujVvdCpfWie5XzAgwmY87NGj/roJ8Fs
34BIySzt3lhYchu6PIx3ybax6+wQuAk+w8LvGyH2JW5yfXxMezg6CPb3fk9fs32v9ofLF9SMbZ2F
NbZJh9M30plJA/7h59ZOphl4QQwvhLpMOhcM9k9mEqW+z9Dq8LfZMO1106uvR/XUjfE0PmFsZU8Z
1vFRrIm2i7acTozHiITMCj72lEmEmagIMJX9gMYWHSNIul4/f+YuXX7Qr7JbIm/0cUIxavRhcvoa
Xh2aTltyJWguqzHn8w6hZRwpLBC+yTQnXn6atmJQ68Z0YHQ71skuaaqigQIxh22/RlexpLFoXL/v
RXpBF1IFA3ldnb0Mgqika0ccmEhjYIufyAJhzZMLOSXH1x2eQ9N4d8caKrvDm1oPvd1S9vD0Zja6
EbVZ2kLzaXXfD0GVhB97yfUTenlcYCjN6w7taLAfULMffHFoThdxUKYPAT7TOBW/d+DFexiJAbUX
UfPXxIaVSh5+yVcWa37bHVrVsaSFJmR4xsp8U4WjwPgcBaYBad7QVtqeSYg9ZudV+1kBjfhbl9KC
aNHLsbD7/qE2VJtR08XXkfGauQHVzdXck5GPGTUgO+VSy91lAafYw0yA5lCJczbmAYek5az7KY6K
iH/W7W/mBma3FxJanQsjFRZxh9cck+k4xPJJRuEoe60GzTpOKrRVib/e9PTbrQGv90gARQWr6jxE
//+5pi6D0H2+8CV01G4BsjAelkqECjKDn8bTLoSX3rR98V4bMqSrGRzfUU/kaGL/qhV7DWq7trTV
dRXegkNXt/QdD1YY13B5dklfHD1J99EYSGCc4efF/tlQHvhe9rGJBK4gR9/fqWvnfO8B1bwcArO6
qOdcer4iad/rVL7MajiwX8X4lqM/4hantlWDGHHuPoLpsLQpe6K769KuPXUCVaZtAifEsZfCF400
unaxuN4lpPAR3cL0xqREM5i2v7K3yeRoa80pfSqguIk54/OdlsSKMB0qE+rQJV336kKu3RUdez8d
XSGK/W+7/McOJ4FpdwnO5kClEfuh89CtyEV+lthhS+9+U11rIcQc2RfsRrF4ajA7IjDoAMMQAi+p
QvEDVoGQUVvKUlB3QtX+y32L/vNdolaR7LLaCJerzVySkBLbIgxNb8Fvki83pghERfAQ3TnM/ccx
MS/kvd6nR6EtW6HUUmC9Ko0adu0V7OL+KWkpCwIIVtfBzEDfg81Ue7q1BNj9XLFkYcDH99pZiukF
jlnWdkM5+URnjSKdOBoW2BuDSEaKQ3wl+/4mUTdUPt8+DaeFJtkFlmsknhxe0tcr0ZtbRTs49/Ib
7PYAR+0pQ5zr0UD8ZSJq3/dc94X2enHmiFAfYV+saOuCzCNdkC1FU0E9dQmkOxkWEgi489opumAx
JF6jR0Hb98gczjFs9Ul3ifVxX2peaBi6h+p4qw8MtHYG22ubqaCfjC1qZs8lMKmDc1UtT1xpQk3r
kqAZs/Y8M5nUNcXx+dJYV2H6E7Zuw9YCHNR6tUy1aEnCLvh1I//B1iD3vHS7wcqX97LTOvJ+Kom6
6LzaKpjvrMFBeWqpIpkHggJm3xxujbJFEuUQ/V2+HanAkBPKhXhr81enqZKQNIrWLrJJxyjjtg2K
SL2WjDnDsOtExxMGIu/ROXRbzJvCItm5B/B0Mp7GDBVDVqhNOAH5lmsvU2MWj1CZbdH5JoK9MZ2B
th8p/VBFyVpwTNAdnO07CaVmF4TuDWt915l5juYGU4wze//ovd1wta2xmFIVd00tXD1TuPJOhxM/
RAMbcH2yM7O3SaqB6MEN+smzHTK00O7gFdR+eEjJLs9namafpsYbS0x+5wHXOTzxunsqdSZVUTEa
/B3CuDfl8DNkjv1aNt+EwIxeP6hh/nefOBqC+8ewEsOh7cj/t8csxC9RBpG9EBUvewgjZUHuOSJy
XSp813WZEUvhQ+AlC9sWor5AXVsv8TCA0Yt2ybm17mju9/dePrEHU/lXMVAsaBJ4sGRwpK0KQXyn
9sCKzINP+dd/ziB50w8ecOUnCssPdGiufJSP63fA9Ltlq0N/VnylaP2lAXrx43aYaWVRaunbPedr
qdeblgWNjwG/RUI19dARD3p621yFVOGC944toIR/8sJ8e3SSqmMMXsx9k7meGHNwImb6boRaU+WB
ZQlVxBU8HWTVLAfWexjvgVHVNny0cULd1i1Ny51CNNWnULEBi/fQL9wQiA4W29kx3uCLSV1R3FOn
giF9on82enAV6e3v2OFbxHXXdIBlXbvlctXAc0QS09v74MJYO4Q4Yp1ilZpYUrfQ0mj/ZMss6EoC
vcfdQmYJZN2lc3/S4dFnAVbrvZdSwBOO2n7FDzKhKkkOIiI8kdqgUxn+h4DpHE1+ReWnRIqoSrKy
Zb0pujM0InRCE5hlzw4l8SPLMNyQJgrEIm/BTu+F/hYO2cTx9ojtx17FxVnZDx53tsMXU4Hwuhmz
8wUrwTCD/bkFkLED3GtdFu01JzD+W6yXrrSJDybCTrH/hsKxe+A3Htia5deheXbdRY9Pi/UQ+glx
BiXiPcWWITsbu7aKvZBNwcHa/iPNt9yaSSGrJ1pfNdVXEk74bXLlcPziRr7U5W+4ecJs6nWHlGXA
doQm4CZdJOqTfDfDwZYgOuH9f8E6SG0IHgyI73eQpfd/5TtpfcPmUzobKoK99lHAJhKJHAMN4zpJ
F/V4zN3qPphmnKbxd8Wj7vZgJGhX+ZAQ1RxKXtG92oLzmv/vyh59jpVRscZn6RL5XFfsmAvfedoS
s1Fh/gby/wXnK4nTdMVUEJWdN0/ztJAYSHHLPZSXP0yuJu6HIhirAnFP2/3/1X7FcIXv/+n42Y5u
TLqkEoM3TyLK7HnakMv/hUiTQy4L2RDfoakZ4XxL2qc8J7XZpPT7eHPQuHgpMzfQS3Y7XRNtUJru
+7gONEOjmpUB/JQT6xsTasmlZbCwwEtdVG6UFZIltKTbTh9Jfc1AkRz44sUyheraty8GcREVVioO
7PONTRpSQSSOqqJaUnKrru2QoMcEB3v6USXYfMa9nUvw78S2PkSDhKqTxs2zMIykLCVBACORLYzg
ZVHlWKCFljlzMiUI4/thUAO0fbjmtNzOGNBY4O6S80j95wGqmH5p2i7T3jwswqLq0sBoThlNT/Nc
gzEP1cMUOtmfdpRCUBUclXM3N55FMpk0kWClEY1FDuhU05wHGXjzSHz4Qwm/c1Y74bBUQNCx8bJU
opPz+uKgz3hMVo4PQQ0OJEMTGIMtIMyYG24DYeuzn3sSxI2ZNFP538khzrjuFkGmkRaCZ235Rvix
I85afHQmI8A8Ez6k+u3iq4zYOW0JKdjzWjdijKq06rjv//FoKDjj/KAOLNuumvE7SeFkKya+msH3
DIF/VKBxLtgyQS5qQ3q3wH4UL3PF4jwIBRTxdX2AzTp7g56qoIdVOhwjgdeJJLjZBZshEtxj9xBd
LMFXw5DC0a65OSk54WZy2vIrG0O6dqS1M/uyJwMoxfgJIEOgZsGjSPMXs3SegGU2jUO29+hQAsJU
wzlVEy1i2jw997gQI6XoBT5GfisF7H7GvEcIAcsRaD9+q2bfNUku33WTuAjzWsuwcOutJy8dKvAD
ywINMX0ZWsooo9hbuVSWlnaKCBu9d9TiPBdwzQqigljXYUhd/0fwCkTizPlbsNigh1JF9gLNQoLV
aFx+GnSdqXoX1GH8lWCrtaFlUuFyl5lcY+kzvxfk+3qMRQ3LdjrqMzjvjRq6HjXnG7eA8VHqdEFA
+10qK25g4C7eRJcpgg6SXLELeHqNfLOEV6oxhWzCdOCjRtkFel1vrAFpJjo6jqPWy52gZqj1mStJ
IReGIQUwEwYeX/R7h669SIkh87IunY2/R/rOBA8SE2iG5djrclM8I5cReg/Iuc3s+Q7vq/eqae2z
97v4YNATGsamSRDfCi7oZrYshKbxqMkA57Gffmq9aWU2J/+KOc7LTn/Y/WSpAT2CSynczndAiWtD
+aoqNJLTlAD/skr3KCk5LIlEuJMUyLBIDC9/QgFKFFzqteEiS1EQWu/14HpSqUVUHa6anHucgxYK
KXSJQIym69Zlz5LjmJzcDhD+Nfs+k3tfW2r9keQXBG15Is/v3/KQZtfzoaxUej21TB827eHvrC1d
Lr5it4L+zYZpUdrigi68w7W49f5DXx1mESO7dvapVC5KgGjxPw3XvVxe5rj+NtZHqgsBZAxurg8H
BdbpLhU0S4EqHXRHICJGBFn/IPs2jHOweQJcDIOWeUKWrUgLzR5vcc7Ra6JNewEZ7EQyLP9ZzZCN
7ZzlaFbTTzWn6+kEfPWzs2yqditmKGrMMNQEarWqQI+IvhwgUWDdqnB/DnLM3Zd4xHcuv41PUT19
a7TUOgSw3Oqwjpuh81suBrEkDK+g1F6VNZM05jbkI+T1c0LaVQ2ATIBVPUJRahM/qqk1sJjgrSXB
hQYiGSSj/uZ9wYkco7YVpdWcgpeyiKK5PqJNQhZDZwlxt9SDQ1G3tIzOYB1tutLcQXmDzxB5TXCd
SPd7nKRPG1+rCO1L9ovrnM5oNxuHSFiBCYJ8ZmSiFCpTMpcVDDHA4u5RiQbI9Z8YE2z9zfHmnudQ
4y28KTS71QEOzaXPx4UvLPQ7e2I2Mk0G3N3VWn0gCUEYv1MG9m3m4FKTvbRvCmAq9cLlT/19OCmo
Sz6XNX0GGmCKyNfOUybNRZqnYGR4M97YPKb/pv9ea1RWb3Jb6d1I28GglqkI3dWMMP3kljwuIuqP
Gwcz9DzyeLmnYA76HSqxpffPDq5reuJnAvgBaJMsBsgxmUVsbJiROIGMmxTd4Obk655/i0RrUkeP
NeqEuZuK4OG4PX1hEmqEUYqhn8OJ195edLuPydkmce4BT6qDamHe9DvXfTNgD2v+BnR7vC7oBqag
9MVpZ6W1OpyxH+OM3YahWeB0qWKI1uxpJ8CbatlVm0C99/9Ph0ekW58jpflgNtlfbMyt2LkGQQp0
jE7sF0dbVCUrtU3g2xteAjr7FEarmGJ5ZwlT29bkL4SJyq+q7tsPr1grEYcWMJ7uq5iyG5J95DqZ
wAdOPUCy/fYj1r4+Wt4RYD9r/1G4xELUp+M0aNS9zseASIy0JhOZSbxVdudR7WGkPvYnsRqY2MMB
PKI1uPVL0gvNEKo3WRQgnyApcYTotzlP2qkcSxuj47Ahncgy1nkKnUXeGLZjZ23M3nFIntCaTz1x
5wksydB9f1GTsXXf8WCKtSW6VANY9r1C7zjy3WS+cFPy6gpag/9l2oJ8iJtb2rzN1g879E+mQ3mH
Tgf+RYDPj6qZo504BL1A/v3h0tDismKbt0BZxep61Flagvr/BmLj6i7ldmc4i9DcGrrPFRdMKQ4E
ktWc0stJksr2OcsIVpbZQo28mkW4jEq6p8409/V2oy24l3mSj4odjNbsXwPWGHt0cJRlrc8IcKUh
KzB3TIDumqRVyfkCBl2CPrxTQtxfSIqRGK/qw9pS86X9eaoRz6+zCWy3Xm+ltmqdlxWz00OzZVi/
6fusXRrmwACgcAV1Kpz4lvje+rrPbGZnvg+anE9tvwC8kCfMYBlyMXFPZudspP0CO9C8rBuV5HF/
0y2m40QKVNIsmJ2lMti/PUFumkopzbgR9jBXLvn/iRLkN20TjD3SPLxnDB+eHJgqXgaIw6p4IvW4
ZpJuFVVxevJZG/0hMbplfr41cDFh+EoPJ2hKBlStvMPP8/z1jVWLSbVZBRWlgDQnbYCm5VfdhHEZ
l3838Yp0ZWu+pbbHNCQFc13qln+tOTYA56n1sgi9itBOvLfwnYxPUPrXsVGEzDFYcm6hjOS01Lap
j3cI2+tvN+M3OkbyJ+de0611zcFR8EAuFWocD0bS+81LrcM4oeuHFV97h6npMjVLYoUDA65ky0FD
XnO0qLS1G0Pe7R7uEePBCTpruSP8hf10o/ZJHnMPznQOBQI1FH/EAaCtsYtsSCVqY80vOobz/20H
SH+fdWn+LduD9gz7QJGS/2rX0LhvdJIfiWPjOFpN3JTKIkYzS/qOyfa+0kpWgLraFN+uXh+OAXBK
M24Tfs7vpM0yW5B61cuTH3MYyTlAlkjLoAS5exB01thEmNYv69zM201QhWKCTq+riNTxOrc9z+t5
jxw4lrHmudgJWWznyzGjSNFW0PMa4n9i/RkZpUjwLO4315UbWBKjavKvKpXHpVvQTvBa1iFsPUJ+
d81N4MM/35JIl5tfT0JmCJU7LxHQOSjgqJkCJouSLcuzSfRV5bH8CLq26Oc74gjBSmKwljeGVwbN
+Q6Aea6IogyCVofkmKsomRp2ca+9H50E1xtGcsYPxqg7N16z6/hrpkoES6TyXm+zOXQME7DGA5LF
+W+Sfoe5wd85XY/aXNU80rEuJY11iUr8+IRSg04WYQpYDDqFFFQgdQqo8nGOr1tvmj8P5MVghHcH
h/kIF6cvw4xwDUEoIX9HC9MZChUFbRy2oqJDeHzkXwvfkNS4L10Rvg4+i35Dl6KWaUN1h+HKYQx0
4q6Iv1i7dK2JXStzMvl7Zod5EQiT1AMm+Qd2fvpsS1Dk9oUNAvyOjoVs5jFKx+yeNpiQi2Ap7EfW
CPenHqwFq+UWXNuBSAbgt3nzaa6UKQGbo9jTTQPFI64mHsEtnxihLHaC43kqYFQWn8+SOk7oCL67
EdmxBB2XK3MARMavFzz/9UtraPqNzVZBDkE3WWf9SLwE22ixpCiW2EFrWbIkkLnKBVto6qZxXO1H
reNNIEGcmkY2EnYGFGpJUsAhmrIUamcfTjLWYDcjRX3FHGLDgiIf3LgQmDx8SMkm/DXsgnkOQ18o
elljP0ue3stnhxLZ+FBZiT4WqAgS2tEPqf8H/KBtt07OSinxcfE5UOuNuk35HVvgFRZ/owZzvnvu
3wOSgMxzNM/9cWcwWsVdCaXAcayrHAQj8cxcD/KXFi1KJP+pV3kMsAxtg5qc8VLZBczc6yWtnNXc
0YGC1udvmEjsXDKHpFiUDnjcavJcq60N7uKjhpuMP5+3DT41Drx9t7bNXJ8n6diqiI7f6+OBjEQA
5GuA7QvDf5Tc1TlE1YayeL1/XlPZuOg60ZMaaUxC3P493Ur5yroOo06+bP8eg2IZiXP0FbNPfISb
LNIqFsaEpGuiaF6dQj8B2tyFv6aNFLFhp3eC9Eew94vYHIG4vyfIySdkRZeNynlq7idnVlMztJ//
+iOL2wvyCHyoDwfbBuplg6QxOup2To8LLWcWmwCDlS8qPeGVZ5FWmzgLMOCnoaxSSMW+ncDVgAow
EjcKA/Kw19+X7gKHGR06yylsdMUzEtFT5E9PU2S3BKGiFHCnoHXBCV2K7RVfbMAL+CJJ/oAnK4te
7lf+PbXmw7rUBu3Cu25lbt8dhIFC3pOgALBfBNeXAmOGSzNKGk9JErO9LJKk+lcouu5G0fc4JDk9
XAV52gjxnlxhK10zIJkOv6NDS3UJZuwKk/QrT+1mDEbExw1Y9lsZKF2xHDYW2XQqUqXQmaSrL3Zi
BsoExfgDKRskvg+hDuKK/roJf3aW3YXuAp+vYNCd+v7jEfmZ5d6UrOPKrWznHDHWKqOkKr5b2teh
pZTJlGvkjwaBqsQ7pRulTdUuQcRp9tQdrmbvXQljWJwq1iFhC/P/SBccAq+/IVdmBHLf43E5ersQ
ImkALT+whYIZLYCkR9axC/Mx2X0Ea1PJ4kQIRNOIHCQWBV6rpHFUrUsh7wMVQgEXOCl1Prod7f8v
2o3ivhcSldhtPb0Sj9a9JPfLzTvwJZL1XGqlcqJc5ztgD+daqCV5B8f1tgnuduGqM2Tm7aUjBNwk
XRqlV5RSAxLLxFvrHndqJIzbgdcrvaRf+4B9In07vAhNCvj2kjvU0OR+k26aYNKVHkX/WY6KOmKo
4Z2ZGgbsbhitfnUuC31wUNLGjL5El09tGwUt+oaR2mT5wk90CuKDo00X20PyQ9Cmr1Tdhs+hSLma
G29/r8myfujVWO3LcwH8vwUAaFfiJeQTIt7IZ1wuad9k7+GA3AgfT5QEYqej2750qEKsDCIaMj3p
CE8hncmwId31x8v8nIFgpxxnrHrmEPizj0lX+/0qTDHrw5YG8XGT9Q0xzJvHIg3Bic3dG77GVWbD
QTs/Ss/vOFDylUq8I45VZQ8I+Iuh8BErfAP/0eYsm4dMCFu0/4K4QvfqD8/BJ27hAZ6MOaydpKSj
mlLNBr+YVhEsm8GyTOvd1qvE6MDGuSHxu5aJuyXuueUlUi+zeyL2NNrA/bwOytynHA0t528sR619
J8sLmXMGUtrutmPh+Y0mDCGcK5z4bMDXfN4Uzq3EKeeZZ7+nlvf5lyIJxbezkBm1700AmwqoZ7/O
w87sSAC+9vZVi+18ve7xDSRUK6wR8JmypS83sEzJaCJ0sfJCWkoAQkw95uI673AhFPU3ocB0g2CR
m+2ywCF5CYPf0X8E07XCOIOMsOKX/BOKpfavYG9PQymgKE36pvbmbXkyBNyPHlZ3OGqZgQ6hjcM9
CmogGm4gVzfGJ7TxD+QespD1A9O/evnWtwRfOPtoGZVwCENJ1t0xLxj1OuiIWopnqUCdjmZ4D1u9
apDAl9tkCg9qiiWk11sSo0bCrJeBpXS+vNmG9qMgb7LCaMZQ0nE01W6QAh9DJyJ4ZWu0b8MZi6sG
nTwSQB4UGI0tVxJkIQSrXNtPLNhFLK1SJI43a7FAlSqj2++QuyC1VAXtX4qGdPPo+H7GLYeCafqs
mrOxqbG35EDJ9v7cpt+/xDISzvv6NHSKfo/1C1bj5CAsUUU+IO9b7rTd0FN7ITKvhwxIOZUv1B7y
3S/Gk6pUnHjZwH/QzLe/ydTAnQ4VrAa9pu+z5Caq8OP6oWqM+MT9wtK2kxE5bceRqQTj8c9gp9gl
F8YaU0w8vxHpELAWD9o0mlCNUsysnYHFb8UOgfLs3ROXzHmQ7hkXtYsz8QwKdG90kPOiJ4O4VQcN
oLL6QNMaoPLp0iAxm3tW9HaEHuwKmn21H4kY056PR5TaoXWV1bGPcMdt9qhcQ5i/I+LHlC0XvTZK
ayqtwfieSAvxZmh4yZrdFsN0bm7O+CFLS6ckp2SzGeDO5rXg7+GLxm2WemIqga5Ntvre4w81Otj3
UAghf1UznSzJWn+PVOSI/n+5oBUWvOz+Ek6hMsJddZIVw2cBjYEE3g46XEjbAxjvFLwOM9UgetpY
FvFZUf/S8VBdRQA/pgzKOxaduM8T0p5SAsqACPgQDWsTBL+grtlKC6mQgPL/YGoglj1qJOuvw+5n
cr93O4As1PsWwW+3BZTwWo+3PkW8pWRtyCROwe4n6RFBSB7Cfv2j4ngSAsfmB1uS1ry/NGRQQua7
+V9Wc7ghWvFBGTSX8uRjP6KW4/ga7eUfwpgeulebWew4eOV+Ozf95Mv3iVJdXsLq+8DyH9A/NtWU
4Dw0/Hns5mPRipX6GBZHP7ZGYb9DjesC8VH+l+5e2fFCsyEay+PKClJZwFuPOQx3rzKI/t2Pdbyz
TLUIN19Wg7zMkIzlSrlxyZ2s5F2IGazHEnfQIHaIr2KhHhMZB1GHNe/yNfbffqtgD95VlTXUqa5V
0lx0mrS4AlCQtrzzuX1efOhN17BSIljxsiOMGKCGlbRVDwoOj6YbjY3mU+dFR3W7HVTyCW7AxLQs
pNuOOlVQfNBi602ND76JDb72HuLNuxotiUpNEjfh+70Pu/ub/wUE9iKtKysTaUYOfXwaFbzzen6X
+pAxA3oDnkUhMS7Ig9SFuul7+Dp2wiombvbH8rTEqzM0GeKkNeolNBDcGhnqp6OgXdbQucsSRDWd
KEsT7lprZB504BoESMpFT2cPQ12oCbaQQbpk8ct7C7dTMCbdQ/1Vhmf0XUUXeHPTDPGjPr+oMoYd
BZyuaQ2ox0cJhQDPOQRFkm09uwzY4Rvgzym+KH9WHSCjOIjnjw8XwGrMfzq/BEomuQtBD9E5x52Q
FTgVTp31KxIc3ZRUfIgj2f135GkMEY8+ZMo7RYF9CSGTNUeuI+uf+OMrWbfZN0nb454Vy5NzAwTM
wqfDyV+Qr9NINOeHkeoScaVFG9oBNRjZGCt3ecAyGCpteCJtFa2y55kVjQqSpxIZxw+qvgG2w9Fo
2UbvyHQfozwXjKnJlxyKLJYkh3BtTSTGhyfLUuCHkO6cu8UbU+eaP3JZC427Yaj0xJZHED5qq/xE
3IGDZAmtaldJ5KFnqIkZ3kgv0O9N1kxehMdtcICp5Qj5uaI1W3dYR9LVTsYGe6BRZThgey+ZgkB2
UXm52BQJU9QVOqZOR2cMhs29MHv0Ii2X4dQcrCVmlBMQ1EMl90BnqgLwL59DSR0QdMTf9Vxe/5ev
Q2UMPTmtB0GP91WF+9SPGrbUatIJlj/GyroNPONU7uXOFs3rUSlbIBQ7+ClmUsRpU3ZAmzh2/P4Z
JheG1hI8r+jkDGXNNF0QvxEt6b7+pjGTWEw2egaSqhaBDcFeXcSMOi7djidBj9HWFLnpJXq9EfdD
aqxVsDA4T2aB+5f92LLBNPQoYtFUGEMVPsr6W9mVsSOMltzcApG8/yicC1h5jivoVSsF+ihmXB86
xu5/A56t9UAmP0e2Zwh2msXQCTWo+uDloEUWw3MjZK5QJ8rwgYun94t0qSkUcMd8w6U4tBFQWa3e
9NCJ/66rTZOF229xEagtUbXKuYCs+WAxXLkVNLeZUp5t811yOp4QcVGgJQOFC38SvAU+X/CY/7ml
uOIIcM0Jt4Ru5zwfPut5ZxfTLPi4dkIhU52Jh1/j9EkdwSnLevlEUnbAQi8MC+R1HnOeAZWBQLRZ
8pw8iI5YIP5pZIvIiKk+8ShmIpgNOEt7n3HviIPQ7Rs9vRV+1L2pqILn/KhhGUGfg8o6oDJ060bt
hbE96/X0n+BoLpI/lNjVRK16wDYLxttp3HBquCeoPAVBxaWothAiEjZFZvjl+OJM/Ga7HdVW9y6g
y1xtpKKJSeLAji9cDyRogwHqd4/6T/EG5lbcGPxFH59+ofDEJV2L1U3YY/iEhG7qzBsbvHGfcwAK
mG6fs2tkSEhzAWvC0un3tNrBydqc+WUturCBTzvpzYpTaGNI/9crwhZEavUIFvnGIgavcDv7zvZU
DyS5dKPcbReZKSqixzbubjoJC4mWcyfE4qJ3KbY5vQq7RFTsBPmJ6wtYWZKc6PUwx9qqW+B/haot
Ele9cPE1vS/Kaj/laUah0v2aZzxaaXztkPMzbq/tbfK47RsVE/5+rpMfN+VSQnsWqjAj94wP4pIs
ARCutAZJOFuoOUIpsgBkxmBx+X5A68OrZki8ZC7rK2Ocu1beUGioWH+rc6NRGvuzCTTPxndpAVW6
KYkZ+IIMyQoe7+NzzLxmSsGI56P39NwQ/KBLRp/zJIwiJRgxI6UTx6NWBoH9ZvotZ0XZb5pil2Dp
1BGUrM0NrpO2KEsrSNIZ22y54ezMNdR5YKSsBlIDkoCfj4Q3gIp+XWQmFiMdvSLl+o4UEsOk7RGT
YWeAdrH9MURI2hNF3bldUb7kc87eju+aX40Hoy/GG0sf96mwA5rOX/vFFo1U0/LhlZPG3WvwJLgx
TffnefDQSJrhkIZndrWlDrU1hFBWkVrnvXC0cAaYdlDskWjQZICxutDzCdl3urVihOL7vXwf0Jpq
h4mEYiZpOjt0/vYnHNHJNqxGPxcJfzkNAV0kzyHE2mvrGeX17C8AvKc6lFsoXQro/XoSqlg+NJsg
dtDypMN4wLxDrfW8TG7fUKGMm+EB8P5KnOWax39PDkvv7HCVvmQed4WfqbzbhVAyGP/f2K2g3sq+
OrUEmd/ZmJa+dd2WmyxeW15ZKG/+4YjHcxup36wBa/0fyFpYrUsynr5Zjgw6mXhvHRU/zfg2rQeq
z8DDYy4wX1aqIy5hNmcQjqdGoClHNBchD8JL0YfhKV1KGvu+qqiwLzyF4jKgpvzo30fpQvsVF+bR
OH0XleG7AfU5q/xAI/W7uBpU5MiM2RjbgRT+UuX7kUBEED2g92XldX3A77TqjUpRqEShR768KROF
jihL6P02dco6NIWjyqLci67/pO8IYRmLHYgc+yCwlJ4LilUB89X4M0/wsoYHo/jFW4w9NR23UVa1
jZFIyvJsZZav2si/Z7qLnRNkevY0nY4+lwl2csQ+2D160fOLfMk+5Zp5cvxiMmGO1WWxoy53tOfJ
DVE1CripIE3kroel5FdIcDVOYItb40pU3sr8Nop8vAlOHG4aXHhiiVtKnd/1hlJnp3B3v6QQ9LZg
hyyWNzGNOZP1tY+bW66xCbwdiJsBuXnNIMuKgl3CpBIkxFEAhLGtnTjTJ+e5WUwW/85OYUit7JfK
FYKrwGLLF0/4aXPa08B6/LmQXh/MqMz5sO8CiELPFEEM2ldwXQlnYev4m2mdZKaXXLqEKITz0TMA
we2Q0OIdpvWFTp5nRTsnlmTd90qWtOERNmPDwVVFWpd744iRvbhpy7z9Ma1RnglSYs1rL7Ae3svu
ya0exjiDsLRbJbL1AxvwsJvANLgfSBlLc4/r8ewk9qLDYU1B4pLHC796fcFC+J5WX58cf3BTzN1b
EZCfR8JZujddxvWqCHhpCZPI3pfObdueiLFixyivFyi0vwA+3qOZu58acr8PMIgHSp88fhIxVst2
kfesQ5gKwyyzDqWER/urG1ZDhOWRXplWFl3bj5cpa4kDKw8YA61f2XKTCu156847U7iybD6UGmXW
Ev1OzjCvbdbiyaObtvGLpRBUACrjdaGjHFz2sHvwEAYCtTbfxlEbXH/mgzT2VhOPwPLII+UoDXuU
lqJWqYvyLRx5kUsCVsBfh0+TBsJBUBD87Hp1BqxK4z9C5HGTS0v9OL89sWfg0VX4yrCZgLFThRB5
idLLtMDgwp+QUDF9yNGcCf3R5IjHXjZJhPYkI3hyYwY/bZGuRuCWnjzrKOS7eByAPr81T4iOEiSL
v3TkEGS6QfdW0ibAwm1XNoX1Vw1+IdaMc5lKUASKP/6AuuoqZY+vIvRMNYMffqfcbVAEx/mk4gk6
sONZ+WTZT00Q+/unZYD9LD6iOkwZ9nZpP0CfgL+1agGmVOjbLHAZXOj/FeAMpu6nnwGAERkaHUrM
kXXD6nYFhb2bi7vViezm8TFkN5/C0pGSiKfmq0lMsxUFkN7tLhhTfQo4+WSGcgmQNMOp/+MVvu/b
UfwsIPwYWOsD7VaXHR4Jof46rM1+Iu19QLXmh4iNXN+hlww5Cv69g+XtdlPqeMuqFDSuPSLhjhts
4/WEpRqTnC+1W0FnL/UT+ZgA2kyK063fc/8BCMO+6la+EUqAi0SPWAhI2wVvaxz3ww5SAoNDdcMg
6KKkoov1oD3B8phz4SV/PV3OubCt5WAbuBSJQeB+vWaoUXVTQulmMOTYxgBllSOMGvKu2mfsU3uS
JTqr10yaHIUllIHZ26rlgzBYLHA3ZiLzFcZBADI5wEIk7TO33IvRJKkm/A5Uteohu3BYa3h8X8cL
5qJM7702tL+T97ImfQSOLftEQdfN1x3pdBF0Y17zvhEJgMQk3D9oZxu4CCbhLEzrG5IAF+hz8RTQ
bMmBYLYvOXMlcuMbc9Bo13dub+T1rNac3oQecSlQIskMZTydtlXeKmSiXL2FXUry6mKCPfOGmJID
zxQOaTN0scYD8nLlxvlkupA2QAo813cK4ng18fXYZshjIxYzwNQJMJV1dmj6nCX8/QspyRSMqnir
z/rI1bxvlSNOFMiuHH89dG87624GhifayuZkVVDrFi1E8h2AHobLLNvhNYeFaQxjTDS3vMceeoAa
0NlOmi710KZ6w8DbmgG1pe760DJy6b9dHnmnzMamX5MmzGXRXSF7yEMmKXl5Ylo+y+Tyz3bq4tfU
JnClu0shOE/NZ15+4UatJd+C/iohpFUSIf+QeJEf+qOpX3E2QgV+E5Yf1km3y19WvSI9PChl0pg3
TGXtTntTWalSBnr9oQnQIPlIrXJHGfBC9Nwty/DPsFOG//a612jTVnLgHlMOvN5JGJfci/gW2ltm
cYqe6xSosIePGfspa3g65kP1hjYC9fUWTahrzxn/za+p0MAjqGu+sr5rdR8HMtNrlbxVV1fv7gDf
uLlLQu2XWsqaB/gxaCCWmLCejECe3wcmv3Dqq7SITanNuNtqqhUVHXUoBK1d2k9JbeozeLDXa8ZW
4SaeH4Tkw7mcgpiz8cyFCSHPQnVaiXB6uVrlgOZi8ZY5r20uMNVeFyXJAnwGu8KcDlvlaMmkHbut
+pDeNw0kVlTSvVKQblJxlavduEwtWO3Js5PJ8hB1WPGk3+bWDnNkRM+25yixFhKN2/auq/kHtWbd
HMFFT6xX/7vfUEgEVuBz58LSwCy1iiW6rWwZomxVcV3GTacL5DTUgSDIH175iuGcBO6l8cUlfJb7
EyPXSZyP7EOPZXkOMWUy14XFBHCLXQFlapUiIS1DuDYpOBvWvsqYwPoIJDQsWfnhBCt8nygYvB+k
f61oc+mteIpwjQRGRSBJaxg3klDXRvEC44+GU3wwgp6ueGb5KrrqhrtYez9P5GaltAE8Y4zLkw7F
UwTubtg1fc+3IrRwRE35FDVhuz3qoQ7Bvm78MfZWCvzEr/Ib9kQada0B+TBdMlM3kradwfhDq0QK
AuLTaamJ7glH2bstrWY5o3uoPBk99HYerDNV6/PZ0fpl+sg1e4pujWbYlol7sWgb8kupyGNrz9Mn
8XL8B5GY7K2qtztOXJ2izN3naW5y5AHPBcF8dl2b+2mbcKc6RrSZso4C4gcAftId2IqEzOze6DJB
fp5TPTA12qWqHbG5l8thiz5YTdVouRgwMNPpIWjZA8bu3gxRf9IWZSoctWwvXHCbUMEL6JXr8eDr
H3sbw+SLkAXB9cQv63TgHi56QvRVbGXfQ6oeppK60JPD3xovz+i0fmOcJ9aohWaT1kRR/rdKp+S3
cosulc6MLKBo3bUqeNovGrkfHd/3xhZlQmwmFaEQHAeWF2alPmXmDL3I/VYCZ42B8WcFM6Bth1w8
NVQf5S5Cox274ADjxTbENPd1VAkQUdyrx1qRHpP8IPvFS/i2fZQsW52MXeamEvJvPxQgy6EKXurs
MninSJUA6Ex2iF70ocNHSR2qncxwIn7wtMPUH+vEjUMZcnSPTlV9E9YaGtWIe9vuC9ZNAptsMGli
iIAQ4IQxt5330Mv0qCQ1RxTiUTenxHn5wnmAGMt/gfU4abaYt2i1eCaPYQxyybHUzSpor8qNDCwH
kgukyVrb19nvvYaV0Xld1NpXFHGGsLl/sXRh50aL05v8l6Xzj1AiCU4bJy/3iHTJy2H4JGERYwjW
nBQZSNtTI+LdKZUus4OOuK02oNJszspxuwPwoDoKfbZvJWlQEQiJuDzukZcSEWyPFJZvuzoJwURt
FXPE+JnYncB0QGWI4wof3G2jEbKH2YTKoOyOezWwISPI9lIztCU/g5IdaZ4i8C3yhoM85hdUvKWC
YVNjOegD+URR69xV9fRxgebnPJhMnrtNpEItB8/u2KXwMstKJdAxPXVukvKtMcTI/CSSnuEmBQ03
grTIf2Zzh6cXc+gJ4jTeq1M+/27R4+TwmAbTsAaFDpezb07ZjmSMdtajhbk/0HfRlYX2Q7ENsany
csIy34Pd1cktblQA+uO4SuOTnm0rilA2d4iRjovAdWiRjZ2YOmOv8QC+PPg1r4PxuCYHcdWOguIr
nL7aYdPqUR1xh3ZGq4mm/UWXY8bQadylAaHQ7WN6YVODlDFEdI5DZCCNIn+eYNnVbNsRmLa+qGjS
0+6rCM4+AK1vP+sktZiXwCeeEWwr/DHmkl7Wyy2tSxyrLpDuNyJ+ezneCOLvYB9swXn6tCtQ5rHh
GDoOrtMnbINt3rXEwjso4J2ENQJkNhLDRhChfzptPKDR54eJYZ9k5pIc0ypUpIqBJRPmkcecL8PM
BOZyr5SvJMF8e3srYTs2/wMqGTbmkqh1HBN1P+LSBHzWS44IbJxYSKjYlj+I5OMMF0blwVxR0OHc
VvtAtdawPa6d4d9SmSSpf9+SJ9c2RI16mG2E2gIQWGwfjnNK8rPUqvcl7TT87PGNJdMjoerBUZ3m
8RU1BFXik0NdhVT5wjF/FaYhkGImKYjBhon8peXMgAiX7ox3Dc2xDYdb9BuCOhPpuvo+XTxrR2Fs
acqFTxFHaTwvaKw9KGL5AjqqrFikGaX6480CFO0t9kNQwmEYaHfTc2ac6t6jKleAXYGeOIY2w1Bn
UN7ns5E5GdXCHS95WZVqpOPQOL1SCig49Zcj2/irfN9VnLn6T5pN13MALhQV8EBx1z3LIevz8LtA
yGLbScKpn0KSxKvGPGDFfMqduRooNCdKCTvY8JueDTX48vP7Xq3U+Zi/w6yTB+H9Pxez6r5i+dM2
mBs0I2tuxhxGRHcT4Se5b8CYoSFufB/pg8cUPSYvpmjUXye+eH5Llgqr2dUe+kROkFaii41Hnq6t
66g9CyWUmQHoH07q+8KDLomgski8nBW5Q3fyApQPC7G6JrXENhjaYjzrfeSlwwPgxUFBuc7gjD50
UNwv4gEfkp/OLUtzSak2jGOi39MT4HQOxwKF4tNkSQRmVvmRf3FM5Bwc/XY4fuBkBTI6+ehhoObI
BlXMJqj1AfTMesUMV23nc+IUTBnQCsZy2t8zcxS7b7bDT5ok3e9KGAcGsGxetSR0GF7HE1iIyvHR
+p3KLLql1hbrbQtreu+e8jSY6EH/a+ogC3ddzuHimxPZat9Nh0M39xlrpiA5exeGVDgDYmEZCvAM
UEC+YG28JFjpE7tnD+Il45zj83laU5t1i3MfmtnvFT9D8+adhVpiL8KJ3xD332Ots4iwEhzQxW/E
UktRGJN439AHmQjT6/gySywzQaCn0slBvTJ3LN+bCUjZmYThUinNPBsFREhUVHP06VqzlsC7qOkx
SfHpdlERQCTCb4NunaQGnSu/BTF5rNtIG1fg/+I8O3hOSSRKz4AEukIgtKJyx90Ah13INKIc7y5y
urUlnJGkAz8d49K0WMkO72HRwuYS5wKJ2SsORiTwjexKcJyS/674XL/bnIP/BFfXk77dGbT/1j+T
v9HaMyvUcwfrvJDV6CxGIBsL3vyRDcBsfnjKJO7wY6bTQwecpz9GjBQorc9GG+TWNM2EI8xd1U/9
VNN9GdaE0kTzYVPJQFEPIj+ilztp2PFdvlModvkFJLaX5m8XHjJ56pUAmkepSXnbfPls1nuBKv93
FPJONkYaI0yxf9maS/UbLVXNvyfZ1wFQxZoPk73+JFzdP7eTO3OnefzKl+SIL0YjgCIfxjZ6duHR
Ll+o5XcOXZccXpoPg0Vlwj93DlRIhDLLjcgTtnFvDmxXidRm5u7bIM3NDFHGS0rBR7rWQzZ+wFMj
YFXJBFOtWUI0NeBUGnNrPv0WT1u2ZgVzdHP6fIyP7Zun6Bz9CX8j3M2S2vwjQd7ubc1ShsIN99q5
aN3Zo+je55UsU6aeCil+8YSmdMxwPTKlfw0OdVLRYfolK7wcdHKmiwPekSbgiJ7ZJU95+avOx0TF
rur3U9TtTTGWnrbKCCjWoEUbQLIPyh/9PiJ5pWSt1vINp3Da8DYgh/ZEhHCs3+DYSJJ8HOCo/KU0
fTyz6M2bS5goh1z6U259mBzKYyFgCX4puGO8aLvD9nJ0tcbh0UKG3ycNYOK2TN1T0gOaOq+mdq5p
fZOGtl8+Hi90BWoe13Cr07kH73D0oI53gp/C7kujorBg5IV1UCjXCiKwTx+Z6oB9+Xbggs5oQiP3
RI/jUnKPJkAExdnFcOGubE0xfIVoWpummm+X5N7Ce76uCCkOt2PjAd7s/vH+TqN+pa7JJLaNY1PX
Ydq2F/AVvF4AzEgJ7xgRxw9cKk43xcq7L4H1MWf0hcCcixzujKajgKBm6k3rryMXLijmYExJ1j+x
InyZ5H8yFTgSrAN+qRjFNhe/PFMfoM7WKE2YomKkPailddE9QdBpoykDY2BO1XxaPYiKlB8UdMFJ
38Xkq7ZymMcH93ggJUACHOUwfL18JQrLCM43lc6Rt5GLiVwmZF9wBZdAxctSnqpIau0+jR0Pio3s
oktSKh+HMYvw1WRDF147IgwVDReVUqgs1JPs9yjNd4OdJEFp56ONfijsq0gU80/KSBjkCR9xqJlx
P2xtIIU96Y9xoDXmoZJGHKgFuKvGeUPF0pUJLdr7Rr5yH5l5nVsf1//OP5vc5gVrXO9apx/lA8SA
c53IvcZ+cPtEC2CmwTPiPZAMV1SrX9WlbCZv0ZvZhfJ/lHs04a/ucZy4qTz8MyceBLXIrSMzNDki
FTWbEMrmJbCAIL/XZJVgZ3+C/S8qQMye0qlfdlWo3pb32IXuJ3xsbRTYrBM7FaBSRZ603Cn4dr93
+x/XZTUvVdGctpselENc/IFWtZmIyNE6GhAnIpNGGllZ4VtbkkSjgV3+8iJCFEuv9uEXIL4yGuro
YyKaQmotgjVGImWtkchDl+7GgWjGlzro4bxH/d4Q5w1sVkxxRimBLHSokD2R5D/ABOIIIfr1s+p/
WIEqkDerKKFHCvfs+kZHhV3vHFzsAhA6rc4mnFJz4vYg5cS7mB8OJ5PUTYek8jqYv1Bf3iXn12z/
1VPBvglYZOhePGX4PsCxgVXNsjPmO5QPnP+Sc/RXR+h/K+94oVPKbTfwbZUjr6sBKSBTHsYwk7/d
uzenix5FS16VI/DhKFYSeCfGvLZM64MLo7Dt8WuwZNBcu6tRlAEIPLmbwRHiy98sNOu7Oj08JCRb
k6f9g4ZOsfJi8vUbHpP0oFgXI890/4envVkaeRPR8ss5lyxdVMjtXrkxZml4e9uDoe3ujgwU/qG9
GVPVywaSIurSd4B3Rci/kehWoDsNx0w9MonwbCif6DqnfN6f4QHxxJih578QV6FByqrr4uex/uat
rkwz11/zTN2fDh5X2sxAx+TOMDXCXFdPsxKzOXSrN504CAM49EM0iU5qiJBxCseutueoFQMr3EkO
l3d/LGjSLXcIQx5pFjTYJh4uwYt72vv2Hl3K5DoZquKdczB3MZt1UjPd9HDUTYXtMAebFP8lgtx1
QcrRVzI3Oz6mzxTdlORJr+ByFSivLoOWncyVLrHJhwjJLI81fhDSTet24FF4tjJ63yDEcIFCAXOv
HZJzPYHZmROSmaFR0BbfL2bY2CXoHIfYh70WwsXQxK9AaXm4kOAvDnrLEdb1WbPl/JqwdEI92sTF
HjLe6egGgVsw2F1IL8cwZwVOeE0h6OzSzc1s4YunMhxC3c7+5tSfn4pKSCto8yzx/gVn65+alQ71
04BzqCC2J3t4bRZyNUACwNXGAsTxtyQPacQpN9MfAONExpb7F3oq3ojydZ4laHF10g0ObJx1suSP
fjM93M6zxOB/BvGI+6XU5K1Z2iN6zRXx5xDSd4TIOm4Zft+e1BU9EXnrKX0PN4lP2q1URiDHP6f2
qmTE0BurINdv6vgqVnzrM8qDuQSNZu5cF81npeDl6X4bqsblFczmq1PtGcLXruLV+UqwD76JHPzq
2wNM9ypHYCtZXaChr5vgWDMUTNcJTMFHmgS27f57Eg7Xf/DAJhK7hu8kElWAKXgEL85l4hhCQuu3
7T3Gcimp49j1HSUSaX2ilAHs9ZIM7tx+vNWa74TGJoyd0+E/KZgkVU0GZpbTN5lxJNQC2fVyFO6t
8+7YY44RQx1j8bMVC7lzVDjCFCFkMFz3BSo3PgC6ZVVivKOiJnKwlS/OLmdVY/DPl3+Ad+DRmgMK
1S+HGpBOf8EUNcqA0o5z8X64A0m2wJv1aYSMu4QMMI9RD2onRxRjgK0Mbs4FsqgGj87Eo15YlmNy
QplB0F0xRcRzNOiYdqGmGqiW19V70whRHpq+Rhy3pLtFRJxkIck5CN2tDrECyNiwO1uxDgOlvsbD
lg3mDL04vspgQVDekRdCn0uOEuT5dBCFuK3EHb4CCXu8gukhklKDJNYlvfK1rYCN2U+sWqigisj2
mafMor08rcLGxckZbY2JIQAfeFiUUM7ICa/oxk4eIWxPXcjSKxPO9Wp5Re3ori4Xdm4E3eeTl01M
WeLbPMiQm8DCIDWlcfrxh2VJmkBWid4beRxGDx8mx65k1SNsYb6E0q6rpkrWoKHEog1tJJ/Fhnjb
Cjg6dtiMvWcK2E30pUdDMquSpTulhPaF6ekyuK65+MwFYmUr85tTJFV2MXqyRL8YGPJ8veyn5+1B
QQEhCuL2z70sQA5f8TwdyCfy9UmqzHn3dx3DXswMzn6yntNvC1H/AbDMSltz24V2MUFBPuRlMl1m
I0wcUNIzphwW5/LJAhoS3EhwCdexPzo+YFkbyKzYIoMRf7kESRNbgP+Q9KwLwn4KD/87c+5tQUB8
vJ1J1I8GLVK4wZNoiLycJUzbSqY/Rzkl8R/AUtLrGha7b7DK0XvZxDoo+o0oQTTXh0fXI+oNI+FW
mOO5jr5tiNumhLiRcq/dLCAXoHtZI/5zAKPMpZIKAmiVaK/IdxF+ghI69UlmnJ6ChmZ2uG5rQl8O
EnEyQNj3RiAvnLeBRmTgQ/Pb2Q/Igo8hqBYMJP8NjUG6x2sNYvQjGU1xGmtNADdP0LuSYlXufuMG
K8eSIdg84Ca37fgwkTMJrQNImruCmeJkpZ4t50X+imSfhB2D8Fas3X2Mln5OO48SrsPMbYSBQ1hv
efkDF94HJNk05BOlRAGo1zStkrXo/QinLr24CYjJzUUBOuK31iAbdW1SwjhUDEXqrBZD6e3EEjcP
1P9XNY/rVs4kyefsdLqVHABvXPzUmVGzwjcXdKyhqDPULkAZLzJT2Nub2ZyWLKylOaaAzGIKvxzF
tWVMCHMqAi7PvUes2f7YSTOvMxy3/DL9rWJMKUahe8oqhJ/ZJ+z1/ZUbK47Tt98Of3nbdkRX0HkT
I3t5PfvZwLIrF4QzV3zlcAsBrxHS5VrsoSS8FlwH/pK6OVjWncEgLoEG8KqUWwKqI7sbWXvJh1UV
bM5UBvc/PtQicR192pR8SOGCf4XZHk6E9cYNLvgKVNx7DVWfogv6Ww606uSwRmhvrXJrX6r6LXRo
1u+fZvAS0FW3b3ifRxjDc27/5qvJ+l6A50E/PIYkGsU+FVOzDKX+Bna0pTSLK5OkzgI8EtZwIpj4
nlzPIiRfVH5CsrNWXIFnAwx726ZayhjlaAeP9llS5cowjt4HFaIFvEmMcMu5ZlCAOtaz7/b6+5fi
ZroZ7hTy50Ef8weX+YLJvtM4wlfAmOeVwcY4p9QNP2V9jhw7m1J0+kS2iy5YhHzBfzqMsgODlE54
RDDw5NPtKIGg6ysJ4ojJhmSg7/BIAL4gvr/vpNtAoyjPUNYCCoi1DWWU7qZjmk/L1FTKh4WpaeQq
vtUkeN7qyRwW1S0nOh0aekdmcZSZygUnnFKuEXPpAhn5WtPV3O8AaxcW4nMojDLXXru0lq4RupYC
DYehoqvheUXSXuq9UY0td8pAadQe5wYKaeStGGJ6Odv2nxlJGv8hWnhXlnrCQ5ywTWhNczPPY30P
AA95lxyQw4fGmSgx2A0lku9THpjhxosCos4/3kHUv2AWHS+H3Io1YEQjOEMIinNjzIgQTy/G8yWw
LwxkT9oYDV8lG1Tg2u/H11RjxaNFMke5mggJ13sEq87I+QfH544Na9yC6GPilxy7lKu6//HH57JP
1AG3QDJIwlRtVmtNxeWTJKEjgCYgvma0/ksJtH848fCADB6N10QT9+BApIYm8qEUoYMpDIaIGbf8
IEy2yzL+C9mHqim6TYH5Ox1ps0ojE5pj4p15e1fnBoLGqzFiGW43RqWFp6gqUi6H3H5HsW4bqy4b
/ESgKcgNpLZ+Yf+lOkaTnO5pXi0kYqd4cBD6ZhgWTAeyB1ocY2Y8DWST/eQorBj7gKfFAxyDB+8k
pa7XUQIYe9hpt63cw7d4qjD0yYaUjAt+JJOSzLgNmM7CIdPt6esKeYwCyE1eDkp0WfnHmS8s6gc2
YHMQek9ySD6/ZyDtMJ1dVq0t0X3j1/vLawHWc5O6MaUcduzPrnr4W6FaSAJBQw2VqoOi45FlPMX/
f8Nl0KRomLjGF1hCJp2y/6GvHStCXlnLQ9G0dly+F8QGGzShy3BMWXPmI5HRPvLdcgNj3AilCXTD
A73WkfPFDezkcJyRV5L8M6jcuriMduQTqi79sZMZqLf+Hd3XiiHZ/tOCQtbLJvRFdy7YJYdW8ozl
hetAjF2tqb3GTSn3kJ/7FHTKiyHOAtreSD8dCv8gwbC/Kipo8OPyTz62BRgIF18ydI3Y67kSDuCj
DLxP3i5LL9SQFhDcNjIR855smVCZkpm6WcK6+25o1mSl32t/E5Fc9pFNMw0aPShkdDt0byDTdE2T
DIim/rFporKmTfKMaUFgqKy8NHR2RM3Z8zVDQEdLgyUAB/4i4wCHgJzHx6oCTFgjS7C7YJTvHMig
55izfQD5Whd7krwEdZx0cfwoq/FAXl/aczjwEGiG79fYxvUejy7qCqwnU3rXEsf5gK8ARWG+CeYi
HI9OYQOEvz8DYbDWGq5xc6BBvJKnYs1SqP4ouZHZwTei3xTE+oW7aj7OUIhfdlMWO1hZEoE1ml2D
Xa0SCu7UUypK2cFFauhHo8zNNfm9uhw0vEdreAUs/f5ohJDbohxGSueY7d5i7tOVw4cfp6oShXJ7
hCaa4eL9/MyMG/KL0gkDlvJQk0WG+JlbigQJB5B702oI/sMtX0a5o+nq72OcZiw2ILtZpYyrmxD0
Vf/XpCkvIL6/wTTsycxDSaQiUUMKQjZhy/jRaNeaawUz8E8ngFsb9eb9ySZg6Zeke02SDBlKKEJr
ygAoukBsY9U9+2Tyz8nTmH5VDSeormGUFghd3rV4/y5IDxt6Iksm0U0nQo1joQV1LdmTU4eLz0jh
lzGnDxQW6Fcqq1AssgPcLz2dldynK+D1RsCYCPEyiIOvN2/HYhHSKaTfHqufin+tSxhmCg+pN6Bx
b4fh2trXrm4EuT8aXJYl7B1yTgBG9gAp8MJpiMXPfTrTyMlbVdutgR1Tw9UqNwS9UgiIuANxn+qB
axVDe+CTtOWieHqRzbPJbKRdBijwa5PpesWPhaT0D7pqQ6RTScxfoGXDuGeMq5izhvpJAM0MDDaM
Uy1r0qlnYuG9HfMx5W4w756XL6ADMPRqFTkWM7HtmLhyfsw0ta2y6ORxpyqljISap2/681rLwMCa
ILAnjJNGxPnQ+6Y5FgU5eAIW/Cut94P08dVlEqNTBJaUFG4DiTVyYKbHE16UwJ/kYZH6S9Pl9j4D
PTDIWSZ6x5Hm5q5MqeHcXDzUzCHrTgGJVAZaB/8oQSK2zWjd131yqxtf/+gFeL/FzGlWCJYdVdFn
84ymc3CjyiwSvv4EkyxAHVCxHLKGqVs9EGzpPrAr9oObeFh4USIGtE27PJ9veU+Jra1CzAnhHRgd
ZBmdYIiu415TkuL0oU5QiEDJbXlApGaRXDjehjdRzibnTSP2V/ODgz7j4oHd/4Ee9dq778mpZQTE
TmOP4y89Yq89YDzneFL0E/pCYtPH2apzX7ElzUvUoGc+VKKmGzlJO6lE0ljvcVbRI1GAJRfGGJNp
cpc0lhRLcOv0R8bd/+yn1xRML9Lbs+ZsNKS9JS+pSUYnOPTobXDl9soU/v2AYJ3U0d4Jn/enpdJc
9SBxwVGcrbUl3XuGoB8SUjmb2OFupcj8J5MbGOShG0D2cerxFXpgTJXoWQI5gHc65J2Rauzj4Uyh
c87KsJ2sTgzjzQ9YByAAuUlm0lNkkz8y4JCJmPvK3YKJopSguxxhbkuqqWNW645KgTv+WHuNuUeU
GaaFAdfZJIXDk2nfAFjUnHwmwbKcit8JDFofi3OduiYH3WaYeE57vlFVOuNT5RbqtxGh2veDFJ/f
lu+WFWlMo1VVLwvdIHIp2mrLSnnMeSyAzHDTRmd0tiJidEJnMH893hkk+yE7phTVLgmq7IhmX3Q2
FmWFo/w/tT4SCYLPTh2/WP3F7AGZHaLNvd9sphYdhX25jgsKOicN1vVRjXBi1SylmVTt7gUy1LHR
LwH7E/k3PlwPkEqY3C5Tn0lsu+RWEQjECu/6UzUoZHggv4/8gCpBJtYFH3JFQtasTPiJUsB+asIv
RUdKuSDx17+geXMraxvdgeDsVN7kwWQ5tJJv7hG/qBNUzP1H/l6yvmi4d0vYO+35VzHwMg6LTL9c
LCWFGoaEg6XbHLixikUaT1flqbnUmxau5mCGuKbkIYNARPFTejanuW+FtuElsr8l4EY0fR3Jf+oO
yGyXAN/ucw91x9Jl/ZPngTnBidLnCFGBUa2yeuiJgfrLYzPzew5KV/nD3w9oazxDn1AX6Bx8RJf+
8Tw862mrgWeSW1DNANbZ85KW4sue10fpPUpR9sDKJA3JS8+d9KlYDRDPPGqs/Ryzg+aZ3syiskyH
pGjc/3J5uZ30BwtdURG7Sr4gXn0BpYH+MaHPScnuEad6aINWMtSkDXWhry6+FEMmR8APYEDnor2B
JEEm2XRebuBk+uFD1YXZmnSLX2ulxPdAfUNH4UYDIObQifk8PjH6kUVqaw7F+bNMXGT7cpJDY8da
1p9uVXFY7F1+jpAWcRlHOoj1UiIrfk/N3vcPhicxJKxPhlWeqP+cbVQ58ThKqaZd5cq+ekVqSJRq
k3np3yqIzFE7XjrBnonLEAMRv+qkn835F+CetzTnC3pM6a8Jt5doVHTHvEw73TgH5vxt3KbmVeL6
NDO7YhWXj1Bk5vftdWRifYgvqceVpC9mKa5DIg6MqvRNuCNRdSkSrshOKfy4KbbeM9qGNudDhPcW
WGGf1Tv+SYVvjNEV32NkAR/TrvrMQUDio331o9VMY90/y5NQy4EMGpezATr1rlXfLitFy07AG/oW
ef944/5qdziCOyU9Dt4KSydZVPBKBJScblUNaWRBIw+FXmi7e/ro4wdkrlBlWBWIpurO2H65B2VK
NLrTIjqokAFy9ueh66A6tHDw+EQq0tGBGZTBppvp8emTosm20R3lCaHu9h8nasQLuPWpm8gi7Ynt
TMFt4pf1yO0kskMeKiKrovpnK1DBvh86SmTBEG+PQG/nOxnUETbYNLwU9x4d5pqoIq9fuLL5RuHz
a909ElD2oZmIt2hj43I0Qr1A76w6KRxZxjmeNEMvUtgAUYnBR55tBWfgr+90iVuhxkVUmtn8RQgL
WPIpVBMT8AJhcvg77s00hKJILQGWE8Y09k561ZN8ybDq5z+hzipo+Szf8zKp4JVE7EloBz2nCt3R
WenumQLTvPxpm+3WOjqlnWEAUkc/wyzVhhTEq3WuSEkZoCua/ubj0yIzVQYf1InXbwg51FfJu4rZ
9CmZIJro0TA7qyg8t9v+YumV3xLteRKXnRApa/7xUV5laT60gnHT5kLVzNs+7v5voF0kKHSC11BM
DTHkEopdtCAGvFfAllgkDppk7b9MQMPtON0tiHJqvcXdyCJH/uMHJS8dpiWL7RSIUGCNNJ3hTpFM
KQPBejb6mSWlMcwoEQps7a8JSrmwxVOLuoQK95/+AM0+FR6rOWtCVSobzJocRjJ1CXYv32PRGYBk
0DaqjnqqMk6NBNTZH1EWTpqoZLC907TAjmWVEp/FtSEZRIQUUrKSng74E+EYdJnbl9tPu3/2qpb+
QeIX14HsdzjsJuZSt2Tr+6AtmLae+kwyURKH2r3+ePLTrwEU3O6khAASpRXQDvDsUB71vI1UW6Tn
90zs7wrmj5LtOssqKCiA9InYzw7BX883w2qIqoPEL8oMj8/ObD/KeI6VOf/ZkBW9MLo0G0lsJF+B
ONILgycE33f/skfYmFb7RRUHdQ2CgduTZNv46PZCwBsHJUF01fi7hTXLQf4Zmove3xZG7KP9kb4d
wD41kB1kRqu4jL8elD3ApZ3PwRIz2noRNNsvsARYksr1KNCZcTM9iaLcMYZlGHjBSZiiYfpFS9nz
AJepSUHgDRnLgC4Buzi2mfqXWINkYFQ2Bd1lI07jID0ZYraltbW2fLd7Qk6rwQ91r4CRkpvceig/
2Lu40ao0f9yswlqG9wHXpothtfWSh4+if80Cp5NH2KY14LfHo6+zTiY2ves2cyH4g/z356FKcXf0
ri54hkG88Le2cqKTvsv7ec5lJEyhBz9Fq9GQkMJor6+dg/55ULABVdi8clK62FlBkFvBS06qcIHX
QKFyw4j1XCT2A3L5n/5AoCU9DKJ/l6WPCHWkzYqatKOy3oToNq0dZT02iNOkqbdh+VHmn8isfES6
CJJ9UMWPDINLdq3rbYscfcy6bvz9hnHnvyA3UVUo9oAFYHRw+RQsyHZcGhb8s6q3Mj+JPPZih4br
VbPk1+X/tVI+aPCbG8CpcSHCDS0KwN+nuQMOkJiJkZjDWxOvtnXPCsL1n8Y5prb37gMCBNtTzCYm
41hB9M7w9GPp4pbkbcz4ldJn/JhsPWxZN5ytmty8LIDrL+qWTqeqHKe1grAh6Lk8JkSB1eR4UX5J
vMhK10Exvj5dlI//SCzEqFRGApRPCDK6/XG2ExT5+iONDQkCxrCwjXsRukW0IDsyTPEoNFt5PZyX
eoyvrqrUmvEwNoF+gyhL9sxW6CKaQIPmDAifooH/EVlQj8zBMZKcQxUSubhECU4X/uvDlfpSmHtP
8ropGt1rhaulfUPmv1k6LV3lP6kI8myk0hisBFWUeozA3UZ/qqd12yDqKEy7yectuOaZJVHKX9Hp
xSp+4Q1rHrv2X4ztEiebsPKzP0gBzDuQxI718UkxMpPM2OftOdydMyzgW80EPAbktohZzWcfhMr9
rz35y+FPw07RR788KR18zmDfShDjxGGJWiUzKW4J9R4vOvASIjObybuNvrTpsW4PM/lRkAjMD+ZE
4TGpQAdrPf9JieTP+/XwM8h3E7vR000DAwetGGZV5x06G7txSWU7u9dVh1Hu5Dk32lW2C0UkAtbi
Mr3JcFzYCdKepHhOwbmUPZrUtjdfMaHpiwGT34oJ292WVtQiNigspRzF65LaP7chDmcxHwE8kcwM
zb7eHPo98IUhTufjLcdF4Rf1mtJ1vcaQ+N99umouwbOCIyVQESyT4RTj961+gnFeyIp3ZTm1QypP
C1aeU/GtkOkWpjcdODgGDR0qmbzV+zuKn3bx/ixw/FiGVLbt8agqxZfbCWi7J45yBge1B5mlKKDP
tzq2QboVhyCoE7PCei32LLYHRg0FL/z5DIndlAup3IHGDFtDWudKLOrcJUQPo1XyW7ox9M1/a14N
bkmJbVjLt1+IZU6ZKZxKYAoUaxLNhXy/kuvaphFuWZBrhacpqH/HOfynBblq79IvB245wkgA40iY
l8U5BvcjG7rZYGX2q04wMWjcwKkGlxfKggR/aKouKG/9Gj0pZAu18X+bo6EkL9yppD6OsT4y18fy
3JLGFBnopkgB+ijpXdgnY/YAr1qljWrkXlrPmefGXhf29QszBtXEk/4EDSmZp/SlWqQr/Rkh/lwO
rYCV6N3e4koVbCeG2RbiD9LXSV7b5O/afD/aNeLzhCBaHmv62J8QKs8DOgO/kGyre0G/otE8I0VW
hDDXK0nRbcx52IBEO/AOxEXFLiDAosyOlnEDHO7xkjrcbJB/UZ8RVY4Mysa73u4zdsmkP+1EkvH6
uHNDYOp95k9+p4nF7HbxbjBElgfFOwE0oQlN7L6JhgalNgcCK/RedXlE+v5f198GhF82/ehnaE2v
teICbBzPAsvlPnlYABt8GYs91z3NLQOZxfqyi/fkzzoS4ccjyzXwcpeRzaVy26ztY0jx4ZXYHi+j
3JXoQrrPFH1HmywZFOTqpA2gs+pnzBCAHxyghrjPhDaw4LHNS+qR1YQKdpEwAGqoyBz8pXdxcKO3
E4stlBikLEhGROqu6cMcU+8cbznWD/VxrTNMOONuYDF8PN9sQjnNdBFdSOwesi/JrKvYtHVs6tJ8
NAyLLjVpVH0mXeYyxkvZ9IhAAUf6jt+oQ170S/4CBfPo4ldvdXOlLVubpjzLj6LEOd2NlV/vbM2w
zFGNiDtBIQ/Yk9bSC/W158sNDdKnpx92Go+ddavnyoZHOTgD2B6ckMIdagUsLEImWbnTM91pvKbE
sDTvX6FhrTyQKgJIIwXAF2OnMuRqvdhU7r8xj48Ub0pUObhIuUwQUrHQ/3k1pxjNIuLf7LQYkJOi
VMBcmGv+DX8qeyyXmJYiN5cozUXlatIKmtfWkDsoc102hJTr6ZGX7TT38A7xge4N4/7Wr7Yg5BNt
Ik9aGF5QWVzHhT08ZTUsGP8pFUok1iSq1wGGORbnaIkBLK1d6up6Y3ohz1ulFQ7pHYdnpUJfv8+T
/FbLGczEXsgmRn/HD6J7UzF64CYgZ3G8fKYppMHvP/BENledQvFqimny5OTrRf0QlUCm5Fi8l4bp
sR/f0e67DGuJUtnzxdIyCqW+UjQSCWhTuPI2MOL71vPtbUuByQxXx06QsfdRlDOTeO03GBC37Bwn
VzI8sFAjNa6f2cKegkp8ZmyBPoOwp2zKjDoQ8iGJZGn2kFiuUvkB+1hr+HgmO7uJQ+9GXkKP8oGC
sj/yt9CqlccObOJOOcgih6Q5ElZRXdVfqH4PMEe6GJbpnBBHmv1PXW9rTbHx5CBoS6jbZPcogKBm
U/4cXasBEqfgdU6Zw5iwdNgi3BXy/ANGdLzR6RS1tBDsH1ing1vfAESeJViXjxpbpIg5hvRoRfyA
iESPYZzwzQDNVDRKye+JQYdn2j5vv5PoV1LcU9fL5ouokYnOwkJKhYFEQOSKI9AxcoyNLfHjUBV8
eEOUpguXg4TrBC5Ix+xREhw0pEBjnDjZUxfuxx3z4F9LUaws8jXwpPYlegl4RvOkzX3BucX6iq4Y
6uHYqHX6CwQ4HKxDCSPTeC/cEJgrNqvtWAzFt46BUpWY+wSRuj2YXfgiJs89RS2t7I3IuEhyR9Rk
YIag+eeSYtz4JRGGt1O4pb9OmzP+f4NY2LWqgX93Vem7WJqnDNHybXyVyBCNCY12g72lw2VNTIcp
sA5T40OJ4k3Vbdjge7mJTEoA6jOQ63LdoNTTiSGzgE/FoQ+GvElFa/Tb95BeLkyT1MSquXimITQX
9mYPRVeM7YLkIra9ipWpHEMoUvlgJyuCbIUTh3x68FGqCrbxipYT/PyQze8HX3QDAI514mpbzGxQ
K3fo047Z6PtLKhPBZo7DoDGPmUTCZA5AzdnA3tqIvMXpluXA0kvic+NtbLJT9vcrkaavXKM/dhpm
U5hPOsDHF4K7od7OlRVWqNvbCLWhnuK93J/M7t5K2aBlEVmsS7h+8nnis85UmNqR0os1MuSXFzjk
e4Kuxim8cd5qM8GOkGJHkXcBHzM5MYoK/2xqKev76FUB1EIKcifii44ukNkPeofS5/zxIsDcRpMF
o+QfUhY7T7Ti/6az2WlPhxx73RRVfpKn5MBXq2ToAP5W3sF09Zrn2D4f8mpJvUMyfE0uDYdzBoWo
DKZ3Rx1jSNb8MtLVgYGlw8MzyLnnMDSY0wRzHgG77t2FzFzM1cMwOWU6lDZ+56fEQfXxyySOBJHJ
aFsjSbn3q1ABMe9BvMnuHrJXkejuq5nL3qLAeKyIEvGh9vtZcUscrhtefd8Dl6a/2u5MBv6ULo1P
VKxw9kmtr3hCuYYaFP/4LMWkU0+keCtFutuneCRIjat6sRaqbXQFR5++HosSTYsi/2N2SqNfYWrQ
Tm0mplhOaGCCH3LC1W2kHUnXQ4LJFFX8J1898eCeEDDHYo/TytHQuz9sfNWnLCGqxHqOJxnmlfSr
JDZKAiIG5JLxQex6WMCRV2uVi1hwkz5lDbkxvl0ic6jPLyLJFvFhWpKro6m7mjkRwWxxmvRL9uY3
Q9tjZEoidF06ae2NHLWuOolDZbcIDqEqj0ydUGXFljm2jDRZXNS8gTPA1sSrJVcNXgzpFTM6rRCY
sixoHepHyLk581GRs7gEI0m6CvuCTE+BfQF10WJCqNsmNFwtru5w6Bezl4/4s8DBW7h9dHlksRaF
soMpHE7uIaFDZ+YMIUWt+YIrpFFik8lXGiWCcBwKfRoGdzLD5jy4qE7aIkatS47sTtjXTwM7Abll
qijUhp/zjDYnu4Y4wh7F1sLU3YYu5dXjeIL/TLRRIJXqTGM3Zrrqhkkuls5dqdwdK8/zlkun5avc
GJkUdNpnJl5hQpRdqhTuZw6bKxxGs5U2i3dY0JvoBeIDArzHELCdaz0RKM2DC/fw26tOVjQ6Gxk7
ngnuyP9BTGx+EYytgPOFVWldC1CrPQSchXJixEfRC0aK5yZxrwceKiwW4Z5QruRAXlt7YgxWrPEX
PewVcdSOCAZ2Z3B70CcbCb9TFkLTiZFyMqCJu+IPEGcBfyIm7sfwTX6xnQc060IxdZO1plV8JGk3
cmbscuYEzQbVys+6o9sv/X51Z9dirxtHGX5XXqer9fArTrFSOP30iHUsL+vjh1MQp4XEV5O5AM+F
DPSZrPojvBoMeCyBOlPvzhHpnlvwkNLm/dwqGmNg9NsNDeK0PDnZXPT5KC9CR43g9zFuFxb81Z6P
qLiD5lMUUtq4ec5pGCRwoTgSZhXFAoRX0YyjAGFxCU5vbn8OH0zb+8J6BooHRlUaehSSwbCPwRsv
cg7VuoYi8cVl0ao8B+rtGYEwG9KdTbi+utmjRZsVn4456d9wv9SJXZgMxlDibiRgPE5O4FMJ/0/K
LtzE7Mos7Dro5jY8Wj3/yGiNoL/SKU5h8EdpJgMYfI65FIQUPTUownQFhs8rY4dr44Ny0VKVMWhz
y7wvh1ezeFGlRgxPS2ECECUHeE15594VtCuYdalJVyS/hGM9r8PsKgoL6x0NSOuS8Vme1H/4UNTL
f/X+ssKrnYUCb2o5UdvwkeR/I9lg+CMsJJg0VNU960Qqmch9e8AdtP1oV23FcpE45egegPNnWCab
l7j7Its18yoIsZg3gLxIzyuprO9I3hlELcsvanSzxiI8gYk56WT7x9MRlRsAEIAY+uoA9CHikZQ8
3rqCLTonJXGiqueN0aUSbLsABQf/5Eaf8LS33nBhq+R0QlUW4+/OXtufeenaL3SxqzPEqjI93h10
hRhHIOdO49XWWuLUdN6FwVl/h3PVNZL/VDnCFnQpxDC2ur2RougYt59X1SJI5iS/LWLTeME/QElk
8s/tAw4rHSFVrjUIKFGbpe4ep5Nc/QGMAZMvPCoc/f1FEEfXYokAxzn2LEr2O+6oiTTfLDo1oR9L
PZsFI/i95mq1Pk+2TeAx+y9u/AYIr9d/Ibf2VExiIyistenKYlWWswq/cb2KN6TC6Pf/ifohygdX
LMAmR1hTo8mmEMcUCXkoKsnqenPMA9VDEkOhxuXEGFNm9H6JKkay7uPUV+S2sjTMhlhK4OHZDabe
IQcF1KwPD89Ka8ulI25jSJX3xauhLiArFfb5S7eeaL0Vfu/zqnNsC9c7zBwMZIoPmvMX41p/J5en
86POsOnDNsa8HZ0eiKRADq2uKG70uN1pO35O12FK9nJbP9uk9BRfUOaKX3QET5vQDOxtYImrns0A
YllpkbOa/6B5/38lMafkIC6biFoFyZkwIwnBd4AgZpwprTohaes7KtMlCEbQlEVx8cVhl5ntwTm1
cl2qv7IyAjGN5Sod3QAxGO7XfazdBs5S+jCfl0RE/JRrEaXl8ulTIpc3PSnXP/FrQx6fwcx8FsSq
b4GAc7e36noGnb4A/xpLK5wvkHRxR/mEwYWSPc7DKO5r3RJY9aFpcTKglbSrgXAs4K8wNk+6cA/6
HP9TiSyCCEKUJMWb7SUQ6SoSrfTAbR4lsxNv0adbSd3mn6nci37MstEtSjdYaKMavWQB/iAgSJOn
YVk5qoH8xvdSjb/a1sMbSWCbtr4DysKq+eJCKb9iYlsUoMqVywJn7+XkIGxKGrKqCyBACFIx6Gb8
N8vV4SZgPoP6rsnQ1k7aev/XqlijCqFTSV7B613p8HTR+i2pamVda0dGFtO44m0vOwxHFujgbuLx
H4yegiPKwaNk0B/kv9bIv3kpy8roYeIpXO4mhZuGG2r3YjVW5L8dPZHxb83UZhfNMbt1Vczbw5C2
ajvx7JgphR8c2QvcAOX3cDfh31tZL6HUBNmQI7W7lBt5ubX88d71FFPwmrRHCC89fouSCaQMhU2a
MCAjV5c9WEngghJiw6ZP084rJvQcGaIHONGvvLUMcsYVbCxqHJ9PHbCQ3PiNOgGcQ7A2DROk1Q5D
62Xf5z+DecrHmoeZmLULhGrK1d7q83hcSPVrP+YseA3ITUg5dge+MPO6OBesdoKLeI0pRe4td6ry
+WQh5KgtWUtrrBnVfDi+Tssoa07Eri/rdinku7eoGrsM5hGXPbb9L27lQggSbajqiSFofrvMHcXS
1XGjh5LggNF0LILkjsUBVkftlnyTezLQnd3y0SM2P4iKUM+huQKb9S1n6t3OthFIhUm5V6EkGAMf
M8zZwE0abdEtdKHSrcRe8UHzfLiIsdm3fccT4im7kbP8cSrrv6g7ZhSu/m9SRizTt9KZK3bYumto
A/vHlG8vOKzWmkpBBuSf7aqukUSmimZy9hTf19EFNKD6bScJde9CvJgjwIS+Djl6VQ4GqLYmfUKa
edTQ0xuFsE4HL4x7lAjxG26UoRdyNWPc00MjlZxIlm/725Nx/ymIQEIHfgw6REeguCtCnN7asvtw
qkkmI2hK8LKUN8bqRxS9D/czh/elAa27uMEqoAeTT9hP7GsRm+3MFwP46T6X5UhkItdqBAVxXPhL
2jtoiWha4d+nYNFoQfn75A/owQKvFthqNdHnde+tY8MA6GWikgNhWmX3uc8+/MjLKsnyVgl8QG2X
bzgvQUKRIhNKehCJNTrbXfRa6eyWh8mPtxAyi87DqJdab6Vk+1wgdzghnTkRv5vxfz4q51j3Bd56
zYrVSmBspbMIz++sqYDVxwi0rQ8z59AIujHKN2Xl5bz18TC/xFYgijieFIx+AFvxWqDd4awxwDgr
VbfTb6IqRhHN8xBwIjmN0NP9QR4yfWc5hJcxr4+VSYrED01pHrVqox9cHyDphUF6L6lCr6ZJHks3
fp79Y64PXzD6VcJbHhxp5zi45q5ptGLZ+pfGyCQZP4eu/yL/zELQwGmOUS9j1g/ituqJD49R/imR
RDItT+gA1/GcBodPfDdfemdE56sv89jMVIGyOEanf91PF1VS2gyCEbnujHGDTqvcHDqo8tCFCUZc
bwxrR+eD9bKeDMsEcl8em61LEgSWDb1J1CZTZ/qNvHSgo24m5Bk/WAPLU9fxKaYaRnx/PzA5/t0I
LrtLhABOwPQhkBVJtstktlE/nwHkqgsjoi6AR4u8SqcNrxKQK4lSkeJIA9y0bwnDYHtlFypScXB6
/2e5J9bK9uF6+gDG3eh/+SrrcEG59rnR2C7Otj/lsijT7qj89LrG9PhPf/8y4dz1Nn8itq46Nttj
9jpnOvUa1A2Z/dpbWpmCKK22ZEeRKJLOFiBHhAia6R+CDS8Y315ck+ws2nEZBp8/8fSxSnDTH9im
3yvifkdq/jwbI66EOfw5YKKfv49JKiNKkha23TODYIwPcgVx4/SwVjixm0mEghFXtkOKtPFfbIq3
BBWmcKtwMIr+4ZN+Vh1wn+t4NcpQx2HI6lxqJXBOiM8awOUX35GGFciYnOyAoZOBqYj5VgyoLMQQ
JU6ns1ojr28R7USQDOigr3ULitnb1rBPYqJp1nbM+KCxY3XtPrpMqX9epRlvkSo3o+pFRe6mxTfU
qmSfF4jFt9xelOcPrLlOwhwPW5iyoSAcEBNvZXenCC2EmLvEymNnTew+XBxOoJAsDA7NveWU3+DH
SsSiXXlkH/9vz0LOZ1/zhh3rAgxjW2JvXHTVbA/E4MCTx210fjr0RLJd7WpAasRzadIUdWtwXc5D
ZBuhuiN5H9aiWKN/WcBHL9ywlxxXtJbUoJO6mJzNzy5ijIzJCTiEr/8u+LO9FIM6iNGchsnNOZb6
pfmbIpOHCCsIgviz/9J3rM8UAV8giP9dB6uou32LBXQ/DHujDGNxFbS8LVfc8OK+wIaEl0RaAWPT
9BgMEh/Wxggt+nRUlImL4Mv0cembuljbfa5a3hOzCiGjYjYGBF7AiQ5WrgaeSMGIw3B6Euo4Gmka
+/bY2pHid6r0H8DZp3KE17sCEFgRtUPwHYy+8UGiqkgVYitzrIIN48wacBq5EqUXJBT9jpcAFUel
kVm3SyUortAEsQYXmM5TKCmSKFDdysUdw/p9aunaTbAoUb1/++FcRK+x2tgRHBwPY1yJAwji+lTG
NdEJQOvR2LlJwhVSvy+lTAgVpjIB4hdR7lrkuuqgcv4k8lSYottoUU7/OOFAmx/mtyNGgtW0wfGb
eFTWswKVpz0rKhTtU0ehgDsiAf23frZUlwcF+RhovtKBuo+haJdXR84yw4Tq3A19sakj/0qbbG8X
F/w1tNc4rRczDczRnJ3RJ4gkrf31FfD0y18dUdDTIvsPPMZjgPJPhN6wEiSICRHsnS2S+MVK3iiK
PliPtBfIM3gfV/x22GEuZfz4ZL1pvxixSI7uxopVLvCNaV/Ir51F24dtkoEKdN9+CpRN6m0Tmd3P
moTs5D0TMQS2FxDXuEIuSV9p0Bk0J8nVWW3+djD5BW6pXWPslTWIMuf1DUlfJcdL1FCMj8xCjX8V
0gSFfNspeSjAg07IQJ6o5HnAXcQxesEDeS6QoYQpzNUOV+2BiCLVkNps/5Q5zuYaIi5a8T9Z73qV
+JqllERRahp4ccLPnZpkqA2CHCaXprC9RvWzCGvr7RDPW90Nlz6sa2O7VGDorwzcAabIpu2E/7HQ
rPqs7tL1UkHUShJLVCwq4HUEGC8ebpAmfqG69ls4fXfss1jlW+ND0YgQaUqR6XTWzCTZOHiR2hHY
6wnssgGUN0aP2Q0QXaG+NBprZy3Z3Ynrf8Q1h2CGJFAnHKkgHT2ehi7oV9QcTqJnyeG7IHRYNTcw
0F/oBZH9H9f7iHGDOT2SrmTE0FG9O0scPe4opNeJhaYJFN4KaW8YdsYMPaJ50KNgLF1ReCCJBcJK
UZxHZhcSl16XooTg0xDdLO6FiwQI+7cPxEgUIy4oTFtKz7wJjnEY4M4aWmltik+n5pTSS6aduIwV
IhngnTggG6V3AnLvA4o6ETO44lrQyA+HV6yflaNpbF4QjajkG+RclAAvnwqJd6Xg1Uwaveyj8gdy
lcoF3dCNccrYm5SiVyEuOUKEmW8HxyyKVO7ScbLXGyPP4Dfz+Joj+F3Ig/c6XCfcKWzGyJnhCpu2
uobtiznxpdujB3l5/3N6oF8z2uM3xL0d84MQxRlm0t4Q3G1voEZMiA4mQ4QY36FvlXWzFTkoFdGA
q92kLSUQ7hfbT2t12/3b5Pq4H9fhumMJJm2LqPpRbtZcdGeYqskp2ZZ3bl/ApB7nnIAx3Eq1zHK2
ysyOuA1qeX1cp/QGmSsjEzolyRQ+nV95oarybuzqb2z/p3fgIIRnTj92gakgNMEDDm3baPvPeanH
vuf82Pb4COqKlN/thuSEdTSHC0gYI1OVqBScWm/ykW8q7gCuRqK7vovaxT65gp2BdrKh53zLTJO9
QEbgsWBQJEa8tiYACT6MJNkmuLNCNT7ybdRhQqGGDn3KCKW/VyLrs3t+JVR4pxNlpQXrxF6PkDHK
ysm8YakScYSbW8KX63sYdfOjgmMNO/r+5VIdOIWMpVg8SD56t3UGVDlK4bYPIT3HBZBgJd8UgjkC
nUOb4mSRaL7H8740gB/3HQVZ2a+LtdizUA309fdk+XvECNdDOkusFB2JkDaaAuWiVRmaO9Elztd2
cqOtnM3mioBQJ2uEkzetY8h0fXq5ArA07M0X0+SevyzKOl0F4lv01zvbhHvFQTCQkWFkRd6Lzg1N
z/f1xnKaU0XSe7oJ8/mOXQ0Q0DfzeSW533Rdkpl7Tb4U57Atf/Bt4XS5wGWl8+EhIqoN7dH1tIOG
n7XsjfjlpPxH1FYgcetsL8eXh9Uj542jPT+kwotzoYqSqkjxqPFEielyyqVFT/JvYHM/tsBxHT+0
mR59RMxAEpj+dhu0yU4e9lc/gL8JwaOhw/d2/A0VzfyK8bz1IZacyhE2ZfIKUhqvaxp1LQ0xmj22
xYxPEbzRhcA37+PM0/ktumxMVfzn+FDaQptbq8vkZ+oERZ84ZqFH/Fcsi4nlkDNY89mB8fijkVuc
p5Jj8n1/zvyIJqmTGji33HyqVyzOVxoH7Nz3GqFkiUEsvqr57acyPdmYcBEWYV7EtpaTwPXV4nCF
xnci8m3bSl6zbYAGXCS5ikPcyBv7L7PEANFGvpwY71TbNqFNSdkIlRaByiBh/5X4GL87pIoZRYF3
kDFFfIu5AFYqFY/t3zz59NB3SSihv8ZqZDKUoYMH01VJiFebDfyT5zsLd2be7+uA43Pok6IbQsAD
NnFIpchlGjTpQTjnyVMO38B4eprAyys/GCXojwfNHIyRXDcse58DQ9ShGf6xuKQ8xkBItEbcdOdT
c5MF16zLNpsn4jNvcVrOpoVQWInG9Znff9OQede2fQB6jV4h0pDo3P3s5q3sytAKvl2m4ej9kIQh
LjDPwT7vBv8yis3gmHPLXlnuNKfALzzU2ebvVX8Q77DVaoUBYHI2TSIf2UYKsxBPcaNm53B/o7Qr
POWUIh35eD8Vyk6OycVmUsp+sf8qe5TNDndBFFdHWJjoo7sYjNnddaBQQ1nnZ2pBXiCA32LD3r78
ofZoVbWhUw6VC7tPYkdgCdRrEeURAk/LoiRS2+dSOPg4RUOT+pvByS8mrH9WZaqMbOYsDtpnk9An
y1P9p68JiAviUcJ3MjkI45YzF4WPeNZVX/GwcJ+q6aeZO2CJShVdgF5bjC9KVQ//1tgTIdkJ8Wne
fmr1PWLTh0h1dY39H9rc4G5fPnVplZIdexZyAUVikNVir7qnL3EtI0PXZR2+ijFmp4kq2IBDoS8s
wG08kJogcswgaAXD2Y/78Z+aU7lAoTP4AvjVOuzxErlbx11lLntDSQSKQABNWWerDH+0azvw4itC
X2oGthnhA1PmUVb8MYaXHPap/BcA4l4TN9v6rU86FGFpl31Ioyo+Kt2Q0YlngeLiHfTbJZ1eTfuu
dQe1KhfFeBD127JYWmSuWlRSeVACouZ1NwkE0LN4AcLiIlDW6i0JCUoNv8W7zpOnITlPLvQTpxnq
WA7Zkd6Chgc0BTsrzG3v7JmMEfo2TdMKNT9zw6884eMC0+kAaV36ml/UhVDcJQJFySCBK4MzD94H
aPGrDoOF/aZC+z5FBtvOXHVcOObGjfndSBRRLikwswxpPJ/lWB+0VNqsxgq2i5vCKi+vKf1+GEwa
GcGHe3kbm12D/kq0HI/5rbV3SHPsnmxWuso3YfzNFWK5mQM6BQnxU4srPCvRZCWRZQZHY2/t+d9B
mbgfATw8seLA2Ad8OYAc/xEvky24CStRZFvbpdLrg70i+SXSANoRIeo1xKHrdnQfDfTI15JjpKas
So677+K6tNzVMMo5pqXq65VE9waD2v3wpZtQlksiOHowjN7epQkLwF0xxozLt/YAzMuVlzDo6R+z
/UT4nXrFNj3/mv7v1R01Hiq82+Zo4tXfIa5GURlnBm17xfSJgLgk5nG5ZnVCGolHEFRRvpob72LK
3kHgEIpVsEFcXRRK2S2GQdXofHD4FaraEEfex2MPFdVdQ7p9Fn58EK0G0Zx/G+qYVYXoIHHHYv6u
UnAyEz8fzKBEnAaqLfpQl6Qa2g0oOhf0YoWPxIWwsgPQHzcdxG7Gn7w5dIVhQR36MSqb6zBmIUa6
05bIEB8xSfVAPEJp4/2w5bK1BxG5bSFw4SR0On0iaC1InMTQsiyBxtFd/pIJ/eRRJMZTxlnALFHs
8KbvLQFzKFJe+cpXV97AW7ty0YU8JZdaMx+2RPlQTvtqdR/GAOADlnVgDUyoJvNW8ozIjDulhlyV
EicYfYzcaI9MmIL1GBFMU76CjPKyaxCday61JURFNrTf+9mR81HNWSVYxpofXcAwhM4bDI+i2Kme
vKqh8wyPdu0ifH6g0N1fM/3jdF7XfBPbyTXKXb/MkhSp6WaaZtUJmHHzd9eSbq+gYqx2qwD32cOU
K+pxCNN2oykRWlFFzKT3kfAt3QgdkV2v/uU/M4+dh6jPUR/4tXNpd/nhE1NMMdziQmL/vqnXQkar
tW0W0Jf+30OIft8JYQNYsHj1NSIRzTMLVjnoKnupihwhNVc6ox3ME32Mp65dWEm5k4uXjl91d9fT
nojcZxglpvYo1PmMjMIdKLKxGq06KZUavH4wbjdmITI3RqPg9/i98XzPZGXtuSeI60t9/VKggCfM
Otm3SOjQel14uDYxXTq3Z5aEZ6+Js0WCvliBRiOsLzES4jXLX2THEmR8IKSi4wjB9iCiQK9DfRGE
ffzq9viwfIoCuQ3hOnsOxZ2IHkj8WBaU2QXJuu1s3+SpLtSYmrfEZmOjXrCNhW9F6LCfei1D2V+R
IOe1k87mzhWgVaymHQIvdQPuykx65pqSdu+WeFrOXIpRVCIfuzCPJIWUxl8P9UySG01VbvrT79RK
vNUwDZ5sBA353EncXNEx7p3DzS8JPmllWXV6wB0abxvY7KbJLRvbcFlfduX95JlWI3Bi5U1U/qp0
cPwpHFBQjx1Mnur6TkXNJ2tRe+7ypJsvf48DiO1YhVgQX6U1VKR2m6HZ6j9H/0soQhgJ2YkXlCFm
ah9ViZ1RVZIIfN77wGgkvvs/pnPRZpXVBLbZuTKxh7jnb9UVYY5SCa75zIAewaxb2gB13NvL4xd+
YOoGWtmA2hBYLj8Hq2g9+s2HIZbCjQnI+qNn0mD7ohiofc/Z9RU+1LVAe7bp8BSZXm+7zplQrACk
GtERTS1won5KhbXhpStyvZBAkDQi76vPmPsuoqiBcHaFFTVVIrsP9XnW1A+59s4Pcjfz3oU4G9Nw
xpMC0EOIi+JpwpFeslHuv0KzPw52AsCl5EtJcgU/9/iorgki6lYk84oAqeIRZSKnuxW5q1ZEnSSN
rSctzis+zgHou00xfkXOCwrswRl9OYHjgpXfZ8gjYglvI8GBpb6g4qV7PMAZlqTSgFTmgQ43YEmb
1vjjoKGnDzv8Y9Tm0rl8x8qpRUk+NoKUz/1ke5Es9AkCU7N8k179bgduAoc//IprxyciMJHR+XHr
sUZ5nKyCLAChIxHOeHfZWoJcBbZTBRRwwKBz5iuc5ITTLYjtaiS/Comgme/xgTC/bfQU5MEhFc6x
SMA/OxMKxXd6v3VtMFABYsvulLLBbKqRzE//0hL2qmzZNmzYsC5f/BrPjR1g0KrBcI6P3bm3w3wc
eSzOGKz+ZRnZO6Xb6ffZ7vb4Eo9kSF1f1IMUT+yrKccEXuHRGQ07povitMz80VE+9R9JY6788ZGv
S73WWAvMU+MrbUrpRIpd04hF34rMYmaYDoUv7Tr+m61B6ZdUkIcNXiRGfa9XzRCQu0s7TwZ6fii5
r0MFFSx5Vh6cGnUFklhmtW+MmYiAg0Iqx2+qLEAKgd+rW6vK3A55w1o2nA7Uf0PFI4hfH4X3o2h+
hE79qmcE9kqAr5Maf3qLDp12e9lhkdUPFa2bI0oGR2WFw0AtzAdOGRGnwa6NxsZOiecNPUmuORoL
ScOlM/BywXAGlcwiHSy/uZwVUV/aHiVEzFpuIqmIrjBu8RVaOt3jQbygzrNockWwkFKVVm5KW7cP
9DMFnT5vSRCylvK6cR6n1+OkZc1yN1MLaiEipDphtLloiJ81DU/OrmBGUEkVDHYiqf1dgX/dVAbb
nYcK72AS+VQ9MdDPelPrg7RsJWYvQeBnyK+4dANlzAkTBc508p55vS+/qOhd5hwcOlXAS5A97Kzq
tbiMs/v53gCbNyoNADdnDVap89tlgolPN/yMF5rZmXZgmpbIUuy/GGBUFqIdqE0z6vMCAmsLjPNy
YQIi8Y/TgOeXWYe2POUWmPxtnh5AxRUHlYS59fAz34n9YgCO+6BXFuZit4j2yYiAy3MJV/MBG9mp
ulSPH3oOdJBczv84feAi48GWTxVD1f4MemVtcVeuhxAl2AwLhQ+Ev8EH4riIEejihDBBl89ruyOx
KoNlHYv/bT+td6EBSsa01eQHjlQ7SwKuI87ux9bmk2dHufdowk+zvhNVgjLewFmrsdBdGcQO2b/7
6/bWQBfjEJYwTK7fwFNxB5oTofJVvZ13AFPFGIYEFh3VkXxGN8Q5kzCzY8dYXWaPngmm6XaSJE01
j89KWF2rWBpNt+8fYF3F+85py81BLvS/898GUTYzxbBeBTqc+WmsbWDc/zvhlxYujOB0LapfQiP/
09nxHRu6Y8EKGQ1SkBdbdwYx3uLnTS7Kd9HE7e7Lqwww3ro2V3CPQZjPiFRm2hWrOvx2uqrhdzSM
tN83HH/PbcD9ZWaFlYwusYqbpnXhJHL4jAp2XzuWppf5yN+mpW0DP+lkzWsk6J8SPPCmo8xaHbMb
160LPLZ1KTQQ2U53mFDSfLHzcPTzKtX72RaKiSbwbVEWY4dFKTNdodh8Chaajch6O44pd+POX5zN
jbz6RBOjR9/aLpytOZ4J/9eqvSvmm8z2Ft86bGd8wLngkXy3Qzah/LwOlBPmHjhhOG3+S9kgMV1z
QOb3EO1tq3lVn2mNdGSQ5+EnbjjH5dHl2AdPzJ/H9s1H1fykfIAnrsnFhIawaCl9xEBKTdyWc1ff
MkGC9kMiRmwsDd2sRdSTwvz3+A6+Dwwyil54om/njSjL4y3GWDbmhboR+/qYpHuO3wzrrOJfTw1x
26FGQik2JGa0CS89ctexk7cztYkAyn830IFjl6ttGyMBlxNdIt0DcHNkAJVykN0v6WHPKeU0BL2Y
lD6L7PpaeqxJmix4cOQ8gqeOxYIo5Q2s2dVbTzn9H5NV0psRIddi+izzGpR0sVXzjKIjLszMvrKU
ksvE9rTqTdexqDOtAhwFCf/inot9ZUIntd21Y3dto4L1qFHel6V5N5HbNaVFnSriwXLt+Ml7esk2
Y2srxaKla0xMVaJh6CIkP4F8a/j05zzNZAKt78XwSCMSSZyicHOZ3Y+MzI04yMnLX9M4G1GTtEMC
DKvPZXTk23ECrFjtVMzl5ZO0bb6gV2EAGipbLybxdn8FYQ3LJzMy9KxiSarMaTEd2G2PV/TifXft
9MzWrTKqs45liGiaeJtEsFU63Apai2fInkNJeuylAACxGjk7y36DWTUjK2T5XkC0/+Tnmcl8yxsP
bH+y4RPdgh+gh43LF6flJdeHIMWN4IVZJqPh2n6LqzveY7gWFJ0W/4vgcjW7GYKm1lK59HGGvF2z
V324/bAAEkTGch76Wxzq8juSL5LndgOfqx9l1gk/aDz/wUnaz1OX3rrsPHMpiJpdqnRB4UfdnrVV
tluaFQzhngAjs44KrYo4lwqHytLvW1bF2Z1z2IDHXpNmmSP8YimMNweEGNSvwbkuXNujjX2icjat
KhcvsOxl085oN/9juVS1365F1dxPYHwJ/pHoKLEdGxwGWF4S7MZQtAnKXZbN7BtMtCTeIXFwaRg0
Rukop8OUCfu/aHx5HkXGEXDRyV+ZCGhvMR50GygfezXEMYiV+Ab/Kc8iiMs+QX5xTQio7nqp0Uns
LoaWxWDNLNZJeA2GrqisAxgCZQc4JTiX1eU077d4POMsmxTW72jd5b08r/9ZI6jSP6IWE81oeKHF
cLfjiI6GZzU5gangvKR5E+vGRNKUN1MLoElUaIFej2QKD6F441ePQgDZl9LlptSHaLD4OVENlEhz
ZtWF/emfTWfyXsWOdT8YCr8tauFi0y0e5a9PJz/gKzZqlsHR5rtDeqHWwzPEohgxY8/1vIA5fBZ9
4M+9Ve6M2xVW2wzsGv03gltQXAFj5K0HYRwnIBcCe9l6GvreA2WO1pGzo/Ctl9E6LfN1bcBI5vME
gz8/WA+GXm1vtY/5v8nvaZUgi17OKKRcC9ZJoq90kv7lAD5kc70OKRLsCWYu7HlDlb83QCEL9rl0
5UoBA6XqKM+SUca+3tISltTTDLyYTNoLn/b18+X/mVzFlFA+0T8td9srtWcX0nyEhZp97VkZlP+W
TYBPd317HffynMGcXHxV5gbGiiJjF7e9du3eBYcmCB60GHvndS9oyCQ3xT2s3RNDQlX/ajsQt1Z3
ZRpbpQlbPZp5KqmhxL2icj8a4ok8WgaQao4IueAfSwddFUTgxDlRwQf2mnAqhBepRYsaqmf99XwL
mJogAqjh6m6gb7yL/U62niYdeuD71G8MVctVHOVhht5o04mHjFb3/xMSXZUMuJvC8y0a8L8nHEz5
ZFOBCQzzStTBbXZMDclN1J5icPqglyQguVB0CgSLa9QWwxvJ/VBASeNSDKZIhn6a9acwrgVebXnP
fdnmq2ieIWtX5pBzMoVoMHCsMVSvwov1qQDxgvBufeVLs4MGJ3nVNIYvlWlkD9qvb82pQ7KNSLRa
CUeHAPQYltHZT3RQ4QbK8Z/RQlRdW6qPrvVUOadH6glKw+hLvHe+wNwjG+QQlYFjFrqdHVaGDhFH
OLkx92Z4VdibX4mZyd0yg0dqa8Lb1WcFpzupg1N8YrkaZtjxJlLf0xLgH16sqOmfj1e8p1tCfF6X
HzSarUW4rFfCvLNEsiKscyoMqAJJklTHWV1QUIESWNDkRvftmxcE5YoJoT5FtCJNr+aEDFceV848
rCmQ6ONqtrK6ZMPgtweEP72p+ctd2E4TyQRGF/bgFdf3PiEPuoVI+IYhTqh5NcrKqR81kWORGndC
hZhtUGybxqWmPRPg4x//1um1MCdJf/7yXc/aiQ5BGxe9O5OcdFObvzAG8zdKsG7x3ztgpAazKhe3
UhSQb3RCf70WpX/rtOGWPALBmWnKbNX0zUEEPNQSvbINYgUQqe5UI3Cqu40r8p7PvKKat2Bc7q02
ZgbGdnFijWAwqOT9f2G4fDnKKpBFYz3N3/cGdgNF6CZumBDNKE1dhIfIWZUtrayoAhH3s+8ISXGM
1PR2o8Q1Fn/6ta2FppD2vFH3JvYITPbrmmpRAu+47wbftbofztiQeM5OCqDICCJMxZA8uYZetII0
wu3CGZm2tRemKvjMbmdkmk6l44nQWBc2LSRgwKV5N+0iAScxl2IYGE2UZkvXh0CQWgmc9aQakAkR
6NBIf90QzBSWmQl0Hhy+Bsf5VfBSIADdsOjka6JZ0W8xcWecuxhIH6Vh9NQREnbTXM8iIFEyXJ1/
BU8dX8vEirqdYdLqbLLF9UkOEGxh+5JSZOVB7Dtk/y/I/vBqOV2Nfjqza7e4Ou9jtQ9++I2cM198
/a0hymuwpcURECcLcaUdpJcStmyzS6cdVjxitXNBSr2aQ1EwL4GZy4rpQi413mxIglxKzn9Nit5V
x+5rtdoMmo8cy/zATvV8Q+BEQgvZEMV+YVvTnrqgSHCvVoiKBSS3PyKCJ12Yvp+YRi68XOWr6aeM
tJXJXgubgC/KBAo7HbINnrWbnRZDA6R0lTLgFkJYa60WEqO6kIAbHpZnf+qo5Xlbp7evtVDxR0wy
AVJ2dVV5kmD0pxruFBnNm67aXGHEoPrE0dlKR5+8Enxlk+sriBp1OHFhzanAQ2dhPZf7p3wegbXN
CTTmN32QOmP7QOqGT+N8UJaDe8Fy7fSXDim/XBgQ+yWtB6zqVwZ3Fzk4O4ubt5NNaiAcJjv9azbk
K3VxdLlEf7+MDg+ai28Pk8rLs2WH3uYtKpZjdwCXnmF3ne3Mpuchnijr52hs1QMfrwy/OhGwFonT
trcWquKToVzvNc95dA8v/gHPZ+Ee0XUEFjKHPzlEfkPYqcCdzn4zZi+Fp/ufOIxFF2AhLYNwM1qu
XAqQhKGgpmecvUfVhGtsfyZZPN1z1SG+ps/sBDN+1sZeLJxr4e0tKAjTCM4Le1bj36te2AMnVqiX
MZ8/CSrxQ9kxC5/xYQneW+VD/EunsP1yO/DifgmY6No/f/fpfQj6vMnp0wP5cs6C2nFpXd1YI1Or
luLBeQmLs5TvqbXuZcYyNFkRYxQIdPv7pAm4o4H3ReGYz6QBR8UOZ8RHO5OR/b10edmExLguesgT
DfcPQyR+oAtODH7cEBGmm+8pDRLjX4e8K4h9KB7GaC6gBGki/kmtcePiu9RwH++KQxYMZ4IQqSGZ
+PP/2jQtci65I7do8HopItdTaGxcPtyXCAUqL456G5ttOiaMJcsUt7lueqhs+yapfTgTYGC1M5AQ
4JsyRKTySAJChrO/7iw1ObX05kpZx5HfyLHyBkbrDhb3bGknLmRyMhME03duFDvryBrZTz3BsaCf
vonU0w0HR6mAdkFZ0tiLgoH/TnIdzt7TGHgfGIqFTuH9coJe10BSTW1W8BHmPTri3bEX4vrXBbVE
jzOvOxb/Sc7Xu8y32xTH3QFbI4ONup/47DHDHo1FBJOo4EOxaL9ZvqiBoLBYCLdoXrHl2aPG15Q1
ElRehWWd8IJ1+ouTK+4fXwnMGIs6aR3EQGTFzaNuWLLkIXhYhTFHd43JQjzp5A5uio75FBnDo21s
tt1rgJBZnvuQbEkKcAAqMy7T3R0Vszg8xYh+uADwxEuJ1N37vY6n+f3hNVN6UQfpW3PvY7OxMwdu
SwGhauQje+QSFupHS/mHsZRQJiKtNoZ4jZZK93W/ql5al2o2a5WpNBu9WD1FZsq0vyyVf9vzHMtV
4nnqSPq6qjnrSCNJgrk4ZVIProD9m/n/o9jhxujbMONnXbYanDeQK1outs0Y5x6xgTyUPlQTcU9d
N/GJ8ZlDCXF1oPN3hRoBLxqptxPk8tewSrFYQpBFx1q8QS9iKW17Tgt52VEf6jNO+ECMzCnzlIZg
7rYJeJDnRuzcWiIQvHYxZR4t67yRQCLp96umyFn8u8wbyhG9pvkQYOw+aFba6gJTJ4O15PPJp/PA
iabGLtuso9pBZDbIvjcb6evcv1gZ6nyYla+3/UTK7COkX/5l9jAc06odxB27tz7B66MHT47MDMit
Se9iYhj/HrW0ekWylaUbxXLeBAXF+l0o3pEJ8edxGGY+cypZ+2+P3hfkc270s8qC2n6WDc9LIomU
6hHt0LTb3O8FmeRHXxfdhP05LMLqC0KL3w4znbYqiQ7CMlsJ0VbWVWmeoJhJ0jhPAaeCjkusEa66
wdBtOQ0sP/NAYzZaMUYNghxpdWx64mUvBn876ig0m0u9X2mPlxmG8uF8yB6W80FwlgprM6WKCNGT
p99GVRxJgDXNFtT/1z3d+T5DFcFwaAaPkcT0jL1yLpZiyNlMtKxoHbNquP8Z/U/r1vjDJJvTy7bp
gxKNZlxenzbFzmaMWxilCCuyrxlEXxFTcQlSvRlPJ/cGkvRUgxwkA6bdr2JXx+lIhS+UH9DPS3rb
Mtt9/EzYnUZG/Ga+0budeipgPL4wbSc6e1Mzy3cFWvgK22ZHv19PfDsjqqJ1My1Mx24fk0YDJ1o9
1YyQOPNkA4pxojpQb5UrlqcrBqd1iFZ3pkMlEmDNl+M1eYrDXz1MlvTSeGaAbTK5kTDGJAPFJvMR
+XXKKByjelYRNY110RoS4Wx9eu9LBHf2vJhvoE8MI0FTygZ2nx1m4s5qAjD6IWD49t1QNQYlSFT4
T/nuEvbLbcYourU6Q1CjT07rTwLPxqozxenQZ/emg9Y8TphT9eDFnjBMIW9yXZ571jdSUMN3fQJe
B+1qWfD0aa9QSalB/oB3qEG13UD/7IUEgoIm7RFmtsCjv+gEFvrcWsSn1/D74f61Do6XGSQ4RFNb
Wwo5ryiFhuNecddX3tH+FSyY3CevX7zgBjhRY5ore/1xvi6Gtnfoy1nHvJg/ow80Z0fyjdn71FTo
2Koym1YnZ9ripk/NOOo4RQXpn4NJ7yJWlUMabKoMWim9zeTAqU2/JP50vj+y7sl3yNGkq5dfKx7X
x0iuBTH9Ls+Cb8QNOJwLcA5E3P9kB0i2rI2yD6E/r5lFxsRAlvP+7t0SOzaJ2CLRjQp0JtuDZDeW
GHdGryY+6y3arMnnkdD8yhurbXCrROA0ChTDZrvgyxIEcbTtbCMkSs7w9zslOIpkNH0PcrZjZ6NB
WJnAOM1fCVVPXdIfe2DbE7RSA8/8KvnhrmUsle6VhYwNyHmDQtZOjOSXWkK3YCzPbEgoBlTNdWCz
8qV/JZN22o8Y346/Q+GrgYErMtFDofP/m3FLpXbynSKSRmLdz1iJsZNrr83+liSX+okoRXYeqPG2
SsGf5FfzoTJlFPkVrN44GKtXlFkdg1+U++gGO5g3Vb6EoG2RO20hWwjtuI1WVv2+SU7Iyphn50hr
ItsIqa2t3HMUcDah9BB4aFuRnAxCB1Y8kopKCu1JH9dRJFvqrnxBhijg8FpedWKCSuo+s8F0qZC0
+jf5GSV1+tdSTFf6B5JxJgepS5pQOGBQPkVnseDHda8Q5615ho9NbO+Ae0WJr1FK0QhVhVhkBlXM
mRsZOEzNfl4Sl9e8BNrMJ5EY2Mt14+FB3V9O6Y0oZvamnxx+23ESaTP0nkm4O24BPu/cGG3xC83h
kubrnPr0nYzxMZpqU/X83ofOXaT4Zw2quHQ3NSRT5JivaQBVXmrYbDeR/hrJDXs5mnKG9zBNCUrd
fuO5n4DesGFMKDbQ7b7hq+56t+DpEW15BQVjzxYONEsXy5RkpAtZvzecc49phTZIChW0y3tlUq4p
RrTgxG+Kxt3YNOs9t3JN2TPKzLCbrvTtbmIeuiJiHdxuw9NATiC1Lw3Qiz+1ZzUp7l2h48nt+W5s
QU5FzPMZyeKgIFCUUJy8Qb9zyR6SKEE+fGAdlXgJxzlFzB8nIWsi9nqOZcPTQ3kcTC5mxNwbsb02
X05rfAiil/b112GHDE6o+DSuxi8GYiPSQXndJDnPvUAm/AAN9QfISWd66X8uL1aYhm1EiuaLzLjz
YEI6GScox/zmbry88CaTsB4KieaoU99oZF9qqyJI8IJNMgfAs42voa+9lRMRPpokua3KkAqjaMWN
KPHy2qGgu7HaLwGElX9MB/nd9Gqvt1Hhi4Se7XxoH2WDwmTukoCvo2zv3bEAFIjaFiekNOLpTIib
cdWXPsTZCL0TmCr+x570rmpBEzDWFhO0CWrfJHK6OkM37r3lmi0DFIq/dGPD2TIwvQw55jYXac45
nN2c5H2CRn2MhchsUmgsfoLBOvEBAWeU4qEURF2dY2igu51ePjKL1+ppIyNmggkpf7qe7VMiYizD
xhWJ3YND90Hx5TWVGzZZuJVzO6SydWfY8LiWcKp8gGmV0wBW4INRrOPe3ZCudSVDTkFTGkKHgZiE
Iog8WVllQQGA0tpMR6soA6iEUtZZqVVmAhDHwSpQC4NfJg6wESegDWUPNi1qDHhD2l9blDemhE22
fdWXgbIEZTI4lpm46b6R18j5sUzXaZX8EKiEMefWBn58OG2NWFr8EDiX3Vpj5gAgg8puIDqyMLep
Kc53mtK8++O9crA9Z5J7bIKkPxFc2gOaobJkp71X0jnUrcBAusvWyBSrSmqyncIEB4rXhuRnGCq7
IBIFh9jfFhYujdUq6NrbaTuDVCKEpZabR0zygyJbpp8s/OPQ2YBcVpcnthIqopMNfUOIEFDtvHEP
E68vMvVPN0CWXaCnGNtLol30USf0XAItzi+SXG2p5j3yiAKvpdjZcxUXbXO2Mroygu+/5N66nhjZ
ASPMBBLHDlMXW2AzL4xFMUrbmJC01mrVk+5OG13JzOdrSz4McwsoRBHm6dJT0y8Iyjw2CC6ISF0H
r2Tcy/J8Xw6yfwpwT7UekxS1r09WshNbT32FLm7u2d1yg/ceLuXSsxNgLbIeeMcGz/XZv3kFxl5r
lWoGBOPt0cckLRZjNsFsqyXqfB45ZiGQ9j2ItlHMnUfy7S5Jv+KTCxHPRzPanpF8D74Lg2LpygML
vB/45jtvcY93HclmUuFxg8rvrnyJeqVsAk/XRieWMTfejYjROqNPFFHkEyYgPm1Zt7dauOW57dK1
FEDQ9/ZP33Gsn+Y/qGW4tQ05Lg8yPezzc5+azk8M5Rza9EluJWweHAjjPRIQxVNh6Vlo+Cv3z3qy
GaH/6O4mfvFWEwuLmt4Ru8RVPW0FaSbyYhD89Gm18nfRlI7IjnQlpAiBaZnUN4KkQWIvBfMOClMa
f/an3PXWdITGz1qoVF1F3jgxu5eKXcCd1305pOWxim7xkLoEpy+1wPlmPeNYaKpzxepCsGlppAtq
To3+ocfysY0z+iYu7FV71KrdKXYvyQWQX8SsowIVRCbWiWWrF1Ot+6uzZ1qSyxqfkIXdc1NrXnUj
u6NCqYJ3Cdgql5A/bAGwtrV2fguOIX9UZ3ep77ikKVS7OoRGB1mNOxqgMVHmITPSYE2cxWOfI+sc
0SdtI8Aqhr3ojaLUbVnQbYaA1huacPcdgmi9wfr04AZ8sEbCDGfhvFn14r11aRQyXL3Xqc/D4ri8
INeFCPgvCfkYzIPWdXoxCNLE3pKXh/B6bHCPOb6NsmGE4D0w8kbWUlrB4SCq0yr/QPuaBM7fJvDK
FLdkRSd7EoADN7zGxDEOPdGpkHWMWn8cx06akznhjTAPi8exTsVRHrFb9Z3ZYO+2P5yCxWXTOggT
Ja/ngFWN2UhY+XdCsNLcwoSeLnHbO4k3moF/l1vIobNW4cBPLeM+av9sib7ZmR/3HcM781LSkTQQ
H49j8LsKSRYziZ5eNANYiWmdpLymQHewlQFuFUv/pjxxTE5hlC60oVTQeqQ8xZKamGoG9ooyqeng
YtEcSWBsuLqUInqwUfWtwNuFAaM4Kqe9m1M69Yt7Jc1DstvTKdlz7sGfj0LYtIAWS8Uf2k6jhv3w
45aozv5XgoQjj2fFID2A9ilk3eR+wOOLaH0gWSOeFTKR2j7QNE3/u43UlWO6mJRD3mBYTNNwkVlS
IAJ5RFQ+X5y2OaQ67soT4/sBRPFcReiLQkcP8q1m4IB/B1q/vorJ8JD7uWFHpKn4IB5bpifYwggP
7XO+7CKoNt2z9WFu2TJkZUQQJlhxcBM7gohzY0zNjb1zQsFO8veV/qkTMhyG55DfVPOcxRvVgRjw
OFTlI7wPvVc+Tb77lgkmRLjbi4xvt4UisFiQzI0YPs08AA4PX84IrvMKawMtB6FC01YF2Bx8dDYo
3Nh6ihZjAjgNeKNpoXHfrDy76b4tyfeuqmBsjeePxtsHVEDbbSvsgoH75T3DCFmVuy5ghGGK5fhT
yy7Yz+Mna/vULi4w9WgHRUs4ORpP+tNoDQG8l+xu4nI7jfRrXPzt0KJr7v2jJkFlmSPCyE1p03uq
p3ndHc2hKDwoAhaYgzHqhGPHB8S5hY7paq77qRGMXKBpYv2htCtge6Lh0wignIIWzOe1iHYX6y2K
hmMlwlfTXGPMLbM8OYLpsHmFQ/aSkUT5Dqk4iRoNAl6aEERhFPjzqQMbXa9K0FecAAPkm7V+u5uP
0TChtlWeYzlBdFBnOi2P5CcClg5gYbAYDp5YNX79F1yX8KNLQucWz52hCdRPFUWRX+DijpoHjAyr
4GtQl6ZgzKiZ8M+BUJ/AQ/q6Af9cuhgpIAHt23l6ctvylEf6SUsxXAFnogi8lWErgsYbLrS7eU4Y
PwLm+j//pZYVGtgKCZrZ96gQo4hhjj+vsxh3gToskjOuPkLzF7uCAlZp5x/FRnY4D4OcKl0cqr3r
TyHCcwjqLW7Bqo7wUc4RGMO6LsvqO7lD7gCTBF9utcxLUPUQ2HeOoU/f3lF9GrQdQevK0IY/aj88
gkVsnE2i06Mi+WlAZR/MNX+iCO6/He3FMgYNIMu9XAerz3B90R/LhzDXq2P6r3Sgzihuep5HoAif
LDMVaN2V5yPmeS+6eZkEMCxwCzMC5O2pG71AyfTg28bvLm/3+rZMFREvOHakmrstdSwfCERykJlB
tbsTF0EO8h8s6GY4LYkmWMeMBFq7T74LuKx7f7xHmu3rZBjIxi6gj6Y6SaB1BFoKxBhe/TpCoGBn
KjlnvFLEONaChxvaFnVIOreJikhTDJTFwufVsvsXY/XkrOw5/hQ3PU2bagYg2qoe2h6mmlVdKZUE
r47B7tqxjw3pX9CSsD/SVbQwwKwheXWy/cFuPU1HmtimfLn4kS0S1Kcm9LZ9gBtEORCpNyxoJRTu
c6MzMzlKaFl8YW1N+wWriifmO49jQ/rtC4wKuIX2kvhDqQGUy1fudOIJScNs0wfmYhnY/78D8ExB
hLLnuT161v6FZxOZD1lKrMzYFCPWF7t1ZE/hxXrsPcoYNn/nC41nJDn/vj+sXhU4OnBB4iclfdzg
qwEE4i/O91fziYG1Mk/jNjcTci10HYEN53FiH7dvfvytfDRvXaORBXDh4bjtNlKyfS5YSoaipzWB
5W8P8n+hLBr/yWG6FM82x77Sr+A2zlFKNtOIQQklnk8rq6ZLLKELxQCwYxQZDqK8me5ut3fG55Rg
4LzDXl+fzBp9bBYCJDw9CwVS0W8R+MYGgJyRmj5naRVe5kiwSblm5LyaH+Klw8TtMibQsrzS8HcF
BBgILWJoy557kK4aStrWV07J/mVoc2dcn4p3ACBF1zalltJXirGvq6QHsSXm1XLre+NKV/PxKLEt
9m1wMjsJik7M5dDO34Aejmju/mwK/Hx+5JiUn77AOU6iZW5uwCrBtS50UhPeLg5D5L25CSKahOVK
DaEisiPxhBPxKCHGmbQv3W7Av7g9OGTZr3StZy4Z4qYC6BkY0CRybG6lQ/mZx6PLx+BQdr6Ruu9V
gkWOrpjTD0iXq+jwwJ45A+ICGoUUK1hiv2lHrDin/Vi2nYaxkEpctT0eP92K0A/vR3jfYJYomtv5
uYHumzhZP14URIv7sIqLNvVSFXynCE3pemGDqKB7w3BSCHKznji0EY4bdUvH0tL5AOiQebLdF4VZ
aBM4/ABauZM2Q+WPLeBoYeD5KMa4zO1n6A8mN59l60OeVzfwytDkytClctd4TGkTB6CzIgm4hnew
aln9bxkxYAZHIYQlZto/9vleqlxdAx3R2eKwOeL13LMn5Ci3D7aSyg8EozCAzIc2S1PL8xehHoZR
HpbklFoVHoZz45NuQ2VQtbuCWr1am/tAvTogVhpYL4xWcQQZSWB6p8nnOtLRSs58l8TknlIf8R6d
prx/LJs7ME5wJfqAJZoK/2G7yuC/ZcsjrRnLU9ygh9NeZfrqLcBTRTGcIvaFMS0Mk5pZEHy35jrv
eitd21owO5ZAEPGNVlNMV9PPHaujpnsj1ihFMkBMR1wxBYMq4NLmu3PwrUQ/XV/JoR6nDLvFE50y
Snld9eJpaJU5dxXj8NVLNdkyLV0hkF6qmJNJCF2SwJ/MQzATT6mguJbe47tsyPFq2bkZ0bzjOCwG
ZRPcU1JBoSWRv8FjJcl5BSWdDGSRhZbGs9nRY4Qqg5A8P3ZjZzrBWeZrJ6u1Kbfc66221fFNKxI4
H3frx4HO3ZwjAD7CU99u/kfx+LK8Oxmp4U10CyXDAXqN+ZtgmMbZVRVNfTpJuo/iyldeE57Npogk
5gBk1/684XA47cUBDWAxeGLjGJe9w5ZFjUweUxI9M6xwUt/wI6QgLoOicuJZ/AUo8v+WogOA9Uwi
5odMOlpUIZdC0yzqfjp8Horci5EBytrRn/o9x/u7QlyNStG0BVgTFXTT3XAQLgASHqmousHWtkYa
UeULOiIZ8Z+nCluagWw5uZk/x5Bbptn3pDk6eB3usJucPostvVtkInfC4BQtW9P3PVyK1bbYkle5
F+yeO7MeOBV8dLxIo3Cl6xMTZxSovDohNJ8EMC9QwDfmGEmqvAxg+Njl0oTStsp07NQnkkrQBgVT
esW+gsCt/Qefz3S+G84SzG17S15Hsb9cbChe2xunc0A3tTLvG6xnlUSQjASa2jkoVhmayAi6g/Ya
0llu/MbXfc/gRlXllFpfAakJXuWNu9DFg4Dsi8oFdNQ+oP5Uyav9B8Rqq67C1LgnVLls7ltTgbVC
b+vIQysZVRvRr0SDlK5BZS6tJuLOKYPjS5YxwLhN2Hb+dMr/lUC5UPqlZsr2R5XeVGEvM6XRnKDX
SaRF4TOTw59ojRUwq6X5fz7ggOcsgA49tQ6aPxfc9v+BNSeJa7ToyJLPty7Phwm4UfnApdQrhPgd
m2hhTsGWXhgBbn593v8hz5q5uzQa83BGWMpzrjiCtaKo180+E6gjXGI8MvGDTLF2wHdTFkSRhLtx
ukC1/McRJCGEmkW5UH83eGD/dmHGTZ1AxcVNU9K027Vjem0i/rzA36fHiPeSM5OEFrnaV7dcd2Wu
O58FThcwZgz4UzFeZfplA2RzciqZTlvBtAlvOS+2peO1tTkQGPRJrmzNTUXeiC8n4xS4c/M6B1wt
tJVxmsickBsSSQ7ZwOGBpFX5ymlwz86ULj+vTH3RQERjrCBZOrhf/MlkPulEENpX2Pm6QgwIKjbC
jUr5fREVQK6tviZPXaR0qX/wRnCQAGthoe+vHh958o98V9ir+1+oHBD2M+Op8dqJD+tKtZgDbywj
Qx611Vu6mexSFUOGZZE3DmUZ1fUGdSEj9hT354ZRxXHshayK2tJ49NkQbzuLN6+iMMLJVO7RYzFC
Bo5DMGv5rPybYH0nWxyuiGpR49LXGFqYJMGs1guXeOUByoR+ajyCPZj6NslATOZorq5usvkdirXE
UxLMreXmBe7HYbzhx/xIPlZjRGwdyZ1GkaK1K1fFRIiYQYqLGlzHHr1l5q26b6LyLXYjsQKlpmla
zstPA+DhhmDH397tYa7VgXs9TYVEglo5W3dIKFk42jED8jXV7PYmPVOgC/UzNa8LSZ9eri4UdDGz
N0M4egyC8kqGOPOF0e8LcUlxJ2MXZYiHyCn2e7DpePOQbVYb0TqcM02ps2COVe7zc6/YJ3gtLhH8
D4/asmkLFkIx01FrwfuxbEG4X137WX4riehl1v4k4JF4l7iRthIHAlkXMyYorLiwCQrgPMUzRXG5
i4ox8ZP0uis0zek+vUoZHfOlgPGCNQn1PyTtbOf8zBKGAnh40aHfiyFOaLJGRSHUCS+7/UKIDU+I
1F29CObfbf8DrMHUPcLEyXI6HeMjy6o8w5j8Od0mSGwQttcRTJqU0aaLQUakBUhSIOQ+xnm/tVl4
XTUrXsNUeDy76XQ+JyUfZzvXKJDgKvYnBUxqnD0UC+K2XjcDXphgMArnxbbBDIx/Tfjo/eqM5VHD
11zTnKnNQjAJI42aiBqb56xpsC7oWH8eitz6thA4q3aPxW71NV7ECuMpZYkU+MWD1kP0/34kPrOh
2tHc0chPvYypIUjJatC/BycBkA97DxhV4BM6jyw2DRbOvxJsLu0FODnR4yHl7hI5gKcGJ27+G9YW
wo3S5f7ZAYaHjsIoTUDEB+J8HkEAI4AT6a1v4wvrl8iRVDLIU3nkKk9o8qOTHK1YMxsEl8ldtnhV
1xkNpxGlJif1Z4lCxymuKeLdtfi2oFoQ1M4yYnaM/4BS0OvKcLXUGI3NTXL9XjxGOx0pxFToH0Rf
pkmpPrHQttzNyWbdVFHpt5VuIUmXKAikjgFD33bbqPO0qOEgZjCEs+tZ35xX4+LyxJGjkogtS17+
P1/jBnsSktwVLNaA5QP0oC1G63N5aDcMixX7heDAexVud8b952isM44+02b9EeS8W5wdGWGGkk9m
QKOlKxhKZ/rPqLwpJsxK/doH10TIGgI3+Pe6Dn0zCLTKQerHeUFTjBO+eTmFkjmnpehrgbq7qWjD
wYXip1icIs1RYiOu9BxY0xC7IL9rYqjAKdAiklx1xNdcxU3iZ9+7ltNcnuyNdFLZnnGHsu4xdIES
JJCriy76cFkVhy1rYnjq/n5cHLzkUkhZWTAfSuMrO3J4nmCpYMIoUsRY39/B4EyKgPGgvx2t+J8P
qtLbpg1iwwEtrkksLjMpUdHbfYzqb0+ZWfXDXNGA2AT+vGRcBGm9b5/GeSyNnPxZLtE/Omzz0Yc6
A4f7f3g11Li1QOfFnaUvdWf2/UIWPNPe6tltQ0p2phmg4FcVdJx9jOlq968X5xTb4xdhDJsoQveo
+LdQgqzmEn3VF9zKChjzppEG1EY9N6kMXO6dmISDZVyt19Wo0nlt/neFpnzkhwLonnNVeW/Min37
OvAQqg0gCSVrng/X4PnMZKA5X2gzy/iwm9uWLGV1cVitTNmecue5zpTOkg2egCLPq1O+guk9bisb
EZYKPNtMMF4uHAsDtFEFOvdkv5jbiz37EcjRZMb/URRbSdW5yt0SctdP0sHU/no8D/cc37IojTn+
WNZS9zs1txTPJYGRc4iBmBF4BKoK/F6G2zRRo+BqyM1sflO+g+dbARNa1o04PlbvY/mlnMuzwxTn
tdFpj+9VxTHZeioyXtCOLtyqVcCz1LQ6c9456BB8Q+tdpSir0mpN+WFaI0SGnJt3znNLeHZucKgT
JhkiY3aYghHgSKSuS5j7iV64nWJjKTCTWx6FkOcM6LLEx+O05EQbpXtmq8ll9s12VfRfdil21tWF
ESDF7YGYBL1AGfXj1lM8qV4ppI8LKynohoXZUhQbGOoxG3V/wP0D6Jq7OjNZxKmK7Q7yuuwjRIjN
ssJP2Rg2cYZKfpahpazTLu49+7R+qCdBhYHkABcQ1ith3kZIeSVAgTtdxD9IAGJpl6v+u4G4L/qB
ZMnfENEAWuNklcdS14rrVQpa+tWTOYDEvF1Lmi/jS2CuecPDAyAIFzdtVX8ir5HWp5U50o+nVjA8
IF2RyfzpZrpthlEo++IKEACwcpk6gOznQcOZM/FNeQcBGMb2xkwwKMebniekym/xZWwht7lkaUA/
PDxMdWMUbbosO9Hj3icehXgpnZloIUisES9Pr5LAMcrlR4WCvNDeiu536WMYU+Spa5XnVaO25M+A
f1UsODGNyiSR/W0MYFRjioS0b/i9Q//KMS355CzNwbjgKTrUTs4TOABSPtVDOOfKe7t1kNyECYsR
+ASA0pGgOv9w/ogXA+FbTuMRCUZwyxiLBa1Fk50innXfOwLPNUi6G8FS96f03Q9fg0GWoYXEroHK
xJrDCHB+Pmedcgi1dWWS+ZKNOXg5yuEEHpj1Pe4zWXcSMflrIFuM5jcq6KDfYbCZOd5X/o/70rwH
jYenjErOc/UIaaTtN/up3WWJfBBwBeOuTL+qLQf2s5dhOgM54tcblEy/BmMX3mi8jRoKGYvrI+bV
DlZF6Kg6QrS3OKbTCAo6WNaD0PdZPDgMlQqs0Xt/e/5jptXGylsV9aOisnF6C2vsp8De/7HmXWsV
ID4tbRfqRiJaIo2/iia2DzCn/KMEa2KVQmOcJfZfDLK2o4DcFpL1QBr8PAoYNRPIJTvZpUA5XkKb
q9NlXHIR/DOjIGfGtjMJ6aDYAOgc/OqfYtE6PllxWEvMuLR5XeAlcGUxt3sZ8/rVQp/R7zKIxwBY
U/JbLzZKOClmo8xJ929kz2KwT9PizzbQfB13Oss7nGJoQDbAmDPvhkXC+4K0mUNfehBes+Z9+CrY
W6QW+lnaWQETDhV1SHVTTuhgkPrxHZl4hJZq+E6mGE7nZUtWVn7Hx0m39lm0oBEhYmG8mT1X8iVN
E2K/zKxVAJobpQmw6xQveMCbRughbG74mgH52wAYdIq7mkDz33aCFPmPPgZDc4vhD4FLPUD/gLZ2
1RTF0DF9lVDIBJb7siFdbb0GI+N+TsiEx1YFvipt2SX1v2YpMYdUuAGyPrQ3aLo/TOo153xIuiVo
lK2+ZIc+b8HS80OP17nUhIuh7uTGPhxnNO+J9MtscMKf+Pmy1IMaZuiLgEnJF7UMbGzQfocXxH6E
7/DCHLD+I/OVOkqdibYUyc/xXmDKZzFxhGKzZUpoWgAmsQd4mK/OPlz8QOqaeR9Rlmygjm1tcP+G
dmXmQSFnyrUbe1yTslJlZ9DtOWO2WscxhI1mlvWnG26YmfSOFHLMPEUjWXNPdcP4Dr3lHTr5fwlA
rEk8hnHjF+f+Xe55e0yzM7pvh45ZHGzBR/DUg6mohFurTxxLyoIQuhh7fl+QxX7fe0gwckevCjzl
z1EgCpBMTFhJdAsko2yseu++yDx+hfg/TAcsjtEUivVVEbz2nbwMJxKAyJZD7btUV0045F0j8Jis
PXUusNoTdBmt+2TuIUfQI/g/IShGARO9u7n/Q0CyQAyDn6C4QdCSjETTdnZtEK8u96kbdfx+wlWT
GLcgd8LqMlktA31SqLHcbshMXyYtzh4zTkDFfITwHJ6Op+GLt030WHlXcm64RRSjPQxLuVkpwioD
Sren6zwwv47Ble9y9wfE5toDoTP/WQu2tpA7+dfMt3uOwWVkOMt5xuzTTMuadwYTdCR36Y4OM//Y
8PonC8t1ZNiHy73JLdeLpu5msjXpD9QUmMyTTAf8v7fToLzqdjoYoEtwoUcNRcO/Nr/KMY8v5gfI
Ajh1KC7DQc6Hl/c5lJDQVMw63d2YyZaOLMOVVbAW0EcYZSIqXEbE1XJjBjcy0N2g1Yip6rfBU8+C
oDrgcGfHfgxT67K+oPrA00lKjxJTkUIKeMpsOVX1Da22o9CModTdO3Gx7G4logjmHo9OOuraqMx5
l7Uuib0152oYjRXwe0P0+BSfEN9zZrgovlc5DJtXtT6dbxPTifpCEBpFSZbIXkI8kfvBeCQppmqy
FFj0Rx0RRD6IMfDwZTbUeUcDjqoVbA3a7AScv+y+mYbACxUfN0ZyHSuhKHSA56sXcUf+dw+PwUpT
cij8eZ6WUiv5//r6YtJGx/lSGtIvdc+L8jRQ/ldwQF1DbdxYC/r8pEe870oEuSnx5z85ze3AhJQ/
DoURKN1KOZWOWATzfMP/D1A6UB9hCAfh8cZ49tRBoKE8N4gFUfiLLSVbi+Uj/qLTWuuRF/i8N58/
VShoYew39iadVyFEjguaftVKs0I3F78r+RNzl3pUUtNR+Q4vO2fDJQqT4l7jTxFAkffQPdClSVfk
penuhugiEvxFpS5691XANrvXBCgbc8e5/YgZsMNt+i21XtgSScuDWFj/Q1gggUo8H9cxW4VzFzL/
ztjt5XZcJz8SXNECLzLBidaqJjiP+YVj52l8D4Wi3Q+/fqQTLvVq5+USn1XWkGHXkGV9OUhzTSB+
OOPp5yJ3jPYT/ppr3/bVy9RIsX5Kauc3cAuE3gVW9KOM7fqaJjiXDB573NoYnUilTuL49xKvZBsF
gxYyEevx6VgrKgi0SJNuGcWFPcOfGMsk6Vx6u20PtXiX/ct6UiK/ixyUR8278JoXxB4MlG8728VF
gdJrO2xjTTOe83ZSB7TVxSe7y92bBBeSz2c2KJk0AMwGSAXq56JHS4ZCsRdbraxnVkMG7JH9v48a
mydxghsEyEZeS46yVf/lwPjTPrcXonjZe5rmb8keNHZDAP6WlPDzXfYAFmCT56fOxaXdVed8uoHv
mwvXHpIybrNTs4YZudCDDocKFINVDefi0NOeZiChsk+WmyPwqHO3ryXgA7JbECLdb9fWS1yoMCey
qSfWOiWHbRLoYXsj6975pyBrTxn84Rt3Mpgxx3j3am+c5MzrgX+J++LhcPGNZhYgkMy4rsI1RYYn
57RMTYKBeebjc4Cl4DwgScUSSGBxfhUv1SBEdeN5L0B2Nnx85dRXXEh+F6bwa6ftgys5BkECBcAr
coySLqyB6q/Rh46ebBe7p68fJpMrhj1cm1vOXpBLcMY659yQDJpGCKbGWUDtFOJppR2hWTK49TRj
Dri53/j7uwef6JwcCvw9aKyLsCaRoXy0jlwhcqxv7mPCYn4sb7TZBOUi/HPEjooZuvMoeLg9fakn
FK8O6sZP6+Ao1cmm/C4t1JaVqShRYN9CWRCwpLUDUOtkdyrT0zE0irArdIHg6lR5AcrFvxXtpLbp
SDgK0NPZ8LIADrREtjHaq/aozy27vt4/5MzgcwqgA4pIsIagb4nGHugSP/p6YNyxeq0v2cEXGqT/
xF54sxYuUZhFb/g2XNviAq1z4xlOQkD1nc1oEwrqfydFpZn6jlWzBkLHJ3k85wrYVfQpqb2J8gmg
I0HJ22Aw5YSfh/Zdo73DViOqp+CVu3kPVfuKTvLDSnUWY0c3j6vkRuI0uUwpVY4VbbUbxcUjfjOi
uxmDkhFHt1s4w2iZxITQQHHp8naIAMJItq49DaYrMF+OAQXXXnsG+CQZRaOaD6/+rwrlP18bQNFR
Q5VCtMAEUA91MVUd0nEARAPCb8MQcxVTI23CP3QUnIo+dMTt+iL0phEFiC2KJA/9LAYpzXBhEEkp
BIosYt//+RmaP9Wl3RiJSStItEDq0A1dgI/1L58Jl5hVDCJ5bfGnVDmDg8xz4aIQqDXeM2OkklRc
wulTKCFy3rQsp0d22opJMGvIg7wpbpcQBcPeHgRin/B9cuDycdXZrH1VZa7uyZ6FX9qscNXkauFD
Br2XW06bmyIBwnoDi/sUxGsxaRm1JeqalT3JlYFiPAUeP6sMrSGsCAy51f+Wb4tUVIZfSG54nTdw
Rgylryx2IJUJory43SjRxy+v5n32JKBopprkmUqdpgaAkP3wz2QIhso7AZ1NiayOD1oOtPqhwcIv
coutH/aBYC0+9EOtyNg1qFAB10abCqDmHZVWG0TqhGlF8lAOv5t0PPhEV76IOVI9qVS9mOW0PUEp
Ki4u+XPbgf63dCRzstwm4fXBir4MQE2jCckcFwx+H1btUizAGKvMlHPWxXqlPE99FKwT6X6JT0fp
6ee7Do93CuPuPEI4MT2jNZ7MomcAVX15Hcg/8fhh2UlEDomZVT/VTefvLoiaMY0ftOtJd2ChpIY/
87C2w9zAgu88UATvTbeFrDNvBjCMx9UR+aUb8Fms5jyVpqxZogvVqtZnJfDvybMihyTbpY7Ew5oB
qi12Q+QuZKybucqsu9N8WEHqbhwh5Fb7fbLX9zfcYXE7UPGow4uXDZv2pB07KObpFT9g3vN8zcVo
+mrAKZtLFd0PTqKMS+OwmjAjwDjugON9z8UCPpsumlmoMFFQiI4i7zMraAIteqixngSYJtS6ZGrN
FAWYWr+Jpz9aLnYptQh9Yfc+XMCXVDiAv3EmC0c6aC1P3WOt99gNoofjZ88WRReB59zTTBhkJokx
WVhtkUaoEK4c8FZiWBb/AxCB7QdV9854SK7kOqol5GZLlBFoall9VQkf6BzA+UeXjrMsQvrX/0E4
xA5TRdZzm0rHslzuE5C+wRhdDmM5CgoEC1lOwMOMpghxq2LxTPtEf4UMBFfu/j5kTSvW7jtwCI/B
t5/AdTynE/jJWEWWxmE4fp/Qhk7EK/y0UxHJLxIm9fMzVUeGzbH6SbppDLWgkDMzn7Anl8LqV8oq
QJgbYSpvQ635Afm8w8FjqKIPOx4BFo2rN7gh43sdgz3lWaJbCOQ6EYtUPC6zLA+dIIHrkp8kq4FK
uGK4Y2dOAya6rMklBhSdvRVq2NEmU4x18c+HCHpTAzpghfY/ddP1t1RSXcAPOH6JclB6fQ7VT+YO
rRtgFV384AG5mQ6+/LhKAE77elmTn2JLLAqnfCkDCYInUGHsTiBYlxmjPsC9nm59rqE3uwnSQlda
uhDAPinHpSdNA5y0fnc2F4LpAsHtt9wQ/MLYTnZTUFthrgjcFzY87T0HjzLCGOkZg5Qo1Ml+/fV+
6Q8KsxvO+NRFqeJrYLye5blZgh+JTuWCxd2hbrSfoSKrykSvbXNHd7zTbQPl8hkQ4SlQPLLcijRF
DgLQNTn1tCqa/3ttHf7tZYdG/d4A7bm4ci887iBCpxjvQK3SI4oqGIbOCsPvXSHVx3ALAp9aBVEW
Kdkhitgu53nZuz5E7Jbg0Jxhfz+e6lIxDdlZgmCqjAYNVMzt0atELNXYqpmTsQqSzJEY11Cuv7C7
JniRNPqNerpdZeZ0hXQ3/r+PqX94N/9FZrNZhTMWhxZuDzBnYmt3+o49UVWX/E/OYdDblNVmJarx
VqraWaka5nNVG/fOrTFeRxM+Dlp2xSfrHq3qRU3E9rV5yv8YCNaLSwV0SxW95aWvjdkOpcnarviG
vOFWl+qZBgaQOJq2hSrP7dy2F5nC2BV0uWlb/YL5DjY/9tgVGCBgXUUY2Ax2iR/KIyU3s2bbv6Qq
6xqFrahbWeROvzcJUiUTIfcUHWWQ9qeTeT06hRQmGoMSNO2DaIU15lH1EAIZZhDu3eT50bD+LDWq
MF5Cmgyr9K1U0j1AC9ZZMk8GtIZoIn/6jeNaczyjGdSsnw6t1bwLTO2Ppt6k+Pcm4KmEztYT6vcW
b7+GmP6+EWB8dKAg0vJOzSnd6We6vAdCW2kPgrIdvkbOkGKRBbACfJoeJ9FHws/P6oxcufNuwjg6
JUFedX4ujgPcCoUWr/MB90MEfyXu59OaOcgInBKkyVIN5yg5CoFdifO0Mgj++wCC/3o1/joTThyE
bsiuk1mpAg6xNR1tICb3Zfheh0FoCqgf1dfUaH6U6Zv6zyzF08uxLiH6JTtJ+4uQ/T8h1R5TBFU7
D3iOsB4EWv2zeeK3dg0huG8MKMb8E1DCS96pzX0xo2wBwwfd/i8ARsXTbKa5FLvymcra/xkqfTbc
YL416IcA51q2J6KLhWhbi9IMD/orF2YqHaRpZ3lW/F1SaX5vDQxJAiS507VKzRIW/4ec/6wIqGmN
tf4rHrKH8W9GcF1pLc9Rjo3REUzRRIvoaeklIGnMuZsHijMCzlj/RgeR9bfeh8flHkAXOoEBFruC
EE8s3r5XM7c8BB5xtQ0R8i2It570UuKDt8xN/NK5wTxtZTSiGsuWqQawUnEPqVmbEuJSPk9cTsps
4ZX0SEY5zwlMAcvGe0VUWU3Y+AtLgWG2tMrZJYR1zxSZTlyvMthvfJ5BWtoUwcD6UBLk1vus8AnJ
5yEoBPLOTRAFMz/WajvjzloNd3z/w3neqJQ/gdWD7F/ZTu0s9/C8Dbk3eY/n4ttsnFqFXf4g9A0A
k9zSbgYdOcSwJf/kKnL8ZXcBO5hJSjdlvv3tFB7GBgQwUbeNkClQhmjV77cDRfU0Iji9dOttBAEH
79LZDwM17SObvnzW+GxKvOzB6sKFhET770PYvxdrOcTCvUi1XlVJNda23PE8zH7dSqSjCHdjuHyH
RUmxxWGBvtxAkpk8kS8SQGndPThRx8puECcweGnW7n17eqRnqQS111a8x7jZgHpWGu9c6oVMQPyV
+d3HwqJdHytcr4OVrWH/Qopr2AJ9TSNU5pw+udFtY5M+vQjivMYXBbFMP66OfMTUeqEqwIJ6taei
nMNIFn2bqbbrqCxv0FECxxOUsOrm2d4j+YOcLk7yT0QJe4+rjiIbReDSpZ96xuwzEpaWlV1xPl7X
3fldMVHxWPYoObdGkpyNeAFlEw2GsN+5rKbKLWHSsc5HvLS4Ea2AKe8qoiwQYGTXs7zxwlgIfOaC
1LtRvMCP5S0czWVO4nlFd6sWgXIjYSzF0ZvXx/1DcNG8Im7RIBmn4nwSlAML9Ol2KirQsJb+xk91
sGrm85+veYXgLgP1F0hEUE1qp5JeyR7hbZjNQtCYdO3r6fDU4Ctihfjry8JGiGUpVZM+BkLGj/Yw
YaaEPCSOrtxYyX2nLiFFV7/K69AsnTkvwYC9lVraOBf2A0oZPqgWAfQ1ziC5LGy+9vegA0mWRkKf
K+DEnigrgsMGBlWpt2izDRghzqhMZO+xIVOzVlh+od2yrfhF72CVunku+Tf7UWM3h4LuEWUqshOd
nhrdAaYcZ3V5wAr+fP3QEPvShQ7+4rL0gSq6m/Gvmmyu1JuG3lcQzG7YA4Kq5gJ7qoMuqSDP95X9
hZlCokGreySl9RiZM6FXDQFtSROtgOrRsEOV6/A7URLffSt/NAMBRPiTCMIO5rS9Zg6Wd98Dp8J6
KfBT0jiTenLT/swBrUTU/uGhdYzsh6weGtMaA/18BC2bCXAlkmJy3Uw3M4UjZ67N3Tfgq/tjArqq
5NshunwlpGnjko51sm/1Fto6LsvrFHJ6XPRAbhicKMSwgp4sorqCpAhrkQ4H1Y5bcyfcxs8hdQPN
yOU198DGxHFcYnoBRqMIqxQLceZIRSYVwN7typAReX6zOgExxkse4evVOwyBc8i/9p1NA7CJddqz
+3a/QOSjKTBkPYsS/8c2GbeeraZiHSvP3nxzkLJ4Xjjn3y5TMHx0XgWwSskPimGFOPCe3Dwf2fT3
lYVrWFbF3Ty5nfR+1iU7BmgoIu75AITpdBq/OpaFQjvaxvvDabjC/3hsJr9QZqGUH5Ya5CjJ0YVh
mTHDNvvRNVDFImPUFnjoSkEaF09UB6QGnDiK5MMT0701r7a3FkF3EuUrLo3qm+uXqZ5D3BFeLS8M
LQtjVC2zUSCxjZp/Uj3JQ3yS8wi/h0cdH0ji4CtJ/HCL7QonAPlA2q+BQTJlgvGy7M5WhnhY/j+f
W10up6a0ZBJRLzfADG6yXQsKZQ02py2qWHDI8/H/2Mt38KGKQpXFAc0R5wwJYwUBW25jmfeSYUmz
qIrSFZpexGg/Hp31thuJQh3DZCaUPsFX5qSOYf36yFPJuSvcJxpF1L/N29jqa2rJXVQkiCvluSzj
hFx6y+Ul9deOvPtn4vJbMvsXqzbj1OR2KlFDnuKeAJW8GQr7zW5MymliGP3chKEKA5EwOS9RNJPr
TN9v599QsUE52eo5fdcvZNJe1fFgzhpk4J9ffUCVqueBaYzsMzw88gTGsQI0froNx3uRf2krJgfl
0WOb/paqcoVqvcsenfhPLKXnfOwMHif7egrxhzssRzfS7NxpZgSonJBSLixBotuCS7LOIf1o374e
zfHZWxN8hI2DimLBMIMMdTjrIg5PzbPjr9hZehVFeXX6Ztuw+1sMZxd9KsC5tLamWmZ6D2HmHY8K
irZZs/KHoBSDxtlTvfaEr/8rDo+xdnnkdbv1ZJC2u/87Y3NYyUqDeY0F50wnrXMTEx8BsbnVBwlg
lOEh3c8sIfJ4LTo1EnHNbEQzjxFHjvL8/ISkC1uC16xShHg6r3GMgu/nUXiywTOhEaRghtloKrN3
gP3R/I5/iLoEJkqyVNAhgt8I20PMi/oCrVSwFrB9SIsu9q57HCmspvGLNweJkiQcy55Mphq8PDoa
UmItnrXTib3Jz9fJPh7TA6l7RJl7SfyBrWgDOfyApyHz3Sh6OueLyuNAR9hA6Sy4R/cZJdRokA6Q
WlLKHuKaBlJYJU09e4RZI4BJoQznr6A1jHnQxOz4u9ajBksIy414rANhxjzZqYysy1aa3jIz9ogv
Gkdg4k8ywqvfdDZkliAFtCpgAhUp1PvM9E14u9be2EZp4MUCk4AXqpdnD9FRsov83ukYikdQv0QS
r8xYa75gLY6nUKwKj19jbDZ3B+6XYwxr+InCq/u/LsIzrKJCbf0FVAH03MTsztOmVmj3JXijQl7r
YdlQZny54rQfdhvnPj02ZcBikh7EqcQjYKn2Sb47hUz37cn+wkZVpE7YzQqp9H7r4bAErkFGw7Pc
TEzi4k7VKjONN/tLGtLxdSjbjclhFAuvV7Li4H1uwKDZpDzN6wN+s5XjGd+Wotvlmpn2ntZKnmn7
ShjfPxrkLNqSoeIBsagmzvbs4MV2DLgDDK6zQQCUFUBdHkrVEEdsZVMhBf09PHMzBtmV1czHiquz
HkmUXyOpz41+3gTrzn1GwuQ7szTCwpTZrAmdNGJtHBi5CARdYEywK+bCCUQZPmUSqVp4K4Uu7HR6
8PLj8455BbCpbDuHawjq9IgLPGVsCkOruAwwj2NNatW8AEQZmbPN+cI5ungHhDc/v5XfyrE/zumM
Qia7oA3G4+pcYupKL/T4mhSeDk9dFXQSZvsMX19B+MQNWQQHNmRAtOwKvcvMnPM1A5BiIHJj1L7C
QIIdTMQ/lecW25gVvdNUesbNGp7YtKUEauV6Gmapfk1zitIPRkFDaFkSrZ4ys0Dw7LUliEryLcM6
WRuMoAZf6eyAVR6DwErHMN6WWTx1CPmseyLqZbNJIueW/PIzrBChzsxxji91Q7OWwcg93714gDRU
fwhuxFEHnvnhlWPgDPCcRmJBnhkY+77bP3Olbkgz0THHstwbsHwsuTk0CR86/9E4MMOQ6C2HEYup
1fmLdg2n9QgZvv6M/fYewX4Z3nm3PlXaQe7yVVtjuKqM9BS75/qUjr8/mkuiBVDH0A9Q/eKzikTa
rxbmk7y/nFyFs/xE7zuJwpmLkyX9Q3LeiT90qq9ojllPXVF3+R7KNy8xlDojSb1Hgei7apw/eOVy
isxHwpSQD+c4AMUkN0DPZbv4xn2gHx9ex3+AICCVphCMflXsErzvC4bBOQBHTqympBLx+TsOe+q2
wVId5fJLoJJnnyDOP/V8z8pLA2Ko1Rng+by6EtwHljcRHnBz1tgCtzJqlRovKKIDpa9BtTy/GP2i
8z7i6vagOz6Amj8SMTghWj3BHLjHQTkmY+zxbm5I2nPvOQ6LitC2KjE39UndDjBlD5GNOBGosqta
omMC6pzAzo/cOuo16haSGyZRybwYnfBh4euDX0gPevxkIMmWO2A2dy8XPQrzM6bXFQ4QBMmU9saB
/mMyplnpERUaC6Vz6YrT+hbTcE23aKIlAy+Qg9HvefXd2Dp2TE5t9/snty4WPaOOGgJpDut69MGk
SGu+Mg+ou8Y2eJl5pfKE7tT8zkzfVRspu2wBlno60IM9nYQZs6NSPxpUebol49AfzXHGLw0MBlQY
yfhGTT+bdnGziKnPUy6iW2+6WSVKhpsFs2+hZ/dlRy2NsY4aJEA+SD4Dx0ZBUY+6G42O6iKOz8SK
+C4tw13WyGk0cru2zBQJjii4TM7K1xb6XSPcdlMIqkhMfjtJfguXHEapSGwXR9UG5A+ftuz+GUDB
ttoCe1PDeJ0ZYddfzT3W1NPWVnRROyh7iZV2dbOywl/uU8I5O2/cOr0JPy3F809TOM/D02ZOUgBM
35bkOZoOI1Ct8cCRUQ+1VPYLlVIw4jjHV+EwMcCdLuoMb5HHsBSFMGLvxccE1WE8p733djubor+E
sF52Gst94Ofqvg42KG8eD+PWCzLBFqfbN3esf3MKiP7kFO9NGy19ni/gdHdyRGcC/fIfuPDqtmcy
YQ2kElcLzUbK+9jjxhmd6uLeJ2mDnJT/EOwx9ISfUlg3lvsNXbGuz/znrJkzBsY6c76IuiiOb0+x
assJKFi5U2tNT7Ygn1rN/FOL7S13EIjee8pqnN+TIKhVGrb7I1LoSnRpJM5351cfKpMG9NGophi/
KfBpQcbmnlhAJpFq+DxhQk0Zn94qcZdKkU8FOEutUYWcejrz8YVKulYVvLGscKAlYi0M2Xi2EaHJ
ZyQLoa/84QAwOuRq6BmRn5BQu4zh6Qa81Tm9/XXJWCrDspVPruF1CsHHWcmYBK/uRtGqwtI8bhTM
evf5MXwJPeV8W7SYdalhGD6BwdGRHoBIN8sXLLkWHe/OnoJra6oNDIAb7DFQziJQgw3NIsBWF2O/
rZ9YdJKcxcEtlJFSA0oxl249zu2VDGQSQJcTu2eyUchY0cqnvgEJ4vzw+LZk46tqX5cW0XqIukVl
HiFmsedtOxpkhIMFyXek9fwTAacZu82P2BhC5Pf3yTkfSOsl2JW4aiFC91bYspGZe9Qtik6g2paH
F4gsUtawBbs0Cw+laX000fkp53vPtL3skL4icKYU7/Aq7gIeryYxsAXbgiHWKlaa7CUksb4rhhNI
0ByU4uFgzVYeIAwge+sVfWMGPwlTtAZlNmjpJkBKWlRb5oaeTVxDLF/7EGdUDmPh78cxGlWgbCHc
iXS5NWCIzCkUQU+mlZ2RXnWq+FGv+dMGR8CI+IZUW0dudXRgNzboGYfaek6rC8v6GH61do/LPZht
rcbZ6Beyd+ToCk167eSU+HKjdVtmXUSVPLCwmc6jDqZx+EzUJ3Y598J2BqI3JU8osd0qsBxQN4K7
IDARFwM6kgyZM6KwxA9YanVeuyNZFARFF9pSBrzryxz8k5PQFgumUYL2T95DlOlH9VlSaogjtl4Z
r/E6c91HLspeHI2BpySGk9FM1xqUBzUtRXA4M5eNTYVXnJrNvJ9eB4qPpymHRYsa0wYYlYgGolM0
uMdcUueKdakhv8YEPsKnf8EOHaCpvo12XzjolW22SOzTV7NzThbnzlntjHSSYYmxy4zksdtuujyY
S8lf4vgQpcFQBpg8YSgIctjN2fE5qfTMlfPcnP3BFWb3HVVV1lq3fzQg/um8OnyZChn3eMXL4okP
DLAbH7yJUM1dkJiPYATHzYnAZi7su2GZj0hSvi1byuuK1sn89ALSBFTh7PlxUdq4OIzxznGm9b8y
OrvcLEojBmfjf/CDr5l0S2SVlDttKBwfc5UO2qIZUy6r3i2ChBkxu9v/KHklhuOX0UUnAr7CPlBB
2bVf+wTwXeUyuFz08eMsuK3o3sYmD5gEfl1/AoRzgYtZbr4juuLxiszp01GtxNGIGXxKxCGVXsjB
YjCiZbOKYcDnwLwxNxFJsPMamuGTmmEk7aBKg7AxwDIIxlmRm/UU1/SrjJmXJjgZYcdwU4C5zaUU
8SokIFh9wm5hjw9+mIy1AferdjS/hoS6Py9uxdWUA8B6K6/RAH/OlBI2051uzsJyuKHNwxNjnnjg
qMOLGzZE/a8Qmu4cG0hu3zKKLRvWTg71Yu2+ePLwg3lrN9MCA++W/IKzfjyS+PfWPD10D6XVxRgF
q9pR/6G3nzQGTR4ZTR5Ayg9x+H4jvB/0eFyzIQ0N0siJG95nfm0cSbIUaGMAR1yMXL0v6uCPfuNO
Mwr9n5DTxYSuo1sSBoExX96Aw/2j8uBHuAdo2/bLQg25N90+N/WxnI0dgYw0w9yodX0ESpq7ZLMn
z1fU0fo60jh2Ove2I0mba9L0oe4mGjD8D/TjksVqNw0CV9juYcFYFHJQ+YES9B/t9e1a00BmZy6A
gthqNCV/NadcTkWLYxLMaaZnCMqY6EiTsnHftjBPRYmC2Wgsyh2AvZ3wcuTNG2s5UElLLT3rwbW3
S9mKms1BUsuh+G6m5rmkGmj24JBZNz3gaZAKrtWpS2jOqN+xUmhNswJEMi4ZmC0c/unM87J3Xts7
PezfQ1uz2wh0+bbgT8+bAJLQ1mFBKEgEbY73aaWT4JqcgUe/1jwsq5xqX7bJcuLNpALgL95iY5HX
9yZ8jQR1yHmn25EtmvrD5hjoq2rcjecu1xZTkvyAjaJVybnPRbQGWvkk7h7OIOhhf+jdSs0mURMO
n3+dOn9GKUIs/JkSErRxfdOiD0M/aH5nYkTteCh6PnsgF0o6dM6btrB0b9VdzyR2ZXGxAiqfpEOq
u5TT/7g19jzWlMGPbS6eDhYSGcO5acXS4eMvu8b7Z1sl17QfOLKPAM9yL4gFOWPeDH5dvLVHdEut
srYxq7XhpiczXDO3EJPBd2kW4AILYs4x1+U0u9+5Adyb2LlVZpm5Fd6hiayQfnHGVWc/are8swTw
Tyxq18AEJTSMoXty0VmyOvU0VrTOGqDlxr8qKWSKCYh3sKbxEs1ZM7xKtvbqsvVtANRlg/XL5Qha
EWoDywimzaWUP8FmUk5XsWWL45qLu5608VzUyJPWv6sRsCDrX0gq3tlnGfBOQsax3r7eM64bWw9x
hkoD5BFBBMdLhgM8gjLG5S9HOBIc4J2EITW40gweXJaVoN6elXiZW57uxh9CEUI9qWnUA2pJCmca
KHkFOVsXdIsFnigB8Zn+UZJduylN0ymprHdULdh9qb3T3RqeEV2m1P57/LO7aDJmIP0re91qOIsI
SEAiPtLXQEaIypH2rKTRUu51PEidrsTGOzVmU25U+AbdUMeqr+0O5RE1KfQ6HFvpoA7qgMyjQw3K
VCOOAo6zYSuBYIbFP+WuQkwl8WDwu8q5f95VARL3Sre93AnEGByMIuoEnoNP/35pYEWs9f3KODG1
/77Z6awfzhauwZk4EeIdjI/uKy/kKjf7L4+OSEOTxYg5Vo5ZIgE69NwQXKhRy1ddJO8PluI2lfb+
RrxSEwcoxKW8kAziKVrO9Ld5ktPb11IEStIv93N3/OlXiHMjpMp0eyaDP+rWqL2nXrJobfxDKo6q
bsX+Ob2bJLjEU3v0r6wPqySMBlzl39fKnEa672m8L0anX6+IVm/zPlFe5+jgS7bZZHBKVxCB4XFV
qtv6s545SRJ5tZrw7g2xPM6JM4R//9K1oY4Wd3m2E72rt81JZufUcA6IHZ0LKnk61Dc/s0alUbeY
BUKg0DwfNYXtrFmc6qKCwodHeKxgy2yn1Xm03kQA1yM5MX68DybQJya5ztCiC0BJRcDYo8ZvSYqM
WMSDhPw29l93i9NPCaEhTbkpvIVbvXRASouBrx9B8gQeQ3iN/JBV5KyfewS8JBeI8PkuLQ0WbTyj
9p//dTOFIlFnuzfN1pPwn3fUpKRlFYkZsxALZ50g76+rMq0gao5P6Cj+gFt5jc4JWD9ohOpWY9/e
bXwVAzjvLnWzSxOlRyD4kJAS8hYyfKmoJpUnhMpTgihiCK7o2AF3iq1dj09ZXj1tUZkM1QHvj99j
q6i00cSCEMNKEkcfJQ22oMKj2K4ufR55dNrn1GGajrnkodNlrCU2JNN7mpKhj5Yo+qTxRMpbBeCr
h1KurVlLTnBcMb4D8qQlNRgKKe7XCSXQ7ByBeL2l9+zHNAa8V8XLKqXuvdikWMhNQ/bIYZwy4AM3
V58iM0Kevh5Ld5JGuvrZPJRGXVJghqG+qG67eBi8ZjYiMItRKe+Aw8JHkRLJchgUQjwsc92ujpdn
qtOTC9hw3R1jk+tZBBL/vKNy2+eq6PvI/V2UXLYQoTMxFAq/bhG3ajG6sFnZrxTdz47fni/MeK9Q
nhKWVghnhLrwyybYCTdpLldh4MZM5CKZNb0S1ipegx444lZBIQM07r4aVHB1iDfcz5dBrTzWh4Xl
fIIYg5tUeoc+Zj7ItkyweswDaB2nKEbS8m14f34PtZlyx0Qtg2/0JQZXIbDBNzHzgdpGPUTvBBuq
jnOTZAz+S7YN3oA328sfhWwpB12JkDlgdvvLz3IXegCP0bNCMhIoDoAyHxNrEuZ2rtdwpWxfv99J
YK8MYsdylS6z6nvtKQgCA1RwYqgBhrM+kj8Upfxqe77rHlczzDE4C3p/IZjyFzchWOlsrfk9fPsM
WaoLtdTvzxF9Wu47wjZ3ghpHbF7VOblzEDybHDejzWXThlXngLQ/1VFlGFtTQBde/669s4tHHC/s
8/5YM556ybxMBZIYdrNh8PU6/EyvcXg/EBcCLVW9XrLK5RH5JPQS1fmrbD9r+HXb7WI+SWU/VA2r
9nhuXtUgR600fSip68cfeSQWHegaKEWdSKNxjjzY7JuHQVAVXcZB83PLiKLVTgRc+FdS2xI6uOVV
dVpVpHwjrcNN7uQ1WtL/yMmDWeN2X1wwvG6bQ66I15SqS/E4T2UALvrJxx2KzMkxUiP3nVyk67Tj
toe0j/hQTSKtEm8ZsVDqny6j6+TVA9fM1oJzPv/CnUdYUiHwT7LFVsKgL4BNz/F77THGMOA318Ia
6IM53e5Qr6iA52jA4rxj7I3527GR/VKRZRQcRlmgGp5k5uq15E2s5V0F1JnyLwUy3R88FDjux93T
BlLZDBon9MRQT/XkoltlZvtIKSVs56cFVHLM21MIlfoNREUp0Fd/NbSm+8FJsnkqx9jLySU2zuoK
CdWM13xZfDZWckXykrJckOBHpVbevDz/dAQmO1ey3NwtgXo+v+osToBV4PxhDVKpSO5a2QrnmG4I
qrbdHMGhAmWAGJfNh62N9Q7qn1m9McPX9Tb8gFX9o8q7Xce3HhG/7JnL3KkF2XsqgqfG4wz1wWr/
W2pn8sBSupLT4iTGNoy0ibffQPB8Dgb+Bb+coY1IoR5kK9UngO6QCm/OApHOjR/Ir3k8aBcy2P03
HptKTgQSDnunCgx2Q6tRe6SzcmC1D95deGct1ju0yhg/h0sBPY1bic2cXkzNfqEY/dj+emFiOhPc
K3AZEz2EvT2dl6PYRfSFD8/9EDzhJLFTTMlPLFT937lxdc+wNVDektxHVl4e3ZeFkHi4FA2pAJ9J
Zd14JSZgixbD+u+I/HFvZbRgIZjWn0DLKTuvn6ZWv2dJi+HbWEVIrz3G09GAzQLe3WXs7lf5TyoI
SNoc1IWytYZf7RQgym5GQpHzKKM/XPNt2Cv97C+C4C9c7oyxzoS+usKOaFbXVFfHFD38n6Pw1DPo
NBrPHOSQEWarKemOp1WiEeD2MEJStNTMZV7awRYH2xr39obQ8Lzbf5wjn51tz5Y1XxKOFp9/4+u/
ZErk4pi2pJX0yAMd9/yymI2CXTm9hI8JfYp/eTwZ6Qi76Nw51uq6GVUONmxUN8geaicGIWqTrP29
bixU6bglUuPcaXuJdERNDGia7xHYnstN3DcTKySvX734UUfsZ+UQceiTJAR6FlX5oN5phMAEagnG
B+eV5jWoz0Unv5dXzVDfdzLpRjnDdCoGMH3d/TZDp2mOG7kcUb0f86kD003zqGQibOfb8kKVk5Iy
o1mTXbKtaI5r5dwJzqg/iUNjsA/K+LFXxEn47nZ8KhXoLLBsuo6LKw15O+BAMYuv5pY1NHUpiq3h
SXcxnnD78WOQMIgqm13ni1scQPx63DEIWsrWPRDXYDAFg0J9faMhDeNzYT+/+Kgo7b0c1gN8XHm7
PBUgH5Jr4sVqn8fYqIwBuP1nl/wNY8q2HylIWRs97bnWAl7fW2Zy6IcgGiosaBWa/3vw6HGdFk1B
dn4vfSMcWCOFd4Rq1Og3B8EF9TW4pAJlZdPDcZswo33BBwL5vV/OgnQ8DLB4DlEwNecPKoJVlbFX
w1HtluugIr/bpc+1tEvRxy/dNK0Ksv8Qq8yLiulqnKkfjAJ/1Xx66zBrwKHfqCiq9ok9o74j1/6H
/fmnpVU8vHbPNgnIQVLoJ1jqmMIOR+jKbcj33diuO6JzEQmuipxPTLxb1CJmigBwOvqMpxSxfHK7
MEXnXXb1OCAVMyTRna53TRqbAJutP8tD43uNL9sfpisf0gWewPzN4xsUHsAdAehzvRew6TziU7fI
hz65cPKDSP2xhUlmAf2bTiKlDX2Ow/IKMsqvPrb6rbOwgD59G4atafynoAJ4JTv9xJgvNJXfz2MK
ZIAV7wC5vIi6JjaLg6qMoyx18yRRPG524YBL0f/QLL+OfT6A4uXHAW9Yp4d1WLwJ67PhbF0gCaqZ
jRnKEEy/I5NnR2UGHCVTCTmat6TX442Ej9idYK6MIIHGxeO4ZuhIEckmQZesgjzMMe5H8Dlf97fi
mhJ8f4lowWieZdMxeEP9HaX1jvnGsbVipqefaTnIhE3opxFpDsbmzQe7x8J8xu4nAgO9MFCA/85k
YxE0asujoxGhxnTdyD7Pr9cUDRh57EkS6aMh2FwC+3q6eLqQ8hyZyHxYPP2l+3zJrVOnlOhB2wvC
6tpZs5C1UzmRRN47iVHPDf/FZC5+tUWrvj89WiGUR50s2T9u5m0kXF+puyki2RfdXMW9n+mNBA1X
VWTEaOV3POXRNhDAhFIzkO39kTeJIcw5xYYncJUJw88YxN1MhSDxv4IU6mrCj/AGs5UoPWCi7WOJ
z6u3jZum92Qi2wl1drKrJ1LnLRv7cYli/N/p/Xx9q7fC9u/JVF3pw621TsH3pBJH2ikv/MKSWh1R
p7Sc5Ue6HdlwPHIbu7B6pqGmW3FocmHwRTaetdvPsOFXqzSxPZTnrXmDO+ZJ3INJ245c+JFyBdCB
TqcS74qBr74R7lG8jUcU1slOCc6ynnkm3sVVTKTqTROj1DAN3kg+ZZKk13qKVgTHuwoFl2IwhSa5
RuNtPUV7YkyeA225Ryt89tJ/abOYrV2NVi+2r/5+rzP4/j2q7YkW8ERmt/ySq6sUkXySO50ETPdk
esaSCKXXvbvUCp2XidqPt/JGttW2wXVX5rpNxXROZ+wAl5NncPM1GoDYdcdUvt6KeNSz1otv+ysG
C1xy8op78S4fth5pru6cwSje6z9jril67yAS1Hv0U5eoGEBZTC2BpETU6vCSdOqJJzlNE4PaQDg5
dLDJaR+hzVzBPmnLjI5fKq/Ces+x4p2f5YI6wAKNzouUIt1Ip9Kk7ZwUNjkwCrDG8AprEw8J8X1N
RCB9EP8qXLSuv5RKeGTw1knBTeFMbMOQ6KBV8A4uJH/RO+0IUHwNlUxoXBIXkPzPkYuuTtl4y+Pr
3lnzvXpsmSu1Nftq76Cif75Meua23gp5gQd0Uo0nSmGS76PsyuLrtM/aM10ZY4xDK6ZCKbWwuisg
3Ca6Ureog+a3uh8Ksuw3WDWTqLcqAxyker4AssdJZEexIkvoRiQSCZZp3WQb4kZNNaIMYcwfs89J
cXUqTgGZ9RYdRuQxePB2WlPuCUyWViRWW/zIySE3859xJqFonAhgH8CsuhZ39jWo5DcroABeNXl0
kWHFYCwpKmNzdCSzHuR2ug+GpKExcHCSKJul0od8jMWttjg3NIQM7fz/E0xiXet2YsmHH45eipcN
W5nWH3f/5gX4c7YPWgJJpeFgjrnacGqOR49s68rtryMgIs8p6zxO/dqk9xJQ3HF2BADlsUHm5XOX
6/CImzKHWDr8W0ht5QylPrPGvqAZKLOZNcxkA5sR6K/FbbvnC7d/jvZ0h9hV4HvlCHXZOsIC/8dH
Cvt8IW124DTSuzvGOPNKYj6429dRcg1pJTpM75bkTnSv68nQqTCyUm2s5VQ5ql3dBHJu6j5b6EUm
SfB7T+xKFVrOsqxPDyq7BuVE0I/ntV+6i7z3cqLTz7qBuFqpmGFD7pNeEVhwLnWjwfvFbn/La035
+4S9zp74JULaORMMGRYvAnCHKFM49QEwjwnCPdrAvosKV8klair4nbRmGRh8Cp4InroOLrfwqBsn
kpoQnNPErZqnrZ29FJbvn4+2IwdSyfqx1H+/SRD6E070EbENXefOY55KcMHfEeEruU/Nq1FWC/T/
XzKVCn02XLsCQici6sLC0cYW3M/0p+RNRPkAwDKatEdYBEJNhblJ2ToRo8GB+N9mVDYM+zWIxs0Q
AMPrYl+3+fqoTfbXb+iDnXtnN11JQD7tbvjEC89nS6gE00POBokUlejaWpdYX9dKffQ+JikcIEEA
wqdg6K1QTjamfPDc010AXiHFu9HHpTI7iEzzzsRsQLHZxlT/y3y7yrsoKoS865/zzjkbh4uItYsT
t1OYx++xtzmHEFHTSnQJRpoXFK/ZWYMdhahirimxG/GUCx6p99ddv5N8nmjwiLxVEu2xz86Rkpor
3UAKBt6yfpmT6/pW/gnCXNyBulQqZI47qFal02/sAzHKfyHnA3qJp1NmQNYkVbuRfYYVvLPoNBKH
C0yoppzRTqFXKaQqcdxJpN9+s1Pz11ci1BE8Jp9VSo9LWgJy0cyz05dtoJ3/XWz8hTXoP7cw1PI1
wEXsmpUP8AJPZusw3HYPJss1SHA4TSCOVbDtAz4YtWKo7FMqDUMMVmATGzgCNUigTj6lMX/WJ7f9
+N0yyPmPxNb6bXlhqOSEi3/yw6qC2A3wH8A5PEDyk4EQ7318OOf/W7ACWQB8UP84bkWshZho4OeU
SH+1G2E+Elta9Lkk3ZgdzZbfww7xDh1thIWfHpl8zKLv+7bSCQlhW95kJ+v2s3/3cyvtAD8agVoq
1mobG3iZoWsFy/6x09qF+IFoK8yma3sM9GchiptWrVj+icR7pS+hl39f+/HtQhaf60mRNQPEXq2a
2uvpEJ+YEEQIP6gNBsJWivW+zt08EAzdIkPC+N4BREDYYYxyGjUuyAzLDTQOtXUtNjpjUY6BesqJ
K92PnDwhRlRbHcamIjFki+EEaGiMb90MLrzb3MM1BgvMkXHWv/SzD9cyMUOxTgwUwezULsHQ0Vms
3ZSrNWryir7ACYbnwNGrXLP0cFDr5Ocx+8kKJVZ1j0l1znvmn+5aP7/n8GtHTZh68xuKZdIExIjc
AwX7FfbSgc6ZNY+UIs/Oeb17VPkyGFyS57qdilkV94SU6mjrixbKSQF4IUvIFz5eKbri+ZBowDwO
Q8z5+HuU10BtqjNjQ5VNuxm9f0wvIKiaqBTSL3idubsq5tOB23rBWo7pBnjzyLPF5u9HFUktbKa4
n+xbx2yldk07dsMofi7e39k5jkwMuKVRktQ3XPDakjlcsJjU6qxTMJxJMfg8v1cYIL1VaUnIMTgF
eK8zyz+Fkdh1tmXKozBtbYdMsBw5OqMoGAiAxfK44fERMAEqyZirWcS+kYsyhN4rXmxrZOd+oWVi
NaORSWZR9CZ6c3q2lknONygoXZ5119Hrk8evhu6W2NiijkUpJf1qU/5gR0lUtYhF+FoBD4tPX33K
mX6XPlYBO+LOqflyLsjofal6FSQ8flAckNlUcGQlZRDYFYHo8B/TS9+CPHuuMQXioi5u6/KecMhG
P5xOM/xGaqA00Wzz8oY4D2cwGSkNIdbeFw+MPZCpoG4k94Ow8A7EcN/yY+6kfgkNUZOBztQqtbsn
TwjJS/DsT07G/wu3BhToijnUeVviWwXChZAO2GX87d84DzPN8Us7A9EHj19jLFrGvYZ2Y1Pi6Sea
dpvsVojAxVEnZaBPInQq/9E2peUPIi1QtMidXFoVz3vPOYv6IsEpUoGfXTJF1RU4cLmKr7d1+0Xm
Jn77jggvH+0dRk9hZpKbTmJtaVYMuJUcqRNV1C1Iv42JN39a2fsFUr4d+XZblv92DwGQ9VAocg7u
afffwGhmLtDeKBt13lwVmlvz2j03kpKK/W8cWuJaYTzRHToF5hfXofVinXQxxQXULSJtSZtWXOOS
NYlA8/I5sBhWnQCszukhDMYVixFTIbMMZ6Xxfa+ldR9jIJJCYFZsyahwq8pOxUPaU7z3JvJWHorn
tziDuq084kQCVFW6mKl2XgGXiqdHnoumQeXgFk/6ohdhS+bvHHdvBiS+FnfEyinDaq8fEQOe1PYu
pEgkGrINO68tjiSet3+N8pGw3pKSs9iyol1/L7EQXGdBuyHXqABv7puKmRnh5Fv5veh361RBPVnh
l0YhYAljqPkcjKQ2xpn5EkdiyW17lVuBMIm3GFuqb5fbUE19cBKEh2xQfvpRS060VZWd1cyxTr9w
QUoWUDObBaFC/pI5mRyGPFou9xmOHAnOkqBuF3gTWnkvPiPmKccb7pPLLMyhS8o6XlmPe8+aQChl
WWNBRFzZ9743RM5suz5SoHqu3XtSc8eyKnEVCC9dpRJOmjA+7CdxkciAoIobgCRYE9kp9/n7etu9
0U47eCNuyv1nLawTdCKSIIRgzsnpu4z+RX+jjsP+q4XUFaKw9IYNiuv0sYmZBFGwSPOYrzvHzOgD
rNaxeCuHFyfEt4DOrpvHxB6fhM2UIXc3L4SobdP3Dnor/Tcx6yAh18phYUVbhHFcUTKphLQbMft5
7NxGzaq+78x88/2RMhfI33/nP2FcLh6I/45qh5N6COhgb79LdyRChIDn3I19YKGt/H6PdJJO5jW/
blvz+jQdfgn5bE5qyiB30w2oMKmGGfBASA8Aq3l+DSnXV2no7UwMdt62KYwJOY04sD6387MvW84W
eTyyk2J3DntG06N0kfRtwnuiyUPAWHdT1J95nnsRy8PL3tWkuuXpkCiwB56hJ708XvDLp8yWyVGk
XzdYM+XZexDNJHZVsbwTjK9Y/Eb0qLFuuIoWv2nfwb8YLfS0fbVdt2dAmB1Hld7uC+TIsGYIhBbe
rAsfirv6RQ1VETg13XwFj13tcTYzLGw57l5bFAEOjIjaGHAQTSzE8yAfqeHUs7H+Oh1igBm5fGiP
W5QJSce7wEyMk6u9ZfZ0GEK1bSV9lS2si0OG9FMe+kDiNZB8PWjnDOeAJQXDqzJdgdngzcDC3bu1
s3ORiyGU9rT7fWGCr7UGT1lItfia9jnapeL08jIUQ27GhVRagDALXtErpnBLUIo6GBsP9FOaYrXW
D5wP6gCzSNvcozt8qU7TAL8Kr9UshMo5DttTnLAUDJ18vXE1yLULTaSCOJ/sfAZr+RomTwzsP867
BT+z9D1gpCvVvhgsqWthCAzrBGUiaBe5uMNTgjb+E8zn6BW7CRAmKMvI7m+QqISeU8iNIzBz72x/
1BycR9zvCkGN18GtRR6Kun3Il/DpT5rUo94N9AY1MtZo9IG5km9zG6MoaLP6KJOP+zqkWGAMZCcc
ygE+TtiwTpw1v1lqyGp1UBoe2HYVI2+67aAYCs6bg4CszbI70GpHwelekdgGnMuBZRszDeEL80xp
ri7B2acxpZB02JktgZp9YKe7AyjTQimWAtBGv92jAC/j1PZR3EMkTOHEl2exUF5n5UPhKR+AIAKL
ibXPzkTZbWRPMv1OzgKHT55VLrRFNMw2dbWh4BQ17rUKKFxxiCxRpLPQ8jjz8/m4HhepzCYPA03C
45uygL9KwuAlROx+DCTLgYeT9lIcw5Pe4ziZq3YPosIxxkxdKOH5/meef6Q2GzzQgdHSldyPsw7k
gH4rqnDezzJhiK9S7lC+6uq0ih/N5yXAa+dEBqCwtACVadMGzSp/AjqjL/FL6XJwF3R1C5ufJVc3
rDVjCe7IHN1kioEggMuhCcwqZiXJEDD8o90uXEwWRDILi4mVQ0FqwzyV0aBK6WQHgAd9QBx+8WTy
QCvxcWrbG6DLZZVuch0bcAC9CbzJhhuYRMfO+sK7OMyb7yVUdd4j2NCc0jAjlKtsu6LI8sb3WVIU
sZ9TJVxVM/W3X70LrUVCbpvDwxmUibaTQROZq4lak/q5Cuf3yeZllDqIt9UEmLx/glvgYDt8MiaX
6XB4v7MgbuAmWWm3pgnpjbFG/benIWIT5tyFYuJ6b3HWHUxTPT450/XSm5+2gqvYr/I3De8VVjTa
woqAfGlPuyIoiAk0N7B/q2drTfGcohSL8t+sF+WXDQ+PX100Rzaw6s18pFVvlKArVroZfoW1hysD
5zVUk7Qo0iIaDnkjj6ejmmjaspzcD+aDg+iYKZWO5V6V81m+xdstZFjiL7YlSn86gyi5iv7PQ7oz
mtYM1JcarM6hzHRkaCzHGOGimWA9IRcaal/NxTztNsgkSl0ZJQa+X8ZRTogn7Xhxty1yK4uOtK6d
3Nl29ibLB6XONY8xBLbNyjZizbkOc6fYqPN8vSexhuezUwLrgDbC5N7baQ8E/7siKzLjdoKfmY1u
tnci79OReovYYOTovwig2VHMLgzZGgtMCMd1THulV7maiWr4HRYOcvi6kIcCrivizu49sxVYWDtv
eIPjPtKz0GZpLXds2orStnfYn5oZK8+NsFF7biqZP1p7V4fcDhiTlc67DZPweDPGB6FvXtekY54G
Ub189gtmIQnox7rakSY0WFlkoV2T11HypZ1aUiwq4M44MP83h4NjCBq50suvUBNUuxZKX+zAlB1d
1vQeIxfh+hOH4XJs8mXzo/TI+ZgjxQhtBmSJ1L9R5xXf+M1POF/lZf8zCw5JYJ8oAYUfqbGcvt5f
ooF7tFyfkIJtRsdZC94u5/FcQxgeYCivamcRanrpBjUmTazb0Mt5w/fQceeTE7uWGS17o3LzRATz
NxLFPZo3rcEdnEwWkiW6NzcaEED5yh7uZYC1Rx+a+azrpfnvyXZHCF0zDdV1tjgjSlWUoZYrXfsa
QNJm71sDs36RRghrRhCXQKesM9CLUcMu4p5wGXmTC4hgS+jaylDBETdJwFEU0AhPBAYInPnvZcFE
C8DuuGAJdKq9LDzR7IT8N6vcbHrtAya4pR74RzUrR8raNt7TgK/KLdtLxbBFfzvQw7rlQ4tznj5b
fCAKaoWGg1aug2MyrkO6VkSth5GJrTUtVhjD7a12j9YhQ4U3NbtjhNH1LZUdSKyCZW1ubrHJ4jZw
8Kcob5mtzNf+tBGwj4npPCM3d50nXv0uESVzvQ2qviIxbpacWLXoWN0Fitxo5Kx2q05SM9EwnMKI
VtlneQsBFnl/3tTtJg+TCmdr4m67tBYfmh4Ix3IStBULOcl1f5ZNevhbbR6KNjKXikh2+xMo50wR
iAie21NKqThRjSlTzfW8TObni9gLAkObZDZSd6OoHUvOxMrWyd96KNh/MTd95ELQ/InPXRUVgjCL
pONp9DiovHiXGrX8K06arqYUzrJak+roAiy/ityd6iCxCBOK7TdekgRZmHlJhdx+MkX39Bj0/KYI
KXfX3HiJeipQA3cFpxdhTrzryGpj20Crm9pGCHB6xAc0ZtUBZkMOds4gJIIIv7MYMgtL0QiutF0l
nSd1DsprbV0xy7Bake82tDtxs7JV2yw9mzA+ShYboYwZZzV7sLn4mL4Ll/eI3j4dANanRMkEss+y
Oe0ovcrkGL02+wpzWoGnxDeoR5+niJ4vCp+8bHFKK3c4WguCTxIL6NuEKH037nY3vIONDJ/HDJPn
KoSdbR+8VB1miaFoA6Ck1pSxk+KzS2xRfFIwmdFcHaukeBIQ2CpLKa3IohbLlQAk+wHoNqSli/dE
cjOXqIIhkNPTRL+LVpVfTq6zR/iiWOwo7nLBUa/dGeIIWdC2H8EEOBeNs13EPTVlVkRrJva4pCr7
CxubZJ60jl/Hpag/eP4ymf+BRaGzCmGiHZy2/iEJNOwu/t/f8Zdw4al8qD8R9ARW9sLJJT57L6uK
4/DCaJzraR2c7RAsw9j1Wg9ZvZRTUMCD2gRJqqukuUaOGeaU+C+dFEl4RDf6KFdWvXgyFpr/r2w8
8jhYhW6Jo/IaDgZeIL2IHqW9rBmDdXdAW+fekN32rAimOt6WFuCk9WBe3r3vMcJ9rCdR56X88Er0
58qZ68hu4EHWYQJbps3jaW/Fn7zcF1F+VpDyloTR9Dk6HWOqkP29fDPDtnQ8l2U0r1gZ8rzvF8AR
NAw9ofK9PnolZfD7EIo/BIbgVqjU/wBvtjNCjPHdwrp6oRnGTFysA0dQyLndxg5hUHtsKUZvXCG/
GaJM9Qu+5eBH5Ymo9+jV8TfLRMMkU2yjCSaLrkjhuIKXkb9XZn8fLdOmGIAlWUsW8X0lbPif3Itw
2GRk7nP7fwHKQpjbzO0sgvLSXsRRFueQdbYC96HhZB5kVlofFbW++Nse3/mILuTEdoiy7slkLY0w
lo5cDU3f1A0joiKtLkWrbx7V1p9X07FBpkyZiaIz+dNVwgr4BZDHWl32WYw+Z0vithSMv9DWXkB5
tOYTPn4imiIFUvagNX2T0rTImjDQasgIp4W7aG86kuTf5dSgyeqokdSCKo8BQqmi3/xL1ekS6WoO
NU3n7yueAhICR2ZldhTme4sUjMQJdJ4ti3GjXcUv8Qk2vnpN32x/1L94stDOGwXY0bO0a/qn96Vh
/4i3JB/qNEATIlpjBVXkDAv32L0crqMySHjeNu6/nhIX01M9vaiNIgH9IrEmEawsy9Wm5HSIdM91
rp8ikOcJrCKrGgYdQwK1hg+2PiYF740BiQL18vwtUjR48gxwLF8YnNujiDryemz7fczMHmo4p2IA
1lvKZDtN4tqjpelkVMgcSEmG387p5WsagaUxglPR/xr4umFiDUzykyRU/enfUvyYofSLEHaSnmW9
0ssaACXyXAD+C80Yr7GLDc6eayN38HXjvf1NukCB0CGy0LRAx8v4orekyHNymHbbY4l8/zkvC/jc
L+jXeByw7k5furXoQRpCy3OxQLONAWiq1UaKa7zepsfnDMz2o9ne+gYzTR9w8E04u4L49Oi5oKmY
gHzGXe5jQ7fPmlCwzl8gaWVud+pOnPOP0Nh+AKrgG0a85D2hU6A+ham8PXVygynEHzto7tmr391S
RGB5UXOp/13reiDa0pnGoG6heJNaKpb6S9M57H7jcWc6xFArHVYoWyIiwdr/87IwnW5dtWjunv8z
/Z/kZLO1lZzNNK/ZG6lLKSujIBKonwM3WZTHHht1eT6lxcdYhrwh6eEmipBTyPqwQB3pOWW2xVN4
5wrOlM+o/Us9RofR8hyio26u7kTodHFbJpziV0nGJctEOoD/FjZMfPp0+FqxOt+27oqAtI6RR17P
yArF+22P08oaob2jZ6a3Cm2eV2K2VcMTAf4WZSiSHqOmokMe2ZUJhv4XFNDwKqm0EMcYdxkzvCdL
tKtbVFlURa/UWblTaScnwldFzKGzP4CaNynBpFUu7dzNbfzAWGUtjdCN39yWaNwHzcrZ+Ka3hRCM
Wvri44KPvz0Mw1eJ+yPEUqwwHG5VHGjLbYLZKvMFOO4y+NXxcVXj8uRVy2ghlOPzGvhOaVXbclue
aRwjTBkv19u+x+lApG1HKOQxG1/tiQtq/a8beCJ5tOg+YL438e3hya1uHGXnPw/2TfLe63A3SymA
PJgDdUa9vyTP4R0Quhjs0NIu71Yr4//E401Pgk7n3pCrG8xcvu0hMdgxJFNsalvVZufptYHcKNpM
6VMEy/OLRUGQEVR5/GViDmLZkmQ1ih+pvkFW6utinGd730V6TuS1PH1c77q5OJYQdiMHbSwlNXpZ
pIRTTZL0PbV9OPQ2XrKymdlSwLO35cAg+Ws+oI1bztTo8PrrSaR7empnL1F0ucDZu+lFmHJmCyUD
PxQoTrF+OPsGb+owqfkIpDKqmN7+M7ULiWyup2JaRayyXy+W5yVaJHhrAA+y6aqkmdonKx6xP5WU
1vMkDrg2pkKMN6/8gnUf8z2BzcOnwAZkLf71T0Pe9ri3VLMg/ZuKI3Y1B30KBjLUDZGdLmvOTNTa
GHHmNVwQymcLbVpuRDkwxaL778rJuPvZfrCA030GgyABdbi1qWpY5Idj8hyRWgbHRIJ4cm/gd97Q
mL3SAs5C7etgyGLb4pwRck1M4NX7fC6OVirhs2zv11df4FjktArri6Ate02TEC6uNOH3Vftq2S8R
8cptxS/mUNhUPFYHV63CnHHIQ05H+WxLsM06Mi3YBY+FHKUBFWVcgNoQXFvFgh4AhO7u7GsYpwyY
tI9e57u6WpWuOEN6ghYkNw9ICb+6zIu+0nfw0Smz5RyYjc0wy7K+f1AFtvOEroR4Tjy0V7sKnY1b
4WJfFArReLcKTzvmSNHtRIgAZImAR4Kh1rCGYPs/9NevYgi97BMU6ySNJHLlVkIQnv+cqFwe9HXR
W5hTJVnxFZAqJkDzXgr8833s8ltBbAiTfYJvoT5tuICojEKMhnfDuoln+iOX5h+Cl+fVvGrvDS03
hEQ31fIgRZhT/Riz5iEB2LghFg4CK3Wd6iD8+zV6N5PCpHC733impVQ+W5uXuwLyJHAvQNma12Ig
zwE08MEUhVBTmP95X1QZDJ3o/v5emo24BaNiYPhZ4KtxsUHfmU+s2TkHL8hvIa4aYwJu1aP+TtJP
zEkJWPj/y0ahO4i7Oj7b7y8ATUFx7b1BUEzm2l0dvLLzdMUOWQ+FwfMcOxf9kjBOqKUrBGRM4gWQ
wXEgd6KWeN/FHyBRl8ku/1KiHK2+ijK/TD3pCDWaB4EjgYcLn2nMtReow74WqRDA7JsXHz4xSfk2
vmnAUjDQ+occHS9iykdWjHd9VLhExfVs2XOjNgP2wt3ZCteN+ZwZqBb0SbZZso3AtKfng3cSdLTA
sNCW/KBEXuZ1NEiLShsgsDMSDDvI3D1m6fL3l4LlD0k4KSPUQb529ctf3Ype28SBuSoY6zU0VHFc
ZHo1PbgetwIfHc4VFUSH6Ul6wZjNUUmlS2Q2Lq24CM+Ef1857zh/hnZCVQgxrfdQcLgHlrKwIquK
xCxldj68gKHGugrO8HgA5dQHCVLthsto3xSzk4UFqRtSnNbcEOqLT5d1ab7eO1hY/56L6drtl+Xn
R42qrBFFFGZ57B/MbTKy6kmButX1NKWSwK9cW1r+xeiy1jPtlk/e+QteFYfCEgwH0nzM0J6QbFtY
It7cV1Nvc8IYUV7jT6fCax6IfSBzXAVkyrIyNOXjW5SePkip9NCf8qzt1SFGUq6alP7n1GyS+/hE
qYp9XawWXRcmx1nkOKI3e8W98hiQCGFs3EgNN+zevj7J6o7RRnTw2RP8NKAMLSEQLNgWnMwux0I7
6uBT2ZXmAKkqEH05y04OmEK56kvyYOb465pVRIl/tdeA8jb3ihZasybhnO0ouR856IiRbe3Dui+U
Y2tW8BMGn4HUvhWU+D3xvXrvSLcfAr5KeHl81CSSr8BlAfHGgLPF2RZaC3rev8Xz3eX2W3thVuAv
z5n8lGHVwAHpr4gmFQkYPcwSnSA9/Q74MJj+XTkclZEQKnDs5NuawhHyBdHWu2cOtYwKiPtjKdeh
MSsr/pEA1wLycA+gFgdlQ86jz3x37NfzHQjfQj3R6VWUHFDnktrJJk5rrfuw3A8S9ev8fWps0EEm
j152bxpSobFizyMtEvsODil5jar6lZJEFmXPULWtlGEz8Xf3kHNpoKJLaPaGmMkxzMxasH0JfZg4
OZgtR1x2YSPr0f2/AjoiTkl90tlxgu7ft5zFN3Kcc6YMbxU8J+1Z1pPLzWqpc+UZHRmh0cIEMg7K
Zv3lLqrdmIXdkDtsADEUeQffQT8jpOFKqw1Ufh8KNcQZAVQHCtiClJ3nbge45LcVbBQGt7QveJDQ
Y5gPK2Iv0/aR2lXGR6qOZXT0OSnilgBniHfAfPMIozLm5OPucbbgjG+c3tckMZ2uVK/xnIcqxwyc
A65ikzHbMIUZHLnWyOQfwNs14HyrtkaZcRMmFLsero0l6fUajuCT9zPmp3+C2VAf0Iiyj6dNWo7Q
6yqwGeD+2Ic97Ll1XOM1zv1vkH1UrkTKT/pyd2k+nYndmzGJdefq+0iZ0weJwYajG9VaSA2ESalG
0xw/fHcJs/gAt0DhlfV0LPp8kyHr0m9HMUKR+mqc3srgw/xBx8EIauG6tgxHA5+oZwwDBGnft5EL
n2D0q+r2/aC2m/B6BYmGPOZ1zkQMqFsDPrYX/uTizQ2O5/6UJKpA0vUpFaGDYnPF93sn2s9eqplW
nk5dzImp3pqXRnSjpWb/Z4jVsk8RbKHIm9wPsX1mV7dAsRlFIRlTphU+l8pz0bjONTVE2NAhIwcb
ih4f+8/1Vkw6TsBL9NfBAAljxtNUh4Vkn7qM3hp6JeZpvYzFDELvkQIoMrFMu7H6QYgcgjz0DYRb
CarBtImtAnoGmtZk+yin+g3c4UadIBBY1qztSm5EWQ978tvrjF/UZG9/Zdy3/oqA/Scq5CbIefje
XWefqF2XMdYJwwG0ck4YPPtUfI2GmfRh4dKX0c3b1jU9tB2GAGEWc5QETBy0gW5GeKIJ5EhlO9Yo
BNYtNtNTUcKWXWmqdOcDdOy2C+RaxukKb9b/RIelRzAr58MUcKuR+aV3s8G3dFAMFnwLuASsVJCq
oHSdSTifkXL8jYU50g4+tL9bEi84ESpZ823V+8DFqQDBig8HasUhzzFzePlP7V+qMDiJa2jRLW0U
mlOuH7p7M4DuHxmFmupRHIit2iRwLW8T8ArK3uK7VZ6Btmh/pVlRV+M/xJDWTchCZAXRjbrwfKCc
vAuHq+oDBnC5kzPgDK6+x2B4hvMoC3+uR3NXekMy5W6oSkKby3j08kseNTadJ3K6U8FxTgwvf+9t
GU2D/p12wUsQaife1kniFYZdErl6HIwFSJNuvafKxLcEFWaAWiVyRVP80o8HULiRDqvyXeliB9V9
NmKBByMuq0W3PljIMGEACvJCG49vSG69hsXNB0p5ktURW338dBtKlABwYmPKVtrTJtTNAPWRYBeo
OkCaEjPtynH+kKxc0wsXKqqOxkwODBD/JxEb9mn/+SiJHJpk3EoIor8jbbR6lSAgp2JSlvU3nBTN
LmGzj/jyVsTwb+NinIjE7s/Xminyb9GHofF4tnVsOlX9DwLTTdWAX/c4SqAt43lU698XVNNbRhTT
oU3Va8rc/iEz8ukdxmgMMX9e+UJYHsyYt5XuEMlGrFenStvIv+WhKzw0PesGtMRBBQo5Zdem4ZGS
cNKI/t9YSrPbDsZjIpgAEAFs+UfMkAtVcUb6y5ycPIZRpFzr5I6ML75Mk6EWBQZnHfPgDOP90UTs
7+a69LrLrm8QU3ZFTFL9Y0V/Ks94krulac2iJS/pxCdNd2qacvXiVzz9gVdhcvHK8CUjtvWrazAJ
UaDKmOa2AKDrzYogApW3vjZvdUlghIiBayhM86WZb+FUznAJIZbl1yVaShqtGi0cHitsiWq/EAco
/VA5MdCDnGDEQbzNiWINEo7a1v8N+yKjCF+a1HIIOfxvo5o8w81bZ165ri9sXQwSJs8hKf6xXFxn
U4HJBcMEBvcNgY4i2fKxwc9nC/c8A8ylatplWTNNdEAPujChIHkH5RoMFoZaqyolLjo5BwAFMfwG
W26o8Vvbq7s+Cj2JAqy03vuoqTxfin9Qn9+AJMvBLdV1Itir+RWK+MjIVKMN/+EKVEbw2MBfwiPa
SmoZVNC4C4S/EzeA3qYQxrdujiMQMhyiZRTiAuU5XfFdpTDKam/+nIa4Db7ZeiJNtIeGcXCmW/UM
54WDvKRdLUrPM0zcTDlqgAJpzd5oyMkJXt2gpgFoe+OlcyGiHLl6Tc6WO6HHhxd94RnX/UWci5tZ
xhTihCqrUFBJHKGYYcTosi0h5m1tKwoCqTqFnd0d9Olw8w9K0tUpu+b1B2mXgCU6RWCSLj6XLFTG
20XS0h19myOZ1EFclf0eJMoQnGCXzrT+oaCkfML6JsZiQZQp9ZkrrVoESytG++J6Gq3w/glE4/BE
0lZTCslNVJ4IeLV8cGtJCYimUUigMwHSfPZ2NXWZRFhTENnKfy7ESsumAdvDNVIyj+oQCPw8QU7z
NVOKQ4rJkQNDlkwFHFe8cF2inG5q4rL2eWfMN2fGs+yD+w0vfJZXmPOrw4nf2urb31vLE072KVvT
v4NM5H7GGwa/W6/Y2N3CT7cXXQRgcRZxnGMDeC5I5ZTef7f094L5HIQFC9s9QsuEyBS1rOnjWwBD
0caPrmnkzr/ek6R2a24vBey/pAlYGaOxu2dBvd+0nXxXal5nTvw4KZ9xwUayGHrI7oeyqi1MnqHY
dWFjlMEU+ZT2YEW5d1aYtvRBaJNpBqCplNKVsT++gGiC9dNX7tCwO/b68JhZCxD3K5rB8Lw2npj9
+5/Sb6ZC50hHzKjqd3BtNJdh9Zxmr++bdMiq7JYUxlSYakzp0l0haaDbB2PWv0bV+C8kQqmQsHxy
tJSjW9/OmeAv9XmHCpsjTp0JkNNNOt505j/SwJl5pYxIAgggM+f+JjI41NmMPX756HvujYZxdqIw
rocOPuflkemMxQmITma4uDAi97Ecu2EvScn3UFav0SE7DU59ghCvsS+4gS+NolrbHYce564fBo8p
TBbaX4ZnHRrh7kD2SApSKe1FT3d8HSIEH1TfwECfg0Aialg3V6Hfd0f2FWZAKc1dKBFazJl0+XvG
rlUn+oRAEOpSm2KcUAW5Kz1jBRrgqzj8ro7U6a6Vtkz4g9MKqCHfJ1kbM/exg05ICQzojqvqNM60
X95DHS1j4YQ8mBdmV3Cui8syPoNP2uOQaWwLPkVZ9h6kNGsCaVuTC9rjEeXXcURVx1h8ENGXO7Eg
lWMyhcO3mbgEWAkUHWktPqeAC5MBlQsA1ywefGExfxZGv3mr0V0y/62VwN1rO9kehRRyxQNm8QLU
NIdGQ+PNqb3/OclW4QXFvQGMqQc+vzIVJ1V+1uIhcyRc5DvVlNvRHdvuonALhHd62NYz9bNAsSg7
lCN0dHDMe2V9t/OyGGqpnbFOgd3a9UcxEfqyrmjIDiz9Cyu/kM1figCgfmH2F3m8pxyUKQukd0BL
EUiPFHtzc/3JPgpFE8omfgiLccV/3zpQ2Jv+OfXkgxfvvs8PWefqX3iiVx4kKhrDqUL57V2e4n2d
B5WD5cyQp57rZVS6cZODGwDhlKHR8O0ctmctQS0UwxjN3ww4sJj2sxPLioOEQlQ7WYA7jmZni5O7
DFdiwbonSbVsXP19yf9HnEOLum/HPxzsXYMx5pObmtU211d5qURbeIn56aOXF4lXD7mFKvDOCWnL
Ydaz05IFrrRoIh6FWrehnEaLXCY4Ad4x56E6mzhccqdzVR2VNlt1Bgsn4kOald5POntAylhEZIc/
TLq3ZrUhKtgWTUU1Vk7/vMpD+OlNlvqS9WwZh/1yRHFHP+G/kp8svFlvNPpXBw37/sOZUa+oQpOt
NDsbVcpu8G4Ooee3qMmMV78gI8long0g2kEHuvQ/r6lhnj4bhXVDM5wqAN6BXB5NfGcnMvWe8Lsc
UUY6otg1Qq8zxeeKGPTLgq9FoUPqfAXri6hGlFgV5pI9go1jwOhJTosAohRrPtUrvKyc5AZHYtPM
+q0u2LlBtx22sjn3RIsVm1avEDkRQyT5VETNXhEPSEU6ZdjxMhjY+NPBVe7eXoSbOyHK84Q8tDih
Czjax826Z9f1t7KsGnol7zDbXpMuE9s2zzxe2Rk6G3t9g/cAfStBDSg+/X7h3kaOjqqn67AbwhCQ
WS9Uwm1dm5nsmbsbziMFULIMT1lDHrtM851I6ORp/ETa1cXfxmcasDJ8W+Q65VvfPVGrjvcq+DP4
1EqIN2jprjhH9H536J8gp2mLsntAX5FtYxoFvUsQNbcKcYRWzjG/JlzyWGqw99uvIM9M160kItHr
mxvsSTctut87BUCrevFQrtUT4/SYThXppKkZ6MZoL0dHzGjjFpttkIMYx6lIg/Uc0h5NU4yi6wUO
reTOiMK39cP6t872/JLy6gZGM9c4YSN6JFdC1vmxXeygCEhIYzKCSDjlCxZCWzpSTPnbIMhilERK
V/bSuvc5BC09/wDBzTNxrKW16r/7aq/0DXw15Fw27mae42qos7c9qqpzlwsSKSc8e6/gpgd1u8+M
wYSv8duxYeEapWJd4nXDOxDjVypIlqu9OSupvx9op8vmGWlApPxlnmBLM08vDOzXzdKUF6Pb1XU/
HIlcWfC4aQbh/dtHgEIfnATNBlteMzqja8uRFRot77ROX5wijzY0sMLH4VVIkvMFQO4apF2M3mdb
/AWvDtw7Aei6b3yO1auBWTGNjYzok/Q1SaFK1ExHTl65DDzmO1ceThgpVGC7Ye7CjMEkGbShMlGY
+2/TP55wwFsTIrEBZYgAr6puVfoQWuPWpKw3E7HJvVuIONR9OmryzKXdpGAvL4nS1Psv3Fd7X1Ul
YYmX2YWPDq6d2fcd990zEUV6y+szGw2B13JWICW2tBcbqnzzPt3CbTb1PlbO037F8/ldB4+YvoPd
QnpbsYWKFxXCBBI7WUlYaE1aMeRUpZj7ewkBfdAirQhmuI2sdBNRHehEvsZaxjl2aaiWNHoI+nmf
xdaYLAVRWwSga97uQ1hhhuUORYj+15iT497mlNDJvlb1JCoi+r3B8N70awctrTlEbYNujZJzA3e3
Vi4IKKHjtl2ZCKkGyQIDQJJtssseayranXD0TdOlMtGIRlK9h7qRVvA3YFi24SNFfu/uD7JPM8Fy
WOQQi7BV8nlbSdfQBefiD2m44fANgQItr8VicDKgXVTpKSFFuaPtnZa/GovWifmwLeoutNMeavdW
JbcXkbeKtAZBesVhLqgEQ1DdHgHCWs0DbdT/UgHoGgk/YLL05LTSiFj5E2397xiE1J4FYxcKmLHZ
lOaVmgFq8qOd3W9eMoCDEgMllYDK8AtPqBO029Xd64iWcAxT1O8OdTtfkclAftinZwGzqxfJvs7U
b+/vCaDKBr+kNIDUZ2ywIuBICFnS5gim/blZFqG9LBWaGBma6KqtXkHUdkvv/ATg9qXPiq2cdY86
Cuz0cfpj9cMIeHZcuccHzlkVf5qmaubaDNbdIGshngw4nPGCtbKxEFh1lpJO/CmbJNJ1sLb7Z1Qb
d2NpEBE9WpPMO/mlzKQmcys5S1DMzuWldlgzBrz5PnQeCpCiGoTq5Vk3v/q+PHfUjHsHaAfF7OJT
Vh6JHd3C2I3ibVr6Y/zO9kXUDDGC5depEVKFuliieFX7gXnKQiRp2g8VU7X9quXkZ5pIFsuQg8ZP
gOK3EkP/11ThZxla4q5ZExI7rflDyzlCl2DRf4F6v5DSI+Mn8fE9gSeQHUcJt03L0mQmFaTckp5N
NAfKrIhtM8NCjeo0uAWMkfn4/YGUUClh0YNEgc5RxI0LtNDPqjjwyIYhR5ne85kZmmuhWhIkURfX
P00fM6Kc7V3yQyXAwCc+ymj7/SDp6STdrfkJH50ORaFwA49dHrKU9vfVOMr8lN/wtKs5hyzMTT4f
2ybtD+dVW0utr5F8eLIi29ahI9lBIoMtTxher8JRSQpdE1qm6DmK2Mnlh3AYo3DW4jajfo7CSKS/
FeAWyoOnzAiO3bcF3EO5oqSofqVOkfDPgnugf/qlHGOw2YTV3ShsXy25BmcbQSogN5FM6oH7fukK
pGwBT6UtZvmv6JwyBhx/Twcd82Hb/VQJluBCdrpJHlNeZZ/+C9U0z0QqCbFsYmWrSWr1Mn19q+SM
i1MJHQOa7pO1+y+e0x8pqmXLhG0RZfg8ciFcS4NVZZx3pK0qGzz7us0W8gXI2meZChnU0j3AEvw/
023BoNrba68mBRFT/NLeEefHD+Oy96dx6/PC2jFSFPHck1EM7h9UTB9iOOTQ22ovkOQky6Mm+xbx
EThdupNpUxiLbZDNlt+T9X5EN8IcFa2hCKW0odW3Bzlvi7+UR64kgIY78qGt+di0NIWt4at0wywn
7H5gHV2tCdjNTC3nCXiWbHfu1g5WmY30Qc47HCulZEUP1E6H/fMBnBG8lFDHfb54C1SZSw1KzJXS
H/DLscPWldajb6vE20MZS/tQnXXDaSvJdJcJ6VlfFRUU1dFhtrIL6oZmnEOsW3hrnErnSe14pcCh
IIaiUOVsOrdyoosEYvJCw0Wcfn2HcRtaS1AkKwlUTgkHUJOYTMuwm+zTIFON/Ttwr6lHNrGln2N9
bjeDwHeqIXFYHepXX6XMrvjgc8bap5Xqjzk7Dx8H4MJsyOTBDegKnQXM+BR3Ki36AEmqWDc6kJMf
h727FKwPtjmop2SBGYwFYbx9Ectf4Ta4BFPLIwCbZkbfFRZj7ht4xkp8UKstkhH+z455IBeaFzJ0
IKEWosAyTFk/pzHyj4hAwme9ReZSuLsKMJkagUcxmDOtFzvwF6eDM9yppUxSZJ3sohOqYPyedOfp
gqoaZPb/qc3w3I5wSXi1ORJ+HTvSPjvWkE2l4gAuq481PEThjxBBGararN7+WcklxhWGjF3Ga/O4
rIIGAxPhmRNo+Q22V1OB0fDy1XX0P2cIvv35j857x+j2llkUCeGjiQJzgFKZNlukBssK0E2q6MUE
jshcWB40E8VTAla71rST89TXL6iWVojfEOJKIUXDMQtnUkizKlN2+aVDnlKcLyisoiI2RZXdhlX9
4amskWD+2OAJp+yDkxr0L6EOilDL0EN/R8EKMeYFo0G857o64SYhgrFlQGOwI46b+8p0EKJXWftY
UzWIptG5ixypNOQuP/Cq+QtABrn4iV7GuqXS1B/DVTBnZNC01vdxLDCzpwz3No8K6fLxXL9OcN4p
RCut/25UV+g+r/mDMBtqB8VGOA+ZljTxNnfD9eBHZbdeSZHENPXo/cc2jiEhCftoZof36V9/pIRN
P8VFhP2n7uykZUvZ1sHY8Tf7F1tTk6oXMnwpFgejA8iBxVQKsl6R4JcxR37Br2nyDNgH0NC0iRtj
uvgheCZQYfv1yNsZN4fFn1Zr5SWxNZDX+WomQ9yjEAzIgLo+uHe+FyzbXzKOztapE/OBwfW2QAvp
R2d5I7372tfuFEKoXKMHSwwwsGVJyCQdj3X4vQPLw4hCOoWavsOm5N24ZN7SBtwClCdN5G046YZw
OrxQkERmn5gPPnYhL6yqP6+hMEMpSLaHEBIRpoPL4f2QfPmhiD94c2NjTHNmkdWq/IRMPyzsi9QJ
qg8BmT/PtC1CA9pDPnxUnuF+lUWWto6//oU7EERRsmsLAPi0KXbTDBgbx8ng4s93kcN8+nthbmbr
Lz8RW3t5pzyKaw3NaO3f2rrKuArN5Oj482NcNKqAL18+DeBtfd97QTM9xGmSImqu2+XyW/mXdZy7
wwmOV3VC1UL3tL7G/QreTjF3TzwzycNdAJnHHOIzA3nfSuKqhLTYriZk1iSVri+t/x5WQy2bRzmt
EVgnHMS0WP7iLAw/bF+ONc99cRO0PwkewfZXInZRI+5PCxQQg8D0uQz49f+I8ECxS0309BlpUoNY
V+Up/Co6yPKw6pYBOSTBEtH16DAnaR9V99Sdc1/ZNKj9Qkv8bTgNNdXM4i1DDNOgpYZrevsPWQo+
mItz7zV2gr88kWFviPuHIAoEBOV7ialedgmeJdinVhtnPztLEAtsoHPmIGlQ4vAS2te5IWCU/yEN
m7N9X3ZD3sndN2H0dgNWTVF57CehtFBb/+mXCI9u5h784ExYX2wwPtvi7vfi7auoLEQivp+ttOPS
e0MtVEyG21wrutDBr78kgLUgdbFDWdkTxT1qP6tlVXKgflBw7ASMXYnSEQDMW1izUjk5RNjQTrpq
LcU4Q34V6Gfy20YnkeRlbR8R+IG54kRe86LsOUrBbacHLbdWaaBqVoB08MVLlzkvoQZQOfZ2iWev
nna69suLDyHgMxL7o6t1NuGfCnTnpMXmsAGCpobUBgTPrcQ2GVJsO87KQ0k+cevPpeKPRCMkauJS
Rb9IMhVfXBxnSOEBUbQplCHsdbJ9zkhQNC1QOY5GlAc4wKPqmZEVC2lVTKhakO+ZsmmynjDp2zMI
eTsKNVS/9YdIPo+VuyX60055sVbGwNxHvwlV/JR7pdCBkpO2jEJRhwdSCigZtCEZAnGr9iae4jMH
Ow/Fm+TwD4ncvTiy2r2/Jz08Kut72UuJ5l0bQEb2puPfvbxceGvNwkltxrE+rl9GPSF2ErFstloe
h3ZXq4klSjZ7dN903Y4oAX0uslvI6db2idR6NmRyXjsKfqKr42Ilryb/LEGrcwT2o2n8/rlgcwr7
cYsggFbMvjxTdHfFZf3vIRk+eHybzk5HRXRmbuEBQWkq53/pvKARCRJ27h3I2cMh+m0UWXh0/Vo0
wVVs/5jCSZBXyS6gNlxE5Eo/ASx+abIBR7VjBQs7xhlyeU2W/KVCrj+tral3XnuKDUl1sbfVEyZ0
GcBrJ5Ko6Ha+j883sZdarPRHfLS9Vu3A8eb88KTYQNOcaWYFg3of/f198MueIsY9sCgFSsVc3hVD
V4nzr/sQcoDcPUNP2b5vF8fDvOrH15ABeTAUIejpFsRzeE6QVfpg/E/rKWR+zEZFf3IJVq6iOZ8y
KRabOcQ4dU0GyZxCvXqijtS3wSNHhnhN9zq+sSMTfPPqh/2xPQ74gJEGKxyGrUDcJZXkmYiYAfIw
JJRXF3O6nsfBxypG+gyYXgG72SJscsGT58DKd0zbzahnGfJNQkCy92ooR7ml1KsnccdrSrRC8v4A
uHcBjX2/h9rllp6OtzdcNhR4FuFc9CuDxKumcRAuBGpVg266jC8c8/RApVCRI1Qj5KOotp0KNkcy
5/xjZGXoVXI+qg78CFy8WNd7lXcgcrbXucsxDov75IOH2e4V7K7ei5dvyG6euRQHR024QyrnAgDy
LJ6IUijmp057tkFBH+VxZCwWZqDd4zE6WseScuHZjtZyxFfwBloeKlmHU4wINEzl0AKrrHOjOhhN
Htdhg2c8n7h9XQ+pF4iW1Twbncc07xPtTVVlXMV7kFkYSBjIZD0P1iXc61JmHvsalzHx20Q+MTGL
91LtHukixKQjXbM314YjPArtOJ2WZc1TnzfmXkf15EdHggUkYin6EuibwidOQdV8UwLoY/Zyr//l
K/TDHO8lJCf0Zq1/vsdoiAbKsHzjB4OrpEKPTpwgUdioAM0UJIffku0CAIzogyExQraXuYmo/A7s
aWdHMOY5KRnKEOWok8uFyBM0NlWvouT0yL6w0YuDJCny7R42pbTziihdgk78LsNX9Q0ZrKvyJPVx
/tOythj/hiK/rZ97bfaAGVD9w1kYiAeVPGAU+Vm4hwUR7yQdXSmDGnFJ0GFjlp3d237uibeoRvpG
WLXDhvWmviLriWSrLw5EmFEz01/wmoXOldMADZT6V1Hob3xAJ9tHltytApcJse6ad4YBqqhSyEdS
24D+Io17GkIdyPw7s0SG11l12+wvloIlkttHl5XtnSvnqht5/InhEsBBtGNaycSiXVrXLwtN8Myw
m27Bun1w5udBMA2ziHKYGrUQhdhQjpTTHIQZqPAYzBZ3pdHp8cfKUJlH4VM8OcciJhogV007Ns0K
gfsTuDQatoGxfdshV142gc7Bx5Nd3mXsKF8NJ4mfFBoAuauzJ0qa83xT7EndlF+yNoizwCNw4RCT
K/mi3/7lkES6E3ZCp2i2eD4rUegiG9u5QNJDvxouaQ8LjyTOMznsddPmHDFtJTyCnCIYa8DPzF4T
1GzX0WTXRcQpuOTfmwAoGLR4Zpznv1ekUJHFDLE0k536VplJhHjpGKAx6tUFgH/eWf/cgR/bZClq
yegwiPO/wp2VQgbydMZCrbBvTpPCiRl82p5G7JElLaScM7HnCYKgz8MqXeaGL28YRLy9HyL9ihQe
giHLq1q7MgJa8yyDSZcqX4O1WNKUasiJso0GZ8GrwDDYKk8cv1dCkCRNqEdcgL+p0+95IarJA6BC
iwnac5YpD4t74b65+BVjDwknl7J9x0grD4TAZdY7hEmlbx4tSKUoPOGl4vXSNeROvYXUTbc5yfxj
pGnGPgzYYUEWxMtlsyzk3O5FYT1OeXwbZTUa39vRysvRiNtI04wtg9I858hiU8IAmnmGFFqT+ffM
VO+jEVFHo3ZWV7KpZqIt3ECn+5RaBvNTlIli2tjCp7ZQWLCqqmSEuIoqNDxSMrYsu2qjXiZACrZs
Gt++nz5JucfcQ4yJeZkl/3VtySm4hTDYM9wLTfkQKyE8S+w3jqhVp/eUcxyniUA9m5axhFp9QexM
TVC4p/yDE9W311kmxqHNUATIr8Bee7kvLPvrS6JQJyyqquUbw+6uk6H2t6ga7TfjyaA/8pwY/XyK
DH+T+puPWWhTKCAUrpys1DLTCX3jdPJIpcmX8+XbYiLJobBIBgqEXTiDm8zt3yz8Z8mpmuvtr5Np
PgkeMnT2Pvg2cM4GhIU9H6/5EK1YitmTz9gZZY5U/ShFdIrKC1t6eKD/b1VNIsuWMDkycbCvOu/F
NcIZDhc0yEP6grFtI7o9Cf38kJgne01P0Bjl9ynZRZz8R2RTo6vTCrHt95Tc4FwbxqtGkMvf4KLQ
ZUpr8KjMi1LjxayW4+AN3kwOEQPaox5CalhgZ3ktwzb3L+sk1DT0lniXLZ3O25dtq4xILEMKoHAq
muwQ4DqT9e+Zd4OYY2NwpKsTZMASiQwYksjUOwGyZrtClR4N84fFa52lGIn/083BgmAqfbb2i1ig
lWmbdJI0+qp/Dus2nQgeUPkg8SxE6K29NeaVlJuGgfWOynn5TT1L/O4Wq8PZsGOMcvWFR+nah0lS
/wFrcYsIL8gU8yxjRmDtKBPMOxg3UAIYkemIrB6Hy/S09yQyiqoI8FM7ekHTMtWUwPWwyjei2pmi
UnawrNxh59epcfTUDhWLW5y1DMCMyGpzcL2RZA+Kr+8IrbP0bsYxn6OVQIHrpH3MTxsrprQrLfNk
hiLMtbl4QA0UhjJX/OSlUVmXOBHQ/felDrLWJpn490XgOMNPwSRVb6247Qd/ntV6dS2Ab5g/V/gZ
Q++2qzSXrSa8/PzXfDsy8S1E+Ru+Nv6Vgtiz8UwC3qsoVLjrbmrOgy4rqj603TqOJNIhOIj/6MuH
hIWQw4LWFtDfh5pSfyeKPpnXZz9ERFr+G7/2iA7nybXahbdKDguU3ZE8L6Te2+n0KnG4nLuJJQBZ
Ip4TjQQDCKXwQ3C1+d4Z6txOddWnHLQIvky4mJWe2GfxLJmCSh7eWpZD9c5WPFapPqpnby8G8ZXE
rcNSi1w8agimcSAn9WOxIRSRV+oXCODP6ZB+FiYo0tEYuAaFgu2QhPkrfeZ2PwLQShYc7Wu67gyA
xebgVTB8kpnrvWZhPQ18cHjHkfdzsEOQEjIsphSbqd7qJA0Qsl+A6iIqgNI16XTyhiDK3ly2bcQt
zFKvHxmhv0TUmvy7ZCINHuFvF25ObLBm/SbUX97Hl04bQvelt1AixaqpvYgfg8N62TQFCxYZXZvX
LkzR6E4cUPNBTJh34XGj39EYjUSOdRx6+wfWrHItrhQd8penxfIhAAd1WAT6aiadO73Hb6Kf9va1
D/WswWAO6G6tYEq17cwgycj4wzDyLYHaNj2xQqXU0jAvQ5+FAm3vj3NFxwDgU1JFsr6J2Dcooieg
l/hUWrLzP40RnK5Y8xdIaYtlFV+VEWmw2yWNTqACpmzQJpNBD+MsWFITXkc/eiW4rYJpJhnQpS1x
ES8JwjyYu3T57SjGa2zbma2xRIQ966NVms4wMIY03hk6qkgcnhXBbwlcWWwFPDTxcMVCSD+hNd4p
EgBjo2PQ3qux6WL29w4JdHjZUKfsjKnFnActB3w8VoIs+xiyo6Lqe+suA1WaM1T8PlQJ6FbcIvJS
tox7ZqL1IAVfdyPGz6JLK6oEEIK39yEfFvUO+hosqSg3yOhAINp5LpHx/lkrxpURMn/twwKdRhlr
SXltTZPLInEddQKs7m44KduEI4fEqIRYUeLhnSEoAFGreqOknIxmO9cxLdA3SUeiXpetWsrPgDX9
+YO6ToW1P9LuDEs8qdyhQej5C4tVnv6ydz90mpwr21DoHMqNJ8fN8YXg3tXN9orjmRJl0zmY7Tws
xjISBsQQZOenlNk3fxvWRa4DsWYwF2JQwxNVkiwsmiRHhWziZ+dFMy8FrYJODGxA/Yow8abJWTeE
oaX/mtNgWflMicdK95S6viA9ooT3DWjGkWoJrwxUJn2byu/P6Frw4R+ncyX9JGTtMw0JzeTN8Nk4
Oyw2KuATPy2sjOWw6a/dmD08P+VwrfmPFuhHUtLdx5kgUzqoAUq2Qozk0LEApPPCSL4+sQJKWymS
dI7Aq5y+kTcgraVi7wDzw5JCsYDY7Gb9kfEuYj0ntBzXlI8G6SqM1tJzbbULjeHayVb62I/Bv4t2
X03qiK/c3y0ub7bvQGttM0NZd5zR6zScvuv0oqwVLRZjktUBkK5pRTEzYvGTTu2ntgA+4YTMbrTs
GO6KqqhNQiEgMvJvckX3Uf9RzMdPj3arDJ5qYYyHqAMUocuUJqT9Bt/EQZcbv1E3gapCZqfj6+rW
Fgw8UXq43SOTWfaz2+GcAefkX7HH87kXp1yxNBeV8NX9sX5p/EvwYxb8j2NAZhYqHT6bw44S4hF2
N4+j9hKllnUGXLra3EUe83fHng/Uj5EFkgFYMN3IRS/+zp3Who97sG6oLDiu8ZUGzSzN8YZQJ54l
l/Wl2lZ0Z0/WYxkAx6caKQqzaxhmn5C/BKsNop+NdTKvdRAGC4XxidPCkrSKvDp/av4T23Ny9+VR
pKYyCQgh9lu5r2PTYvQTZGfMY468yo3fTK4Vqx+pOH6rZ3neM+l20+9SDWqOaryWOg3Ey9cRt8dY
5S0t6lBwvKTe2oXhLNNV6ILtOgmO3MLzukMNQVikdfY0zyG8Glib1gPQ7sI7RdDzshZWAmcbRd21
iv9hxDx5R/2lXS5qHrb7BzsbSBFx+R7utF3314+0/U0ocKmfM9KUg7/UFBFnSYeYsXvt5xg6riNP
WP1y9mhEUKTGtwFiJfSrcS4UqEpMpr14K41Yqnast0J+1ewfxEdQGEVthvhzkvwYm+RpZSXjM1hh
McMxNYeJ9TtpFNseIF+7D330c84cLC8JcjJJJwGs1aBLaSjgKYrcRDIt14iP4+61ffOib6gg1cTs
jt6uQiG78FtlJCZrd9ZSZ93YE1EShmfBviJ0CLEL/nVpW0s3trgLgA2oCumofli73OWAL0KlVJY/
In6Kw6OZvA9v6CmFNsucfXkITXJt2+JRk2NvwabDutFL3CQ93J3B9x5gVl6RpYrydTGOhaKg/qED
4GPzdbsYYxCN82/Ke68UcKMkdNO7136/EZn8+sKeAa1t4WSd9BArQbILmO2cF/t+KywN5vf7Wlq7
GyQcQJR8yTM2+cjeET7m7b2e2PYimU5zAGdWu4VbbaEfOLt6i7l/uFzG8VwiCoEcqy8HOFy9Aeq6
kitbpagk16R8WDrVoWbdK2PlkUpJgBzUFVQTlF07BrUTTEb67o+8aX4wG2C8+hHIXwnG7tdw8PeJ
TKArswUWUMmD7vaAL9DoX5w13LC/UpByvzWJ2hxwh4OCFpTZnHVvSNCOEhl/WWVc3nSB0q43Pcac
0nMUuPdPssSGM5SSzrJOAgc/bERjpQFSM1uf2+8CJUUwve20FU3Fijjcfr6ghPgKUEzBo9kWh3hk
u1QmUoqDMYxj84WA8uM212lAbSOvU2K2sl+u9p28CJutn79WpiqAoryQ94na+SsExYRyaGt5xElx
0G8UtgZdWR1llvQvQdf2PBShGyp0ILzgXmcXk756NI+XWlyIIC2SpHgyohpzY3ntl+qer31l+Rg7
jTgBIbxOC/tAc4ZBF67PDEm93/LuA325/Bh77+Gs7jF2u9zDVqwFCipJs/arQTdQtwHijjfgcrFg
QTlJDqEKM42V9dci6uEEaOlPO2A69Nf+gzF6lSsMx4zBvQtqSAUZh+TRC+WH4Q9cML0BtGw0hTBP
DlQpnkAVkW4H3or+kxpq7WkwwszDgYefOznTfAZIjYl7dDvxYYGxTtkMjPZkvRtS9YvQz9fwbADQ
03oqpMJGCEykHwl69kGCXnkbGUjfr8HN9a3elEZRsI4SIh1Z3pGZDMWtVQkSWT1JEG1L6YR/GUHX
4gu5U9DhLWs2lolkrTVKbtoHmOvVxbmBeWdS2K9BIBPtbBBz3wqbT1jmSoLM4J6+w+7c9/ueVElw
GHmZAWvrbS6zm10vqJMKko3C3YlCTWC5/USY0orKx9e/kwrXBdhjlXVm4Ed5S3d8AvlWLqcMkf8A
B58h8AdyTAE6bxQy02P4Hz4FhmCKUJC1MYjqDSW3heE00pIT5Rz4EqvX6bMVEbvwTxZWnB1XXw23
P4wMxFHBwRX2Z3xU4PlK4PiVftzdzTBoULITJ/OZEP0FcaWbk1ilIMH1KzYNexZn1AgDFC0kZaoe
evMUUpDzH2XsN/6EpZXNZrQNR2FIZkec6NxwcyZCDwcZ6PK8CWXEwy4czomeal8PXq3JhU+Fg/oz
swzalFi7B+lY1N4IeMs0F1+rATxPOHCRRPWS+ySoDOE5zgo6Zf9hjLHGq5aIxLQnbTabuorbLnob
asRdxqhyZPe0ZzqJWg2E07rxecodZN08ChKHzObNwNu0nzdKBkhimJoBm7tLnnEB4gsoD6ebrj0c
EjeNoagugXwvIkNCRImvQw6DedeUtiaIQb+wHp+Lp1Hqw6nN5h7B30TBFGn1RnQnYXCiDSjz6NC7
vxVN3655QJOWyVqAx2EG5G8QgqDxVzxpPIcsHh/v3Dkf7gE8vfmNgjCb6K7cfHrh69i5aOqGgpxb
B/GHFS1m435/yDO+fyGSVjdelNZ3riUzQjSrAQ03aWgMjAMXdTr7tRV0QM+sRZEruOOo5Jtjem26
SLpyZL1ccVUa+uM/8mHtDOiexromf9RPzRsYMW6blxanVA6W8S5EAQuy+twOwqP+647WkRT/Ge+7
1QczXzen0MBZbMb5+hYejWRb4EPWr5UYUJ999/W7PAxOtp4dhS02W+FLY/+HvXNAbhdekh0zoM3m
fqxScaeVqtDsfKOQzdLpl5dLhcqvEOZJ+ZYkXh+FLjxD+5sT5ht1PXxTU9WIG7hYZF0PfTMHkalD
PuSLIgJw5faDurSt6ILd6gJcz/IWhMW655ARkAOBZHTkxAJ188NnDHEjV4zsXEdwKnQ80tPPFaYw
XU/a50nBbB3qR78QHK8XLn7jJYGQuf1rLbELzOxI3PXqo94439h77+SOs/c3D3hYwe4JwxkjIP+4
NYtIuC1AU2BJIwjY+a6BJovne9uCZ/nrUIuj1ij4c/wJitCI+a4Lhl7uGXX6oShfuGZRCFueytkZ
6cLc15yHQOBkrC8RdNQg9uiFC2fLVfeHHcB0viD+MOXaAS7eaT3i71p0uGB80lQI5w3KmWVBIY4b
3Zd9tMSmaxw4/mC6AEZdgAqXD7AUkcPZpYLdXRuRUoMhHeqRrHR4pstErPokLt9/7XtawJ5IiN3K
Yewxdtt6qyb2+ab94x7casSIhkF9mr0qgX3QYO2qa3RQir4BUtew4FQLL8Vg8fr71AzSrUYTUPnT
0kky1N6x0rzKtXIEfXpcmM1oAZxt1F7OdYuXj/YfQbt/LI618mk9UlLj8WTZd8AZmsOjEf+hMd1T
PKwsGv09fq4NP1IqEVa5eNLz5DC0foeELkf4n3fELRL/ExNemoMYGj3UfMZbBGih5cK6LLFIepv5
yIzS39kT/qndCNX6VK3D/izKm3JOqRnsKq2jS/tLhgB3jdn3q+lA0m+S/WZJfmz4/qEm4iFE5JGu
V15yq3g0OgEWSgOf6devErugsZ3FjQ14l0DHmZGK8VRvFgbgAIfj9AN0MJEJP/7/XHx0L4Ay1yAe
8bFkCmNpnz5HCAz7/9Pz8/Y1uIMDN8i679ljuq/6TCnmxf7rc9tQwpgXtL3UtUMHf6Q7p8iBoZMG
yXmrh/RUVLe7FoIF1Y63XwYNj8qoWY72l3Vi+vDsdeE5D3qZDLnWEJOSViIt0Epqe0EyCpSlcvjr
wUHKGP4MSsW1gSv++WzvQiNc5Ev88y9COUJcCs/ieItH28P72IxhZSDsRmLEKC71+prjNlUMyPZ2
q5u3aV97kmPwEBQZc7KDwGlKZpVrZjZ4DS8B5zkuSNZMVkxpfpJ2RmyF3t6jnHOqStdeX/MPaplB
MpI2n4O5rFQCf9cQf4IDkUiF9YrQQBwHl33domuQUMD03eUoEDlO5kdVZ65sSmlIMla4RMxhMN/G
3Z+yXGuz6qnBhZ/IJApjF2xCcenyvCrmo15IswMN4MPXbQJvRdwdMw/3gMTQIcnB+Ws3NG/cKJHq
HHcDA5W1H3VkBazsunqAQdY/Io0wcJA9fRqprDRiupYH8G8QSBxbzi5nmoJsLUhlUtIuhHIkAGDR
ZAkX74iPBSNBpl0WJ+84gQWUYX/k90fHFPCgNbJdjrhpkjee19ynLUtRVkCg3V/vJKhgzRyoPxiw
Lnj/ajVBaXi0c4WIhfyeoHiiry+kPpOntz4HbPbi+nCrjnvaRiPJp8D8ULErywXfNVN9cOhgWQDu
mPoUdeIPfii5cvSkVDmZOhG/2LTob62VrGMXoE7ODGc+4/rqydJuq9yornT2e1fDA1CmZvj2i0XH
UjWsxB8E/keHa3L21HOykwLXjosANxgkMXmL7xy+SdNJoS7Cx9pQuxWS5ksVyil40NbcK8XmVFWH
Tdd3um7zOigHZbeISjNEzH/alq7bYGmeF23FrqWQglJdUUupYVp32eviuHhas2Uh3oxoVbnh62rD
+itSCwP6PBOQ2/SMRChzqB2SEpcm0y2uuPHd2CdrjOI4BiU3SE8nvhb1ya8hb77OXb9Dq8R2OqAD
StF0Na0ho+EMzurPjP2qWp9VV3FWeBa1h7N056H4lgwe4pPzF2c7k6XIOrvDPhYdc/LwixBiDv8N
Dgrj3tVo5ec9gcwOKsN66SLKQqlncviWkLFqs4Rib6oN16/j2eqYzdEssSoKV5Lf787d0DyOEhxv
384bqrTbWXE7i18v6s4HGqswhe5uys6H9PiLEVyswCFWJY1PcA7dxWlNp9ExogBzK7kFeN7PuTcO
dpWRV3VOKTZOaEfREtiyQG/Nneou7iAW44RFfCzyUlGKXSW9gSoEwjGD/Uf5H/kfEqAXZF+CMqyo
QZFA+HDWVtTeJJLSxrDGkg3B5jRJLVATugHRzX0pMu2gMyjkFH90LLq4X1pzDHJ6/ow1KDr/VXGN
2fd3pfWb+0FDT4u3mHncdY4OavSuS4KJgl8AB/dSJtvcCvVPQqbzaRXnDNxAOicJRUPbJSVZ8Tdb
jCSsUxXCsc0NvbrF880Nd0kFja0wQSrQMrs9uUyc4kG97IIByF3muWnmdV6gTL9NGpAKeNJOHv4s
KRXinlGTk8hP83rXXe0qdrtk6AaL+OvxT7AHIY0mgQUMkPegqzbOStNWxCr5HGCbK/8u1MiQ94ve
SnAS1Evw0NuM79lWfTiTyB2ax6ifdJmIh5605dL5vTronKaYYmyqfZ6E6RcqgWB88/EI0lSW8iwN
wLJencY9ctL5d3ayAMxACUd72VyndlVW6O9NB+/eRmLMUYdw06zhV91LhjuTafsFjmXMz3N/z99y
qDbtUW9l6i/Jq0Rlfuoj5kfeGcBJdWm/ZCnTMPEQU1gtoKp3zaAw8rTUysFKooy+StwXB8icCexa
M8REo4p/lM6rfELwMSQloYOpid4jgOvhHAg7kvoXUsaKKLQMyQ5IFOiQGjwqKHJJmI1p35nBzy2F
hskSkPbxEBz4KjH29CBUBv2FEUH7quIfS3WRYZKwhUWrgE+qUnOd2i9jPW7lbXEEFPqMj26cfkWS
CLq8acKgemCHWK2cS6bP7c+a5/oaacA+lYdZqhpRuLnP5AJR8Mo+9BBM+JUMJkSRmx3X7Ke43IoP
0pAOFoRNq5RBfh5sLH3NEagTV3TyJMaZ8UWUSJPvXyYCG6l+ae8gRqB0DF56uNGFwcfyVYIOqf/4
B4gNpYbBUeZBM2SuoyZnC61aY0BBSYooUA4UXuWCJRyqzqort1hjchGdc0xjAntTHTylXqRdZYsh
5B43gL6pMr/TAPwWX7eCIjXYPerv87X0LtAEaIcsGWnV0duRIZOq4aqAXD31IYEb5Aj6mwbCpGzO
I3uo3YfiO+AQpLtOHmYGVTVCjRjEAOnN4NJ3q59TuYkSYgbd2vd9Xo835JyuriTVTMppz9mByUVO
e39oFryjnyPXfZUvsQfDpXJt7CtJVoNkW5D6lRI3+PMDekpLN+TehK1FSO7E1417OjOICuWSQE20
MeSSzro9dxGuXhfUn/m4ZOhvqCBlR4BfhDXVTqXqJdyBP7meNI5A4bj8KGsxQoIFAP8XvlIx0d9b
8S8fcJ1KQ+XR1Ab07/9uoYU2r6hyHy+jH/X+euOyU1UYJ75uHZPwrEhrsblnaeEseIF2e4XPzWYK
t8MBd6Yajz9QcbHosd7D9MZijee3Saj4/wx7ypg8pRl7JvZN6FeXgvtjTbvDsdUIkzCUuhGHTzAn
rTZuLfnZ5uZiorzWPLroi+UtzWKPNdz2a3b+iE/X2D/79nfD/U4ZdY17svFjhHJmiGGQ9sfdlPlA
jmrmmUESGWquZrV/njLDItZuGUVo1VZxfQtoDGy7K02Z89U+QIIkzx4fnXsHXJlUSui/vat4JDT2
zR08wXpfxEz8zOkoHhv9kZVB5EV3LvO2HLV0PiHWx6V36SQJERKRDeTskO2rzj7+hSzgHTWsi9pL
R/wV/uS2qzc/MNj9vxsqqNxC4YkcvuD08rXh6sTQgl4a0xAem9jmHLv9AW+h03Zx9GQI9uH9HjaL
RvinamWpQiGYh3LbSHnALZ7jiZIwUxz0AjTTLw7tMVp+ZlgZ0aVHyENwQc460ENTlkKMCB4ZqHy2
9abYvG1eSEQTVzKIFRIkE42mHXLeHGvztaAbR3HILu0qxiiXAXCstZdHqoASGtxZ01288r3fTKdZ
NDIARURMOEXCbyDhmcnBNd6hrqDeAVl75+ZMXSgs3Rd1KsQU2yzddw+SfvzHPA4U+fFNZcsuhjpl
th8atDB5nziBq1EgnRJW2OtTT390pncnuPyPAYQm42f0DS8Mt3nE/nj2nWkFxwRYBcS8Tn8fwvBj
SewPpzUCmytUySSVvCVwzCDLUb3pRHnxDsnqYaq6ESnkXghmLBQ70UsPvOemiWiCcUh40tz2szQr
HZxQWNpHT5p84OW/SOZz7BDD5sGZwQKjW+gihHBpCpHpNmhGIrfFlJPEqisPVzHErWYjrqz0LTun
MO72UqX/rhodPYomrGagfhBMzPEr3aZKEZPk9xbNweDJD8fP36hM97UClaj2AuD0yUz8d/z7gBT4
O1/uyg/cwViCTm8ao2irmFWpqli18zOKz3Lp3RxnEAZOI8fZyBYf2OFlA5RyQlZei7h3HO2+CONU
Sc3gV7vjt0csUIU/qUU4E3J7RqhS9SYvjk96eoW+Gooulei2mcOxvZ7VJdbECNdQpLKjfTUuovT5
GkYUC9AzTxmBu2fcPpzyl3e2P8VMhpKhl0ivUiRMgq+Iza7Nqtbsuiy5a+Df/LecoOeO7FyjzHfu
p3Cc1pXvfLPoRZnJj/xJp1SuKI3UoIT5c7A6AadmuJVRp6PjNpB8aXlTsVMrQbgRLjtLx5new7To
Xz85Pk5sn23tHMHMiiyDqbuo70PNqHKdZyi8DRrwzSfaBJ2dWc4UYjH2CvGfy0qfvVYyngEzMOUq
kxGRT7oYWR3vZOSN9GyYk+UWvfftC9QacpMJCFzdWTHPWNYgUiOYOPwRfv8PdAxToVDn4NV8FV0Q
Lj91632GmqQn/c20HUq4kx7NKpoZIXSqPY7CxJYgyiP9gFTWD+Bjwu3saXG+49EF84+ghL7FDKTH
B/yCaoq0gT4C3rawjgJ1D5NPGxgCm9DaDZVFX/vVxIxNCTGEQA+57LHD8JgFZ4ip/cGCvp1hpe1/
6FtkCBgwRhw7xUZT9vWKzi5ok8XG90hUdYhUEN58fTep/cjXG4K0hYvz/GMMpwbWevjomEB51JTq
x63ahUyEkiVxQC4oFJxDtOILVjvb8RQ4Mlu8pZ+wVCEQqegKowm3rWu+LPgtv66b3HfVdgn51bTS
9TJrllG8VK5XGYVtz6zT0PNGYf+z3i0uZdB2yNMCrFZEXIQBN4krVF/FF3n7AXuiTDvj5ZrjwMgG
L/tPyIT878fyfOHmy3GX4QCyc5phUe5vL43o2EBdYrtEBNxjzL9OPeqt/+YTxxV3l5T85hTamtN1
PxxTLszKuhv4KXOq/OcO0nbVvNzV9IS242+JKkKFLCmQMnXXUSI3SpV/hlBSQ0HuLcqpZzbH/gPN
WXOGm5u7k32T8f4MX3HuIuSZMQHGL6Yihn3brF7RinGxd0OI7cbehQf+kmJhwavTUgujXcJRoHQ4
fP9Htbn2kj23XxGAtbHmJbwO0vfFmHXiYzl2W33aNTwN2BLgtsykReAq5dZCHuezDLuH6Ot6tZrk
AiE08YU3mTVS3gpKKlBmMs4SBNFD+NFCvTUmzeAkCMqdGV1UAYZm+jXHfyjsvf41ReAIxb3JZ/kB
2R85AbeVQorQg6aw4YEO8SWiYjnLAurhHfFhJbtHkRCUGPn6BR/KSA+mqhFf59jHe4E3g941vjir
oFaiW+v9zVYCXdxvIr76BAuIooYuLrC9EK102WoJ00XB8t4ZfG0bbS/Yy9Ts4yhwNq/P2QeFUGYE
DF6lD9nD9tn91WGdQCnGyegdvOBA0pJATcOignLyxeaXyATVQM2+SmB0ECrPY7jUHcwOkW7YFdKL
0J5IWeMHG77cW9oC9rdf1flysrFEE7WmuxaIuP2phb3w6paWULrmOzA8KVOm2g1nFxNgo40gEjfB
7Kos99j7zMvi+G5FahQgVwo6BZPfxJiFgg+mZYC6gjhMDZJiJRIsQdQnM7zXg0+fvPDuSQ1xyjXU
eoA1Hd7KsfaeWOCiGyfsOL3ZxFElxywRWL+K/96giuJ4lkCRbb6QTPR0geFMa3oDSNwl59hLchmR
GFXyYA6ybnhdpvNouankLlqirQZn56fY82hPZYarHsAB2njruD5X/4SBaX2//8EJ5bRMKpgAO3dH
Cj5xg6SGR7dSLkrrcntlTVJ9vuq+Ze+ybFEbnVWjNutsypZWe8SEG5LodYc3Nqp2rw0xDN6S7DIf
EvmJt0FLlruZBfrG9wBLwF1XHfmmymqP3rat3pM19RpvFukpUCR4MdMFrl+rEqAmLKNfqx2hpDwT
YjysFBSgW78q7UIHyDDYhIez/P4PQ8ytmOVbM785+dW+xMAlCVyQRXyG5kVLjehe59cLreLGdLzU
9ExPtYe+sxHXl5WYrLDsMbbeBD2y7ejX3WHN0LD1x0XdVT9x4/3GE6wO8GSJnE3AoBsmdkWrmd0c
OKC9bt/yWeiHB0vv6QtHBvE1vd6lisla4+uOg2OElsDeeVc+JaULM9GbWZY4M9BunUhgYiDPoRxe
VE4XbT/ISmXIx3sZrEzGcnMwQ9ukpk3hVApVXYPOTxN3hv56cKyb9h7/NiWUtWBYN4niYlNjGJkK
qnBU29NstZD8FbMp5gCJ8W7fv5w3nBWyOhi6uLLTfjslppBXVJls8Iir1Bt9l9DXTL9PSyjjYXVT
McdPUEiIhvcYwAvmf10X0ppWeAvQW93GgCWT6EsFF3jjOmu9a1TLh6j0zieZY/4lD4UBouvkH2DG
GV8QkiKS6TXPNlK5q1EvtddCenKRwT3nkwDLunrYutGia/NIfFWHcAFJIZlOrI2782lK2nuFhoyl
hFBkbiIihj5QeNLRnA/sd1lHyRozHJ/R+WedUspuwlS5h5R8HFdbyhkCs98PUoApo2Vu3mje4q31
p0NISiz0YKoZVKRRG7zVG/pDo8XzQgz6hiMc+OCPlVODR3eudhA+8wOeVAvNu7OM7uIn++8VfJhF
sWaXQAK/knm0BBeeQIEYElwd2JZOv5tDw8OY77NMd+8vjHOgzx6jYid+la0drckZVStkc28vnj3h
kN9r7RqIehqJIIXDs3olRgJURqHCOgJkcAtMCkjG5p7e/libnuAo2nKfziV4wf9DJpQj+Agjv+X/
+S82RK1WPNFXJQlp/Ix2NUinL0zvLK2QqZq7t+k6ovWPzvzW1GC97NJWdVTx8XMQ78NuwlSEetV2
6UNQiGHmblTg+QnQrjyGrImI1DnHUWX2LpZOGIifVGdPrCpKHrr3pz1C8uH76aBylOh/AWSWBZwX
R3LNG2NlA2XDs1f6VXcYqJuW7wstaP+5ApPCSz+aWTpWmgXCCAAnHz3yCGA0BqMJfH93bndF+oQa
h9z/QayHENuJ4z8o1R8t3BaE6Ymj8wZikBdni8MOFpfIYhM/YFUUy/nTRnarVNmpyTe9rzmKoUiw
KP2OwRitKFcJ+a4qKyAE85CAR/p0ibhzW5PUv0AkOd2eOQ7hWu3VimRs2SOns79CYuGVwtiTrpeI
pch7Mqi2i+eMVTaMI2owNSt3lWI9IkDzbbF7ONtVf2KAFBDVMoaaz83dxG5zB0TL2espCLbd8BDb
uPM/LuzOJhI44CCuyuXeP715sVo/D0mBPDw7fByRpVL7PYeE9E5qazLtJ77vlf+u/+oY3v9dlHBI
Bo6Td4U59mCT55SMiQOR5indwzOARID7TGyjb5YDHZNQ7u+NqKMBRfKv1xnZe5RUJT6jL/hb6dUk
Fv1kBn7Wj7se5eyQfomtCN97cpbKqZeI6V4IF64asHMVCdToEo5tbpvgG6yD37oGSwBE5z4phMcA
tY40vtc/eT4/4swOuZYruLRVJIBAXJ2Cagv2FNThaVLzA2RLlDS3fK0fdQRo+cfDVo+Q1hfYSmg4
zde+29X9FX5t1tbDEYFUk78MbcxAJidlKHW6eWg0bBST2ha4Lsohg0xBtf3Zj7OJzHp0Y7Sa7eda
+RVYIOpWrv/qk576VOnTfoZmvhFyyUCCCStKVcTwf+moDvmkHK4fx1tn6hz+yXgPlhaUso2FzEkK
yoaSjMUxt82sHl+oAsblx0XyPskQi7ZF44xlR+fXYeMhHWa5SIGJNbYhgO989sH5BjsKvKhWrlVM
i0lmI03Csra5i6qrh6Aju2qKxp1Qux/Jz2hGZTw7HSajybXE9R1QT756ulb1hWdze/LvDF8q1COn
rw9JTPLrXwP1rk2Ot22VVk/Om3o+Y586SGnaIUMWWbDFu4aE6oQSAiG8wzTddJ/UCb5mBDWWyelW
+SbZh3+iR4OIX5CbIUv/Stjd3thU2wwPAg4UvYmtVLc7ywRRUHi9n3F92JxuO2qdHu8SbBvlaG5C
8xC2e+4ZcZqZZiMOxcuAe4l+4+69b1Kow1OdpSVAQoNpozsOC4LtkwJRF5x3H8xML2UNB6pLbYTw
sP/nRUWUU1LFzgEUJy26qRbHMb+S79U3+TdwULOFDyLvLFDAgbGWNRMLTukX/DeWVZBewhxYLNyg
TPxZl2v52zkExPiOZ1dQGSXhX4v15vYL9idzzp90dKBuUuBxzHWb2SMoRFrJpOc2H+LClb1b40Do
ctqKfu2DYasz4wy/yatPI1GKErkxYx/0noc+YNEDPsltBBsx7KHQBzuI7TaNjPBLrgtRxbdBxUwG
oO6p1RVTkxmO9KnAiGFu1xI33GerSJoer1tad6diWr/85YZ90/mwdNEn9l+ajCPhZQCP/KxCtpjf
GGusMjX+0KUme8eoLzHe4nDEUVQnL27jst4e1Am1+M17TlkroEpi+7wZPgkEdkR3fZK0UAYjcLVB
wOXK/cp9RpwEvLt4tS0QdPor3jH7QnxaSqNPq8XvyLKtN7tjkd2y4FxPuCXqIyq1AGi79iRQAt89
sfprcf/8vQYmgfWT9BB64D00064+47xOCewS7Y4HarDwALpUm9TmVtpI6qMEav1sQYF7ayzsKqN7
713iMO53fnEBsyXROGSfS1rz9nLGGfXPIfu03+HQUgVP0+KTWrTuIqxSXzHbH/25IE1c5Sot5+hu
49u/pq7/UjnllcalyMiu+zfIo7S5KuAuZvpK1rW/TuuYkSbVOl557wvDd4kFb1fLAinjUyE3i8g3
UD2E1pqT0IoviWgPzWUKTNTOHGBmNAYJ9o+qssEt55kR1Dbgj4hyJF8XySmQAHtNAbCmg2a9vhOT
7F+ovNSMRBf8fTMC6Hf9viaDWvS3OAQGlRLVaB1VdDqMyPu9yGaP3vQoD+4c2s9JrzdBY7CkRT9B
B4p2mZNxrqPk4HaN1sGQhLk2ety8fxsczlM0QpjzztnXgEcOGeqNKeNQVF7ksurdqc52eQvyklIt
IQPwn37za5qwg7WFSm+ri+8On3WeJbx7p5fuaZQypdKUGi8t5NhSFLTKZM0JogirQzGEJXDPb/Sq
9AeN4ucY0S05x03cGrAUGp+ypAGSYgZXHeQkJm/aCnYFxQAPra6LD/mygPEHD6ec2r4sRNhTB8SL
RMIdbyPTWbI9fwduFwPWzZ9G223nLWDYqtkn1Biksuvxka2GMOyAQCDwYZWYHNk+59M0zO6BSkP+
f5VxEjqKklWYnZrl1mLysVwENnAU9B461RyPO1hNpuT/tEcCbe/1TBRoKMLF28LoosJmuYH9v6pC
twd1877cPx8mbQS5R25tj7Qs99ak+82Cn1sezU4c+esmu121LJI5x9luPM2GgOltS9JTAoVYjCj7
FKM1NaCXENip0wMt15n1CS1SGqXQ3URvyt5neJ8QDcuB2UOWKu3bo66pjWbffC0sqTirhuqkpg64
HiMjeCOPZoCUOYoG2nPASIc6F6cOD80pGoD0O9PUrvb+Nus5sHdbpPYxIfoO/A4fJCIuNTQ3Yp4v
f/8gknrHPq7cmtdQ8uFdggOJv51OXT8w3HrmvZPc8N7UGw459SV6xjibyhgNM9qjB443+nkGA595
Y3xlQZnWnFveYnEfgpm1AWfg4NAxPdZkDwJtSms7QtRjTxop+NVAgB6VYq7Nf1yxumjH8wFAn0Ms
uWGT45Jk881n7mYEQRd3naOnxG22msS1zSZLFwkIInwOgciqTNbYAAI2jcW/Vyn7aFSbZ2DqLzJH
IhcSvphdt97v/berO4yizibCwCLFMSESRh57pOUA2DS/jOYxIcleuX5DDO1qh/+m4CuULMBaW3Fd
o2EpeX8AUGfCfUQOTOEQc+SXTij4vkJ2dOY+YFGWnvZGO87a/5qoIzW7jfJlep9591fD5Jfovyu9
1fV/NqLnPSWLBJZI23dR5QdRRkrQAd3GHlxx7048ZGsDxGzIAqleCRpDO3u56j8xEvczR5CjLA5h
uBshT2hlAM/UdNxM/Sycb/x3gePw+Ha2VGGeHeFx+PRbBnYO3OzOE+CyHEtkmf7NrxNtPTpZ4shn
aucJakessYzwS/bl7Pmorl6w0WtWInXabJCtSyOpl4o7txg4x7rF4A9OvHLoEj1PfOnlWiBCQRnI
A06paxxrsEiH4vpJmGfeA4YffZlOeke/MSkUmTed5n5Bq9aBgY0XZvpOa+T34v11nRuVeix/bIYH
u+iF2xbxdMQTbYVGvsJ0d7n1BcczF82JhCSFPMzwowCR5rPRXaQKYpHplISttT/dfw60V34RCWmI
DtTN/6ExRxrYe+DKegph+hh5/So51GQ3+BhdNMMxhR5OldDCQVztkIT9k+U6Wl1MYa9I/g/w8WHX
VsQxLlksHyaTD8fBrgqsW8EkESCm3n95id9Z5BUFLR2av0l+nQlsfL90LiH+HPAnEgJIx6aa1il8
SrsuegxeitODmfuKo1tcWXTcy8+fHGgcEPOZVTgr+puuugYVc+p/EU8P9iIyqPkgnYn36knse8YI
WE3GU8J5mYoCYraiyabQiYENkj8tudyJClhsomC/A/YPcf+ydPtehWsXpekFEsiIVuAeplgdm2GF
su2mTerWOO5C6fQajJgL8TKtPPBGrl39CmBYuLvH7EXM8JREMmbbL6O6a0H7zsxSaImuoOMDbujg
ZsHPyEGRmucYDoFBYs5vowJcZ8OVUy9fg/XkAbyHDxankPX6wSdX3J8tJy9p3rjK4SEYRpMjoGsa
tYvEdlRX0QZybsIRsjkaxcyInLYeDJTDG3s/4T0dDAwSOqf07mQ74MYcneOJJYum8pimS1c54jWu
kGdKCS3wN44nprNlpe4OXMidoEpZM5bgDg5kc4XsR4wQisP5ntakafhAIAX3lgADuHTzwMKfkfs9
H5G70NtGh0LwmcWI4J7tsCkIqAWiVoCpQgmUnrO3NHYG5K8NVAofzXLhNCxCpRDwu5YefAyEiygu
OLMhB/Mem+L3OsnZsEppnL9rdyzrcOmC17r1KH1kjkxs2Ho1C3LtgB6e2Unb4sG4fZiQory6j8gb
+v+NxWcWOlKaJ6oyTrEmW6cg25IJSZWE72OfJeYhDiAErgQkYs0FSCqJ2v8KOirZMCvpX93Bg4sa
N0jJmXIeNJAGJx3TmK7i52OyoX3NEvGf7+bT+ihE/wWb6378mx8KMAw8w80e28gFS20rq/zEi12S
WXNzHvaRrPppWIgS6yr3xsMgA3V1QAqykdxyR2xFlQVoK9hJ7kZbQ0/HCrJcvS+dunvTfshj5EFY
MMx6Stk+c7TZOpGiZ50V6LDLQZo+8AUUrrS97FOrKaxnm/Vrq6jjxI3QuGx3YP9/OWGAxHpAPuci
OY8COEBN6K4ZIV+s7npfuJveWzi4Uap22TU5qv80UiybMXdtTbcVsJ3e6Yj2ArUuFkCney5o5sTg
Pnlj25l5w7m1xJnEEsWJpWk6t9fMPom55NWh7yADLBHdnw4/8xFXlCet7zoyt4K1F/wJoqg3nPD/
7cQB4XVRjOuIW37OMDzBaOj3lyl945td2efmhOxbWHF/9d/iW3/sOWGNuw+8mNDgdg436xyarZQw
/Ilaxfeb0vEyupi/vOcexqNO5o6x91l6QO4W0DSaCHATKs4Bx3Ltg0KQppZa4JtXTGaJbOPwuNVN
HzSaDxVtMvhpN49LvY/2bgHhs85OK76P835BB27JubXpdq9CtRQANHmnvO0yb0naxtg9NEvO5+bd
lMbtchZBDnpD4/RUfDmlS8OtU6IPOqrI21VzppbdZ5y1Z5xXu+96fD0aTKBEfAz22vcOSRAc8jcK
QnIm4GNpeCjtpkRav0APhozMdnWvMqQUkxFecSG3a7GhyyTUaPLyBZMo9Hb6rf2sP2pKaZn/ECH0
/9n5MW1EWbdHe9UHlFTZmhA1CD4Z5PAb29d9muJc9cPGoiUcXiqz9S+cwF61qiW68Bo1NbtTDZhA
xUpIQPT9Z3ZPj4sFO/VhnHOxYNbObrJi8jT+dVzV2DB6VkGIK9h+bTJ+T0H2j7t7zTjgk+Jz9O0M
66Z+y9ybWopDAaVNAbq1oJ1zGbAtQgRHA6wXZDPhl73Z8M3brJ7ftYBrt7HrGKr55EYQjoqUVqjh
0eQ7JeGEJIAmxrp1yLUecoaY5o/zoz6YnThxdJe60xEkY+oa/A2FG7RXpmYrFj7mwUnx2oOJ4K6M
Kjt6AnQSRNdrlSOl89HFvwxbxt7IiCyX4+zjrQbvw7dK7R/6B2Asp/fT8QMKYGZ+6Q2i1Xj2PvvI
LkUCn1QRfgZ5ZbQ40Bec6lBIGvYT/lJqjkCXYVF6avKI1saZU8VX04MUp6qvUoUKCeDwq/dBHZuX
aRyclikPvjdhrb5pH/bFbHafJeSJ0A+5n5W+QWS8g0TQVSmT3GPcD2MyL+anKPWR85UNH1tr1/9+
WH2+U6ONGKW4HZiWnSNxdj+/QK22GyexkyipVeYOqFA4EggRqAPj65ljEM53aKEsUEa7WUaOHCub
D3/9CLKyKZVGlkD9sU/eVOPSkNeeHB5pEbywni7f10dZX/7ayJp+V3Df8EJxgX7XOkTJA6Uf3kLy
6+bPygiugxpS/xAMW4lYjsjm3PFYbkOZB0YkkGB1xBxZNnfzRtGh/5iZvVb+GPrB2ZqxM+pPlSuM
vW5jqZHArwMughn8V/n8K50Rnkh8KHA0K2FcA5WBA7/LE5yUepmdLRRtiWwvS7riSNU+xrXoKBZj
0iy9V7iuA06q9y9ukl29QH+7Lkt8rbswgtJ83uEie1iYTlpI+FQyShmyDEvZjDLS3Tk03eJirj19
PI8h09J3oGto4JfTCXzXiTiH9PU8bKJOFZkTR4HGd1UU3X5dIQHPq9gjUn9mUSfPtmSE3+kEDmFT
VPlAD9ge84h/AsG3pyfmfXDpXsc6YTtPf5K6HhzIv5yXfhBNAnwiYoQwAxshQ41VbMEB0UkdRqzf
gn6f0b9ZBaPT/Yu8Tjf99CfwlBajZvWLfM3+Wq8u7tdrh7+KZSWJ+sSrRaLHu8DwiU7V/MTPi1j5
JbB2/2DTLTNCWHJ4OXUSehSLhXPJso7f4ohR++mH+5UAE5Ymy4KGTNVR6dR3UHeLK6LoBLEG3ao8
WhzZbZWUOYnXXdKxo9oycIHOb0PqmStWDgdbFBMeAaSeVGRvwGqtqmgDNpFjp49l75SFkuqiKCdh
aCtqE5gz+yqi7f2dHONNQ8pLlnumsupnEwXi/5Fb2YGwPnRMa6U4O8+YCHTKNsv1O4yvugcbQCDO
W7Yf37E2SD1bPqRqFetlFc+HyfCWkUcUi37Lk3+mO1T9YZc/t9DnDPwKALDSlkOLqV5exppljO+w
b5erYU5A5hfDH28OI/JttmdYfmAQHPvLhDvxPBbZk97LRdByGEPOPF9YYIzgUZ+k9XqmKi47mVWH
HimlDd+6JCm+G8/+gt2BYcjsPIAEA6yD1fH4LOx/BRw+CAI/usXTDqIHBMH13Yp3mUOMT1tjaxql
BzvJZrJKm5TD5HQhqGMdGHhk/ESSftGBSOA7OB4pizkkNJPhfgOMvGQ9Q0BrzfYUbJyZHfT0PEM1
+tgNF53qjT0rEqdiu/jNgxhGF2LaDm53XLBozsqGDCUwJxdsZ2LgKVccZvHJSiQWAE95C0vCI4JE
MGdRHhes+LsAd6k5zzX1BI2Rx/uoxES0E6EFy7NbzdMkb81agthDy/kunfnuZu/4Ua5QW0sE23b3
JH07usZ/zt/AWHXUwNMenOzr06IL5trOWQrWddn+uGOc+2Cn4mh3gU3wOiDazwXNfrFsaK3VHFTD
xG+G0/+io7CSqi941tE3RFgnKV0zQ50vV906B8a7YumPTMV67udUT8cEq7hY8kIlUVcFXXmaIY5c
PkTuiBnRAColcsQNagymvNMLtfR45G97Y5i9SScCE79ipEqOGOpIcJ9ZJfvN6ACNvdCTMh9v8dK6
PwdR8huvvRYaWM0DT1tcbkV2BTF4mYiLnIP2K/pi3qN0BRT0f26s9v+rbm/hbq+imVCSpjdr9gfD
43sFmYvqHNdVBeIaXDUGI/q082Zy4J8O7OiwrbUW0p7fQ7akQ3umu1EJqd6SqjRVQ2MKdb0Z46Xc
cR38nARxTt9smfrGgCmSlQnQNpk4LuK/u3Fgg0c0NewKpVwmA11e8ibfiyXVP6us+FKvh8mqRVYm
C69brn4trsBPdwi86K2JFLEm52LB7sH0OvJiGRpRrmfiOSG3mcsqyRAXOZrg16Egv3DS/sYy1INP
ARYaBCWSNtDlcyirnsCnTnjZlJASiDBYVaShk3XHUhcAZTCYV7G/5F06d/acaUHyx+33OFxXnTQb
sxDv1bQ4BfLoYe3IH2t8mgkSJB3ccCSFOYV5+XdcmgzpMPWMpqZly1UnqPQjrtdSRmHd3zwlhy9t
QixiU15zlhAAkRc/0NM7rXHvFHXL6KEO5pNizYmVpzdUKQOGnRYsVxgWKfNGKdQHk1V7uUXqAv1o
Dw6u0YkoWBlUBZrWLp8lONpa3wdQA/imgORkMWChVRAUkD6HLfQ6CnIceFLPpcCRKe43abkLmeya
CnZFdeFt/kpFkwg/7SNoxui3akH5+0n0tcTkOATad0UIWIv5fe78E9n2gBLkymFRN9E+/d2nP/A/
D4+MY/ksgmBfjE5wI0/3v00b5lHNFdZg9erdGEn9gqNacaK4wM1AgPMqXB9hBtchhHHcQ6dx1JfD
EogbqMVIhT5eY17xHnxqIrnfAX1N5LQ1Ym2dFVuv81bDQAkTMdjD7z92c7UWviAwNTxVzL763bga
TSCRjIDpM9QyVDwxdNzkIOwlm7G7mSxzZXEDs9DEuV8rvanW/WhxoZXoAJpU9BSRzHrspLUY6AfX
IS9D22BgxQgCHMqDOBiPtYQIHHJBK68FCQDetnU0lTqzQY9dGzere6KDnbjEncaBEh8YkQJdzYV5
UVaV8ilmW4TkkzgPotQzTORLFE4Ee3eoT6HlMse+4OtNmoN+EqGi0yV6iwmxu4ppWN0SIXSE2Duj
gSyLE2nplc0kCODMeA8MJi24TX6KkiqsPESRoEZuIKDLJxwYJ8TErX27NBrOAryzSa63M8zplwkE
9BSyDod4H+ivnI3CY9670HHBT+YwMdbvro9JmIWUO06zjhZYQNqZpt5SdRpHWxV4UV64XQWZ7UTE
oupn5jk1gKwSa/sWzeL+f+3QKa+6WOhvFBEaSlmhkEBMnTDDIkb44F0TCQM6qZob8YIMkPCRX56X
WdRBk2YGgCwXL2qWIGAYISM3qCwu4oz9rpHBrvLudFhYGeizLYQbAh5ln7WFmyFYqHhzF7iqRzbu
VW1Rsc0PmKq6d5UHi0/Kq5wAHw/dEgYy/4iRYBhCi6QgIsnTQtwT31ZGjvVcyYDiE+usRlnOKwV+
XDs5NgEb+HunXgLk9qDzJfRhzs83mKYxbhvucgEqdZsoAtz3Oos0GcbLoPIEYBp8NtiaFs8w02kv
BfUQWTk5+KqLXthwZzCE4aLdt7hv2IETMqi3CbT+QSqensjDf90X/5uvXGpqr69WmgF1IpXCIrC3
MZwprW04l+ifq7Q1BdGgf2gROcxBwSyJBmiw0P1DHlqDpZMZ3azbdN2N9E+AB/U7qmt94jWcnMfP
A8uoIIyhdSUrrPDcpzBWc8DXE5DmEsl/Y6Ht4fRgkXyo3oSnx1ysWj1SWiErhmyhuf2co0dRwgj+
2aQ1mxuHGQIDPgdJVb3kDdcOzSkUKH4VeDPbxeMxW1rPXTZvjbpXTpmE2zsQHrLqkkDoELWcxabq
pKk1fAbKWIvEDBDQvOvN/OhSoWxrA6YQl8CoksovSzacMAIzicz9ehtcPNl5a0Z9QHOVgSkiykz0
/rn4lzgD0cUsZnxkJTOxxaZOAUOTKzd3UllwTByAnLmnYOqN3/RzumsB9uJM/9KriBCzpffPOU7W
QjGHb7AMgV/pcYlSbruBv7/ickyD5Y5fArzXkoO/69yonhIa3WLG9UeRozwZwCPBlxRHeVvsPfeh
l1P1vrkK/IXi2zzqRDJN/A9NvnkfEoAz7vl8dk4igiAN2x6999ioxjVl2vRuvyTl+7+0ysmhmFPx
1Gpu071zLJrDFbwbQxzBMJVvQV0ITDGQl7dJt4EUkj8RMN1ZTK3kppO+NVtqKdFJwUYY6+cawxMF
ag1SB6uDL61m/FB8asfpbL2wvzIvZLFa0F5DUHGvo0b97wBasGzKh12qC6F2sZt2Jrn6UqnxawAR
S7Z+C3b2wLCLKH5cvFr1TSe65Ybspy/VE9/ZtyQY3fWNKtoMxrwsUy1DAt7NpnnOOoLHFvBIMjUO
zq2/hS55tMwkGuEhtJDciZsQq3dJSEyfbmK3+v0FGo516rMNJIgMPAw8FgK3TYls0LTXwtsltDFg
Ipt/MMAc3XS0wF8Q6+r0Ai+Vl+Qpy5o5Q8/izzRpeW5TxN/zwJSo478I18gztXYZ34JH+guPDUzk
37VvjFJ7B0CpeVdAQYdJlONKLxYVwdB1OvIuumhBGB5xKUvZuqNyu8nQYWv0o+zq6RJWeEGoNZKx
RTtpl203fThdhRZcR5uXk/nZcxACZowfO5qKpyDJJizc/i0dHunvyRG2pUPu2mj8/wdcx4X2Mcum
5makfmBKfEzI2vLVjNfhl5c4Om7QqVCH6x5gDVKYzvV/7NyazF8GIlpdCzGfvf4gOAYOhd4+M6nv
SWXui8+8a3+cj/vrxZSqXDZ73lxy1X36OVHbW0W7r+lDac+SmYhY6D1JwD9KhhJGrdxw36/fj2Cg
1HS/DhXAwbjDzCQDYHYhivP7WqaG3HEojPIByUuziOFd33f6pOVPfdrPrp9IpUgF1ZpzP6ZaM7IK
mt2EmcgAyMHYZBIyrWb3iq0OLUszCp7ZstXzo7jtWcp+2UcbbfQJ5YUtpcv223ex+0H23FSX3GW4
SEMjnbgwvPtF8XIKc1kKkWLLzkwYGEDG5GgbJUt5TK6Mss+43AW6ugAjX6OyPsMpU7Wt6TtcgNpX
9XSyokzOak9doP5Zsb8MwdMNURbsMp1KcEMOXJqG5fklk/VK69iXY4dscN6O/NG5BMdjRz93VJTP
FCyCksksKFDc8ko1PUrnpusoSA/Lf6HeWHUFW+J4Ia9Q9ujcq1z12ZQRJmv1UvPf36Nr8DxY8Uni
Z1zDEb58CIdogNkisC64B2WD+hQHeW24iEPvfbfjaFn6p1ihB7jr+siByihEWJpymXJ0nobYtjUS
LyauG44Nl6puVswdPRlMg4ogTnqpJjdpH5HBr8ILrjJSYXdcuF+MTBmklgSPLxsjFx88PAqenQ4y
+VNXPhYz247p0B7tKnAMyMi80d8URU8keqk6lHhxR1Ui586GLltci84/fsYetCSTVYa75tub1tph
SnhiO3EKl8+wH51fAOpsHxMxi/uls22JuBBGsKDp5YBXrBz9Jb4kHT/vkdsNRpi8cvPp7INwL6xJ
xXV+Dj6VZ4EFC7LZGflsbUmXsv+lzgnO4t6ebkR9wnok5x+icPv3bHjacaZJQvhC95dPVYR6rStV
9+7cU1ai2YcIFpUtSBRAEJ4Ti+hiv53VNYrtlDa0+hec/4vVLYolyEd8/NUThJC+RM/PQwI0d43E
qjIkB0NGsqwiyI6+mA/NeSoePCuEqgAvRcO8OwTdIxouZ5lSC8PUKCubM/8YPJImv064POKPfUSA
FUAAmBWjTeBr9B1jgARcqgHepAo3cPvMyhx5YiObRFaWlBFU2SSH/oFbpVMAfEXJUiw0hWj4utmW
0AqW5kG+yBNEvbTN/RAe03ZYFltDB0sZZRmyLWqEC+iORtHF/LSql876OOsyfwHEwVtfuT+qU1rf
wmMWHBpWqNLX5w9JzYi6wHzVjbeNfABK19WGsUWyW48XviIGpO1rpe8DU3mSwc3Z3+XKFrAPHohB
g0WzcEsPpWj9l1IRMsfxE/xqC0PRb7TE9dczLO8orXZiIbBx+6rhp3+r69hTAXmdCh4fBnWXpouA
StVb8/Ca/4x6+Bq6nVfRNyC7K66fLz+NJGhkTu9AE1ZCzWsa4YdZK8dJ7Sf/T6KSI5ziVqDw5ZZJ
R2vO5nctxceHcZ9OstR3aBuIdvkLehoPYSgkrz/1W75HdJT9oWuAZ6dFqMUbyzlJfgoEf9it9taa
oNKMHzk0HMZgYIjtHAcH0UTnS4tDk7WdhyEKfohEdCu7vhPPkB32piMXpYEOtO0ngOSMfWOlOXcP
flqzAWrtM9Kx8ynKeXgXWCkyljvb+RYNVnAy1dUbZiimstMZhHlyYDAcWPhgxnVXnmSJr02lytID
ENk44kjZegqfUpokO/EbFDylOfmrGw9WrTuP4C783e68jz3znz85zceLawPKT9oZYuG53Oaf4sEX
IebHZnXV7CVC9idHRVduP59fwOD2zseir4YJ9C9nFxGZy/0rop98mI8hipriCGB51zJFBtE7zKjn
/mNOOXJLt1q4avgAoRmxbci+SRDn7hvhdWwcXQkC19gnC93Yy8NrkQZvOZ2yxvqoFxBIRzxUDH74
tpoJ2E+SMK737VQsjrWc+TEwbq/JgWYpNnCkzm1cJS2NkspuDLGw4f2ywJi+6ubDie/mBR3MW1vL
UlVtzRXAwKulTwsklLIOFUuQJOEtWWFMdBaxhmeKqD6sX+WOgBNEAi6VIKcjB6djJB1S2v5EbF6d
e6PgLJaOsGjMREi9+YeLYED8fq2up5JUKf7Oam/hbIRmYhip4q89CLQKDcRXCP4gdCGYVfo1QJKm
1yzRlSfbT7b0FVLTla7OyEtNvOOQ3z0/+Wj1kD3iF/IAXP3oL0ewlTFunGATtOzoV3C6NVdR9AvX
r6+wawIznz4zSpBcWCQ802SuuQRcEkMf643F6WHoWQeXlfnycUf+darTCkSDNLQP3PFCXQsC4RmC
XDR/56qCgPx+DWQaqLw4Forgg1wganWzAGiYDBbT/hcf027/ttnY23YN2OqRiMKdPoi/kAsyG6P/
lEzNcZxM/yarbv2gFCXDSIqGAVx3auymL+k48AkSw65F1nlof56ZGy4HFPtGUQo71Ji1ivZ6+ibW
O69WMkXEnN9/rjc5QSTFtgKw04ITniPVRigs8vjRjbCIZPWb1Z/Gx8C4L+yBkc1hMlLB2leqoUFP
gR5i97kRJYpl7y1e02WAYwPSXA9zTTu6iipk7ANkNfM3ssRHhK0hGlBNX9mpTF1+Lp5rniH84oK7
G+ZEAdas3P/QJEwcxSoVIkaeXtbAvwTCn0o1MiK0BBILEcQm0t6qE2kC8NFm2MORvZWPDAuws2kw
yTK/3N0aq45UWgk1vfl5oOBxhbLvogLXkwKJs4VuKwpbBgXxdbJGiVWlV0Sc1DQ4jmtSCubz9ky2
zSSfG0nE05MPnSussBqfcvOkdR0pAeQLbaZew8hPycdEIDbtHJPd4xZg+YtXBc44v8ON3uh5wQ0d
ZWK30g5m9JHRUQyINlysaxNpF0FRVQtArDEvKUzzfNb4zgJsiSUpUyYgBMUrAa/a5Dtosxw+GItT
WFadjxFfHOgL2Bdc0QQ1dhd/lMky6uDUhKgyyqoPdxBoWayx9X/gMjo/DMQmpdIHd0uM0ARva7nm
6ARg57HyZWP/hCUnCNke58LCKEGGO2yKxOSvuwh0XXVPjE/dpnN/S2LW5MMaRqcrdiJwUJn/GZdI
KO2BBZXLFfBf1a0fgdvCNrp3qAMf6S4bGhA7UiIBJA/jUiFCslhBZa/iBQddfeeGJQDAR+oK/+nX
daUCGv1QrO9YLJcg8C/dPEOZliY3aucdMkubPrl2DDe6BMU+CHRMlIli6/K+Gf549JvbemLsTwFx
ZUwY28/d2GCXsrn+ZKymjWy5pZtDnUBxtNh1vAbKUvE8ZUW6ZOOht7KfsZH5M/iazP+5s7JvkSe0
hom2kibJqlkEMerAxNolHF65feYjS4USWFLMvd+kX4mnPOPdURl1aMZWPKwRcEbzocy+gpbQAdB7
ushBLIhEszkDt6KNGCt6opOnuqMR7O7S0W/jhPxk94EfsQ4xyDt3Hdq+0u0W1QdPz+LRftdj2KSB
hS6jk6HiuSIoGQFXv9/SOJd3ecwLzZ00A3Wh4tzlsxaBWPQNbsy10085FQoA84FXnwMQa4/uvTB8
u0AMAyIVtLz/DlphUd0tzlWG8pfASOwZuTc8NOcvcB0cH54g17uYh7VHZpBTzEHxxpsha5gNRu6w
70nIE9Yb8dwtbZhyR9RzP89dRUXCebAM8INFC6HZzHxa+k6FU3iaFaxbeWfLPkG+8ev8aQqnj0fF
xrzrHIN19pYDa9KW24bmdj5ZUhKiJqWqp+JORylDxoZBRdiq5XKYp5HaxcknzDiCR/tX8OYQOxDJ
37ttcWvmYHFZVH7mOevnjvsM62y4pQ9zxVgflT0o8++g57rkziYuaGOrOVbauxDy34iyV5Pn3qm+
FeuUwrfgNSk9ovKFDL4fr/Pq1PPt7wqxND/hv7pPJIWOyJz9p9iCjqwZn3BrkZfzpAhvwjkttbRb
Ylpud6owycRwV3ffvha57V5Ux7GWvOz1xwuoEaCvJVdei6Rlcz78WUryQkwSnSPxjsFYxBQQ0x86
fzMOmwNcEyjF5UIwZaky3ZMxi3XlmAMBD0QEy0Zx5aie3lURrVkuycYWnEk+A8SHK+Z+9OgTwkR0
h+wX9CBz1+aG5DUOBKuJfQFrpz1PRozHYUhFH/oARdIWRK2e2IiM21lyLLld8qYT12GClJtjYLpg
XHtcN8khP6aGT+AYdewjwuyvF45fOtYrqbQW1cBB7r7HIrz34PlUow7Zg+YDUNtm3bdUkZRauOtL
wv5Q+zgwDWcqO8uNkjXXOTqiFlpTjZhuvfm3oVj7P66IS0EwAm8v+uEtDp3pVHrTMLbLLWjCEqgg
IQYky7mOItpbc6fjY7cdPXYsdoyJQqVc+cEEAymrUP6rrQryJxBJUK9ehUiFOZtrHKBrUAZETYcR
TqFhtPs/1n/LJ6fMgY1CT0kDT34fSLUuQTua5kRSG8ow3gmUR6V9aX4Uwj9dwdEr558EPfnI6RkB
q/UbP30AxFmXc/36kOM/0KXpUHhPgU/1yCoQCId5WBmaH9CqMl8rHmMyI96MlvJi1s4RkCUUIJ+2
Q5Cu0XoUTLF3UpkOwrrNHjlutC0sxIn2y6xI8xouxminzsoawYk2xA9wBEpdoonjqbUskF2wPL30
MnMlfvNarz4RgoZhK0uzrotqnq4u2eXruWnLyK2MiksrEJ5z38h3FeaiTasszP3nR/CGEg2SxxLj
Z7r/nexZyN9BF3pkD1fj8IHevfi2QWeoycQ9OHUJTs2TVUgs3N0p/L3xJkTTGebasEf4YxCcBFvM
3iO60PeDJztZNch8bQmUREbGHau+vjZoP++DnC/Pg3V1lBE/yw1K7fQnBxiMQI8evzF5++AjiwjP
mUAQR3p8BBkxkZ7UnJ9pSEIaF+rpWU2dKkx9+YcUWigaAfJzco0YnMHN7frT635xGS/wcamQE51F
B0OhKtmByBabGtdVV3idTBu+8Mt+lmSPpKj8KkhL2n9XYuxUj4A0/nSwub8EE32vFxJlqy8HI0Ml
pwFQrCudfPsUdE2jDf3BLv+jv29uxiBZWApZwwhVVMhh6WD52MkjyT0SAY+QanEukSkqUqPnZjir
mKxOOR5vC05jJBEk6iz9MGdulx7WooU1tr9OebfK0MIzVYPqGpBZhf3NAdoh1KLm50v3FNcHWGQp
UrZ117g0Nlf4qcoTeTjBChb1djGvRCkbBFFTOF+Mt2p8zOCrsNYAhHeh5NmAAQsR9Iapi5j4JM89
lUYYuX/tk568djEpSJFI74YNNMmCMVYEhQIDmD0mSwCoA0n/gcmNO1/z+nv/fiNkKGZCbKBAP58b
YHz8SwsXSsRaisC7SK9obfaZbm2flBhfKr8l1xH07oK1IiSja7/J5UNQFwvw17q2Io8lyYkJERLr
Cu73WGOG/RJhwibBvwELZ7vZfZnsbh+/1CEFMYalw/udKES7xmULsLMZM3kU8MyzijEw3Wb0ClvY
HowwCg5P8yp7lZe6dvfIhhL8juTmGz5OGOT8CrHYcz0rsPNbb5FWobTRCKno274bNdRQpIVY8jko
Slu9wxdLCNS7MJlZZ9mfV3EFLyKT+ISVoMlWyW/hi1ve/Lv7QU4Dnm4saP/CWTjVfCEdsyrM7lDX
lUbv5JAWTXckxoZCltAXkUJsUNWGIqjmmD5RgQOEndWH5Jn1TPY6ydyzLD8eqIJ1SGFqlBivs2Y4
OZIuvC0iRYfj9WyUq0G9G9lsAJxw+jFYgPNZNvxZN2BqUuEsBlRNXs81pT70CvmRMo76XtScCVO9
UlnJUvnzpZu1+VkPFMDr+3LVnjP3m5fbyhrG8kzpIcZbyuJMEQaB5fIgaWAUrd5AJAC2xeRLE4IR
IbPOoTt7rMRS09U7D9WECFmi8GfeTWBt4a/wHYYpXvZ7hhtfr35G8ewmddQHBZammZOPi4kN9i9T
UZ2H/SpW6A2+7AJIaiRdAtwJruNDO7odZGJiB98o6/hoGh+Cvt+JldApTJJTvBw0L+MnmE1ICY57
kjpiWDHFFsvJ0rtSXimrTeFIwMm6FaF7w/Yxvg4voHcCO+Z9Z4r+CHRKjRNXTsQpUdWtph94KUIp
IvOMdkxkJ5HGMwJo7KD2VQEpSa7XzGyPZU4/LHvFlkN659bXbpJBawVJiX56HPcGTRmD1HNVsMZA
r1hjPKrNUjDBhB6/aURyVwyM7kKhR6C090RES/5Tu3dygYrOkK3Tqmq3UERmAXqR/e7OkA1pxa2q
zGIpPtB1/Sw6Xzkbcsu/cwaY0ud+ej297XQAOoqjtkJ5M+2zxg1eoXU+Y/DkyqbTZBvmCk7xnqD3
0oEeVkk6qet9RSlbqEeiS7hIYcyEZsm+MzihUlnHBGyRc2n91LerClUJnGzbuL+QX2h7eRw3cj/v
2RCg3OZBp0LezgPOXOBGrIosbBfHrfLulLKjGYsF0b6k9Amk558/5CU+3o5pVELGzi8aKQiLxtXx
tnFCla2VOthy3au7YmhiHQ6fuGe+QzvJ0zhIC3ry8qwbW3h8oIsoHnjbtwiF5kDa9qX27iCtxP87
vl683K6jqR4I1Nu/F6HilqTKdMFOWVJChuzVmXE/FHMq3h4gqJX4avhtenxjGJMfye2f3KFqntva
JkCwNcphI7vo6cemQKqoT0q+ENdYXr38XhefnH7TKd4wP+j0rCpJ+S1unwl6NJCjaDXF0174kIjT
CjEORtNcXJY+oaRfaXkMOz65kGl0HXA+9QSZaWXbDBI19XNG7TlJR6m86aFrFCHi4pxat44CxvIR
nJ0wqy8WtxtPJqxRanZNWTQwvFD9PJbTYKhPdOcn76YVW0fq4xAxXKLOyDQT0Kq+nscYml7vxdgn
HajQCzGXXQnXahlajZxWp4ZkXMlXnuUYnsJzGLZqqw5AVNl3wLxqib+J6D3WOVkKmLcU9VfL+0Ww
Wq7gy79jh1GDHC+g85kTV4GyRR3PkruHh+CoHIX2WqbtyfxGOmhttKO26W8NXjMmhKiqrDyTr6el
t3YFITRqDJmMbNXcfzZfvLxH40JJF8qVFDDTt1xMhoG1AxGvF6oerFSf1nVf5RgS65A1wBviRBGW
Pp6Iz0mDarOWzdb/8sYxIhHzE5oHTqYFvfBxON4/2H4s4DBQQ4PXczhyCDo4fAbcinq9tWwf/3BO
bMzIo4FcCetLsgcnnb6hnhGEYbN6D2BGM2s2k1f4EBB7caUKX95BBJ6307zMDZVxyJPnoImetUYy
/s67NvvYfWKG90Et289GIPMd62mtjQ0AAWYfQxLpDkiWOMW50tZh6YMNSK1gOqGNTKJ+/EMT7M9K
uICwrLuPZGSQz/tfEUBkpGKno2vOP68HMQpofWimo/7XTRB503b3xpVpUuUhbbceWrg6zQb/dft1
VX2EaDPLa4z38P8ZLUGpNixHz1gELz6GyyuWL7ksSFruQIO5S+zIAls2jzIPCY/EEkFTesD+qFHb
J+021xJHohmHNbehvanky8AAmb/vefrgbHegBemxnZ0wU+sR7PsQsoYM5x8GmfGbhvvyvrM+69Ii
5OGBvML2TuvUmzAUzqDcq8qoYHsdbcBal+PPat/YyX8Ew56kzwBJDAs7zWs1O0xlyhdajXQxJDiR
KTfGy0Gw3cHYdnu6RGKcOmYCj/3eg0rw7D8eK68BBK2Z7xBETb/pssDZM6UEYp6Lra2dMLtODgsN
bSr7LtpWcZQGM2uhq13w0GSuJhBPl+V1Mv8OwuvnJnVbfA+0hodsZ30N3k9Dj+lFsq9O3W3BAzbp
5lWe6Zqs7cbyap3uchaFMux8WWLibBP5TbLZ9dZwfCrpkRwkEE//+l5xyJRKCALlEIIdwe/MmOwx
5U5DGIpmHWRgaCl6o5YDRk/e+fRink0BdQ0xuZAg7lJgmxB9dxQNDb31gug3XBpoREzl+eclMDrp
g5FArHZOYfpwE4KZFpRWBrTifuxWMHCe/0/jXePZKnId83OF+2+0NiT+8sd3JI30w5/Bj+kf6hrS
UdM2ibihi72/iZbJiCywG4KDxjO4Pg7Elh7wYED89Hm4Zn7YAK4WNPlMeO2kep3ba6n3iWRHj/2e
dtMuDLrYfnjIGPtgpf5NJY5Oa0PRYb02MBHec50DcMx07byZ0+YLnAzZtyl+gvUa3/ZaF3YxTDoh
ZH2eTonMzdwLprzz+63PNjC9OkkTB7Mwu8T4QQcP3lqAZJBuHvA/47oLTrX2IJ3brTCpp53TPyAP
uGlqziEyX3BQDeLVtZRjKExyny3bKIsKSr+oI+2rJ4miMg+M6lstJJfyqWuLYAo8oh3qB7++2D9W
SvhoYN6dXYyN4lCLfkbjRGMPw8+TvFYA0JF+bViOPxdSeYrWrUr6HzPzYvhJrL84e1bCPLnbZxzb
H3e/Wc0s9eXKjIWI3kWbUGbUSLzjIeuckR5hB7nVR/O80OGqwmaQrYUN9eJ+y/4RDEejXvDjB1+m
PYfKoaESP9Kg3LyHLLebod7A/MMSZRMgIMrJI8bioaWMyJMG433+v1zGlsJ6iySlArQPz6UZsNLi
/0WWcj8vWhyLP86S5FnWLWQzrNkGQMSTSq95bSSZVOPfxVNV70V3j7jcLsn8PABnnYYayEwjp8U3
UKYrdoaVQ8YJG0t2H2ny3py6KOhg19+csoo4phjfNAazo6vnvARv20dPMb6et0PDN4ndEM/R3KVq
yUikq+f7tUO1nFcv0KEU6ZsqJsQerRE+5m+/Oa5pyrxH9JFxN3msFqeHa2G+Zg0o5CKsf5fJxXM2
CHqm7Ywjh8mBEchJFRdXU0giy3byQJo+ts1854Ui/ZBRD6kxIyeJ5Of/sWixRymhSyDcJBsv5EgE
+tBGDT9TNC0FSx3zasaF7u34jaPIJtfmwvX5eVg6mPTsPNhshZmesl7FNcfptwrF6Q19F/qD0s8Y
CWCZsUaBwfKlow3lZfPLFKZJxoMrmELod3FPNKXvGLFt/9kiQWB0iMqzc46Jht3wm9q7LSWVSyJF
DEQfbPAtKJFnxs0Eq6qFX4Hr1J3IFNUGAjzd61fm2gVBupR5ZRFaHwLsHmV6uFD8S1m+06bVMvzM
Mg5ezODUhcLbEtcgdwKcN4hy/uGmVSzGVga2UkzzoC8Fqzh8/r68Hn5AaNmEpX8OIwg+s3R35/Wq
khbtmCDF2JtFefhwUWXW8/pKuKaujoLqg/5a93P8RZ1pSh46Q6XexXlF2OlmLM3qFy3cdMwTb5+s
ozdLZOZalAwF4wlBlRPHf4D31xedSLo81lTeTB9I3VEFpQBQ7bgXnsLDKLuZdQkjqG6rkNuk6VUg
IUifCHk0jdS4TJTZJCr8RyqtJ8Kc3TnxXQ+ahNo9N9EM8aFSZ3ZgQxCTH6ydHe4oiNBGSJOtaQwN
FXfs2yflc84Ut3hHPJlr1hVlBQEwNYFf7HtbCcDKDQaNQwNpeRCfJ58H+Oy1l/udZPtS8Cig3z2a
EZwFKmOIpHJyEKIEXl6D1REToCIUUrD4cLIiThxAje+AmNUC1TTLu9CaxcluZrp7pz8loE1gQUxa
OV7CGNhASzZGpRr330cUFQxVGsAipZyFcWPtbD32IGgooz2US5xeVghiXz24NsLMCuOBjD8nGjIt
pDqt+obeSASI5D/XUHcE3uwVSSxzN/Y4c9PDYZd2K8sIl7CKeocU5Ed7N6Hgydo+3kjz7w/2XuRH
94ruX2pLOs1nijHaCT/VpchuEm1nIOivlnqaDjDQIMVn65BoZPa5meUkQCafRHCmnnbd65E2/Lq0
DQGjQ2kAOTAH73SUdAAuoaxXSusNB8ZmdHY2cHF/rtHeg2t+DeJuXgC+FgORI58GvAoHe/noCCUk
E8ydUV93iVaNKOYS9sgcHLoLvOwSW+TMxzp1gIS6J/ma/G5xFBWnfhRUED6iHVx2aIyhYtTYQeR0
8g/DL/W7/ABkpPqi/G1krAXUw6k8Fs32V4KLSr4rATS01BM/2Yz4q8IcIseLCnLH9GW0QlrKi7ue
OcF99xks59R3WIoY98gzMvbKprFdMPNvkSl1TmNXDI6Nq871WVbJItO18i8ORUQWFwZc8owdS2at
/K1prnCZFdjTirH31j/ocEocBRK26BZVn6QeLWB0jNXRLlbSV9Meoymi1IyleoWTuOSvrOiuX/4N
xUx1MYwACLRljiSi5tJyObm4rmQ82IUHIvrY+AALNXl1FTKkdUkgESoCyasVQ0MTOI4fWLa3dMgv
VUS8EAdOKrsx3LdQDPT81wbrPOLc+gVVadKM4oGQcZK4MLgEHpMiY1wIIH2v8a13xXVwiyPtxu6S
8llL+mFTOA+axo/1cKlYOEBp7pnRttE/qSDZrAkb83PiAU/7ytgKLba3EJAlatagSbX15hgUIPkL
9LcEGp7g3ZZNXF7ernsFkT4L0GkdzRN7Pt//Tm1l7BlJZnYV3fG/zAV/HA7ZWVWCDuTaQkqKr6yQ
lQF7sPFUMGmsHv5j2ZHXJP5//mYKS5XC8TNdgAyX6WPPSRy5WbmbkiI2g3+K9DxVObq9IwDqQCJf
zp66hHXqPHC6Pkzr0FXdbzW7MGXs0STg3yVn1QBaHKg0cVF4gQ4+w65UlMOOdJCj0A+tXphIMq02
fcmbtT2pQiqCV028DLj0PJvqfAk0A8Tc3Nbro8GuDjMA8VbOBSZoZR2FC3vS3vSUGPZXB1QI0LMp
fgg9DwR8mNjn/0koXvju+AaSxIuwioHVWwzjN9sNwQKvqZEmNy7iM+sLE0F2IvjTMXmialp3KbCQ
Cs7Ukc/HARf/zcp5aHP5+dMxfd31+mWrcgb4lfBaepFame9wZSgLaD+Fyn3wSHXzdAr8i2qCByFD
45DOP10fkrm6hq8jMfv6U8VKVJHbt9FjPlLfeLEVuLCViESRMVMdbylg5qPolCS4P4l2bUdk2XA4
oLdkrF9PjJJKtCkM3xB7H4Athr1u9EBQbf27r2GMY5TGmXG8v/uyJQF3d/DKIcRfRJ/XM4autEBb
52j9q94NuViCHHs4bbPX0nRmWuIvMYkm5g+X2KNxQtKRAI7mYY7OOYcchynmzrTDx9Lfi2pWqfz3
4aZ+hfDzLgaUu0zK95Ongq1AiQE27F3IcLNuE9FUApDRCT+Oo5Cxs5A30xMI3YPeQXJoPpdblc2s
aFlKQlN1hYGRxcnKWq0zeAV8G3e2+doTZAZEM0FI6a3bz+ne2/V7mlkBJMXgYsdzrLCjZTco1jKh
0t/QESd7m2r/xMcLRHGhitD55FAjHDHObGWp/f5NopLjViUblfAKXyl4Iw672Ci0d5fri7TzLH1o
K1WQkQbZBXbxjZmgI/BZFA/JVw9wK0pYAqjUpTy4EaezMOQc63nKHjUqlzkZfq4ZvSVY+QeIaVm3
uHoTXd+kzaO2f/BkH2D0tUmNga/nnRx3wGydAa7dj4aATFJpLNdF3bisNuVASyQGUAS9qMb4ZP1S
dcc9Vr/WXnnpMw9z82ADVrt45DO99+oPzC4igfVhHiKbPYhRu2znU2tCpKpyMLlA79sIb7SVWYCi
MmzY8uONV1ZWlEAJiBjWPkD2IVxg4cmFcVCuVtaHSDSWQ43S9cpZdbBBzj/fY056p7HW90Dw5t3Z
p/OX1BCxKiIPwXeNQIOcu3Rb3mOwZ08xwVEY4piSsN+Rg3EoqG9GaDfObf0bdwQI2DsngjEPSVCd
0Qy8JmAJYvqoChNVc/fCnLnRx91UTGKrvXz1yRQ1ZGC9Q7OMEkWpaCLcBJ/TrdUF8h35QrHYpIV8
UJsD/vNwaiO5e7BB1bPB3LZvsWBoyoRD683/FvXpqYoekNXHIaREGe2hCfAaolU43Tx+dQtsVIRd
0R7+lO6dTh4aie7Abo/m5ZsfgbXgeMvWWGhBGbLS0HJ+HU7NJ/3j15x4WhJqBx7HFMH9zspFPJY5
v3ESjFT8KsdnAINw95cC9HrYmtKJmeEdwxkLIyxI2ngy3xeSI/r61R0FAKu064qrjz23OJAqLccs
VQhmG+9Qn3XtiMxmizf1iv5dNDhnB0Jg2WENYmyaFzu+nQ9jgEDsyZA2A+95IeBwGhgsu3JUDtu6
7jzATyG0I5qG8/mVQdrM4vHltj69NnIN0hW9d7XV5W4IGmXhy77Kmxf+3vAY1IyM1z08A/SV+BQ2
3pFM3HiKTyUNyupjuTEX5vNkxhvFoAyDirEwTs7ouBcDy9njg3N9hPoa9PqtIfKZ0DDW4U1sFtEL
zH3rz1Wg1VN/junMDrCx5wE527sBgHHMdx1mhBx4iCgPROE6u303KsMTbxz3UZYRqAD48Fb64rJZ
QmsmpZwJUk1MOgpWdWnEDjVHT8iF3unXqVUyLdpnWsdwbDrDigV2G9A19ChATp0w9QBa1pPv4BWS
tYIstLhfINR0kRgjWp+c+lsQvpcc/J3PjlAiPhEnz2/TnLUWgQ1J137nWxxz1267p74rAhjuxM/A
uFQJszf+9aFpia3ChfA5RubAF/2UFew7O+x/hcCPMn+StbCIz+QVtOrzlOzLkm43GEeN8Q4RzGSv
ItmZnwQZzC1mUSCmGMEkL77N91HKBdgLcj0Op0Uabm0T2KTmkc0eMaBwOzCQVRz6Hf5jtoA9wlRc
yxVqXMnLZGoMBbtOFSsL/d1nOQhPtr17ZKkCauQHyNUwOym1lL5Mwy8YLnLCgvvyggWFkItn48II
MNGcGR/Pw6+RSGvi8dxbsG8SBAkb4UmaDSEnEES1+38E8rNM698pVvoyaWr/IP+iB2o094pzpYjg
cnqqPpnpuzZAuUuMGZokJ/8qtn+4hjdOg1KsJM/+1ZLLz7yKki0WXeNi68QS3NO2ZnTw+FbjD95W
qWYJoXg8aBB/t0VaajSecjix+iTIB1siwPzUsfNq5rRdMz5MFi6onwC7Ejfdvz3sUb7lMw2GdSC1
ml3Ye4ADUzP2X/yUZ+eE1dyCykA1L8702GohtaeLr46MnorLf+aujZp+yJwGrxckh+7VhkrU3hJV
RNhmVxbn0Vvml+taEVoFV6caALL+5i57sy5jjdjpLIEn/SHCrS/ZzvJ4TVEu3IiOzIzluZKMRiog
CyRVaF/qNxM/dlUhIlZ98PIzqiSu3vcS3HlgExlqHTd5OiBj1EbIiv1gNyXW13/C1KBnb7UzWs57
2q5yOQQbNwhy+MEuAOAI/NlcsWHIirPXAT3hGjOSox9n+kHoxJPeTzvW2b3buCb4RjlVLB+pHekV
oLoM6y7ZfYdwnwCfkRsi0lahZjX0CgR64s+4PYRQr8J5bXE/saRUSve1+5SLTOuY+tyFye6xRZzg
miF7Gs4lmopm+AxADODH8vJZBQH/3mGPnmFasAyZLIBgIMh/UD/zdk/Aa5oxa4wwW5BDOypattVc
LtUd10hpYKsklQyIkaq3NT/BqsNJGYyaUrGM8HaaEvig6FRcqgCYG+nw35UEmraNz/wslk1do5GW
ibES8YTOzzwSaFt1Nuecife5YiDc24/ghYIbjolF3Ry5FquZO6nnmffQ4XWuMs9XXpeAXYZgXpAY
i3qSqE/PvR7vrefsaHqYCIGdpAopCoRk6UBqseAeShb1FVienCqepVero9WU7VpMuaLsN3hu2cHs
s3MRiYAMFpak2jR0uQmALfvTvjEbGbbK8RGnKr9oIhCUcYb/GjnwzbDlZW3jyDoJI4mveC+ygCvY
K3KiHH8/+tF6GdKbeeGK2HQfrskN8DhXfH4k7HhcS5Zo+uFdZFEbsX+4B7TEkFfxKaZLMZZt5Nlx
ITjGEJxIvCZLF5PbIvcEd55nAmFYnxr47r1eJcrTzS9Wc11jBMOuWDXU5uYyXYvt2OquZiUbQ22q
rxP53UTpmdwXJPL0EfjHjQw3ZYR7Yg8fthAW/TDhGvFrjq3DljBBk6k07168ngTxjsze9hXv2SLq
IPW1IyVPV/AoXRdOLsH0lilxz9cSBOTB46CaVq550aUFgd0iYYlyot/W75R4TjwL+9p1jxBccoVI
yEk2pNeSStYU0Y8nlYZv28ITmGbmzFGnXDnaSf7xwLTUZZWMjVuJAtws7myDm0O1t9vysPO7Pgbb
X4Ram7Q6KkgmY6JEbX+hiDTMScvqTxFGtq1icXRZe0cIxEBCH/dWHPcRnYduRTIMb+GJeq2gbMe1
KSKVHonMPtDNww5KyMRTEWDNShW5bfnJtX12H6d2PkBDgHi6Ua3W7JnbD+EVmNtSWExyBnHRcU6l
ZkzTxXcu/fIVloJB4CbcesOF+JU4wgGUuqOgv9UIUEDbAysrJ9s3R4Lh43aJrTaFY6fr2F79JVfG
DT8rVIr3D8hbWsuBS2mGd9zzz5Y7uj17IoCD9NQnKRIuZRPrumSQnzkd2vsFV3e5B6SrvPLpH41w
5m9IkVkDI+yfFbIp9OyYJ3VjBwhC9rQ2cx5jNciL0weWVEZ4yyWMckfOguyuU83ux9bHrUmDo4wY
4gsS6dOKRUUT8wFYdYgHhOmKcWT86jkaSq2KvN/c8VpkS3nuBnAwgsTAqvo/4WePGYBsCfOjeftJ
2EWQVKaoFYB66rBa7qumhGXQY6VWz0S3MofrCBsgbuU63Fgos5yzX/nc/KM7Jf7oGbvkSGi5Pyr0
z3/6hVE2eoKx62cJpU10cfKUIOPVenyKvbefFrTT2AeKtQ94dma2XNJjDkNDZIvE/uyuoHoxwUXK
3car7PndVL4VuyWAEXFh5/ypL/xjcpWyvJbVQidhnK+m0Aohl3CBaHQCJNioPDv8XPZW3+nAmmEx
GbIOKA9YrhmYHSX+P4jE2ouFp3OHwsSVt9GcqvRf1sT6yskb3OCwPycsskRVbmG1gbiWf28U8T6e
4vXU35t4zm/gJo5punpPFCuNoBkON+Nr3TZG4sA7OZJ7ZBPEJKFWk/MfARqOwrekDfsydheja2Ay
neYPgrBn4AMFMqxVv0ZwNw2Kz9dXFujq9fwbgpbysv4RYMOFc+FsgB7O5MyJbnHknQaa4dfTwEXn
06Il6S+c6mqWEDAc7tXqvTJYqEhY7oan7Yh2x/98RP109vwU9vqkZigmgfv5JH7LV4iqLDCmcmTD
zuA3BCVf99oxmk266hJAQbvawip2YJk7mB7HdA+KYd6tJSrLMFBwRbjjCXfESWvKM+AXjRZo7p7Y
/uAvZ88UuSlPSE72Lo84UdYGNm4jbjdZHuPrnHPrLmKTbp23OguI7PBEq2uSddi3J5ZmfA0iJjvD
QxAiIWQUyCFKbkQJp208bn9dR/gC0zddjsAIFKqLnaRQTLGOglGCRE7nPqKqU3sWZiXiw0hGYhCe
V6kHJCRmilmIZzkA6cJQ2Zf+sP0zGjZYDWDYigNkUqG+hySjAzCXES8qmUtgBEAkAc3AZEsSTlln
wkwJb2Ld7is+eHK9wxBjpr9z9SWle4RuH8vuEe53LNXoznCGmwLZjw70PJXjIAurQcS6bSAyKfRL
5kPl6KC630P+fbGUR67pz6Rdz7MLAzfIy4OlV+YZHdUSwJU3R7zJE1X0bwTxhBlreBSj5ruvY+ZX
PmS9tJW4W1Qw/l5wF5FP0238IINNij8oZJEH1G1A9QjeKGFon/Yytnj09hp0ivDUivfF96isUIHo
IHwmz/foBV0kzQTwlvpQ3uYXXJJDtCJBlU3B7ihN8l8Q/e56zjoS2GLFdvljUDOIFPfZIYFSzVZO
/ObSoudtCTTuYXa8EO22jm6FE3nzjNMTuRF+5hhe5uUk2OE8d7R1SIdt2dWorbWBpxZZjw3kMthg
eBuC6oCkDPk7cx3hbnwRnF7ipKvyBP18ttb+ObGZY4TWfoz+A1b1tzwGvyWh+QhzVmiLBXFm2Ab4
FrDs8Xq1Ipb7BjIhxUKkclK3XlwXApJcTOo1in/8+uYsJ2zkoXAPjBHjpL3aiT98POpL8gJj8haK
dYwYppyLvWKoQcYMPWJcUEIEbqDb7NmKiS3l7l04YCYk8SnZCIixCE8JjptZxzZvU5Pvd3P72OyQ
iZ9Zp6EnPILvbDUApTpwhYdTuw0l+oh/IZ4Vbc5tnPHpjKGqCmAyIkiB1w4SqaCXKBo4Xwd90Pyd
soB7cKCqsDexQQI+T5Kd94eles0N7NAyUSMQ0qDuoFgR5g++7qpalnJaEHL6AwQum65I07VK93mF
S5lH1IuZleucnpcWZ9KxhpuyQY5a1GGCCIFo5CCO1BGLix5QrdS2Chgt4szj1q1Smgcy55Q2Rxal
rcmGlOFlOUufvNNUelLpcCz1i5Nul0DjEulModmtEF4uL0Vs5jMrE13cE5KUeJ48uR2IqcszBQhu
vw633AYkiGqBd0B2KWw/W0R5320Y5Q5x+KR0lXuFfNCn4mPbLamA4C4bxufJ+CFFUeTxmjuYxazQ
1eicCZb48/SC5Eyi/4Qc1KdY5927y4BhsQ/gn2aMRmblbbOO6lYl5pbCZlcU1xkFC67o9tU/6Dcz
dV4Nawz+R9XrEZak4rsuAMGDp2hw3dDeUAUMHtAZ8a5FbDSfx2uIm5jOW2OBusnBiPjfGfyqcaC3
D+G50fcl6OIuujRMQ9kEO7a6n3T2L/HveKWbhOe/it+ADNpMb26b/HWSeb6k7b2F9FC6HLA0Oj0s
ZLuEZQLx+TZe5qMWnXWGZSGz1P3WA5+7ksF4vSQGUBU0lzH+U2IWsjWJQ5VdzLYMhiB3FKmd3eZ/
2I8ERYEieuN4DqUDW5W7LjnFmtSSHxEnKS2NaJ9N7Hx8WfGQWX0Lm6UXAsIX5aAr6cFOCERMjn8w
J2+STWnHj/EkXiF7TjEeqCGiUgiLSn2A14x7RW01aUk7SFbi2Ow+spsH+5sb+LeFGwdaRItHN4Ur
rDhCpLSvR3qPLqzGjtoYVyswTBtgXUVZwlfwka5HJTr2E3/5HpTACA0F3fsr+MuFhCDaxe5sooBu
1z8z0mpkovY4Boo1WRPBTceLalq8bMI//2agCAKSWjZYg11f5jalywX3ITvnw2eeBTQsNvbNNhbZ
UhyWNY/98ud9EEONAVEa4ObAcQKvpRmSZP79ofgj6m4snedLm+WlqfSX25T7PX7m2u+B89URNqr2
9XNc9zVISow756wAHxuiSh0J6gixXLpc3k6jk8lMy0WkvMw6K0UQgv0w6PBBc0de45VVaurx49Rz
NuABJGd9+Nvy+4IQbtgqVt/UZha+cxsUMgNr0f9LC8rYoHAjBdhd3w28m3lBh7xc8tMELV1nEuF5
C5B0pbd5goHyjh/2/j+rEyTZ5pv5LjfKzSXeF0bSj1P9AHsiS/+JScKbFwu5k2cFdVSqz1/n0t4T
D60RhD+JId4dxlKhSatYitQzgWIA701yszvOhP4QbPQ2z+FTTS+MuzB/y8Q5PZjnQtq9Snw7y8q9
wudfii46AQNYFKakLDQMUq/dQBI7ePCGOxBcUB0DZBMqrObvp87UDYiXYA7gIRH61S/3iRJsQQPT
sRFPygkKGlMiVq+qiByyDjoAmMs0qNE2Y3xxHzHvjU4rq/IctwS2X+2YSyOeZuA8i2X03eNnWvL2
Qwjj/8JvBkSN1swlh1QyGQKnx1eVfCM9xZsTB3RY72iPhFW59iHSc7x3a/EXYhVHcMQURww/HSyE
T0AiHBI9blYaSjPSdFiOjBtsTP+1Rr8LVVsoiAzhC8CYUmNiQLXF5pPbPxKOragik6AH9Bqt2bck
LqWqQtcElUlvBE573ffYmZEXeQGslnvb9MLE95GvLN1qLeLzUr2LCKS9nQte/8BCIaTrybukn6Ss
keByHAZwFPImkpQLlwrQzm7wZvsIc327VhGyW4IJ5Q/i1U7o6sZayrFB9Na7R1T1aFnM1xAwyeXJ
dSLHbgsuUF9MoeWe7UCqspHXp/NTSZzSFYx7y0xdtK9PVsH2zc27rQe3K50ozfqwfVxUsMKLlDme
v0Fh+OUn3re65VjLYovH5Nae0lISx+D79YGvNdMdtgaBi5hiWhYUE3ULbv8+/Zg+aPRzulR0Bh/d
9M4O0nFAtM2tDOJDUuxee+mxwfUiCuo4scFntys4CPLnUNzS2nmObeUj/y+g8eT5CU90+zvbSGSu
mRksip8OStjOfpvFEsLXEeCMB064RhQQoFxSAqAq8OSdGDFwW8KERi6lj584wqTLUCc7LmbGEJIy
MjlbY0C+eXJHNr/VJCmzA9ROZo/7eXBGsbW6CXu1z3xysViEKB7V5v7A+Xdi2ZUnUZay9MHqkuu2
uakM726v5vuvanu+BGBlN0IGVsUypNvlRk6jvBZQ67xfKWyGZ3yoExGQmVvbsL/Jk0yblXdJZAkC
X+N/D9ju9k8Hl2d3vCEkxNPB66Cj2YwGl3m8YA2mDBLl6YLRPL78qmodoHTi+ji9I8ugupxKOg4V
Q3J/sIHaPgx/wstljv14BUlpRNGoB5buWE+Zx/uN1IoIARSU5A3HJmK427WLg8T/xIvHXxjDBcIi
LY6r5NUNl2dHAMwoynJU3kkbjYbj8+IrYkdJXrSxxIU4ZRpTe9B+Tu3pieyUxGSR42fvg3dNacQQ
nMjg5FfuQtVzPy6O4JRGrkGYz9L0bRNaJ+iPrqSHx7JfgupiMLVwNLiSGMxJh6WlcL5R/qweLACP
TNNopa0hRqe2LSKPutS6QEjsbm9UBbmfG4VmW0lB1UcidjWvIY5ueJ4wANKOMloQtwtYseIMJI5O
btF0OO98hOvlU4xEFYvygbRs8srJQAd+WnsbdYZm9niwpf/hcr12rWFCNymeyvq+xgMwPNMXcRfI
b6JBy1Bo4Ch2fIz8b3/H7Qu95X3uJeTucxRLQTOmrxVfLOkM03Wyszd+4sX4/eB/ILlsEbP4g4iu
dziXZr58UfQlK6Q8K59TpqWXmrwSPX30XBctPl8m1/7yVH4etvyjU6GYVmgc4VlgtSMI3Sn8E0uO
pBXvlzm4Rm751TSH1yo8hfTHZIb1bT5opmOJ5+fNpJQDfL0t7M+Q8Rk2E8gs6nr9q4xP5A2POEye
OX11olC4rbb0CpWVaU1dGSw43W/aN86CGLkhv8Z8j8OtQg46qlAXsWNTkLAXvIzHyJsFmb6qFTN5
cqj/FqKwlAX0GGytppIitQ0h6+EgHEDF+spcg4NHQczGo6MJpFNECf31UjZNnXoVLMY0Blk/FQGp
83dOLgTkle195iQxGugwmnhCSYJZYueJnwg/6IPIt9SJCveoN/3u94EZ8/vK5j+9Jxi5zkXLGuHO
o81STT5b71YJtArZnyzysbxedjDRtwS466rHYZHcrkbY0w9dm78K3o8HldfJ9a7TXkYHvyjg78bm
vXcdWQVTWGVQcEQ5yzwPx6ba9vR1/e8KA+Lx38a2NZs7HZPjRTPTos49W/rgh3XaNJvzBZZZbGpF
t/a51uv63QlzIOuz9EC/ZHXyUBXUOaSHoYzkBvt+5+cn54TcaTZTQMAWIDKUiJ02xZ0Ag2Qr5dzz
GmZv/2T0h+uu0/FJEQbPjPVaeUMnX8g9x3JZep087SzwnVtAsPneacAAbmdoAqM5UF+pcLxR1m/G
AN4YOOylxCHzCUXC9t8EfkIEJSxmK/PDSJ2QZzIGeFm3ClqKgsyWIT6GgPdZG2iFkJqpxoiVhK6E
eBywpJ1mH/5kwrWCKd+JH9fozsDzixmJ4qOF1zX1jfH/E4MCq5K8QLy8isKb9Mvu87dfE11AfwTS
VawTA5QAIhcTiKzb5fTIjD/ELuzL90ccBnRHY6yyUR5tE6L6Td88+VJvikrCcOMQ5EhuhXfgjfIh
JIYLTdYQaJpdlI7Wf2iPjnYJwrIbUH+CzIQUaazEgjmirbPPmACvfvGg7a2elEJR63LMUd1au0+3
V01dysCSiMvpXIR8Qv9d/MRShoNYroKwp7jx6Bf0TUjjvGJ49sCOQoMDZRc0jhuq97869xyYVQcx
GHbNstyYbv28H+tYyEk7MUTY+NN0kk7Qa2h2NWTojuNXXAKvWjN2NZD2Fj7e80JaEax48LM0w1tD
g35UFhgndupIxbpB9TK8lQcw/s7L0Jr23r6Q/abrNK6Xu0emKsZN37Zt1FklTbGPOA9AVfHX98Pt
n9zRr9hjtaNFZrq7OC1lZOEYrLoO+1mohqL19zefTWFNRH+xijQuBaZwHWw5By6Jtyk6SWlpNl9F
Xlj9Eaysjkeu6D+g+IREDRbGcVmUEztCUJRYc7Wqqn83d0X//G+tCwu8zrv4+dHD21n26O5jHtDB
KVUwqTKq8YD87rJKJ6LlkniofM5NdxAVBp1JNgb3mjpJHblGUosrb6iw7oIZs423yEjwPaanCWc1
uRBI8wTi9fm5BRwqfQK10Cxz9TIbEDS0qIFs6A8ZY/DQKqeQZIZyFkYTcOq7i/8iBfzOn9KZAhgl
3cdCniANSiTzF+9nkBZRjajHJvAHOjkOIv20MEm6DLsPL2sZhTzWnK0eu5uD2yYxyC9KWd4/7v32
FvSAAY7vmxoFGv/d1EWtCnU7maoQw2E2A3Y3IKRsv/AQGA8GHvv2HDbZ7gbQEjxGciZJGLkkf0lD
kSGwY20hFHDlslh29hKpC9M2U7sA6zbTi7e+aCyZDnagv8VO4DnJWtO7tT7LjzybhFirdBpByiY3
qY+ykcYizs++rpeogfyVJzqfWs7tREEjvh9diqGt7bt51GDby6euqaqHnBAhfODMaR9bb2nchffT
TxbcOH470cGYdjx/71ShNJCD39KqorKLc8Chal+41YZkD6k/Im7gtp/RyWIGFz8k2kv8XJSlqekP
4jHuGdDAOU5cw0UygdmNF67T3WGa7YeexoANcKxvO1ZWOntVpaRZwC6iuMCS7TmIEoemSSLQTfms
AuhrRHPOlu3Q/Px4z0vwc+GNuMpbPcUsFn44gbRi9pffuGcGI2ZgjK93p0RcZIf/taSKiRTs5K3+
GSUCGw5uo+fyXXehZjW0DP+Dlj4eK8onpQ/qoV45hHuqO5pM88+YcwgZfSxtxVNGUdZZ0E33Cghf
XbcLiNuguCX+tkZK6mfmcj2WUnZOhA4zfTgjkq1NAdTQaXF1AUzEBJBw4hoSzZkS40hebwZQqXTI
027qKN1FvQvSLgh9SiLxJCoa9mRMO4lGo2pK9+I0DddnefizrJOegpZKZwLvMk1RdIYXtc/z0ZDU
6l3c8u/LB4aX+Itx8fhTPSVSkBkGQtQnvqBZXU452d1HevXjolUFfBauUrQl521G918KhbvHsYeh
1hi6oed0bhLOikh+xZWGMoAIHxjYVr9Pik6PE82T/1FNouA8TrZ1MON+mA2NIrC4P19PLSsa3WVn
bqGgCS12Nig3PtO7fFfK5QKRJ3ikRkMNhsct7OI6r+dzIpb0J4eAeDu4gQE9bDYjgRv56Yc7TVJD
6KSBfVfC/QpkwXOBkPV5KG7lPjPXRoGYF1sJVGjceQrqgIwjArqFbljxs1ILytSd9wdXcgS52Ycn
HYlEazWW5arJl1WnKjqds7KnCpmvsqUkg/Jan0B509N8ZUD32PNjSra5EiQyZ0crmTBHmYYcg+vV
0fesP8sQli0kYsBisiqJYKEhu8V3sYzMxMy6YyCXVIDy4Pqa2qs2rmM3SUjaruOwcP6nMdyAKGtw
chSrGqylWiAfVaew3PRT18t4cX6udoymW3eYLSPjUsd+cJipyu25qAJd4oaSKcy9JpjoE75DNfPo
GwRPUoTrJBeIylCENxFQE2S5Wjlas5IFaMIP2S3K3nuEQhm5+w9cKXieF5BgpHX8dyALlI3aDirK
XhxVNPGBFvLlUgKes4PIXqfIPXYDGrxvoIQWFvzFdflTvYwOsnp+gmdzqT/bB8BL9YlIP/uh7s4+
weQX0NJx/BRRmFIOVYr3rNUuuB4VAldiifLN1C0qY16ZYgWuAp5/OR25R6If5qRcin8Hsqi2t2Nq
kNSfbmumxoEDeJcKtcS3YXNybU1HJ35jkMYrHe7qJENXNZpuLBqhKTqqndQdhwKedw/zkgtTm1A2
g5ptPtgNHfDcQrWodgvqoVxOOFnSZszE0j59/QrxgjJmCOvG1JUDuOOcbGNwIXVdm7gJQZbd3fU3
OtTltkEt0hG1Oo2OUnt2Y5JRo/Dm+DxfUwfL+2bx30WMKgpZ/pEpPH/wG2x6ysXDmYnDZEnnLhCc
Hg3Onbbqdg/wL1SWVCKLXkG0uztvgflIv4N/n5P53zuC9SLUskdXY1cfW4LIi8taqF66MKb9T9hy
Q16PH0QemJjctNZwsAKBQHmRtIF+S5WPwMWMzrRcspbPfButGBAIZar0b0IrmpjFrOe816ikbyQn
ZYlFnLiy9O5alKA9AdezXLSIgOMQmdb9tTfRjTavfDjTB3XxglaZotlWtCqzEFfQ/atsOhFX2yJf
yfTXLsw85KZoBtxHcXsZmOmM9axScFzcZgOK0nQ9pSj57d7jgC+q3vCbCUQOJ35ddCAran9eqqia
neDP+Z4N/9ruavv4abVMNiKVx+OFS5cgq93Kgvac9VV5kyk8RCO6En6mLVibJrc6RWxNKosujzCj
q87aLJ0EcDiqN3vA3Z4l4S55bzH9ce/iMse2oEfVLASqJZPne+R2abyiE9JaS7ZowIXhTlJWSYoD
NAnskrTtQODfbB6dCCmk3TEj/o9adL/QFV6obUep2uShd5H/1lMWOR4gfktRKDB/ExTf0UaAC4KG
zMlLqOLQ+AlvkEdPPmR9Mm04+Kzf48qWJUb8StPavQB6rMMNq5GTD6Cs0tQiBcfMcNqFgcVNij1l
HWb6d/JwdghWoIYCA9V/rQXSg713aGW333laDPcgGTlFDWLynrurAU4D9XgpxgiE7EGVOKWjerI0
/aSSVbmsUWbJTstL/WRWMDbDE72zL/jLeK/tm1edLvxeJzXCGfhY3IhmAzgbYNJkdA7eWX3I5fx3
+K6Dw1toFEtchJ0jZbPg+zFhP/R7PI0O69ORC1u5LtmwjQ3CSdFzlCCKsyJDHHY2dP5nvdHjx3Do
meGUHtHqblgNYc+CaAT6Ue7pG3o3VeGb//m9akWxmQj2C5WKSKnfcYmkPKblGlupyD3YqJD5K9pH
V7WC+58hyhBJawNHHQJJMxhSsSbIMTbKhZ1/sVWlGqayUDTzGGkcjRDDeu5/3XEBaI777jlIMlfe
QxdsJ7g9uh8OnEe8ojLEUJ2hAS1Ye/vgCSekd904ICsZB1rWnlPS6zWyQGbip0bE4skV8Z9a2siv
n1S+ANP9NfHvh6kcE+lSEjFNzVf47I7NxqGylBtUXYAx9KS/lY73tCdU1t7BN/ssMey/EuGTP54A
KhtQWwj0qUd3KhGif14sG3Ev6c3eeqNlsiNuHv/TJAYvAPaNSmZjb+pso/oKG6o935iYLXJbquWq
JgKnTKFlIK6XVEl3fDx6+3LI6GPjvlosBjgmmmYqE0UMv5tSsW00nXHchh0ZSWbXVaxPPS06zgLr
Q18lfRodRNsnlVTbtfwuz9itWtPkoGcSWDcujsx/6R1BSEVXgAjr/JyC/ovp4ZLnL3DrJIgPZeYy
R2C5NEf6y6jKYnU+jHKDEucQ9YglMTRci+dAexoHPwxPGMV9fN6ntEVr5IaW9uiwzXo7E+boBYmP
/XYCEd3Fh2/W78HdoSgZU0NoobcW9nzQPueUmHg1rnFRcC8rf+q08xxR25WpIDbzPfL00GOa//M6
6SAk+VnJQlE5ZNsqlrh8MUC7HZ3WGE4bh2Iwqv9DYAD4iKdyhU/S34jfBnXiPY6X2EfURXEtcqXl
F3R/RQZWalDUcQ0aJ2LKEh7vw+m6xIbREHmU59sian+mLXOlpFlQEelbUoaES4yKJXj0byViDCqR
HmlzhXEf2RF+0GlrsMAD43Kfdo5++mG5OgXhq6CEFnGI7V7Wtd3XtYSCYIsb2SPng7lNacoUFkLP
Q1ClNYsn28vq63V+eAmA4VljCjV5CWKW+n+SRvn9SGCH+JvgWfCRM2DS2f6imMPvfMgFVDVnbJo+
i2TPaVqfaRE8UA6Xkz31LaNu7F4jNM8ccf0BGdIaXqbK61NBkTwRKjJQcYKUMdmzdMnHoFDDDIJu
Hm1o784g036LKGrAGX+rfcGQcqNZtJ5s0ipy3wTEE/0vUxiRnMtOgD8tcv2g45jaFbQosGYpmifw
JfVzTd4PuHPARRlcqYDBNuK0SRb4brR9PfRlkAMA0A0KHm/32b2P2Q+mmcdGerhQ7CcCnqcnI0kY
aPVPdDM7BHrot2uXExmw8V/3jB2W0OkxVVzXwkE2FIEwvcDEkns6M8l0Xvj80OL8TaGNj+xmFr+u
/Mqgp8H5+xE43M4BOKH+JJZq1fHFyenIbBDjYKLsMvD54/EE1qqqEuR7/eHb9xTNiMxPLkYjHRnf
YUx1Dod6/FNKYaWoLhM3iy9WI8Qu4x2a5BC4gqanMtPm+n2Y41gbVeI6PJT4AT+HGNHp7Kw/8FwD
nlw4axAe9RP+fpEAeLSfhYoX6FAkFFM2XCyIF8t5FMvLkuvTYFFFbhcSpFWADinq2e59snAFrs8n
dj7IyPCAK3qyfcg9PogPvB+kaNho/oAbcR6uAZrZmFXfFtq3G57KldtNtML5Na/ILYtGKSFjV7XC
X2Z6KUKnYnc7GMODaZ+u/1iq40d5nqt0rKnTEW3advMpxr5j8LxVw81+HMrmo8D/D/jRspz1Ogx+
v9jHeyUsNl4pR9tSelB/rUuYxlvo+JC48+zhKWWJ4m/Q/znr+SqvF3F07Lxz7BuFKri9Ajin81jE
adIZTDjTPbpX0BWh6WfYC8a1JAeyH7b7PvFLGHStvV14qqyp5arwgnAqrwuBQpvOP000zZ0NMsGC
MSa5/yeUwCEvd73wDtHDmDEcEm+IofgGdVlxSLYm/CB8iDYdBqTvE1Xzja7iOJnPJ0mWwz4gaDGT
8cZDKn6Qbmy+Nxx3+ujEYahKj6YlB6ELPMzeNHNQLtIHwJtQEVhlMhLX03OdtPF4VA/sm89x7uAN
B9F6ExhxGWDOmumvQ0221F0ouajrg7M8vdWNKMacJrBY4bL0xTIv08DP1u0oU4xIXEyupnOXdqE2
B1PgAMia09jY7Crj5Uv1iNBUuklcW8x4LzRh1jvjQ4RxBaQKW+wUiEU5tpVXG51puMfxDldW6ye5
U0U7RA3mpji1kZiFDBEd8S5sKvApRx9XM86qqe+dhklEzB6DpoJoWI9yJkn7hMmPO0sSdDuMyMcV
STAKKPyUJeI7vS6iNwA6QOCdgREeXUJcmcM7GqSrSMe6Y3yUOysueD86++Ctm2Yq7UyHuwbmqzeA
UzMKg8pSoegy1WYqJKGLzVJQZfPga/iDOW/ofcNbQ/xgz/CaU5vCQM4CUJ79/G2B0enLoM8b6GMJ
SqLEL5UxDh3wio/cWEGHGGtM+4QbjuJ53p0zUWkc3sML18DoCPns4tacwnofqwCG5NFsFGmQ55Kq
CEz8ut6/vyK3tItpX5pCtdQrdt6Ef3Tu9CJpKVU+KFJYGt5+F9jXGYBXnVnRSzfZDjlMFCtrkHzk
T2C8MQlJpe3dWKSbbGxZbebisvL/1mhvWUyqdfbRVCzrQUvbayLledDzJK8DR205NK/L5ObGpHU1
dUjQP5svj0i8UDnJBEDSU1Z0oLylEZYv4bhSGivqNWx8IZTQqusORcjtDsmR4o+BOvAZE3ELvzjX
jzr0tKcSD4aNmjEqm+38qp4sEoK3NfWdijUursFZQsSc9cPMOtEsM4EmqHi3tj7uZ94pKS4/JGFh
7eOpwvsR6YpSQttxNGFV9Anqkxcc9qdumUmRpSjvlVpF+JiqOFwlm+irC12t/R4w/k+Z9CvdEULR
bWmNunHXxe4Tapm2FKEGdfs+qXJ03Ar9/vX3x5REkJyA5zfqYG2RB+gwxPSV3xURjJtlWA+xpqiQ
YRWmKU9VC+s++/bKMrdVgyAGDeaq9W/3DNXe4O4P/ahIhY5SY56IDpB3+66KrDyp+NjHAZG9mjlQ
Omr+4MJ6JasPyhyhZGXxN/b4EWc9EE2TBLPkqC8dGj72JDLonmyHYoddyZWwfX8imRSeOQkvV098
jITehcrbvJBwzMN4Ru8YKaurDOYDxbfxEpP5Bc8HZ1IEgEI5m/jUPPXY/PWj4u5fgUVLpueRAuyu
+M9mhp0iBGvctkhsCyraUQxJlz0kZFY+00e0zlyB83HcBf/3mPWr5e7NL/mMSwg75wds1JL7g1v6
Kii7GrRPZM9VB3b/yDyWjuUoZYKU5v4nDLzzFTvJ0HotkoX67tLWUplF1dN9WUTrPMlRndYpjOkZ
lkx2NbQhC4ea8//vQ4wO5rRiQDEHLyNkIPmcz/0NvZl8ao9UNiEHzVvbReo/QIZg7e08TCY4/T5O
ywQuXEdN2N8OHQO5hzKF1qK7kkFQuxOkLqt6GcGoHRQOW8sdFrGq33m8Z7eEjdal1Ibp9ZqWxp0r
LjhHoKbSxKaorHfcvGcWwWhJhuP8OKJc0SvLQ74waOHtBJO50xxyQxfahu6zhyws/Mc6nRv6Kpc/
kAznKSRN9QiVf4SiVbIPYL0V6wSjlskCHt5qRcx2YikV/Ahn8I4S6Zdqvk9GZt507vq6zooCJeLb
+wjoy/TK+RBP/LQznaq2VzYL5WYx3XMSp9ezvhvjloZ99x1G8sz3Si2mhdWs60lEtjcLMkNXtzlZ
AkDmD0OsG7XPRTBWEUt0GcrgS62UIbeBULOjEuRHJfw7sV15w9zwrrnuEcGpx8jIqmWp/Rrpw26H
b2phkePfnBIQNzOotEkVK4vp6nIT4HVacBMyEE/dc0OavOkOP5VotBGJcbYgnEM0Rm7+0kWa8gdh
y15gJK0e+5QKpIEzjRxcyX1u3eaNFUMAY3tW1922xFURYMag3/MvduCPWVPKp6DwKmskfa5VhPgT
oQ6491pstkjdZ0Wb0og/ygPhG4HWH2jxjqkNrVL/g57QM2W/u1baK5q8uK/g7CWNLBdVwEbm7nBQ
Tv+9XX0YVQj2PF89t+4adYnJc51s35MkGksiVA9HzcuPnkFpV2z32ZEde+LswFbslFjtacgVu6iL
97rlONPwUvuYQbxw/x1OjnP+P9bXWx4CBcLy+Qq1PRB+6aLiQfCkeA/3MgJ3WsGWDSvPb+P6t5xo
qTsk6HDmrFIEiCGtQ+nD18B5NJbUMrUR6cO1Kam66k4lsoeXfElSjblDgyDx3cxFe7sD9rInRiRt
zO9by+t1NQBbeh0hJ5C8oY39Bv4G25c9YQn4q3DWboHemJRnm+5KsRA+ehlJrbEQhLF8ThjS6azA
7yFgTHPiqcBGoV6+TjkJnF8X7+rBn0CkInfr5eHnZ7HdoTTVZ4Wt35mrZdOjXbZ0CqdGH0Cfxw3+
uiaY5c+kt2Uhzwp1h1rAhRMUqWToeyKdR1PsUPnnYWFugBszDBma5O2U+lBAIfpsITfkyl2M9v/u
2yZMV8TKDsX5bDFbb+sBtBYsM8herSBeyLnbmEja2Acg8/u7pAWOrVRc3Ma+FqZsPmbgaQJ1OT+2
1OouD3vKBI4SIY44QuI062KhBBy5Qti8XOWY3kWWxRocgBDxF67d9HZ+CRS1pReIHIFTI32F0V0y
+Nx1/os2E29YzrwHRIkjvuHZEBWjL8TYAdJLZC7rhrLnlBredh93+myQmgXS29QvefOHHqqAltql
DmgdxE3CKnc04N6h3GDw1Q4lSWhfC6D16aspvB/QvRmSCCRz7KQGBwvUSC/E6wKHiKEX2C/rWdd4
6yfbA1r9t1pKFXdGLKrBybhR9zLcrSI4KQo/929TWWe2XAB/t7iHphKFYkBZklALPVbRu5J0yu6e
jo5lwJJ3IIpdIez8s7At6YUMaAS1FMhxJXoqOrrCE1ZDJW6XXnv1g6JwqXuMUYtbHXI1Fh/kgq+0
2F0f4jT/sIU/Zej93Sgw0ajCrI80U0fVJ5ZH1n2+DBZ0tW+NUECFdBIjuex2qPiJIQzPJCKmFld4
MY0EhkihpeDEP8ayqaTNota8m5KLga7BvvPDf3HeW60nP5y3GLlbfMEg072g+ySLx0X5Z3GzTO3i
0dHFO8FZ44YWYFvYecdF9fMLvmRWmBNhBhG069Gdfp8TX/KKnPBiXiBdI+IRPJFwZ4tt5BBg66Va
iRW22Nq8pvOzDcUVXEpUYw4w2LwkBgubnF2XMOw+//XFZyZnV4w3S4bOryVKGdarfx0rdmyU5cMV
X86Owa4yEZDrXi/KZrRSWp8QHWVBvi0PQQoEw/3TZVoNAapFQjjldLNjtLsFtiVir3VeZAzbMaIk
eSaC0SWe941hAgEiJeToiPbl2Sk5Apkn08m3LstZvQe1P79kxXffTuNyDdlu5QLb4Nc3vNVe0yUs
lN5T4HxL+PcqW/x1Z79EdcCY4govpKEQGAr2Lo/loX9xP1O7h5HJAxr0DVHst3FkM9UEKrFEOoUT
HLT8RF3/ywqC68gE8X48ShxozGkZHeZY7mrSkF8UcsBu3jmJ5+/rRMMzE8qeakBzCmMAyv0BHGwu
bsaREjPOkNKJcP7GNG40Khs92WjZvvNHYvkWKY3qk768ke+9dtISxi6AlDJwG/LBVN4TsuixpWZ+
qyim9N5p40HutBBIQrr0VXYIk9aWOmw76uxjCHl/zgIdhnPaqen9rgqhnBnGrXP6ON+KoeMddJRr
CKmb42wNRCJmgLvm4TUI+Je7PGAjj0t2jkWmk+4XCaFxvtrrhZMXLqpBJUddYi32iVi58b9RtAcX
7jrvNSJ4eTguiB2RWO6yoPzJ5pOLhl2uAWDEHs3WHkNYN0jtP98L0tj0jyJ91kvT4Yh0ViN1UdCj
5wAiV4AWBwcvUt0d+l8po3QcE0Ioe1GJqZty0qTvBkf3jDdYLCVPt19KMFiM4os3grWrBoeRkkwC
A/PGfahOUmV3WpBjZMWnqYPzJze8ELvXX7BUGQetQGiGy4+LyLTPfZLUsA3tz1/R6F9tBZmSTq6D
lpDidbmvd/aMhIMUnZvHi6KhBKq8xZ9AHTqhdjTP2mak8aIiz9NvvHYUJFUoMOoJaoFUub0DSJnW
1KahWrgYTZn2YJ/SwtPfEvTjDHtyQ0t3gI04RgmhaX+JNJuHV2vwBbsSjYFNwcBJWxZuMbRTlmAf
Xkfdr3lSSVKqdq9KzbBaaTRKTpCSWha/PmIlYiJOv6oGPsGCrfyisL0KQKHQWEuS0/NNGfq3JZ0L
Sc6e9dh0tSSDR1cm3p4NycB6lRGZPW69nWI8noi8DF0kUfriPoT04GCbmVd1RIcod5H/hfaYcsFu
ejDpm5cgonKCR2p+lXMYxGTSOgp9ezKphTd8NzoxQJir5zzINvLRjQG9GU8tYUkw0nNtGaH4InR/
qjLseILvnzosC2vh/O3VYcThOUjk6UFb79Eac7l4SshOwGszlh5aDLtnWM3M4Sn8//zxTRVKrWTK
gOunjeGvI9X2FAidvDD4ZXACcYDFzBA1LjR+/t0dRE6QgQ9ZBFCj7U/5eXJ88TXFn+f6RJyf/dNF
JWy+uQ0Un1LWgGktgWMaeV6uLGKlCeuDWClRgo3XdKoJkPpv3V4lILuuPE9Hog6sCV+PwCzIFIxR
0YtOZBm2p9QiW4lAtox5vAs1Om0xDHHA4MGk/OsZJbhTsp0wZ6u1z6W8npQoXedV+cLn9HnIqCaH
JPaai8cZr41FoM3GR3hRtTHYqSVQW1jMzg39/y5yKTZEyY+QOFo9VWDVui+p1zf3VK0EabAdv7qZ
0HBLPipnCV8McF0eJvFOWvjQ/otq5PPPe5s8Tub2ILNe2gr5jUcG9SevNDnCAZTRujlOlw6u+/b8
Gca5VrMXNbCpHMe1Zc1o8SGgUx17dClInRaQh+dODtWSc6Kg/dSRmG5Aq0IAB6yiHuo+BOK9bYH9
CEJk25IAbXPOVPyZMklmsNzIYBlkfqKUBc6WFZdpNuh2P6V6hsPVk8IDLz0PREjUbyPVKGXWnBrl
7NIjHzxSJgwptR9b1gx6wVPKGZhUxnldojvi+ojpvAQod3Dra5TCkBanDjtZOmEXpyg1BfguHcOv
8IUT1ZS1hLWdUpq/D5rvtGMLyAstnb2CIhl66BH5xSD/iVV9xK8f4dRuUPdlHY84kcm0ItaIeYSK
meaySkcWuv668d1F1YsQbfvCIM/H9TVqLDTaFFrQV/eMwjsNmsYIT6ALH6mrHrndPacp24leFTj/
V9EXV0WjcQ29843edHJOIczgIbfy8hH6RTItb14TmEGdARGv5JhjzhRye5YSZjDBn7QPKo3+TqBG
Vfc7/W9b/+ekeNpjDO/ozoKYzm0DK6B0QaLFsIQFXAbxaXSid3641nNNMlswip8fCf2M+XODSLnl
ZSEsSORx5ajVf/7RNn3GFZMRAYyxuBIREekjs+JFKQS7HVhk0ZyKBBKo6QhshKOoNWIN8c5scPyX
VPjbCm9TKURofZmSKcMaD+rCs0g435Cj+pwiZIEHaMsWhcNOEhwMTPncdisQCKTMLPwFyAgXLHP5
YWvyk/pv+2Gn0mwqmDTaTkXRlWQc8FGoMrcZmY5+zKs6NLt1QdhonubQVAO/QwGe7SfkYeE572qh
icBaHMMOoXj9/rhYDTFprc30XIa7uS2PZTBXEpLdY9Jv4Znooh4ir+PBMDhg+dyVcmhIBauWRqEk
qG7W9etEiTMunYrNXx7l6lVM3ce8ysAg1qXpUNTJNGG3kyJF3BCZYZgyZwf3TgkOVsxRRB2jXBxU
tEv+5oqiIXjuVRJIZlElIlb9AdXlnk3MI5iqeBX15XOSIYZULo0VG6EzkbGoTWgAvpTJNjODSvZT
8rcPLDscMOiVok09NR7PK72NHO3vX46Se9aTY/1OVXTAC5di8YjG1ar9SThPb5JypSxFSqgD7BQN
RF6ugFRdN+Qg8t+Y5Y4RMwymY5U0r/0GvToCb9+wFhlFAzHMJF0h/2ta7tygIPkCyUvw6e4ADe04
TZ+CMZnPFcvMcjf1hpyfCRpjeSa0Z58BM0eiuONjlG36G0rJyR9N7l7699mD8gh1+6DMFVvWhsXE
ntG8EQ44eExNBp7SL7oIpAwICkP0e7QVQmcN3tigeCR4ztQFBYoTFao/WmGRhXwdZawZA00UFxVZ
wl4fhIimS9qsNOu9Ocf2SHpVAeDbS0kUZtwxVbor8mOD26S0zBGcV5beWB1KjxKf5h0RLBM45SVQ
VmaefUtlzu6p1Z0U7mE8waCenpAjsOURFSCDF8tndWGVtBVXibh4iEUT6GoU67zQjOhHl6Dg9lrk
92zhGoyNgvOvA8UHzTjJPr0NgPXhewoz06WNaq7E4rjwWdkcdA4Q2m6QDGS2GA3DE0/M/+uXwORV
nPVsKUKzOxQ7AvMX/Kg40D4gRs4T6gknpfHsZ1wGSdGlFIZMoJR91yN+LAkK6RHEZQwi5b+JWZKN
G6OrAr/m0+yg04Aiw+Mr2cBb0z59BMCwLjOLUIb8c28WqC7XYAoxTwyx2Lc1cboYxJsjQnYLV498
+k37O43B6Tqjk/kcM6Kofp8C0r9x5N3k1VNC9bk3oHVrXa1ntKXXBMdsxo4FUSM7oa50ENpAOWRO
N3hVlhxCyymg+uwoz2BpUeeJ8evwjSyE6bpxzn2GRo9XMiqn5WgqOnaAnG+WVJQiywlUIU0vMpO2
DuKQgVTbNibHAJnl+FYYUL/x/GevyTjiEN6I6/KD1RiSaQNYHZGwlNqUhp2wPS0fHRcmi4UQ1T/t
poicavNlrzjU/sueSMMFPJIeRexDi3k3lQWcBe3UIsRuhN8daJE9lVGJn1BzHmyvRMHEk84QDOzI
xtQbG4UVRgG/pVDfGf2+rkpzmsuiIAUPkAeSLRJwLWspIz2gWbnGpZ/mIIv2wTsw8OR/tXMScVUu
SN4jGwI5qnYrzqhIARlJQaWWIsJKc4pj7jL4hpHQHImdBS9Qb+1JAD/qfHQ9k1E34zH/1KXoCXcz
DCVoyHu7N4VN0e282odbMFUjsYGo/hlkDtpz/PIrg9P8WpIImLAUtOx796t8RCxUTVhI8nepYMVO
smU6qT3Jv4nBA2IFEcIbCJloS4+Uo+X4RS94VOUfvY6FSItLyyjzJo83NbiI65zkHBKef+g9WUJY
jhqyP0UY+M4lmvC8S4l4Tj31KcE+4wPB+ZjmtItmeAqyxnu2zYN4/iT2DJ8Dd6mlZWeQk3FuPWPN
pLEdQ5opGCoPEQ+Qih2YZsbo62rNhzX5ctCyP47vV6T4JGicDq1cLP8AJ1Mg9PImsA9oNNre2hzh
LE1jquSftxHUwwz8Oi+Vt/K7UinE0fe8VF94U6BbUyGKtKuA/au7l84LL38Ma4GyJqb49rMFws7x
EyZ1lWvhsowGi4GWEIgzU0SDls9fKeTvbQo59l+uVJwNebsaVsKCwzfnWvpWrHwkQvmi70ixxK4l
VGGUzJGNvYbDHrdsnVUrjkVV9tDtM+bzYK4XDcJjTyGVP1HZdqIwdvqwV+q1FsH+5YQtGZuKNzA1
4q451VHuOSl8O2YNBAbmxn5FVlZRzsj2Zh0mQk77lyTr+n8TBoRZnY7PfpCTu6WNUbRXlMCTdBRc
nIo5HELc6/8vOB62OYDkpI7owwaoFHleHgbkDaH72E0DXDOxl/EQ3Wn4gc7LJ2IVDgXRxOMElIsM
Xw8mU1R8LqWv+D8nuSbDvy7dZRgAVBE/U6mRphdCSdA40hr4uzmbnVTeA8UuiPyUat/ie2TmRpFM
BUXmKnDQKzSPVasmsUU1xEVYZiyukesdXmBgAP5+8XoNcls8P+JkbqAz9mfjdKDB4r3Fka+DU9Lc
MBoa9g77ET9dX/VJoYmLCn7iXhOUKqUrN/VZiKkyGiR9f/ldwFeUX9+iDngcRBrjTZQKDHn9Z4GF
tTc4EAVM8VDew92rQGV+Q2vZPLbpilI9cTcfMsEHdNIi00j66HyvpKYKclr3z4vVaqACZzEDpAtM
G43+hPywK3CHwgaBfkEQ/NWXSB0SrjdSpo8nrw4ubivv9DU0wvbSVZbrj7/8FUURM4rdOQflJFpw
wBKe57ETohAHf3UIfCy5ahzdyh3RmI1NOmap805xnuy5+2s7Ur7bkbM/0CALD0zDKyAqsO/4qrTn
pSuAcBfZSX9NIbRn610cY066hszVsMk5U9PscH2V81sGHdsijPoMKOPY7gM4qFP0CDIsppznLTsX
FNOzPCbEocr0BFSitzkdDjE1OAWps4MXF+kXN+Kc/gCIt6HxKZSACqnI9u73HbAkdoyRk5YXsiU9
uSROKFaUfviDw2v5HGOc6Bya9VyGqHrsJ9CBbDcKykL5NunGID1nHxzVdHvA1G2B/eEipEcd6a2o
eCnl+F7/NYKRVvzbtY/SPtPyutxFBZ2XO8s1lYmAvtY8h2d5l1tz9UEzcN6glpd9wow4rGwzUPX6
2QxSEl+Ll+9tI6eXRKGQf06J/0/2asUuMxfSf3DxxuzKIXhM54+Qpu6TxuZxDeZ1WxC/XUcjbC0r
88bRvKQfTg71ZxyMBMbcB5pbWoYC8GeJzlN//Oc53ZoHyS41qg9rJV7DVcHdCI21CyJItZTv/mYA
jcu7E3s9vcALL1h6z9EFWLrW504yMMPPuJAuIGFTXI4FDwhAjznJHLjSX7Ew9qgvem6MqHdl6S0/
1HhhKTVqm8pF4Z5I5aQV1cN17toxzIlU9IXf8GNkzbDKkzf+Y7A9x26SrHVGgUMI5CvHUuULX4u4
ZGPNZ77Iv9sX3aDoF6kjuE3PuJyzcNsD1B5uKQa0G6ir677SkCIg96LzoN5Kt1JD86joqsRPL6d8
ss4nNt84m7i9KyvVKDIvWaRPm24Y4Ijxz9pTBHifHYxwO6mdDLJ12Xit+JoxJHD+2m7HxB+OytSP
nNCwRnwyycrN5LbARPtYLVzZffNsba9eYZfbhGxHBxdyeuTFCTNtvQDuIv9YFkM2AmFZRQdXsmG6
VXNAf40G7V0ZcTp5MXkYbILXmOLAYSSLMbGoQAbl11ad1oxe6GI57Ey4QCvcB0pKmVZXcLv+QPYG
APVoYvlg9BrMHvd/Xt+Gi6hEcYiq5hTJUa1sMiZ/EtRNvIkKrdIxnsJxFXHq8sBxmmG6Qo8g44Zs
oDig2SlrkwDTMw/9txMxQy4tyWgTVPI3k7/WaheaRrS1BEkEEQGT6m8FYvdM9nHGhMy1IrjIbfXA
dRxbGF8UHI92pd23k11b3DUvi45FhMwiNT3tHj9Q3JxEztufFg0Uw3PSqKlGjalnCI3Erih8HjNV
IYzFkc2kx+CReoEJX30PmyBY9MQU/gyTKywI0trtQsnxuNYpbs/7CTaabOvgJK2WNTJYkX3fd6C4
1VxzJuEl6cYIx3GEQC4HRKXYOXlSlBam1CVJPYk2sC2pKOsDAZqj0rlJK0dNV0GREaX7+JjcY0KB
M8TEy0JlEoLHhOATzliCe4bt4Ike8fBG6kRY8mopa37HZ5YGi0xmES+YFR39SBfcZGdFTuZZ2BFE
/hTsJ2TUChuSZPadZyvAF+UUEcBVxw+jJ+ihlJLoaisgISgCcD8HNa0ccfUbdq06EMow0lhFtQm6
FYwbPiL56RuX2CvCKUY7qFXRn8M9f6X2zaCrZVjmSpACBfEROs2MmjOeTno7rvhw4MHYIBp207j4
s+WSVNAw1xGKkKH07v7QYKJqfAEglFW3ZVgYGMqcQcXoO/GZ51bxU8LSMOFR8DzA/2VC95LDEpUd
x/3wVfNx4l2at+jm0V3gybZoEJ+BlTu9IW21fwWE5z6qO3Vyjyw2oGCLWA2XGFzDrqdW7/vMoiP2
I/7oXCAllW0AmHwnxBMNFIu3bGjDMKsLeITD6a+hom3BnWzuWxp+1LF1tMbws/UlGtBNQ9bAF7mC
485jxfMy34tAmDNh6ISaGSHp1dW9qnZ6Zaua8Chhi5nXZU6nlGKAVEhFO4H1WnOqNRL2gSF7St2W
RSi5WHG0nUVJyVwx0IY3VO3zGnNN2I/7VjUbm/dula5Jhf06tXhLiNj3G52K0JesEQlLE8K2+UUQ
Mj0W5piRyj5gpcxZcOQOLd/h22mtdTWxikMt4LPUrM7ZM7HJ6XU6sLk6QxhpIpV4iz6Cdvk7Us84
SPRVK7Tvk0dKIzOmXb/p2GFBVNgZtwi+3pCccxcyMhdLIvjRnqTpNtt8lLgJi3XH9yc7fYVJRBC/
8+XqMOzV+Ur9GP0+gPN5e99wSNf6MkT7WnGyqnZ5i0KwJE22RqOOu6Du9jisON6Gnigs8Ku5PXoM
MDiseDhzbHR8J9/kLp9Jeo9T51InD+PI1HwoMkb5ZsA3Sfnu4TxrXTlvD94HcJsGQeI8EVAEOMBD
IItdnFsvbKM31kaE0Nwh+2XT0NRW8TfF+Y95GWi2yAj1FvOQXsQJCJoNQ23rhxRp0IHFdmPBpB4I
vMR7Zb+YRG0NLzhfyPBKkqQg+fyWWikwROsSTuAkMpnFsaK1Xn2eSN3y8yszNyqqS4m2QmYgQVii
GlJqXBocaDrWfwG+nQ2DoiORm3Zza+ff3IuAruhaTFM2DGw6l6C9vBaZl8g30+Tj6Hv9rNheYsxV
RnTKNTvXB+s7Faa02D7nsjI+loclgoctrF+gg9hWiLxDD/AvQfiVUZpC1VdDGUH7aeonQHAHpykg
d/JBNXAf10P9w8gqmxMXAK6xGbmhLIKSEsYnVMTaqU0R2k0mK29joiC2FknDJtb4JdhqjaNbzc/M
bOTObfJbsJan986923hO+gp80h3T9GqGpZkXixlHbHpdj6NZAtBzl74yNWcZ4jkjip372RkJhs79
6HPD5gMWR1QUx2rp7d2H3OCLR984i7jRJQyfQXTdITXfcJDRZ03ZNG1LgfHae6Uc86/8TTTe/ncP
OCzVqFlK2RjZ78BQao3a3canhL5fmIaobbTrL8PQ/AJx4zvxXLTG8f+3q76xH0rhClWDnSZM8uIx
ZJarJwRQiKmwmJDsPMPuTvGHGUxM6IpsQTDKpVnpdsgT/eS9mN8ei3FMj8/ARa3xyO//TcHgJgWt
On/XvUYEK2RswxL4nmavgmO1iQrpSsmnXXf3H+vO7+xf90uKx+8ePsujMY1TWVzmx+mPuAZ8qj0h
8z7IF8KFt4G9nixetqapOGp1fhwAD4zMMFeGHcsWu0GMdTpRhYU60nTKMOMmf2sD5eeTg7Sk7b5w
nJEw8TO+wZnuF8c9Wk0pKuWsRU3sftQsF10aGH9Hve7LBS/fwrjgO+j4sz6KPwK5nxtG6YzrnAr6
6Hw12qkw3gXh8bJNX4Er8tuXhQ/9Vj3PiF8uZDwxPNrWIfEA04Ni27tX/0f8l3MhbYKGq+BSeCBo
L2AdPaJJp4MRahOnErOfaLQ+nuuqhjXHdwN/l9xoPWYFrVm+L9v/eLkdyGiB+kJdyAera/6UCI0/
i379Uk+Lg6eOTGnktlWqMsKZu06+/wzxxJyTQJaikVEPNwro2UtOSFHsTyLJF4PDBB1AGO3h5o1I
/UWdoKolLECFwvIrXF2fnppAZ21mghbl9pKwXGu7ZXGglkqLhWGS7bKq902kdKrFT+azxdMPLnyK
EANFZUNVETxpKPZQ+30bxs53oSkBVKvtPrkBkhcT0+bZ6qZ6tsuVcQ2EChT8nuXHiv/LpCVkZVtA
bs55P5tIjmA1Q48RRKw1XjViaW+XZEeRUxsxp8fNIzDx5jwepNgBFox4muUUfRwgOkC2SwGQ2OsC
zvQdgBh8/V8LMZ6K/6xn+MMaexVQoQKslPCQSvo1AtklX0miwbhn144mNdMnsJmu155xlGozl8lp
ekm8CZd8u6Qbmyu4dQ6Ull9UrDJ5QbmnK2gisOHuDvlr3ZRXLqs00bUoFtfI/CW/p4ETHvxRU5m1
QXQWGX9uhDfLFGJan9McMhdHSKjT/NFV4zJCrLqpAA2b+dDkNP16R9XVR2upImhZK5iv/PrvM4MD
4RbID3GKi2xOHVg+TawbUXwkIOfcDWHuvQGKYB4lrP+iM1Z/CjFSkR8XNRZ6Rxb1F2obZ+F2/0s4
87X5TvNXlq7ZN3UUTjjGt2TjliOm6yvsJis9k1znobmuzQME9jTvtXJIUANGjBG4nZViVR2erjmo
kPtQH0dJZ+8tKE47c4Qbe3xFIeFDTNWw/jo59OY5uOuQQwEB4s9hmbpmGqTua9SoEYtt76sglOGZ
2kqoO/C+ZShyNkfnGWRbXv8Sn1e3c/TRUBSaLo9cefPpdfH+TgwtazpZlz+2tbr2rhCwVle8cNGr
+ZC06a/KLAMCSWzZmd0q8+CmZtc1AbmT04KOpAWoA3zWdj06teutU/fjDTVX1snDrOnJu2rZgqS4
ZY8mnUbSUxPHEdOsRPilFZTuiXmg2p0dneFyZ7702mLRvvU7IUz60P0HEugvkw357XqjBrfCghak
gjstpDYHN6sLuQyM93TJwTIEmnAyRympz7Y8LWkWlr/Oa23hC90VUzbIEa2K33/rNnccQKyI+6Lv
5NPYz0gIn3qM361pkcQjROMMVxsyR7CrwIPuKMLawfcuFFnR+OVfcNDfPbCSdpaFRefrVYafqIkU
PEMtrTBktcsVbA/eZcLUtDTCSpy4n8U0aPHakI5lla2e8fw5OcgDQ2YJhUFV5uqKJ0q8V4bNRnvB
SwdxVALbsJDRjh6Yuo5FvOogMfJp64qz21XcZtW3qyORFD8mkACN2IizV2LgQZBCtM0vzlMHXU82
nn7JK+dCfxnINJVPdKAt+aR8ZSGIgLpeOSX/S84z4f7POsrNa3VzdUbrRM9GTQ+yW58swgtnzLt7
owdek7YLCRyTOM7/vb/4PgU7P4VfIuXvuir5NcEQqVClc98FlYBCuNmKFS44cskbLFzbZG0F03TN
Ct+eVlhyL8UgZOBQPdt1A1VCtjWujgjMJ+U1YSwxs9XOdEH4bJuycdjW26mCeJOzzgiKN7aWLsMC
kY4O4ryfk5UgWSRQbSLw3xBYXIeOvG/dUL2jz1yDT3XYjwWAgXhVw176WnGhdr7mrwi45/F1tPF9
oZzLRiSsIYhWuNkgcokJEVgitgusNsv8+FawEVOjIgjgxMiREWJX6S1tKqOT3Qjje11amMc0MBx/
U5/hi6mROv1lPSUP2LhfgxllKcRFeEMAFlP2EcTHMgsQks7TwVMYlVwa5SkV0Zas1yUGqeS6kqFB
bymv6kr+NMy8O5uZXHyQDBjWGuFrXWE12Y8epKR2UeMcuX5F0lw5DQIvElkQj7vz6AgKqPt4PysQ
VQb4TXY0en0HnUhBtGKq0iXBt5F7AiXF0Ob3SkeAI2m4tMh34OrbhjuRF6t59DoMUc3uVkAjrfWH
az9Y86b0GsXOLxmEwUt20m6vnQIlnvatYg7NiDnGn7qDKLcdE0Pe1CVJNNtNs5kdLNHR0w1jbVN5
Y5CBQPIz92GgzCkpZf8aZOVSmS6IHoDwkSUpfQHFJxzRUc3A8zxi7jQ2+elVH5pO4z+LomhIZcHv
N27EkaveBFY6YmymlGyT6aISPo7LSp7xQKS3v7a+Mbh0KUc/89bjT0wU6TBOeXHfKDsCsoqzpAhT
CeM8WRDC2TqW2iRZvUNSixiM9/dVhtUrgkNuIODrPpK6yLx/rOBUH4eDEceINB8URf5V2E3la+ck
VCCj4e+s9KsB+w2PQF2TcwuLHJQ0Lo2Fsd1Cds6hDnmqJtdFV2a784M2rFMXeWqLA4OW50o5zgLP
VKCyPemBzV2/xHKRn7nQSyLS4hgNoa/rYO0SeFAI/9AFY3Ol7y6954ct+FezF/hI6ZPI2B6ZFAS2
TOapbxUh4juKRlbI+7ApOBagh9XaDAYzZwPS1eiuUTda8PxBFd+MqX4A4V2fbfEauYsCn7e0s3hc
ra0YPDOIovJZWX9zoO/CRW+em5npIvzrdCGiDfJhYs/bc3LlzTqAysUxBRizz0IyUg7HlfpKKjLg
+ZxJ1p5GcNYxy7/YrFzEt8jSD3Ext23JJp/y6v3hfDl2J+M2X+Kth2TM+tkEORw1U1N+eq5dIjn4
aL7DAYLlXSv1YBzzYWIPN/WMvwh/8BSzTQ+8TKVeLa0qh5iNCT2WdpsQfPnpK8kiDTdx7oaXMIUS
tgLHX5MojTd6mNqSIEsQfLKD7uRMzim699WIcuXxzCHBTcTJO54w4nDhz7gb8GL83N73yP+G7JwB
5jtA718sdjvQTk0gCyMNIrISjHE4GU+TIJ7L06muZQcIFCKs1O3Nfot4/1uQV6gr+Gn6XMEg2lSw
twieTllumS2ygYbAc/X5tXfDbLNnOOKCl0hl7y9EmwxftWtZ7rrtRJACTbaj8IzXBDqWYjSEBSwR
YsouvpRRwpeLBCnL3eWW25a5WIvqGGX+huJsrwOnuPihkQ2cxlj3RxQhh29tQQkACEkIE+WngMlX
eDqD/KFVVm4D5dN3IsUki6kQ9CP+yj//Hle2UEvv+0woBBCVRj4sRrHeFiPBrP/oj+4xj4yZN3Q6
vXYGJYJnO0ThAOFeTzQ3/Y2uggq5LiXBVy9JpKzznQSIrPcIXDPx9aGQjs6t1zvo/I7xLHlqGsJE
m2vgKeeAH8t5ukPGBgvc0eHJ/rvDt4Qc9EIGvtKKKwoth3rUjbjvW0I7E051BYQm6bFugFxxII8F
9H7AbjF7ZjZbgJljtaV2SIA3q9UxYinw14LfRUyFxjCzrBMHa7lc1QDtIM2B87LxgAd8pAxjNgfi
hP5EF33fMdOdAul1mdcbBPCN5cjMeCVGg5ZL9x9z25bfXDfhbm4uryBLgD9Uem/LPxowM+e3LLFj
ETDnE8Wf0z2+Xe0PeRQRX1xRAQ4HwwY6n9CHsQXM6ZVqe54BRbkkqbQXS0Ea66SU1PIksmlMb3og
kLpNst1bDXb3MYstVn0xGWXzUGwBDEmmH0RH8jIV6OxAuMnSwmsHigJz61FZ27ZbWKklX1ig8pjS
2xFPUTzuyWoHrr6X5h8zIyqqHTMyjh1yy6ieLQtvandf6KMmbZlV2T79MNRgzHPuWHyD1UQFigLT
+sJYLr9HGbkmQU+p67inSNeNIqnOfyZWp6egxStbcQe70BW9R2/PyAgQNj5kBevGkNhBDBA9OrE7
DSEvY9zno9W4FAoXvrmFQq8XY1M4X2cE+H5izOsQboXNOUkoCi4jCkAtfGoxmD3KcQ7++MigKwQH
JyKDfBX8Cq+e7QJPDXqZMKqHRc5ktwgJuitjuja1a7YpVn2yWSA5AqnbPgpU/EumjePvzGCyE6iK
hMUpLOTNg5egd4tAEzsHtNb+wxGrIoeQe9FG9+aY9lAJfCDdZAl13cs2lb0lyQuGJh2ZkwXbNrIC
qmRMI1XmLJJWuzYdmQWkAaQ7wuoxMw+9jvpP7SZkUhmyVn8YaG8uOUL4LQxXSDZBbuq/vcdl5wDs
zxV/x8v2+90PmsMT5PsHsDmHVOTrk4s4p3V6yQrbKMqdmlexGA3VZLGG1CDL98qjsTTjOzvkd6hP
8388ha60hfqSNM3IFk5D6KXyIY0p1NIK/68dB4GrmJ1JZkTEZ1CBTGe2r2+nCLWyGhKIMkXVCJBm
WDscnUV7+bHoryRQ9Fqr5DhDSC75lyCR3AmG8ml1nW5FqsYdJNEejfWvzWOWcVA5ytXjDIwLwzt6
IguBRuuvTmW+07N1PNojTQs194kGGaP7Dn590qIEdLs7PXpFrQIYyiJSjgNppO/kak07nV6vGiQI
7f+gpgdt5DF8UtXHmeI8iIiY9DEiaZQBBmzHmgfPV4w4yvrGAgXPM/q0uXfxjVLvV9UMD6IwHzh7
IRL+xL5wD743dIaLX/nSqyub4e259G5hJvJMwM6So1abGMRTbrJbD5ilEVz0U98CP9prk+JcPmDp
fXOBMzM8xqDTI5vJOb4EktJqO/IabZ8MxpATvntVpUA/V2wZKNvs3Y4k8jMYySYZb7ZI50NQhiYC
s7MbsXHzbbpuKELFH3QePoKALHgiASP5DujGLbD7FKLn/vZjROSgnWCjvqMIkQ7+nsPhkmByVN1v
9DKy+JaGQhawUZBh4HTpMaRlsQdO6FvwgFpamvGsI64m2Q7qqr6njQSuSUsjStXORx/WetsESwuh
WXONqtJDzYAeCyDSG8mWECxMnm3EBR9xTQ67gRUXszOXJrsQMDH8xNpZ32uDndzDehnvBnKxOKxh
pvlhuzzViTPX3wCDXw2KYEeMwtQ9mWly4BdZrLAeiQJ36xmN8xv1y50PO6ObIc16laSOwZDIV/0d
0COa2Rhevtk5983oVV46cKYd1ogTgkLUjwvVdNzXKq+B4rUK6UapK/sAR2ZRuHFQqhf3DRjqk0dy
tUnqiEjfWjbJuafOihS5b6VwgTkCQWPnlqNWkEb3AfH26gMfU50EmsnLwYsmoZiHL183Bd36kO6f
ZFWiG5yrlYd0pKVM2uxGQmkeZ4nQe2soNrTW3CY/WC/t/I7hDm6duIxFimVuG1l8BMZrk6MAKf72
HJZnB7ZzuXr0fEQQ6Qcn0Eimygx/IZR4LoiQGNoFG9qYEsQESVDP8O6Vs3o6eVvPWRHoSakJRk7k
vxzDx6WBj5DzE15QWkww7YtbyCdL7ft0RsxkUnjn5jSq8RvNzU2ebwGC/1iGTIRgH/BVA9lu3HhT
RjKklOQW8kzrQWUiHd+nGyvtxFEsryWJ4YfMV+HtSWjgX4THjeaGVM/0Fh/TCMiuyg6318WTs7Xj
qRMDFLhHSpRNzs9LUZOw7Xb42VMMIQ4/Sl4v42dxxYcfXmC/OHTaBHqjAnZHxVxg5g6TWDkjmT9a
6rxzOjAHEKcROKsQ079oBUk3ym7UAUZHZklujowbS5F7ObEKf/fudImhCwex9CHPH3rBFeZj5vwd
UHrWRbY8JhHd62V5xeDEEwgNGRTCANm6vdNvrrYdP8nf1kZy5Czx0qD8jPXbwm+Kb5nlB2IS11Kn
/MzsLPOnCS1ZkZzCvsFGWESLBhV3fG7ZSg8pzq5z2swRXHPvmRmbDAdRVufORVDfQcUYekGp8vQo
lzIJ/XZjQRVAOC0V4Jtmt/eDh8gwIu4JcBsKPKzcV7GfHcq41BxXHFhvlw+m/RXMl1rYYjwGIOtp
Xft95yObtSa7BZpxmBBQAIV/EhWFXEER0WWNcfVf3h2Y31+Q5VEZspqYooTs1swjF0X3l/j7DPYi
l6wMx4L+GT63WuemcF5z6Iy2TTY6BxUvRdQ0lNxx+U0dwQoqVrF0jDSPltNg3wrTMw3mDikBTPsC
8VWcpdX+HpT+ytDvVbQF3It8ysvt7nIKP/Hmhr6dxQYthTriDO32KI/YGmkzof65GyNJLsqI2Sva
6YKQCaO8POXq6RPlI1u7ux6XRwZsF0zIFLIioa0ydZmVx5YH/dBS171EIqkEOf9mf/kj626CX4b/
zObgkskQC6fhCcFW1r28nk6kcfRRffbiCgkguZcu3/wEygJIhMLgeIgMDwZ1tY3ybuOE3yPlUcJv
Ko14Aj23aRvCcdHm4Fki/Eyze/2yKMicig6YyG2MLhoQuHOuyGGs44AQOd0C/pt99e1YfUjGswKE
qkdHCK5p4yX31Av9/sjFDkA/H34VwaalsgWN0IBGDOEQOpuUw1FQjTSVYhmhXh1u9AsyipPNgMsI
1hMJ9FYBjnszn3wJC8d21erjz8BGLJZJ6wVSBq2KV2Ypmi7O3hbpbNmHUCDdifzESuilzDSlIbrh
VpkygGkhsY+W8aHUjCCtn6uv6Wy745KWgxI1xu7r96BZeq2ElFxyIkRSx4jg7pIJ5iQe//uqWIvm
s/pMLYX25kbulG5oIhoAM5UPArRtnE9VRajCaZrSwhoVoiGH0I87dyLgbTpJ1YjefyNTRQzlbK8z
OKAZe1RWz1ahxUKc09emBepuHLQ7R6AS86hcLhpXjaYHwbECrz4OHsTSwg9sjs8ypywgNjrDlUsV
SNIjFwtf0t3MVC5RkE7kbrTh8LDQlWZSq1s6XjMgGEOgq9CXDTzXSaplxI/tqMsXWhm1Kz5HGDWy
XbkqbewC9+iTmFHhxvQ6SVQKClr/MRBJA0UHa5e2BjEc9saTnxOS5Id8xo1On2uqiVTol4g6tQpp
wDKiXhtEshPrexGfRnYKw4va6Lv1y2H1unXP/pkfi/Vt6X3GuLQ+nkiMHmkfjKImDX6fYoi7Gwu9
bl37oAu2flEJBVn4O3lNkt4dzCaBzOuSd/HMX3L8sb//PLJJkQuyQskLT8LfnqWIeEwAFUWm0jkH
9vCx5FkiH7Wbn5sUSKlMDQyK5iSmdQRXQ++7HSoWzCvDSJ/v6AbTyZhWhw/0H7arML16eUPmZf49
Sh8sQZVHdVGeMmWvnR+PIZRqT1q9SaHHT3IO6VgSju8ioHMjqRi6zevQ0BVA4mdrurUZRzl7sP1o
2j198ZA9H3zV2t0RUkJdNHgNc7JpuI8AFUVCWC1Zmh3MmYgPtSTYl1jraPbC93yoT1kvv3mRVvDi
Putnqsb9EVGwC9cSWNeRGUOAXvR4ZPzUnYvPHTn+CTlrKRVF0Alt0vJQmkxTrnGUfq95fWSjeX0Y
2cq4bD6LZdVGIXU6bbMZDl5ti6dBwxAzLmRuTch1O8w6Qx24oxcEc+/vBiuw9TCK2xM8Fr591hz5
sMHhtQJ9rgRznwjUs1nvws4u6jWR4rhSfV/EHLBrK9/0AW0o9KH/VfWIVUYQBm/yWZQhIof4hXOn
a95UEDEhODls+PZtmROj/I6pB5+orbsaG0fnLJbgwHHEonWq7GejLOqsQc2wBvk1qVi4K+YTW14M
v9oCcdQ33C/AkWZPh8whDk3zzQDxwczg0TpIahqOWaE86n/Lgwgut083CPiSU7YJAP2RyFK0+0gO
urtj429DYG8F4Rre+OHeHt01kRCt3mi55wnOhUqUPzgmJ3MxTG9CXkYchpu7Wad2cZKvCVQdVQbL
nDry/Etvt/IwE7hNr1XJ1YAKLYugGT6/59vl9y5CL3zB4F+ifyGkSaSsW6sgAW5RRLGV2tLE7zbU
SfZULdHeK2inNVxdFpGUGWT5zMkaK6hth5IBohWpHFFB4RY9tfo5uoPktm/BBLSE2h0ev1us8d4+
zzwJ7YirNyB2/SczWMNnxeD0RuGPpOh9Y2cCIoHHMY9Zy1qcaTMoXboe2S43x52X7sDpLAWs9rR7
BBp+CQ92yCVkBSkkdP4kK5mFITbY0w4dmBPcRWFB8TZBigdeDWoOY7m0gi6XukgVMkSyCni03Arn
yYaolGtJRSvUurybNFFGgLQNkQ7SW4R71bUOuARaFj2H9qw19IjCnW/bSDIgXPFKCMOpD3BC9Mbc
vIftEjmFM6X0txmFWx6CZvYmLrhLjYk+zlodqkCjR4zQKDc0HAnXStrE3d5yLt0tH984JPVhjkp6
05Ln7HI7V4L0HBp60M5k+cBWjo1Fql/5KwmlXqa0k078GMcFrMggKya95tKPruuwMrH+W8ZeHTN1
HdorBuZcvWXH5oqyoO8SdyWZXey2nnX1u+WURy96dmboavM/JYsBlfjNvk8L5Eu3Kza5mbx8zqD9
oyV6UQhdYITQOR6mOAUZShrzp7MY97JmFMx73t8uPD+9LOv02kylFO2ZZmRHrk1uiKXL8kwLd+Fw
1eEmWk94+yhqY49pwGwQooVmS+UksGc0q+SIDmF0mKSRtTxkczjXCFbtR16GXEiA4jZf+bcx+0wb
QJjmcgXuT1FHjMzP5MQ6ioKF0PKtQ0RKilr/CgwYBusO0HvVIpVOW/KpW9irXfdZBNPMMtHYh0+J
oCIjlDafj8ZLCSGt4gNlXK3OXdZo//zWn5iGD4xgMpmbmg9Dg1xYu1S0xqWAuMAQc/qibLb5TAIH
q3+z63bLdzzA6+dBUcgZyCv1C22+SBkvWZFJqnQ3vGKp0u/h1sdmsYIp8/7B/qTJIx8nI7lUPbJV
nNeJmnV7kKGyBFiOW6ojI4gmKI2uursvTPCS/ce+0RN+4r/6Y/yQtCG2riSJ1yktGWC8WzbKIBfX
XXJGUYJNl8dOxVmOe+Aj0eQ7oYIJuQloNzDBieIosrtQikMj0QYCOuUQ1oqUGNLfe0gA/3ORfX1k
RCdyS1+mnHAr1850+nk6+otOVY6MXYbB7+Bcojk39y/GFg62RqkEdID/JW52osJPlHsqCHfaFg9I
yCmv0WuiupbPFX2lQ7H7FpIgf4FHwB+m81Kric5pDeLXYxKN+4OPU6USlon/qVLCPjlIc9s1QvY6
Tn9JHD+iSzFHeLCibfz3Nx2lBdXb5KOxC3QJIMx+zdGXwQgqo72wks6s0oF7x+stzNAaGIIQ9XUs
/TtKMBrD6EFpMf0dVo2nEURSgWLtmuvbb5agQcuPeREnWn83jPdcnOqCt5VfegwaBBef7SX3BQbG
H9vXzhsnnitqlO81+fn/hQjAhb5VNbRmsAue0MD5tV+nlaTw5RO/5/434c50PTcNbI2rTggu7Q0q
MQzLYlPksJAKs8IPO/gNZeVQHlkgPyWUdZnGxf8SCudtWwC0Hfuqn4M+2ZEF9+kWJO/rm2WZclB2
cZ5uUROMponGxY416Mqt36BdxTqApgKbkh3tWGsGdyJHdARa+6zWSdnVDyg93OL3SbyK35JLVJaY
AOpXUYPXimNGhGc5/z3mfqO23VQNmvPLgLy0xdZGNlnv9voSZA/1aZ2DXtozf8zQRwFmOICO6LDT
3NqzW2f2G5ueXPZm9Hz1CAzeebvMP+kIuJxmaxMqME6+QZyEugxA6vBBvgXHBSADYIfB8jNxnsjX
BEOVyWNJLPquWyrAdTdgjTlreI7I0+YB20k47U6rienOkZkOvUIqGgwu6mLQeu5k63Shu6iS4igh
x/cHz7sqnBvyquKS4/SKEPPfrKvYeBGEdeRTMe/A16MKQoPxUa9OPP3T7K77q4RmM33vnzm4+nBb
kX40N4BHN5NlTHQWme6Ya7We2Y9DhbmKtcW1jSFHgsbIQKc4BjRX/yus3wNTFd4sxNOtvufb8fcS
0nTstRsYsuPdCRKe6693tQVYXNO6TJJw6wZ8rGYt+Zuea2n1SEvKkA6VvsftPcplyMGZZhBwhni9
H8pG8RXG6i69ZNOeeUuPyEdtepv7f+v/B06dVXXshcby52u+Gg/o6ppsQy0i1LVf3d7aQEvRHV2r
3bBp8P9op2vGA95AfGJAUrnL8QpsW7KZlvlyK5N8Eq4L1LCFHMTFWHL60Q8x7R4sw3C1KU8wdCPy
YT4KCuPkIbmCu+/DEelUh8wh/lqxwgSZIbRB0dswdnMcXmh+Bx5LXbaeeyyfT9r57FoNwHJTwrGU
c5vdKeUyOM85IHPQXQcOJwx3/Dj8Lm5UNyFRwunoXUEADuNNR6ZbBkU+Qj22P8xkEwLNdTHd7080
MdqrXzHiGU7C9jX8KgVjUlSFLV+7VcbJskRQcZTjuKwnpwzGjUW9eFyLGf5F926cMy3qEG6ZP5YZ
4/dk091c7Yp902Dr7ytVGJk4UEJYFO/0u2jA/20GgchFsHn9oQo54ApDpfAZnY2YXtSEZLWxd2q+
rqFQDrYyspv0q/SSgIGfWw2fK2gdrrHeTZ59xsT2WUcOV6f3ydKibiehH5mtWTtLPnUl+uOcC6av
OaIbC/187k87kJjeouJNrNNE2ZZ9i6zqgwIQIGQVPrvkNOLVPBrefIWWiQVulN/3C0Cn0IJvxXQ4
tyoivEFKgNlu0USlG8yArG25PhcMMUsWWtjxmBDryj7vHgnrVPaZY+3bdFKuS1ZeFQ1XXzrBD7vs
zmHIZf1MITr3u1Q+ktXt/ALntpmlBNK6/BjMzJ4M0Sfp2L3b4MCIaXudwvJBzDTRt0gx5nrvZsCo
qnlETJ27wGjhL8yehyBjy+4zrgcYI1dt0V/UC/xI05jWCBejsLBfolCsgqPyDnaDOvjE9pd0stp/
GBeiQyI1vV1b4dyUoj8ZFWM2eIZ2Cf3yz+nH/on6E+N/fw7h0emf4Ts77aN65bB97j4iecB310I6
icRdfK0yawiXrTL73XM6NBjVk20uOqonxQ84yzC82+sknmqNe8O0e1wzvgoPyUBduaw7voOGUVE3
PPtzJARZdsBKyTuAIe8bg/doYKrNjhl2iK4IkPnfJrz6dRyQSSX3Ot01nzbk0ua1iXK0CvbLxp3F
6zz8lP9eeK1xbhpglCHCd/yKT2/INH5LmezflqvMr8dBC6Fhh7iWiGu0kh/OjWG8CZh1G/30mUVX
xPh/dLXoeUzynjE65OKLxQ+KWUI6TMDh3xASuGRYRZYFeL3f2qjiutk+FYK1gTxVpcxctqCiXJKn
5lWYNHSZQDqLLFyNsPZDhrhJOlOuiXzm17bMQQc71c04G3jWfklCwrLPjQfrqbeDUbumyuIwhMAi
gfJ6TudSothuOOeTzIfgyD7IVDI81T42LaCqFUA9BscZ4DT96GLwG1GkwY+PWhlHj0PlN2zZITCe
uRZOeJIpkSmLLdXmWwr1h3QTbayEWFNTX9fnNq6stDdJ3KgCD125B6TGY+HP72FG1UoMRRFObXDi
dH0BcJ68dhOXeJ8eVN0xQLb1ybahSeTHn/s/0LoHmjhOhXnAKU9dSdZJRLLmE6vGN8DQqmuuNIHV
iTqTA2EA0bE1FU0FHknX/+irtLgoVdxLfVzRdUDskoiS7FM1z7HhXMsOObRSBJH811kzUXw+LB0o
1UCDpEghvwf1cgbN4NVDHhNwAzuKLUaI6cRvf8AKrlyZ2b5+wv7Dp/PHs4Cv7O3lSnzcIIKSGpqC
DcbVAwB/jXrxNkqClciV5N92a+rXbRI3pfynYZvJGy6SJhNZxk7Y6aUzyi26J8vKTZqEwr0DILff
DroL1Lf7w65qsXSo9VNYxUrjTQQHaVTaR9Rtbs/qBi8wkR1mfqwSQ6DzyvBoJ/eZd1UIht/xAzJU
tiC1EHZND2m2T1IC9NGPDmBKkXtn5uvhodbmwXRT9vLN13/RTXfhMj4g7PF/Bl8E+Cjgo4Xf4KIA
LjcVBNJZzX1X+oTv2MilNqY8kgN4nmD/SLK6IoZ/6ZYQV5dP++Ma8P0l61J5ggL+Atus95uRccH7
7oHMGd/BCnHPnnkcTUZKfy+nQWfn0WXwgIkZckKKgRAPRPbnuNKquGmWh0r0EZ70W8np0hnpkCXb
+1DUr4+NIXzMYP+KbYO/qzF2oIGjoTMzx9RRkX+/7uJbfp356QzWUzm+yRag4/iTM1CMt2H8mJEm
M4bRXRnsWgQJgui/4R5ZlsTVMQjUT61Wn51696uhRypZzgOJ0EtC2fFcYwgYRnPFTvXJ5X/OxJ9j
DWut8OEdEkvdNxAFe3MnB6YKRrZDitw9K+7Odj3tfjnFHU/gH9OdRWOlgxldbnVTU0tHRLWjzsNa
00GPPf//ZgzS9Vb/iZYEhQ18cpwRF9XjsqOXxVUgdKHxmW5HLJgAHx1IcURzbuzXcbsMWRmolNzX
MKwbWQ3b+Klu1TpWlwwaUfatNY8croIoXs4Bh0wzgqLorSJ+Ro6KUN9+IVYc4RLtDzJYxtfTuFKB
BzcjmoWRVldPO2LjX2Oe6LOtu+30YHNZrnw7LwruRRLKrEaG9SIbv4DIcHNh+KsWl2fmvMIEMUKS
w7vm3qD9a8CLesXi7AnBrJW8PUeL6uwbDrk1SN3Mt1HsCgbgPHQY4a6wk0gzdNoZ1Ry9P8b6/ag0
MvY+7yb/edl5Th+bdXQrldbuwMwXC/WJMNCofKGAlaRls303mC6lw0b/5GfK0Y22DSFDF7KPBxQd
QTjYOQusvzZuM+YU3CnGvYOGJ/xiuPpQ1xOmuiumbrWbpPAyIHzxqupNq8L8yJWiFCk6aqwUr/JZ
u80B1SBMBCfeFeV6hW75cZtMuKGbGHMEjswHVRG/lUyAsYLglwVwPNeo8TTHs9S3f2QfVA2LOnJf
XSaZJIj6ofWB3qIgVxSkjdsmUPURcpTpx7jToIgXgqC1nVFXrYJJ8zVpzOq1NFUkROMVA67X7XPc
q36GgCJSo8edoM/chMReODJqQS2wksshsmVm+JWaUyKZMC7AI4AInr2Hq+O1dg7JEWFZPChxKmCx
Fd6JtAQRBIwvWkzWvf8RzXBgGEgnkF6LhJV8lKYSy3vxgBnUaYf3Z/6AH8UJ7eKkUb2pPf+VKwCv
34ixJarASoQrwS6vC7Wl28B/5mnPTK1mgjg832AcPBSEm0TiIQGtvRDpZZXVMngvf6R+9TVs2jqr
LQtNzwcbDby+cvuH1ZPNQ5eBzc4MSw387vO65G1b/JmL9rfcZZ5SoQQ7oc+Z+emLmFZej+AFxbY7
uIR6y1KSIpcK7Z3++h48+wUkb/LUshlCE4NrirMDQM6Bi7SEU9JpJcqwfpAOqMaQ9NHDiZQ13I1v
i3uJ/Btxhzt8FCAjkwKaWu2HmlSQNWiwFFesVU9XtLbSZOh/nVhebhcT/LMFclbrc84tpgayuIxl
h7h7sUZrMvwZeMQCq+3xjawmYKRQvujVwZKwAl/qZtpLXg0I7AE3XjnmFvhrZg3z/vUs+D6zwDWB
buw+IklKe1NC7Z6lM0g0FQIDaxN/wetBPm/gyfA//X/WdNzbZI1M0iopJypfPnjVuSLAbZ8s2sS1
ATsGaZ/5sOQ0AD/pslRObkvZnViYOdXIMHzwkxVdMSD8WO9At6Iri/qHCBlS7bA2rfy+spa0Sr/a
fOUNovTNA+TQWF/8WGHB9WSCLOqv7SMZCJcmwlF+s2S90lpJfVJHjoDFrLmgjzlWifmF6WWCn7+T
pom00Ir1cwn4PdVuy23ZbJ8YlDZqL1ouorh3PHx58u/2o0vd8BVZ206SekxVYNc01AFeC3sqRPXl
0mGSlqxDRYKm3r83/jJ7qcVQYYse9B8k3/DD9BpGOEkHPSDwoOAqHc7MDC3SSVBSHQ67vLhn8Sqy
zi8XLZaduGTiuBUXMvH1hFddoEqncG/w8wP36k6zvN/VYF/TcVCkbYY+LLriIhY+frrols6YEMAB
UY8lP7Lk6XWskTbs3cdQ9mvsKgcfcyuNAW7afNOboRCyKsGQ4UuT1DMOVraIVgB1/6ZOcIuPcdJp
aZWvHaFNbuWsTsBhIwmVTiKFbns+KRcG3FuRc8hSrb9xD5kpqvqQ0fxfkbRfQ2954oPTEihSQNK6
/8EwQlwEkvYqUchslu7kCgYgdGSNzongPoA4MYvJ4iT5YyC8Mdi/8B+LB0MBaUtaj8gOsdzQ94ZN
3639/C0i9PbrzfeGZNLEVCdUPQRMQSrqY6Q3cuJ8QadRoQ0uhniUp2+3IM6KdTsulU5v1kacDkkM
tDk1bJbM21PVwpgIOEjZbXw8Yf8N7NNdV2q+tt7CejFexXAUE60kRQDCMN50e1JOI2p+BZzjTCV4
RoVRY9NEP5WdLuvddkNkHnSp7CcYyEhVgNEUfmRW/1f9nu43hadOE8O/Q2pytTizo7yER/GTWJ1w
3G7T+fEVGyD4NM05X5MZ07v2MYm6gJ0LHTFp0pgyRFLzADk6tKlcUzupv++c3KiX1AFGQWUKzlej
IN+ZsvTpyxOE/tGVx3pPJj9Z8AVSf/uMnT6XKLelVZE/UpomGcjqNZcq+rOI61nu9vFejIs8bDxm
nm5dLBN/wWk4wUIHrMwtsIahGsOyqs6UhU15DrJ+c8xcBIZYD3xqWnFVul/fL96O8syj/BQTRZ+p
ACi/w/LdkDjwYLviDGEeRgpZbk2Wg+rrE138sI9g7KerlSnx6Cz6I0TPTz7J2YIRDDAKYBn4gHBa
omoTz+V9PT5bvf7FF9Uij8e0736wWvARGN3KTCdsgSdvsr+aLdiWyIklLpnUt2VU0YFvg8YmePgg
cwZPIzAe/u20MZTS423LXd6xHqH+69NQLSNQxn839gN+Sh3f3ZNiaXlyGbixDmaSOoAxeUuzeF8m
e5Z2OzMhgonZqgRgQoSZ8+ditNlI7K6is6f5UZURFw1zL8DwfHNPkVQ9M6j34yqRT6I3Ww11AUX8
K4yUPBCgBEFtrs/W9YIaQ+0Du0J6a1Kw5ile3LjE0T8kd/XBJQdlZLIoCA1F2gAY/ZAPfPpWW4mu
alDuICCNExdzkY/KjNsGkJ35IwZp9yaYINmWiGxXisNyRgWZwk6R0E54u0zgAG02p58Xhk4njurp
94/Ldqi3LtkLB0vNcvddqSQ4aM3LLfL6/mrwPUAur55P8GtznobRMkrGZ5NF8drlLhpW4Th6pTwa
BSWM0NMGfwutWQCFowJHbmaahowJLEORL/QiP8yka+U/MI0YdfhSHYIF7qUjtsMMQg26uRlBGV6w
IuG8FGWurMErQKxypz3aCFDJLxicuHeejxL9Gqw6n9/7Z+jO9wVFAP6vU1BgV/xQ5yah29QoiM0A
wMtGKbe1SnXgID7PwNz8maEy97P/HxDdUgkXYAL9flCRqHMFLb4iFYBrdplgWVpqBd0fnn6r81xn
Mn8L5NsxAe270ZaSr2jkCBUlZbwr2fYPyLUG01mij8wO8zQGIlDVEYpHKgzkvnWayZRfbIgG+I9w
RTLsFP2hpWoNt3amYM8mhr0jMzZq6M4SBXhylYejvr3lqebdYfbZbTktcYmo7iax4rmLSuu/nLwa
1KeefAQFHch2hwnSnFg3MxPXuywJn3eZzi2O2wQ0XlRoJ2hzDvV3+S6ikyyeohOmKJ7tzoX1UVnX
VRqZTsM8o/mZRVIE9jnOrKoVsWeZzOpM1RnMQ9Wu3XP3x97sqlS5W+2jnEManZUqytc+fQJ+YzOG
1N+OUaI68i9MQ+xxc1EVwcC81+ab4A1wifSp3/Jt3qqcCmPfmulD7kRl8yXWgxVLTdrMbrm0nGGI
D80Pjds0z6UGv17D+bWoVli7qQl1/noPDVQIJQVYGtxLAyl5/Q/pHViya+uwWboWvKDnY5B5xRPY
EwQjcBE9347j/Zy9ERK+PHKkzNSPuuoKqIEaYgzcbN7mAlLv6TomKJIAwuktdMOmKH7WwjoovN4g
0HTlYO+GR6+MuFoU8Cos87dMjzY/rCdliGhBbRe5UnQYYdGNP0M8GW4UodRuqrwgKDKGM2nNC0Hs
RcmZmBwLVIHXQmcVta1MnclMH8rAnAu/gGk5wS2gFOh+MrmDwAEERZXAF2tj5VbllA1BDVUIzrKO
i8EUTzLJB5n0FftB/7FdPIydOjD0o6HSu2WxiU4+gPWWbY2wu98yDrIUoxcTUtqs+BB6n2XLYcKF
yaEBG+coS4zZwlkaa9vvaQMWXkPDDg9HRThS0zB8j+4AJWdZhT6HPiXdS+HXLydA8oZU1X63rrRR
x6rNDnxPSSnNkcjnuqKZtL9MzcIqdayfWagEhJM0W1DxpPdXjtmYnCGCSC+grnLpXITpEYj/gGHh
H4y1H6JgewtIxw/mND2YCgYaxdRkLCEQabS339z/01Go431NfECMq01LOPtk5zk7Org8wNMp+fAs
p90QQcG5UGKwi8227mYv3w6T/9NPFIAYPoYv61EDXX3vY/TY4HBrsmSuKpFVo+BJPkCJP4bb10PA
IYtD0bRTYZOyB6/1+GfvL70jYfUSbyzjo+zrdSqXJQflLxC9p+f1kOoJejgcb/tOk5vALmO7BegL
k5XPf+S1Q9+GnKWAi0SrMMc4KlQFJPUZl6Is00jqyfmAmWUZ1qpuNlVHbgUSP/6h18fZ31IrFhgw
WxjsAkPYtE8NOwfZBGJcohrKXu6nnSRoS2jC7cDWLK+6nFonZxsVKGjFPrzGrAkvcZ8Newmw/ZXg
bCrOYTMNo6d4d6re8aw2LMtP1ZDTGcDmwBYMmBWn1X1sd8lz7HWxMsjb8IC/WydBSyCVIrap4pcW
UL1BwtXYmGZmX/TnG7HBYgOqdvkaNMjOEbzkpYgju4BLdXuQECwQg/QkqdBIg6lq0TUlSMcDE31k
CZDHxTob9HyFLPzDn/VJ/wvF+D4546ApJsq4Ur73xCQQ55zFnSUSz3QTuLWwrRAEnguklGL/VtMb
3tevhM0BDjtWsxfieG52p50c58R/8PLffw6ita3Kkym/9sgMx1PskrKpJS0r2YTaPsHJTc9TwjO3
1huGIf49cBRC98uPtxkAU93hscZUm7E8yA488VTpRn+NwkPSXPfDyfCUZ/ZUtsTywEn43dN6d1Xv
Fg4mE3QcOIo9oF7Unb4cRbQFJJcegnHsCIMwfSxEiSpT9vL7Z3as8/TwC1t6ZLr46ALjpPRdgz45
eUza46R9hqz0+RQD5y0K4qS9nmnqtgF21BBi6I6exm392Yr6x2Yz/FhQGUeN6Ho0IqQYdjgxUK8D
evVW1XJ4tqTwFXtmN31lFylU1e4+xkF+HSwrBftPvMVlYxNsAq1bUlmj38I3eJuZsnuuB5yTSK76
Ztk1H6Nc8KOxStG0k6kGh21zuxhYZX6U1C4ZsUcz0CUAVvUnLi4f9SZP6d6PaREAL2/snKeZ7v22
8zVa8LNeT0/wpNMHHZMx3QQS/G39jZaaXcO1isWq49uhjzL/qrV5fXeOvWQgYc77/wdOhWOTGFg5
12tjSBdxCJ8ERASPVEe7XJ2q5YnHS8VFFxjT/HRLf6kTdiCcsItw0YSe1tipZ8tW+1IpLEexalFw
8VgNxZx4F5cgB8cltsJTzbkgZn5yX0uutngmlxkXeBDvzG5YV0X+g+OFak4yqIqwNcbMYDQ81Yik
vI9rJs694Q5iRvwWbOkx2edbxNExbo7Kndbcm7MzdsHveGD5NAHkpsmBRoSYyGx1u5jRN5r/EaL9
5AU3581kADJ8qH0w57GfCKeopPO47yJBKTi56u6YmsHoFVpOMWHIqJ+ZKOMQEe44RuAzF2lj+v/D
Ga1RwvkaxXdlFdF54nUUMf7W+ECWYFY4B1sJJHDbfg6oHOTc7XLjZkNxkzqddGL/jd66oazYGBh3
FCzIs9So/Qj9DlsgcSpiWg2JuRFS5hiDlrG2djPVJRNFgjWJn/OjxhlyYISQPXAbAqkpLEPagxOZ
ur6YhEMA7wHeWhPOgJSmortVOlbTIl11sgU7gvZ8jzFIM0LnInxnV6qtxkgw5M/50D1sQwEKfy3Z
qQLd8UbBMrg4vcWJrbPe0dHSru6qPSG2RyIT7USDjXQHLAu0Q4qNi/CEF1Hijh4lHeV3nO8pckNU
u86b77mPAHQsINny4fVQyQcG+FVAa4AXolgVx/2cPXoe4cs7SCX9cRsFawsZP6TG3oOx5ltYoLf4
eF7n6FjlXXP5Vt2XQJwrUYUIger7i/ZFjQT4DHgJc8p0xUVBvnF92WkdybLFOPPfphI7GScr7Z8r
MgaU1Gd6YR+Trre6BQddSWP3T1k3rv9/42WofCNiy7kc8gKNxEHSd6tdIddiaPbj65mhpeFRsBAV
jV2ZwqWYDEOv/R6nyK/Q65vENxHzLze7EFKSVXQWtDIV/l3GAv2Vcx82elInP/vzm5OLs20IC0ed
fHugzTPVgNyuU2vbTc+K2+Dj9y6Hi4BR40wiD6c3U9+jsemgfQ53h+azEQELJFHrcN+YxZpANyUd
/RRzE9Z1FUYpMUZjVxfXNwYp+YyWyOG6NtU4KY4cGHckNeGUcn2UTOMZjigoKArRWGb5/IMROQgG
KVDYS8X1PzBOoolnOOfRIGm5C5dpYVr3J/272MR1VbupFHBFuefhaoV19bjpppfIe1KtIZB3dc9u
GIJiwt9YHGn/JTfhcv5jYcwJxcQDc/BzAQhiEjIt8LJ0W44V79489qK5ijLksaRUW2UC6DxDGr1Z
S2Ig5+1MkEkzB2/9a+rX9qD8ptW0v6Zr+oXDNOopbGJYF8KyhyXXjmgxzLmo4hU5q0u4qaFN6Ihl
2HD0k2cONlMu3Z54OxTjFG+vqs24AYAd2AaW/iVEfMeGWuASPpaoktK7+7BsALDbC+wsRjWDoTmB
XA4/jYG/pXA6+yx8HRKmKwuFwGymSIFl2S8XLOGjp6FzDWSJpzVGROpLPs/dOfkZVP0mvsFRn7/P
y1LdWonKfYQmnx5e0MZ19rMar1KYSXQ3ZWJNfa+mWA8ZwPh29ca/eOUFKMdRgelqkEK0z4R8bQ0M
H9Ksg5t65MQyyGTXp0OzchYq7gD/9NHxrIFGzXyBOCTNVyCw4tioseJEgzua1hWWtf8DUhlZNMYZ
/gqGLLMmN9xENsjiTkgRCOp8sHf18PO/XJZpJ9VKooITzngB3y7vNnFKdlXQubmAhaD/BOWXCcnw
oKKGHKsg3FKG3aMRRCvtcoF+b1iEbTVlmMuThD5Ef848HZJw/GOj80VSYEk9PV9uDpxdVpz4Hhsh
J4lKDFG6JE2ziHk6eKLsUKICAmNHC8ZwQi6Ij9WL2guqwpTp/6A0CwugK2GehatHShTNdRo9dnxV
pcSPpPwtbaMZ4G5H0mi9PcYsbH80A6ujdUttYAUbgrs5fSzWFofGNCUqwWKtX09RYjmFtpAmCXyE
QqYfNYIn0NAkFh9tebcH0K0kD957QUXp7DIMxsYuuE7shGWAzEga7wxelRaqJfqbcra5yaDdQBhq
X8RwDVREJ2BRV75tfGiTKr0bjkY4n0GT1uUk/A1a34ZrEBPAQ4R+pPvrVUNNZejJ+bhd9iniHYWH
dPshgQQVaJBEoF6cAPgegNC76LjOxfdCOP+CXhOQlIBoPjmisYQ16h0RWHWO/+tq4YQ38NhQ0TxT
sTg8acs9c76Bh4NKUMEHM0czr1xo9mJ/3NihWiXJsfBr+Ckc4thpKOfiV1SzGR3FzxrORDJZp1Xg
pKBehQISyY+UQO5QfMbkQZN5BXYEvCmrE32DhEi0BXrrRp2W3M2Jg38PntOdvvrNLxqBEp9GtqZR
2vT/KS6rlrQjfjleULMasb2gySYG8p354b4HGeWmDPBE4q30cmjM8sa3w+ckFiZtsJfy/ru/TnmR
rDpQ6/sCyglRTRr9qLHo3iq7tC2aG3hybFPqFGPn/WllpfqcBKpVOSbR6VFT/KssHTvKKRt2E8+/
hHgdKgyvR0q9y6mwLnALwRkGfO7I5gCsUIbP2ng9kr1Wp0OMCE1hq+UujhjENcizMqdLqaoYaJQG
Id8+A2ZTN04FLyHPshmJZk4FZ+0+cgWp/9+4MP04ONz3tCppYNHrbwigvQnvTXN1hCQnF2A4HaYE
cU9p5r+GpebgjWJ46w2DugOQJKi9LcImJdUZfL8HgBY/dcCezIEs5uHAgQmyvg4Sm8Bebj0uqlu0
e7A8euDOz9ut5Pr/zu/dGIeH4nHf/BYjuFa5aykw0Qa79MBkw0nUp6T73EMtnrv+Th18dBnskfoD
k4q2g3igP0+/qpYR/tEV9LxAysp9SVn95r6LlfWvvLbulAB0Gni6Hn0k8lHpOLeU+K5rXq6/7uAP
w3buXyYDoJJ05xGfOMiPDs6luqsUXZfqxh3FGFq+A29sVpmIjG6Yhca7hsbjPWJkucds40fcVzoQ
ZFjLO08fOjirTb12uVRj9Fn4fPtuEsH8rgOTLQrb/TNAdoWZ9MA8BR4yo30xufNGNaB+Q+Y77EcR
oILxfb6oR23tXTR/mRxB+wZfKX6IA0LyQCruakqAIWqUDXA48SSYWA61e4Q/fl+QLAB+jjqg3onq
L7Fp2yudjZwDuXX3uy2dXLQmAMwqVXXmF0SkDxrSEeD7fP8O8tqB9DTFmy8PCsAZLrskkyVd3iaG
MfNVR1g9L9JVvRE2pFYwVmd1s1zPMtROwyJepJ0/ZrTSK8DUJI0wtgOQH58OymoBFKwV9/j77CsH
vcT6bQC+ypf8sr3uDE98+cQKGxLRNgGZpE6n7rZ0FImTFjMOcsm7W4fUOKqg/HQgOCsm2VwkhO+t
JRntB6YSngbzr+p8Xa3MWVbpAgSdxr/+zCSiFO4Wb84ECQ2YrjCBXn+xgNX9cat+l6yOFw6SLTe5
q7cqWeillsuC5GNo9vv1pYd2dVvR5Sk4X3UJ+t4rz4s624oH5MZEwSvn8L3oORrzQ9/uRLhKy/6w
Cd9Yu3DaqOcdRQhglwBClwexle65t9e6YhzhZqeU2+Nz9pLwUOB2I50pkSINa4Q+1/ybEwwbFLO+
fK4Dt2mCRa2ZgIJ+2tYSxygXeW+Z8Xv4oWxgNLb4WBNu/4ruZV8sy9YUfMX2D17tsxxvDA96dBDZ
xrKYL1M3MZmHkvTrpUEFhkwjbHQ834ls4TlzaQpPNY1t6TzH7I40yPBVBwBVBAkXNSch+iRrTWMp
nkCucc5xyBsuUPlUGkzkWuPaevwk9NmYXge4WM3e5C2Mb6G3nIXh4401Q8LCc5hLWa/azRQjb8i8
DK9As4oM2V4tFmZJmSKQKtAltOuLc6fykwYgBaUqasQNxh+8YmxeKiSp+Yb60u3J1klxAyv3zHW8
GGX7aRzI/b2KIV1h+f7HThvegQnA/s2FBhDXU0vRxELWAYM8qli04oMLh98dnDvpVsPq0rvAT9UM
kXJ157gcttfQVshJ7c/LXJgQ/eOZYjHp/bPGRhlrib1Wn5ix86DW6svqBqOfNFGBWjPSPh7+qkwZ
Fp0Op9ReJFj9/RBYeojHEsHeULJlrI3qRe6a4HYH/FBqJIddnYCHrfVcun8CBtoMNm8Is3TIF46g
I7X081lVcR+KScTWVlndco9oG0dUGiYQ+SN7q3IQg3ppVNGtZaY4/k4uLqnsMwXvq882UummMIoz
wwAxwtkOpYFRDFupbVqUmsnzFtofuQtpjRagUdojFfYHbtFCd8+xuFaeNVxFL0+5ICqGLEQbBBHQ
BKZFNoty7QdqgtNXnZ4z2c/a+wxDYyhegguuG6lwArbVgSZcepswcIEzQmzzSi/YHS3+TEtgUFoT
LKUkal+TtUkN3qTZnKDaPSOsS7aMy6WIUr8hxkxUdDeE1MeLQySDif43XKw0J5V5PB2OtQofSpSp
HbI1dLg9a7OpQok9Ol7Gg+QiTt8wtUhtSUAB/zULnqm/RaokxiM1xmA5ULcb9GOCRkLJlQccPJJT
po5+eBE93td3gY0FcJtWxChxDKIWQLnoFE4HNqNlA9nS8kvaf74tY8s1D+pZMs17e/8ccYh/RTvg
6QwszJEtc3wixoAOCZcpBiQdu80VImRQsyDNwJAMlmI1TBwzZiayOy7uzPesykuTc9UQmKGAlriV
DRn7vkd/tRBY0xryChqJushyzqf9lBgjYl3bL6RhkJEUKuz/qYBmNcJrZFU80KNpVqmoQ68UChfj
20d58upTLcRltaG/6hhd8IMHjH/5WaepU7FVzxmsl/hKwuLnb6GUqKPQLzytnxKrayKUhdmUcNtP
hlb5SN5XUsCEtvg6UZChOuingeAjqxYepCXXnScw3oDsT2kcwfGjF2zVgRRAcXPWjgB9Rb9ecG/Y
3q/HHXD4kqBPczfEGtOyDKG40uCvCLy3+VWClOuzqGnFx73YffEl2HuRpqMB+V/0nNfJ0tAeXxEQ
NrkS7jSOO+VSuWyLnrg0+0EoUTj1mIQSqwDTmA+ULYm9AMI5SG8gBXbrjmFNS2erg1/JsMOgLVN7
LALceRR5Cf4Uc59ne6Bq0Ik4Ic2x+SxlcCpHGnlRqiTwgCiDJ+j4VHYQy+d0OOVLL20TJRYeKz4q
9frReV6RCKQLS+FmobcrHZ1JuaSjjpzUWxiiWcyl313gXbRS8ZOuHVXkmAMxpK3KomSHquhx0Sab
2uWmtRvK3KG+h7hwr4eqPSQtpf+69KNyMe2hmugMBO1/s6au1kGKcknck7ei8Oka/Eml0z49VS8I
sv200mbH0e/KQhaP4kMkf6RoPffmRhKdIl+5k6Xzj8RRckaEpU66NBqOGNTCHN8dH2xUHAWttsQM
ZV8u2sR0F6xjseazajgk4a5GKMqsr/02K7LLfckrLbyuD2veFcB0LH5zvErydT2+b5+s2FgAzSfl
rVDTPrjHC0oWvRa/LkKFNizRKqgqErc3lwsLzaMTtPHPO/L8o8Nr8YYpiMk6T69sOeSPJBzUamG9
yaLk81b4mKFcCnJcPsiCktwGrvEozoa/Uzx080GXugi+BQm5KTvNyNsA2XE5LbAiayNnOyiJ74+s
GXxZF+piY+Vu+wuCi3Y2PqcqIGP3nX640niygDM0SeRvA0h33jBvUIlpF1/hp+0XaKqknUwZyUMR
k2e/9NIwp3M6bwCY5RqsRPIhDfMF0lZXZVhHBqA5Y5TAsF/Ev0ayGMymBp26V6n3qAU/NPtdzpgR
Cxpi65IkiLBsPjC0VnbTnyE8DjjMzEwQqgcDWUtxA+w7TjwftT2JrJGwZVYUD8AeoDPECfft1phf
SvM0zYBvSCLpiPNl/RVXvnwPoLEH8kZRWqlhRhCi0VgdtGbtwiJzpXGGz1IP3Qb7WCumbGzzPdW4
eTn4irIShU94VlUTkS6ur2OBrlJcCG5KcNQAv+FSKlWR4hRqlL7nSFT/3Q9iInnWQ9v1+Cv/1LR8
qkyY5AYKNQrxlC9aAsf1FdpqF6vdUrizImIbwmdYEWh1BOlBk55KKTPl6pyjBPRcQol3j62CoYlx
k1r6qVdNBwJDyTTpgfm31weUxAsCYdAQiUo+EgAkqeXqCESoZWm/qVALEcpxNJfZ9k3kNcKpwQS3
woJaVdjGWG2xlF5lZNyd8j7PV+Id7d+dM7ilBP1dcgI1ofD4hoeGMV9N/6heSgOWDCiwj7IdMTr7
dDKOyQnczfDvkyiAyVLGHrs6JfwTpihj504SOniGgSZTVQPOKAt10zfD7GFQnznGP268z5ryPxdd
L1GZfFDavrg01eitHaMtK5BmecZbNAHtESB1rLJPExbdf6d+a4++EZmdCLUWt0bT/eGBvjGiAnbu
5HEkc7LDNPjSs4+kxPbrKafgyggCY8NGx4JkPPfbzZ+2Ks97PVEoJhQPI2VQz/0Fsea1p/DS3pzM
H3lXK8TUZpLJqZyuUYBFsV37qNB4eqsQkQ0hYAxLOWObD9KHPTgekd+yddXK5/HNU0HwOfzhAudE
uJ7rbP/OKnm3ncvhyA+8Y35mW9wEa7k68Wk3dz45r3cRMtsMod2/RvqxQ1HovRN1v0APTcoAPQom
NY7CF6uoD/2pIwnaaFW4coqKt4pzlGJ8GFQkmfNvUKKy7QJpc4UXaYJYEYqllj/cFUgC/NyQlg4m
Ce7+iUKyZ6CNjpEwdhTwaEK2u1zJ5MxZWgsZPyKqNaLE/T2JMQceExH75VAnTkIQSnpJLr21h0Fd
k42nmNMmKNjTuKZIVOmK7UmW63wp6Sxi1EaCV3SEc8vgADMqPL9f7izhQg/SwpY+oWn2T+tvP+os
I+eN6rN0Zkm7i8rRB/K/YGczB3EHZI0PXeKDzQvnFcEqqhelxXGvwvVVWX9fR6+lHXbDWFSVwFZa
IHn93BkrK+UQJrTcXXmBtmbTYme3wby+9asB+uyHX6eXefnMAIBEBDrApZAKOW02P5SoTtaomk2y
SamhJY41f4Af9VxJFfhcJqyan9hkB/5d1Qe9DrEkvoMIbjiNigEJ2IIXzqzTSVAeRmhxt4KX5tM8
gqQDReduOV2Wa36LB7OroXn+PtPnh1tlT9jtdTVZKOx2CqdYDXnr0AY6gzKmbUyv4NwCcYh6MSe8
vbxKkb/9zrXNYxQbG7bgXxtn4/NG4PDQ2JUolRb5Ux9jWVFuJTrCoZ+QdlSu92uAn+e8euia6s3y
9BrVSCutPU3whrT4043LN2MHckpJikz04bqH5gtubwzh51LthUE8j5fLZV6YqLcV9Z5ZhS3YSVTC
KU6olBrLD2+jCi6SGxvpnXowmrJqywYVef7L7cSAPM55taERCl8LHPeKo9lPQ+6ZLvEK4jIHZsv+
lm4hGmOzMCxwT/DoSJi1DrQN27O/2EIeV9npRVz8ze9JeH5OlBj4CnAQulYlzWZMLzXpoRJDV02A
0yW6rGDhT1/yi8UBcNeb67eoJmC+pkpn28r4f+FQJ9T2Nwwec6FfWlDmZSUYAee3Tl5jFDfuXteD
684cdQsE1U6ewgl8NEke2f6ucZ/REYkLUsHyhymvfNOvujNTCiD2a3WA+9g4YOdiRWX4+TlhIF3i
gntyLaP6O8ZJkTLCU9nfJbS/1s2IPb6WHCB7/TcHPmWBxYtIOqI4BPmmcC0SwCO3A0iju3HJDxyu
vduzp1kKRXMt1q9JH8FA56FPA+JcNLfOFJ9gF0jG/ULn85D7qGPVkeRUIljAPxI8vlMXobbtwPrL
ECpd2hSMnb/Z2o6CvXTWUBYPLMuXvMN25f+1WPuiQgA20QCAfztLN4+ndOLZKi0/7B5m8G4MZBq3
8IqKct+q2OhjqCW3SVfFx7tuQq04kaA+Kk4CmIep0oGbU0bZvLeaY+VDYbx7MMlrK3o26pBl+N+0
j8gdlQNX8PCV8GwMaoERGDv3DC7qjL0DGRPkaq/9ita+kd5Hbc0rIXG3PI+xCjGANZWXscalRt3L
BHQYP60BzTyJHfgIP2yBfkHWApZVp4UN9Gvj9GS0TDx0+hHdSqRLFq4cUDnCIckdJoqOIdK6SqWT
xVo3IUzD7OmXuOAVXOrMSwSJgocq2JPz8bjmfUUdEyuAcPfyzvrkSmfoc290AVzpp8PzA5FXMjxP
6CE2Nq1CHOJqQ/91dYHOcAwZh9S9bLchie833dUCqkj4CG/LTbaffFfHU6cmiU/BAXS2WM6TT3ss
Vk8iOuFWxXCEqTjoSXB+lo1/XchG7cxrcPkvD1yDFFtbVwvGm2WoscRxUOeXNeB8yR07+DaRoTYJ
DYgBOLElAKyhgMr4nh0H1Xg9j19xJWKchtdD8rFc8MMjnCvoqLgqRu5/tdF9v7U3cFnGiYln4e8d
+b1x0w+M5IvulTNtsMjxUf2R1ZlaUEpcMjNsf0RpgEa4l8ekUiAQ5PrglLPhamwY0zwgGK5qNjzk
IUAiHZCGxncsUR4j5oe8xcz1ZkXmWixn0uUOrE8xfrnYxuM6aw4JUccewQ7WKGCH5LaB1oc315W7
1RvG0EUfoP89SXWQ7wgdrhAssHgH5M1utHIdijwA1mUtBQ5OlL2ld+8fWmBNaVWj9Zhq47Xp+x8+
qhEzOVQFZex/ZAWZfFAxh8EGoJtxy/Wbe68ciXKzm4uVrbEdQeZ20/3y6MON41bKqxqqPj1uEV2m
ZG5vlE+in+w3MB0lN32ZiJ5dfj0fxOy7Rxvc2mbuvz+76wMDQuDZDE0Jj3h4HSVR0Qim5/CEHg3P
arWVvXHeZU1J5dvY2C6d6WaWJ3CYCVtO2+iAB5eR7RlAfaBmMEGTjWAnOcMoT5ciz9dcwJ3q9fu5
Jv5Idb5T3uiITerb2SAKj40IK0ZFU/qsvtdTXswYOiQmj6ZJzSs/pcDzof32jnKczumd1FUlO1qh
QEHiufjF6Cswi4Rm+6kgY9pmqVOeblWkMsCCSrtsJWuwdnvHYr18nYjcZr566r9sKK7WFygJIdI8
BTdyvrWoWOiADm4CxH0tQnR1E6+SdDtRvzr1QhzU3sJzKbmtdRU7e3RjFjpltynz+4Tw2Ml3pUSa
79sK+fGR2WTb0ZKEiXu8KzbN8bG33Z0b65SjAtpWlH1oTT2sB6dLPPi7l2MtHya3zsk0qMvwsziR
2ttORKHWDdj/6zbyJPaYtAUZTOwZ28+xAm1+c8rcKE1gNtczjEsgLmu+piSuPULQJFAG6nPxx19o
GHurQ5rt2rbql+NemY3mHrFn2ydr+nJTNYhndrlkNz500D/ZtqX5c0MQQyZaPgQ39VbJcmguX4iI
+8gEUDaAmH8x/4Ldl7WwjSVFZoT4KyyKsUoE6i5T0nFpD01SsQTO5tV0zQer0fbWSZJypmP5CU0b
TqlEM4HfF1Pacqz5KkvgJs/06Q4vXQp2WEx9ZRycWqL6fvUYm6GuOcIXChHOj113RNCI1m5N4L+F
UPnpVbEIVioBMzBdyh5xdGt0edWt9dWHTVwFFCA3z/yIg/Ju4T5JYwtYyh37wfYZcxXH0UHs4NY7
S3GXdrLx1sfGpSfuYqKmjO3wGV6jtlYOHhd2aCH1Ni0vgvxV4yJGeQ5WgZGGgDkpnf0CPOmby43L
RqO2MzqeJQdItUsLG3wCBJYvYe/+YuxQAcYGExYhstm2pWOWhMVg0FFP5fIODITbv3wdDAg1RVeD
i11ecRdmYqUxQYZfnlxYbZjWJF7SFl7momx5tscxJP7Hj8MXIC8t0Y+Zzw0+ELIzJsOiR3cCXM+9
EJ14/dp5QY0TjyZa7j365GJJ4we8xM+iFhEeLGfB91vj/maXe4si+idL66bKeg5603lKSdpFSZwN
zafAFm+/R1tz/9oByKltX8DvajTeMrYKmf047sbHf82Gdj3wRzOKI596XAPHby/QbASnWzHel1qB
fgEo10LqnWIBDbA+xd04DBDFywi0IRLmuzP11cxkZcaFWq19fY0xZsbzjh5qomdRUtRD2DGKKjcZ
//2XOGu1OOXXiyuES7OaJ3UoWcJzWx/SKao5GiLXBtpyGDjT4HDQW75QeOU/noIvRuHjRkG1J8s6
WP5hVNpCaB8Ta0JCFSUm0sX1QfjUECOrTdd9+AFaHWPXGxB3cs2fXblu0EZql3ArPrATfkS1osnP
nGgAAqbyxdyTnoFd5pS43lTULy49w3JxF9IGbtiauAdTUw5WN/oWEhCY/JxGWZ4zmdfW/BaeEP1Q
vInkpjzS9fL5x992bMouhwiFcjINniDfTAr6WC8/vJ79eSdBZB4y10C60QDou5cyjnxjepjPMOmt
+Bvr7GeXc193scljGPvx4Bdjzol38UaIGUAvdYST0u33BzaRKebBpdqxICLeVxNlHWe5oF3e7NmX
rmBPP490oGkNg4cGuaoWmOltaseaNwzMQR/6z9qm8bQhAysd9OD8++ZLYSX2DLjZY4hfU2c1lra/
9I3gkaQd+/Pnnu5SkW6b2h4RqMXRDsjMg+P0+5O0GtQGl7I/bEIARj7su+FGD3m5DvtDjGfvEsQF
RNRoUJ8BQcUg65WjMrUTgpUR11bj2g6TL91wLNwHgiMgG4vn9O1u0CrSUlakYpla0QSrLe9eHxxe
hpnxYW0toXJOgnltLVYwmzfVC3+p7s5vTY2AhwLgcdHUGVc9zMeJD977t+viDNLukfkHzbG48X+j
/1Kq+Z6b94RsO77ooN0J2gfoVojK/U+xFpDYubRjlGPeBOzvQ1uxG0KwMa5U4wZYKcUiG7ojrsYG
bfX/6/ED/59UD2qs6mm0Xw/KR0igt53oyjyAjaTXRb+iFLAfel5Vewdi11jiygGnsYdaJNhGK8Dy
GUS3AGHsDf2NT6cxh/n7dnWiph1zboOvLK/HlF5DAl7IQ+PiNbTyzCMjwlMCpxofb3sSdww/P1jS
ZQ2qWyI9E+umLco2xqWKyrlQSKUgpwma5gPx16WjCemrywRl0R5GQ+1qZ/KeVeSKxPp2UeMsqlhJ
5XKMONfw0jTrwgEwOl2/sRIxn9t60Fih7NKGgNoDoO6R5O6gnubO2BEz8rQMnxNGAPP44v9zV6zi
0IRzkHU9b/OYaXAb4bPlr1ZG/wUldWHZT8ypqBjnb7v5IGuz4hAtkArIbdRYjGSFCuW2n8tVhzJ3
wZjlXkSnAQG77tIgWCVAlyDUiNPsfs4nKzTDLrcVmRkEAhrWU9RZ+JusPV0eG7lSYZcw1EldPLB7
EmoIgjJHyNtThy3hharqXmJ2L+ZVdne7W2HYVAxiwfOY/kApq8pVH3nLqjXiYaKgnYW3TtQ11qiI
6hDVmACX01U78loZllEfvwEe2DrNRdK2HAVHhYrmdVS5Ri5aBrJPm/zkKq+O6gpzchbiz5auw69P
oux35xC1vT1nHCIm0UdZv+AVJkLTgusqpYP7tnaegjtFDLpT4IKJ1E1M5quznlfRnGE5F19Pdni2
TRc4CPkQcarDZTTa9SVokaa7p2JECRUWfZWzyeWIYRjG8PT7aX9EDkKVA+s7/d0mJiBrUAVppx5i
P7wceMEoes29R2jdQwYXfua2HrRfGuEgzSZjjt5pKHbZTdtyVs00huGHqs+bgHpfMJcfnK6PtZ3j
bZB1eVSOJJkGVMt+Xq6UHkESGfXy1gKBu0aQoNCYEJBn8X65jbGZKNqHuqg0QpRVhA+/E/DbQeXg
qiRHdw0TAsnW9bq8sHnmiOXvgd/sH0g4/TlnVkIKH8HUbZbqVJoADGJuPQZEmfxdaUltpGW+JZU7
thWkP8KJ2BSktxu+qm72KPA2/PTRBDc/TQgQ9nO3K+LUpbeMGhK7pBkbASBkI0dK1bTc23HjfV17
VET9YvEpuU/oyKk9853H9HkhyESlFgQ/zDow722Q4x0GZl0hZ2hnFXb/7HB7meh4N3MxmMtkEm86
cVhpkecnHkXbgxYmoctgzkIlZpASFFdFB/ZEuOWM5szsdLABpIw2QX2Y7QL/pa4NbTjJ5borUECy
+RimXKhzsg1Dw9tHt0xyOLVjcTCuRXCq6tRdis+0y7sIoGTPKEa8F5L1v116hBXGtMpct5NhpJMT
7SvoeBwH/eaSY4oYPZpgc0Vah2M+DfkDgjtMRBIi3berCTPPzyYkoflpQNsPexSMOOWNLeWuexLE
B6eaOCTOjJ4o+W0qgLpNLke10KzqJZWZa5jnzieMlvF8IlGn6I6JsySEH0cEY3YIX4E/ekeD8VsB
XtBcuU+huLVpjjzKbk8g1tBE8rd/pTNF6SoGdA4cB6dxoxYPzW4jbwX3Q0OVMCxeojKgwVDt/Vbm
g+lZ7QGgNSnNprPaotdkt8FVZEI6bWM+4ied8cQsdcjZOZ02Wmjuj/TEhA95mJDbTlBT3LaWURwj
TTwsVrvkzaX29eXWOMikdbNAgLAR4U9FosX6XT1e/OMDiuSEjdXeHjdqdOkvTfcZQY93kvwnD/Qj
Sbu/AIXlKpm+tzvwfAhe1MlzivO7iFaGFjPdvH9kjjkaVtI3K+57CxgctnyFJQGLFx4nNxtDMB3J
KEjBUO8EVjwhomfNpHvarrHut7TwxFmsmWjAa+/P+QUj9svLd/laCK6qZkXmu5rU9vF1p8b0l/Mr
QoNGnh9fhHxZsbu1l2ShV+NZ4ihUfetEd6Y4rDGi0gP4jzK2eoNnXKrTHIn2i2/nQ/85JXsAAVl5
lpICtp7cqCS3Ut60gNQmtZW6p+JtweZhYmJqu/lM6s6GERgC/xbc6RmxIyhgwbSs8wP6FxPrLhld
rXvNVbzDNhQJBfk6aa4gIbkTy3cDLoM+qAeaG4wxiyaHF1b//eKB2b4rQirqM9vNyaD7gqLwwpQG
EdU5LPDy5///5MqwwCKGOT9ByGr54FDMy9B7XjQavnYJxNe9M5DHCUVrtaS5H9jeR0OrLq5ZF9b0
jW3Lk9vHWbGiKRN2IMi9qvhryOUjmfiXMHNzBbu+5RXs+FMJ1us0DNjEDewXMQa63h5nbRvos2XH
GK/XlYmKIlFuwV4ZNYN41Uy7FDaTmEi6n103XfXzf/5v558kgP/OlAffsnCrfRa4ak5GeCDW45X+
d8NHHbWEVLP3v/KfnAhi9ZIVpFfi8KlY8R9n4e4ovNmduZ03rC05DGwRBuzTdHIsbiwdf0kPyI8t
Hv2zzcxDq6xs1f9KLNsGkJ+yDlxaqZxGhlevPUYWz/ryJd1vK/PjzHhlNo04DhwQxyef/NYfPdDx
R3BI56svgdY9zEc+6AcQ0kzqsTsNlJQwY3OB6HSGQf+gGeXLnf6Pek4xZeI9U7/heQaoWI5hR5Ur
o+NgNAsuxIYXC3QJRVdklsvx/afSJpKQQuTCUEpwsynwpWdnLglwl4+eGAzQpCHa6yWQHHCqOpSB
kdehwTIQdnS6AuB3vOGnVTCsRbVKsHD0DtkZ8IiT2fEjzT+K4gC10DbZFCHZ0ltpKbLJ5lF0hEti
AggC5+2Zw809LXzWU/tYktZ5J1bty6xfZNQ0oye1l3YSGzVKmlcZjfTs4UdM8c+u+TFiVy0QeeDy
zeSWTi/7VS0uiZcBmDRQKuOblZ3Vk5sPdeet3AKyv4RYzGFCbkFhT36a6oHwLu9aWVWhmZq0cLMG
6YOj4cFoFj4CwoHI/5TPLI2OeYqR0HL8mj/2I0JjlJqTg+1sL6blaAjxIidlSm52TJCbMkKl4FXu
985vxYElZ88EIKSHTgo8FQOfHtyb6tBMEMmEEnrdIeDLaCHsOLFtyuT0ZMh9P4o33mljLNtcAfnO
E6pMT0RnFFh3PaE/vTKStqKsGV4RJ34/hLBAQwsTYrV8WMxstMi5zaNIKE56f1bmMLdthqFbbIYY
32e84sLA5vxRVPuqZpLYXZetUvvADt0FhVJnILmhDD/UuGtVW6yJsGkv/OA/qspUu7zBrnOSlPvu
oGmD8rZfAKBjvg/HrIRnxsEa8qx6pRL/YUTQtU2YtYWSigISyvQp2jzOG7tvcO1grQMDCmDqxEaH
HlNtaATJKztv++91mM+ecYqSMYrNGO0UFdbD5gM3BOcCrXMuCAwBtMuLsKY7lmFsE2UdmLVVcAys
n+DO3JInq9rRMriomx5b9fsaCbDONTb0kZWNz9kOSu92mmV4c7zP83LvtKbSnoPh33iMwlT5X2DF
9WduEBwX3JbxPzp46R8hdae6Lu48Q8TQlWWf7H7AI9z0OMKB54QF99xoi6xwDTFNELkXx3VipOaB
OBtYNkRysEfCkIqmP1/J+ggpD4UCE+O9erlgxerdg+kPWbwtTo0nh6SWMIdvpwGUz9W997u+pkLS
vi1SoO4s6K21KLAUZF5NgYhT309RHGPBvUZNk9xGV/RnBdCCDGrYIenqUaMng7jKSEkfkA4NoEj4
UunTXOD1hJi2NZETi5jM4jp5ynEhoW5YIT07/8ffs0KLKPGlLsQUAtlBcRbj4pQdLeaRj1vffXoe
C8SeHC75si8qeMhk2dcL+4s4T+Ehurest7AzDmOMV0dVW/R/bEyLNDpgnkwTxUbCj0bvExHP1qX3
xWelzIVXTDfgJ2SwiOoeTcYPeDZvvpo8qZYSu9Y4xmEp8EQG39zyVU74IcOCHFE/huu7N2/2j7Jg
k5ieOrmlN4/ZN9DmPGCfsskrBtKQSIvc5jgD6vEmTHnAVv+A654+SVuCXknKXhcnPc1eqEPtPIhB
yDLrAmtQ8nNloc2JJwZCMUu08QB9aDhVyzgeYBsRGaO4BiHCOegerQNQTky0A6CAldK64nGgk9bU
URdjBnroxtwwsxMmwyjQRfJmrsyRbaL1FMdM8+hm81ArHHddJ51r4EZWLZ+20fGadgUxAp2tbLsl
CN/QlFAmf+RZb+d5cGA65dOkYF6RNp80dhIj5yfKHu23PCAQyGnCQTylzaIsMjUmAq2r13hXu++6
m8sLNezsIPNYsJmcHm58HSMIuzJVORpxHj90nZoxrhAe3fymcQIf8m1CbPWVGQyQDjgF+j/JvsZy
/4YW5cQ2ijRj+6VH/VXAxtfkMK+xhxTo1IWOwwv898BBh3oMI0MPvDrno0hToEYOCtMTw2RwtAEu
waG7z7Y567G3cWZTH0kQPJbxSVmd7B7aYIEE9gkW41sbKZWY6pOSMTv93QWqz+L8riauUjZPKyyC
pzvuMC3Wb1ZN+qkkIC0X62ydniAjCnc8o0WNgxp83d0dfpUbDYS3QNH4s8mRR5zNzaKCry8Ku92n
4q5zBfTlwmLSzSm94KU7zAXntt0Hq4jjTUdhFG895VD+id7qO1E8MbqmuP9mMTbW8T6u5ypKHume
GnYf6DqQ/r5CUcjD6n3DcLZ322bgQkT8i4HN+A9zyNXjiw9qFRtambgpi+WSO9rEnHDSqiLhIt04
Iw61O3473TDWEYlJ8/iH7Vw6LHIjYmbRQBpAAGQe2Cc1c1KTirjEm7XJcAfbHdSzCipS4pReVP+x
nweiZiNp8Sj7fpSyhYPGVH0v0pWJBOBr2qcK9etdz3UqmQwzOlNiPAM0pauYL5CinGBUWhDaH7RJ
uvQC4RXzKmnP6SNx4BmC5S6x41VxsLubdPiD+ruoigPT7CrmT/tr3zmDj7DqJAAlkcV/VlDv9WMv
K0kg96MhLfsaWoLv4VVdmnB591jGQHd1X6oYilFq8yPeGAOHxTNbZAU6OV+Y/7RQuyYU8kOzl7lT
txjtwo8+wbQ3fADG96KsoqVPfna/ZPKOvbgUjBzqeYO1ZJtFUg+XQTYs+5vZF2VGHQP5wP/GYM0K
XdMiaGDdkRWXhjA7L/GasvTDjZDf/ae8MU6MObwZtCjscCaGokQshfP4FvAPPi5yniwKMiV/NV0u
PUBzLMoNI8HfjrABmdcH9N2Wrme8qH05LfcqM7W9DWv3yuhFn/L6a3d4oBmBTF913Ix+3OxEdhEA
mMu6G1V+uMbwu77CJwnrhiitABLTzwvl/BpwF0tYq0mqiUBu6KGuJpCBjXkFsR+1vsbBB1UAWtwJ
2sCGvV8YtCX24kVJ68oA+CwlHrI2OGxGa8dlQmrbKTc+xM1JuYU2C1m7Qid20hrONvyX1dDf34QX
kuKW+tSp2J3OleziVH8Bubgbxu+3HU8vcpCNGB2D0yY+5ZqORjM2CYLo1INarGdChhXrFZY7hMVv
2trHB21jhiECbpYm5FErC0Ms6iojPIqUvBqI6qgo3JY6PKHG+JZRPPN9PaPMsVFezEGMc1Yq/hAJ
88agXkhUq862s8w1wQkee7QjDtNHZemxdbzaBn22MjDrtOCOKLbHzl9qXH5ysMi8R0g0QfDPFL0M
hw5peFpMLAA0t3HwkXnYmd2j2EOYLTF832h6DQ3VogWHsbYHjnGIdpM30dxwr7YEg/wtFv8Z1IeT
ntnxnlB/qYFvPUodUOn2hQsFSQDbjQogxbWQ3bDzMWG9/PSjlc+7161gnP1IDPcjRhSuo3dKeF8H
7hkGcZ3t4WL0estnNFCpbf7uYUv6xEjvKMoYc5c5OLgC936tUG7J5ZAExMQJhjPGE/oq+QXHXa2C
ajeqX23hmkr81Osu0HLwLrQcTjjbIw8/UQzIq1eXErFVL+UPEnVm8ot1Xw364WsIYxf0juRzQlQh
75BF9UTvNbcebFn0KxQFLyjKhwrbbBmFKUO+J97unMu0andXDNM/gmslsbAR1fAW4P1D5C0JYdy+
ghpPOHKdGMulb3krg+D09C3rJl9/itIAlobCwZjAcYNmaFUYOuS1tT4gXIU0YrLKd5tliVOspB+n
3kB92cyEhMMlXwMj2rSCNCLmvHJPufFyrZ/aHTuMqB0ijZz10p6+Rlt4At4PQDBuHNrJfGxP1spw
ZoyXqbebLKbdqv4QzCgqvV6bp3xgqROVI6b5Eh/QeYLsfI3b9KpJrStTPj4cmO0ebgWaHwfS/ZwY
XgtkUY/9ZFG849J8HOIg6ly6WyHe5qSOBiUY/ERP9IdkVEMNDYedaNFtpPu9+HviicflVuI+76++
SEFGbo1Xn1Fk/Z8wGLiQtTrVK71kAIlG8pD7IZ2vjSAWiV4KI46k5bAsYWKMYeYudp6JYLxLTPqU
S2raZc8weTx/ZZb1IGmyN7APRxjO1EmRJll1zhQnmIaKbSFjn02Vk7lWT2RuwGvygPohdwdP/zcU
OSNEfigus7rg4MxPRzx3fZqDhpW5P5IxV6aBhm+h9pKCR9XP6UQ0MbFxJZwcngIzKa63IET53oEx
YhyW1qvmaxICM8NJ2cecsKU/2JeO8+0bfyJr5/YDQKHocwG9OL18JkmLhhJEiVWmNr8HJjg0qy6J
JDDRMmDLblwtav8WTc2Z8gze2HfG6AilcqcSq7QL/dBKWE15xy4lZQTv+eGO4Bph4v/Kf9DobaUi
v1qfh0XGPGjq4zf2oGLwx1Jf8eDC6VQiSMGDc/EMzAdPjyXz8km/wUM3G9KDDT8j5p0N1MM6JeZE
UP5AfiJPflqAuL/g0NBA4ZLnO6muofaUJHpKkojLWj0PDs57unMZjCFfcLxLP9uYrLVJ/tlE+KCP
mcgKhe/nbmXnKEumCO+Jou4WxD0ER5MD5qifsWPY2VTZLAmhO6rk6kAivVzekwHUsEqqgi7cZPtz
w5pq0wt90Cp0vxZpNwTx2/8MWRJqxAO9+ZlknCX+Ad1S/Fov+O/8uy5UgpYdtVC4Xqovs/Q7nauH
mL7gVaokP30ARpgy0fvamidOifsSK4weOeersN3lOuMAO5PStC8I37JA2ROXePCvjH3i5mit2EOY
abdQxAoD+Muv8vAw9a0vcY5muCQYpt+MeJ/gVOwOwwd4F3LbHhCLoCdBFnq2XUrPTz1Rxs1ODoHC
JaoaEsYCgpjAgSttvEH3N7ReWpXXHLPs5kUfO+lcaKOMGrMWlEj6mwfJTsy4j/7ZEUM5xQxbtPDf
b+ImhWn/Rr+5lzYxjHCVMmC2bg4kSTzz4/OTu062RLcXDJFampkd5uu35iXfPrwo92Kuo49x7iqn
HOeOQS7Fo4CPAkgCFsAI0bkYlb6xDbLLlesnaoNPqmYeyPHw2wd90h0yK9H/dxD43no10Z3xD3mP
V/BK3zfxKq0dEDXxssPwMjwEEORIVbx4eTsr+3ftor8w2fwxh9WwjzYhHJX0bunU4aZu2tWWhpwa
8s5aGFufomvl6ABHsN8thq9bnCeCRWaQiZy06Doe5ww7x60d7ROY+T+AFCeVCjFDwCcETPAsaRb2
dpbfwb3BCrhuaocEMV2c9+oor/iys1UvpWmjlyESgV4ZBLfrqwtmOSF0Lt220yjyMuh8mkvrl7s0
mptGfISJOItV37sLRUHhuiM8rBDttE2qTzJCKq8Fkb9U54bOCZqsSfMGY+1EbtHQ/+QTUf7VZHMy
LgrZhCps9d1Gi5i8Ye06f3IpOZ0xP+1vVs/o2oX3y4z7RKM/LE6OpOf6yfkttDie78LUuOYZYsv0
V+rxYZPhLIS6iqJvpK8sDC2y8cQlVDBnSsx86CBMpAsYyEkaifnrVUbWYMPFN9SA9VFCzr8QfqBS
oOAgvHU97k+OYowbhs8RjHD4mlEsSIV8B59SRkS7EL1IjyA8GVqH5dqPB461ycaAZ4MEiFrEPNpn
yc0QL8C9NaBBCJL+kx4wG+1b6Rp6xwbm9TG0elM3NoGYztAO+EFGRkrcuVYQrnvqjNmaWuuChnHj
Aj/k11LmOwhFop8grnDXaq7G4wIqDPu8CUDikFBXqzSdSBF+bxxnbKnEVvS2XBVwWhweR7RNSiqm
H+T/MGHfnsM7pIH1nknmXOCw6CMrPgkpLBcRdpqUynYtJGCJbcxt+H8kg+exLHQwlt4g/leGmmcP
z42UININJx9vFKGJwzQMcc3cNDAo5c6bm4oDHVh0xsiRd/3UlNCVlqcZHFz0MPKzi545+y8AJ/Ku
Ilc1OZNNQS+YNb89sv1nkHI7qd+YiGuODyLgR12mhdytwR6ldtpd/AmnmmV8pHCknyhG+Qyw3onm
EHYmH/XmUQp1Oh4LHGrKM23nLC17tE3MWVa7xuW18TsdwSzpJEIPl2/szdyuguu5IRzWBm/Kmf5b
QkaAtMTAfjLU77PJvYq5WdOu+yqpCNqeC0phHgKfI+BNx4eaPPKE/1Pf5o4rNdZ9D41s3/s/vccW
Ra6tgY7CyOyv4tWqfWruIxfztBZ3MI9h/8lvEwEzzAiVAgFkwpZ4dK74L9GgsD5slsE0q+T3rkdW
x8uPQwHbcd6nbmkub0Wgjugr83zJ4zTFQaRXn+O86Ouq358zsU4E9RaDFoxddzu6h4tiuoZVs1TO
NjZBNIz58evv7U4nEJM+YtbVzb7Iv3CUb5obJzKgE5q89pQnr/jbuUV5aQMzvhsKGMkNBf5QEFZE
M4NAx1JFwZTKghebJIPjZsF9zE4/SLYtWshgEzYh6zxO78N2zOyYRFZxLcwvGWezIqkMzZD03gY7
I0DYrGUb0FJa4Yo0kLC08atPfeXH/AUYSqAsGmaiROprE7+p+xp9v8TyArEDkpFwPb3FJwqqxCA5
Eoui9YPoPt9l//aFSlZG9k/kkJQtCXLr3V6YdfFA/rBmdotGT+UmMg4G7c8KvDTUobmRwCKSikuD
odEVuGP6d/1YBk7qzQvmzuohbLLYJ23mY20FeT1NkZQnGyjpt9zeDA+U5ZLsz4UBJ0OLrjZ++CTm
KBFK+6XR27dNXs2LTLrKKQKb7VivL0oq4dq9CcTALp+p2jVyZAqJcWEmL4tjfxT3VNAJkxLQES1p
iORkP12O8ccTPvYdVr4YViIu6BoIrEZFWiW34xSmE88CD3btOgE9jM05+WSgoiq96afrlUnC2bfL
NvD0SNnUotE1ipheySrTd/V667UfKnfn+cr9B4UDTDHZTNgoKpmlSic+UE+3w8ztyDRqxJEPwszC
CsoWlit02QlW+pXMFbfEMY10nhNOk2sho+FuEh0yqDlydz885fh2eD7zM8Gdb1/jZ7Q2yTu/pjnd
a6yX8schjvsmP9gRG5dZVEOH5YZn/SeMudMv01hghWAz+0L/zdZTWx5LUN9Hpr/I+lyf/B5RWlvJ
d2wQ3ETvPawmMPWTWLKMXV0TkG+4oTuXOwHb6uRFLAJm2Z71eSqqjYLfDyKBu+VtZ7xr6tGFa5Wu
paQ2QvJzeft/FPQLiQvNe0kJJTSdfr4DvzBgEUUf44Fkjj3EzOaKYGRp8XeukxLSXBDPAAbrmwGx
MJ7rA4r2o/q9iz7HBEojUlh4yHpALKXIFfmKTp7YZ6VpKbmsEicZGpCAHM4Nu4+YMzu6QUV08228
Ost+XZ/A0Y18gj9wWkTVLap+t/IktJQMRHfGSKXJvq/SA7RD7IIMo36KQ6+8U0AE5AAYihNlmEkQ
iDuVQbpk/E3CrbCrDM5e7gDxWQglrsfccBcouuv5FuIhz4dwYV4ukfIrk4ru4YYyixoQYMhdzMer
IXlEcODpns//xExwK9n/8qVDeYdRlKnaPHehEkxmKxvSGKjeXLCs9X6JRDme/YKKHQw84HJGy4jW
rlyKwScJAmPSHE8gQJiqLcnI4qmGW08dVmmSF242cGD3DQIYQt7eLf48DIQVwi3mx8S8IYJReIGq
OyBrq1G1PXuFdZZHiV+jt3WFdIoyhqovJhnFLJZwjN4CKa/bgJIwaQivescUwSg4jUHdx9ubf3Px
+IA4D0DDXg0iiBB3wWlvAiUztTmWj7cuGy4tb6CqLnGK9uGtL2d3KwFMPbCXipvwBQBvkAkUfS07
aDc3DEKQSjO6IdP0NOhpObgIsvpi+n1O/UJUwKg+M9tsQvYVETBLvgQ3Go+leZiqkTgVLZEzurFg
j8GoudqYxkMa4lRi0RHnUYpBK7C2FuF/GoZtvOiNCa1hrJDkt/cQTAnyza50PLStP051dHN51dhw
+IyYd6kMGw54BJqX9hj3qHOQ72TljWwshluU/dZ9J+uZjaR5nfAKgztAaStHfFFMNyq5JALoehU7
8gPUGkFXvcj4K6yWpjravQEed/VayMzzYmnRYak9qPNKHybVuv1TLDCeCuqMOXEOoN2VcOkonMqo
kc1iOLw4vDxxuq5882FggxMLGoLOlB1nvVLGhW17cGmzmJAB12d4jjGjHxybMfyOjFfiKSd+ZFBr
9Os9Hw3rIHhJI/0eGKcXGlF2acCZyVvdYqBcKgs+L4JfzUSK2CMlmk6ilDEqp5hY1VWibqTZhslO
U4FETd8e2L9FA76bMfxzsD6XGe+TxFraxnZCEWiz8E24lUeSUHUWqlHbnZDkfXrSqQSJ/iXZq1OW
D2nXlFSn0oB8W2fnR2v+u4MaAhS2qSJO/oM4dqWApDfcN6i4N2R9dsL01jjtCuu6CbSb2ot9BDhZ
Z8ad9R1iEMCOQK1lcYBbVOKKJkiCtPgLWjbYLX+dcnIJXq9nE3C4DLb3icxacry6MRZdSJJfBtSe
ACxq3dg3ixFihgh5y4nY/Mzp6AgxHd7/Dmwn9I5I0x5TGq2SlUtr7OVeKmLzoDPFEdUU0rzzMwKj
0eF4fD5ceNAcFrfJUtT1Io73ce61ORnKlOYpQ6dLpDqmBdSpJw4iSijTpND5KDfsm2z3flhT29cG
UeiqvwgSiopbZxUBP0zQvsbUNe9jUiGUdv3o67GCMwopQGSJ5MONq2FvPRrefqZIChYpFPZXmPyM
HYA8StVpUKdzfDLIDmezQTGS1aerWbAqbGHxsRLrVmtk6kkF8+9Ec7M6aIXQl8SPwdvOXx1tJaWj
EpemqReLBtYpmQO7+il7dnAfhMujckuQIdYSib3j5sONcaEX95bHRbP5SXw8Pq0C5Mn8bM0U/nFZ
rPWi9UZnbkiefkHZmm4pI4T+DvA9LNltWg7NvCDr5iQd5HzXDNvUmLI8+3HxN86B9DuQ2McItTvW
gz+WPSbJq8OMuhXDXQSlWByJTlvk6+5+284J7y2SculKLoe/0usXiU/gETPq3nNSMWuhRgI/8Rf6
XCXvln2/K3xn5CB2WcWW/2Z+EEqHZeD8xNXoBY7G7Vkh3t1OYlBHIdO4HjJ9/QCKumji5YUAMPJb
E9kXDpGQGA9Gm1NQaDBXuRS37M+6ckP1u4cD4VF06NPVNXseF3aHpY6a+wAcs9bLPJ5HZyyyH9Xg
72DYExsRewphpkKnYO11ieKpRUURDE1U7IBRR+kwkHno3l1/+T9zvTvE7ub1HgQexDrywZSGm184
a8UnfvLRTmL2sqrrd4UN1Y5O4ByzidVJgnNCdiq59FnHwq1GnK3MU1Dmlesl3MOIyLP/NcXHKS3G
auRAMl2w8vdP8v9JSwMQ6fvLs8bi721C7dXgMLIkGglZ6qC0UPWQrS/5kEK2jvBgtJymIFrO9Frl
BKZJyUg1v82Wj3/WxOIV1MTmE2i6RRYgi8EZD1J2n91O823EPlz3Bzpk+ROo8oq544hlkzIBTpuy
LBeCSx1YipCcLP+57esTqsAzb2wu8ay0bzUL64CP24nlZ0+LNq44Q7e4C9MfGxnlXpOGf/thzLpq
YmmLTsMChpxVhQVdO9rMDTj+1IjYgWXK9ESKevtxQq3uDaotvMptv1qOgfLvG7gfqx/6JXcPduEJ
ihAcs5NidFgHdwEBv3uroubUPeFkQh7+x0plMls56gyJftToNoGjX+q6AxAhZP+yRHUBoj54P0Tg
Unp3p1uByd8/7z30BM2c64Uu9E3KlEmsAtKLPtMKxv5kNbElaARWzaGKJUu5GVTPb39NKegMyGAN
NEn9ARtSqfk3awB1CpD2JoaQrYVr4hi142J6xOtzgXRLzCnzNaLZ3DDY3CGKSJLrNjqYftROKIkQ
rKy7AcgzxlOkiJUDXzubb7kmBsguh6Sw5Xn/orosbpH3V+ttlWkYyHDL4qBwDZIK2jL63jkEKEg2
7MThzz9DVYSoToY0Hz1eo+MoIrcMeAxOqRSrFJsgLxZex4OKNaicLjTay/nAYwuum+79ir59rwEC
94Wx4iTRNso2BAggLDpmlBy7Yv1/X94hsc6NcswKQqS5FSMtpJuSOBgLHRrTN5cOR25mjUE6OHFe
UWAQQ2hK5mlXoAZdgiWfKXhZgLao40n97N8YbfUGjkrsaiiMDBEXh9/sRHFywXF9KHccNXydlx/l
NZdpnjDK019x/WRJvLTb/wiLIsZczyfBM6ATSc1dsA2KE114S8vzpA3tvzkCG/EJtUxCDygY5fEK
7AMvHFUe9/nIARtGCUOBBTOHb+g1DUH/ClcWs1sH+fR85WLU8iiMROz8C5ya/d6uYovm9gEwsWqj
S4uyzjhSeC0rHjWn5lXsks5pTQfn/zpSWpNVSs537Xe10PBja4JuKK4hw/FJZJq5IIz8ah6UASy+
2UD3vmkWOnuqTxtYDLEPZcgyyXq7i+gotDwaKWMFyT4zt/UMGmq4b/30CaqDu/FPBNp8Q9LFSLl5
KIr1QBVSHBlQcACnPVVsicW7uEMGa26m6TqKcFK63fkVFDzF6RFjkGmLVc8D3Glp5UJkQA7/5ffD
O3Yqw/wc3bZ61irL32oyUtvYwNpvFd58yWIk4FhcV9ZraouGpq44UTVY5fBksTMbsdbIbHnuIafH
nLcwdADd6DT25rvtlD3tFPjaK/WuRDeUBR8ZlNdZJ3FahJmvH/EQn4f1JEW8UMLl0z62njFczsW5
gwnEFsFadAslFY9JWXzFQ31514nu4CrD/MZ/TPteRT1S81kURAHbOpZpyVlKFtzy/5+FclhQfqt2
8eH5HpMc0O3xZFPiojvxTa5L5hpSRRwMWWG+8OfIbEeIlbqVEJGxdVvysUPMFwTGFeNC5clyNqU6
QVVxOMilZFtriPqmXBLWQG32qFuJNQUBoENPQmysu8oG5nUzbGfc8kWopws/byDbO7n96d2ZaWU4
gVpHfmBNnYzKSLC+JS1WFiML0+lSthrTLwS6uoUoQGTwOde+MBEpcdjr4oW1XgSFHoxAB6hvoI7L
LhSlGdu5uqWS7lESYYQeCYWX8sy/NTkV9bGuTUeMa10pfbYix3PEmwOm2HUb06/zGeI0+4BjnZ96
uKm0NRuUX+KEmJlVCA0xV9PhJiEwGLFGj8acpcplX1qiLlfABwtt2tyNC3LAovPMHg7mg/PvoyTW
eFwS1ZtFbPmOO5WYHxUslLNFrcU+yfWjDK6huL2n2trcLOw2aGUtm++Ws+QFztYfdzYTvvbviiPO
9jcZnf9WiqzAU3iyMYbJ2Nw/ujVVuSUdaZPtA3ZtM6H5oykbK1mPDCy1GDHJbrTYNXei/6hWMeEb
tZDzbFj5a2z/QzVcq6La3LxnWQPbMNPg7xmMoH9EoQ40sPAOsm5G+Z7li8N0vS67Bnrz7yNsRlo/
XD6QR9gIBaD7UPaXxCDPLdwSm/7uaOyAvWEGrPbXXxrJfJ5weBpi8XjxOeFQ0GIB8OL/my7tiism
WDRt0cBSI6OXZApCjL4SBa2qpUOziOtsw4oNqway1IRQVaBk/3wZ6D+bdHfRwFMZtiBbGnS2Gy1n
ZXvf/QU1J8cpscr2Riv6hh4Txv4FQFVCt7IyhkFaXA79crapJiBF/6j8CbWsps/VvnRjeYIUeVzg
OcejaVhTmSjcDSmq74mGhFnoM+WVtnOdZ2kmKIjoTzxFPhrszO+K0bToT25q8FRi3IDKHZnIJfON
jHAkzp/zRxvZjR4Dxns8j9gfDtxLbcJEjpOiqukWp6H3ydUp52hLSsjwyCYTMDzje6HPCsF2f4XM
clYL0owxAsgLFyKXp8kBDP1+94z6KtYSD6ycRBtyCjYmPf0BNcz0c3ndUynQDFARxiEVuzDyjW89
t5BkmX5c+RCPQpCdF3ZRq/NrrMRdEQ1R6XKSQVtOK4TuPMT9dHnuMHuWpY0+UO8NX/bvMaqI2zLQ
mcqUBRjFEWsq9pya3S+Ff2EWARpWyNk38OLruMPYzC65Vg2VwNgkZIJkYXdjIQ5Aqhqg6M997LUd
TMpBNcDGYQsfEBQR7pusZaFl1+/JFUx3nrKVnvUsNRX6u2etl0pos44dKW03wyOl4SotLcYNO/aL
kLOsR5G4l6NA7fdeIaE5ri+jIzVzF/6/NhN1z7qtSRVLtJkpVqmEOHQcK1zn6qeUDED1GrCpahT6
8ngzmH9vzWLVOxsd0wSf5qmaZFlBenkRtypmCwHQ1JgsWM+dJam0GTKBUZkkjV0VjBTZBTKaiuP+
EcpCBBKv5Kfaw0XvEW4+6wHrWwYdhU9rIBeB6qso0CnLOPs+fv5Y0MkG9Kht7UZUBGz0/SR2jwtj
lv9oSnVguL+VNWzxTtIf99HXDM/PheNPL3O4K+q7bSCj7YzOJKmmP+wl9VjmGFIk1TAuTX5NQg/0
6Act/e1OGNH7k/Zpg+zxWGSOxBCghD3hPFCwH79d86F5pWgl92SB6LR0enZsqGhs9k40oi75IK7K
RCTASQGjeR6sDTRopOoVoXqmoNAHkPKwdbGjMJY4xpGEkkBN6ekE6bK709ajS/se1Hq5iNXgdCWe
Up2ZcSpLZcsGp2lDPAlMmBi6HB7VAcSpdKqltju5KobFq2gI/ELiFy2OxSD7AeOKL7DMtyuSEBBW
Gb86BKfg1pP4215SsPN7loL401qbEuyLPmF6sCX0Ru/cUkYdZUHoLHu4jr6B1OOAvsC0FkCW4fRz
L6r2iTB1Ji61ETFB9MTI3svmQzlIXWg8V5XzVZzAJryY6h+MuMkQ9eFseSUXXIVY/F3Ha8SjfNF6
fpkNg1ST0sp7e1pJTktt77/Ywn9ePstQldQQha3Thvg5RzU9SJdn+9n5a77053mCUpcDdivKCRJX
/qcy3XDj5e8Ww1e9Ai4JjV/Sx0DUYlTiBwKTLO/HwRkFcBLvEl77/bOmctRKz4OTi3YdL9+003H6
8DaeqSbId843CIU3fw8OrdSiOen9RXX8VHip8cXm6iXK13OZ4W3QNhfsx0/fsU7KirZ0uFq9k/AC
hD6OL1sJeYr+xe4psye6wGqsw1k1XtCVqrRzERufdxu7VisAKO70PON1PLx6IYfZHGU9306k1dq+
vUEpTXgrEClSqKy2wiMd8E76Wtl50KCfeVKyJP4Fbu3sgrLIOIlKlCROVacH9TwvPZ6+6GFwAbnQ
kvZLpPcxqIkrB6U9/qjVGel4uESoDwzdWa63NwSlqNNOrEaUfxtx/UXpeto6jZtE988HvT3v22W3
WyF7zJT5+KzXRuhVlgJjHZqEjNMbwSnqELNbSsP0KRXi5vI1vM1FkuBKosi7sMRbRio/HoNOm8sk
5p0QUwXI5EfxocZy7QS1RcjMr3fafbOG7PrRN0j+9vpFY5ZXBtXXExIHiLyb8cx5jPvQF7kWT6Mc
3IyoLhj94l5LVJFG1meaQ9dU5mi0ORuabW6LzBgo5QyCICgTDJ8E3pk77XBVmMu0PtKqCIkmwIZK
2p2Y0wgNKlfhlDHn2wlsO62upscc5CwrW4WAXdb6OuKZ8rLsQLcb9q2MpNNZB817tNO4L/W8WZdO
KWEXg0v4QVgS2wcE2wa8i/Q7hsnZ4CclEBFs//9yu/9KCqsretcbL2ouYMrAEUjgqKfkaHuqFh0x
5CpzA+C+C/xYocunOdj/R8Yo82yFW+C0OSUMaXCS+PTOjYDA50uSh1GWJUFM0c1sI+8HGiOXkPUj
OeEcvSeFZUPypDzxNVlS43vW4ZWDdKOQozqgRXAiK/rW+CvDnMdC7e07PMdoUpAqvSwOrLso9CB4
QO4rsCHBJKz0E2Aq80V4vWAyeNKo6oRETcDFY4Xhs/IJnLhQxe0TbFuiggO5PhHTWCIZzppIPtmN
oJHAAmCV1sVf3M08V3BYVm6iUP15j3OmFGy/0v0g1KmlkA8i6IiccMChegwclPclikkvlzjeIRmW
16Sw4T49hsKC+XfZTUpXwkhHzW7WjF4TY4v+wd+kNEbPI61fN/YpZVdO6DfSiXRDQtkcyLfwcSh7
smWTCfdxtXoZODD5q25l0e0xC761tchtrNRnRQVDCe8XI640RdMsgUCgCaIdRymwaYDSnOxbD/zN
ezelu/JHCX9bHbyJDC5ZomYUE63XsRmWy4NxBj15b1ipRbOEbYhf2n3gHfBlSG/GYRWHrqPAYTkQ
QxFcTEew/k7DQ/OSTxTQHrI9iusL/yNnXAZlBdte8G/zwRryyIUzXW7zI56VCPCNDqqjgTCkT4+o
SVtPSlAlZrdRHQsLik5q0ATT47Mgm/+W4ccWZVz1eN3ReaoWUyCoz2blpe0a3rvbkrPZBUmMTrHL
CaUb4v1Lm3lTJ71NoiKLdmGrqUwWiUNWm1/hM8i31vuHSUZYG8983yoVYUz0fWcMJRmmeWrlt3X+
RWvZiyaZ1SIg77ZnYu3uVVghQZBm0v3KPcoM2WoBW9Gzeku9sHydAnG6EoOdQZAktIsqk7qcMo51
mq9QQ3cQi8KfFRhyPteJkCIC9pRwX0pHg8eNznAud0lLwFCXjQBWgCxIFytHKZt9WuHU3ZMhKv07
jZcS4vxkjTLQMjE9TQOkyQ8HDLMYHFsJlN7S2RXCG+iusJA5rnAINlFATqeBqaDvH2nnIIExEQnV
bEu2HpNKp38FL7w3GC6CaB0+8524U+tMalBQ2aQO3uytPuUn4uw9tjv+UvJUXw8fvIkNDpacMWrU
vceShhTNg22nTY6ddo414KPS3XS/jkiKu/G329ljvi9Pq408gOcTZBGg60xD0Wh4hA8DAFZ8n/jx
aGRg9F4PZEjZPEHJoTqUS5PXYwyugTv+lF0Vorz9mflwxlDUdKCzOHLrYXJPlXncE7ATX8j5MO9T
0V+oLgmnlUmQk7IliImUO1NRXMC6atcucFqidnNnVHpPzPBKexF2/cokpzsqUPgo7k/09T44ldyq
aZpw7/n1TvXs2Sa3cT0rzfmtB5a0qf8KKbH1HAkYOrbAJ0qyhS6U3yRjb/rTdxxRctFmpeSRlo2e
XODUP8jXtXeyDekP4t95L9qG5MmYIT2Jz2Z8P6UAYjSY4vp0yuqrgje/URDGuBra5wITjO1y4Qy+
gvCXrjry67wwayYLOYpRof4XAOu9Ovb0IU8rgYu+oxI9HSsrSDiiIRHMfFVNVim9YooM5cZQlghn
2zlD8OzYndkU1MR+eEhK0I4BZ0O5dgJvlNjWOVlNjPw3Jxqt/+hVzruoMqS8LBtrdcGcSWRoBpP5
7qLNQ2IaMXSW09uZEqr0QiV7ZIaSDUqPNMuvrLa7TXmtSM090W/r5nGGQ9dEyDC+d2s9bfTBToCn
bBpdX9d6y4PSlWeFsY8n6OpEo90S32gvxikprbiqAldSKUPQZgBjuQS/KRQiPMMr+FN2LwDBhL1v
7c5KGrldO9WDBmn9WGqFJyw/poYN2C10NB0flDdSHPHVtv+swMobTsUo2s1Exb1x2rR5cnRsqv5E
MFecV64kgxdvjU/tTlkEbz0fwyE3TVAQAOKNyQUxb+pEtWkNUKtSX5uVmBwsdv0JGyZVdsBV6I81
dbDKOxbi2hFuQymlmMkGemmLCXAEklFD3aj4VDlGeW/PE7TAZmJuHf+KwZfl+w/aYO6ZEW1gxrH1
EtODun/xCSrhTWlRr2HVM+hjUcWR2zv6q77awciuhG4PLH1+8bqKLnQOth6xqBvyBYPPtpyqorK/
UFSuBS4pkBx4FpBXbmHkvBjfmdMklI7dicZ/+wSPb0zYfHkRoUk0C3p75zgopj+9B7MfTKi9rbAf
1efse4Poj/1T9FVYC2r2J12WfeIk3O7RC0X+VxHy/iaSPsji56gJ7dAvk/wm6syGd70YGUAUOlRH
21MPzzg3A/+Oi/6qt0ktdAsepzwR+PRCS/9BCrHoeybLFxVCoJ9pFlNh2jsFaJgnGxdAEWcqOWjp
b4NDqysGDanhv5p44SWFk1f/LE8JX4LZBw1M062lXsfdIlgAYeTIAPPJOoPWzAQWW/Wvff697iZj
L6S6UPyJmlxRSok1nmR4FbeekS/TRUVNr3/XUV0P4UM0Wgu7YQnj1THoIy/oJiC4TT2ZzeqSUkG0
4FxerK3osEvthectrXfXchzMpTq+LJNKrFb8e1Iyc3iCGXlWtPSjKn4FDuMREhNXNUrPppP7/igM
SHgQsL/RmCnhJSmP32/LwMgVNu5wk/tvWSa9sBC/WrYSeCw20l1HlY3dvijZ4Prw/JpyGP25bU3+
K7SpVgrjhhMziRI/897CYSs14Izn6ogO/wLpoOyqgZ43/iXmoaBlX8d8kIuS6swKXR9HJjGK6h4Q
vQfgQLb2PGFWrPlfgmMqzO8OsOdCgSZNpMwpQZOWNoKj0GR0giaSWS2QQqYqiOuhsAwxoegcbfEb
1YiuCwhedl6VQxVLiXO3Msc5GsFANiepJDB+Yh6iB5pWcw7itYv42skvQyHdiVOsrnrw07d3tKM2
UIGpCmEFxGoSLoInbYrrBHFF8S1lbMrp6UnQuRczEkKhvj1+JjGq+olGA/ojbzl4lfwl1ImYpUMr
AeDiOQeyMTT2phpcr0pyASfz/Q1hLaWnaamRDTxfGicIe9rrbVQVpxuqzFR48mN7KqvNJ2LF8TSt
wCSI82tr9xT/EaQfP1V9+841nEm27e5LIpTogP1alsuUUX+H7+WxtU65pooP6DtHMEaSKnZIUpoY
V0MZx4o5In4nWrOUAHY46TMv4LcE6Fpd9D+T0LydHPfxK6MC4jQ26rOVV3Qu/SbKd7HYiKOU5y7m
3B2AAWTx6eiScQZnc4h4FcPLJvodLfukhBEiOzEeU5T5vNgUTfJTOuxBY2+eyvX9Syi9SOuL8yZ4
Z7yiwjBYIb/+VRbT+EGkTePdBnvVuWSa2AsrjTKCGTVGpjKo/EQkID/rCkRkLnPkdt06BRqUlMUp
qifIoyxUXkLxZuFn9pSw2TQXZqMo687n+U+V234RAg428hcp6eGnXqDmlzIs2YM4EQqHjUCa3zRP
lx45feMY2yZleuQ0xfZxKBbo/l64yJDRP9KIbRCr69Zzsc13oraFsrAcYvcNS06ci6kGvYamKlnp
PNrIapZGwamgVOOQeCwVECAEzu1Yif21GV9ioZJNnjy/L2kmJzZ+ZR8Gw0dlVR+YcvtayMI+gqjn
/hacTZH8DWK7oNUMkw9Ntj6IaTwLVFkHExj3iU9pZ93/ZKzfEbY9M9C4g/mSIzaJQcjP+l9h96LO
DVC55pVGXU62B5FxhOgmQREIvALyRMvg6aoX6sMPuPAqlJgY6Fol2LwP49lLmooOHKXEzqjoHiq8
kZFpUmyPfx3UpA/3PXDdO7Uc+BnO27XrODh8UkRjjXHR7dAjrqTpVNvHbydcbXvvP0JzlxEDiu5i
5qjruTKDu8+OI0NzYb7G0J1TWpv6MUDclfviuIRf0mms6l9LKceuARmSjsunCPOYUoVMo43/qWra
mhtlj3+NjJ4N+nh/rJswNNEKOp4jiW8qSV6RAxQCL/Dbcv/8hVoVP9IreCTpwiYt2FqHpBCyT2xA
LHowL+6TiDbCYLXMMV/M1iJZEHvN6sX7PrHkcW3AQVn81lMi+rcYcBLD5TUS3QvpUI1ULsiQN0SM
qgjw4Kcm1CRlJxoJsQFWtfpmifFzgtLSvTpX0VshzyHEOycpJn6i+qa9GepF1xRjlnMTH66s66gT
akl89cMTzODJSYlbE7QOVvJDbaLBgx8wCG8EuRyJSBMW7v8mYjSEdD9vvcU24AlLR42+VpUDMKhC
x0Ltv2oZ1yIvTUZAj2aHIaH7tLEpu+4cQyUx7t7DKXEGl74zw8pyZ5zJWAzHj3UvyK+3S1sqp3uP
j/UDmXEQ00qf7W0xuYthZ5G+lmmA5oixUxsKvkRTChqQsLeoiqx5as5RhBDU8n8yGb6Ft4yDipvz
iC1odZyWOJQ6HGJYm0v+0QJj1t+5oN0BNGbDO3RsHW+8CyllyXe3rsCVT5nwUB1vYrRrXTu4VphL
ffthtZbow2merYO5PjlFFtz4XET2dwpFcVqEIGFUAlyBi85nXB7I5cR1NU0sQnjmQ0kbJ+hgfEli
iyvNqqiMCLLX6fv74Zawgr4uSE9zBVr94q8PzN0eKnOcyLGjuiOpjp0QuVOeaGdER9xxOGxRXdUi
u/vu9KFiw2ch4H0myp2ZL/uaLkpzKZVP2HP6yxRGljge6BJF4vZwpS7rqWfqZIEFyYVwxyRn9G/X
DWvTFYad56pDoGWQDbldDvAk4WCiIUr4HNcd2KJwHFACddDZ1q6NeeE7fW4sf/FtIL0PoTdJpVQe
36mAJ818iQMFnvJYqlNFWqYVLSmsCnLDjqqUwjZnWzNUcDdDHNq2iCs5HNXDnxVDAWHwe9z4h2iY
Cn6eOUl6+m8+aSNwmCg6TemxQ2GYrFkst8vA7Ay2Lv2gYlC8wUAgUzs3eYQjZ+BHz8dpwxuwFED8
0G6eRWRIjIeomYFk0Jut5CZ5KjRp9M0YnA4lJ8yfVtMVReqefWnFD2W4YDvWlxU3esnhJCqPiAH3
rodX1LOfKqavoHDZeXN8x2CqZi7p36A0wBMF8eW75OiTLfqrcwHn33l8AyiaukZ31AiBbtust6SL
0EhJMZWzhIY35Ap/6REyoP6wKDQhCQRkrFs7sXswrq0ce11d29P7usHXH0Q5ChVvoJowcqlZvhPI
EFRnADeG8CDu+Duvba0Oc4PEm800eXnIev7rV1HXGiW/OY4FqRubR8dkhD+wAaqW/I/NgUqzvxAU
XoLYj+kpxlgKR/tgukN7csCSYPlJdagTVgEdCmQ5bmB3VZ5LHV8JXyNLuDBRzjz4vk7tKF6Fo8bj
LKF1eiJzmORJyRjju6TeRjCVh+lqwX5JCfH2swD83Y6rqTCaWnseqomeCnLF89D4nW+K+xjHbrsB
dK48H+AKYrsgfP3CSq7MKlQBxOpAlKswvyobbikG5ym9KoDpYXZzL/IABSv/jOxHYWyJbCl45iuB
2m7AcD0ggtqTbLHulLP6RCFOou8xIh3ZQBHW1rPmHTLl8Ce7586EHQj0dIibAW/EAU/iJYQslhzl
e9F93Np3PiaZkBuPLxfdsc+sLQSlMoEnSE2a5yy973aOPna5HJyWpfXRSP3ta+a8+l6CHUHcmq87
o9V5PdbfUiS2huiolD1aFRxxV/EIwv/nm1ofCiR2a3YPLioUe/ghyDhBemLtPfu7NRCal/5eEf6s
mMwXXd87NpI00lhHY9ZaON6TN2jAB+wKUvwYm2hqDdWL9ZhmWaCga4vF9r1Z3L1H7w01ZUvZI+jI
eFb1xKbaa/7B1vUbeXWaBRiiY1RvwRFLrqkrJq4g3AsvG7ODwB0Tmu4bZ+38xDHH8QifaGP2M7W/
bWWw1WvEXIMp+dZEQN54oHnwVCq8yHe2NA8Y+LIUCduJQmRIXl1+ZzMLZUqhSOjrVibqAe8Tl+15
BAWNBpsRTpkHxzYe6wD+ExGdC87U3SgLRwImYHL6/2OSFbes+wx2d4BfZmg8SWCmD4tcpz1x7bMO
mWEF6c7giePQxdWTYLV1CNaNrQr1Q/m587YvPLuwCXaoq2zEZzcyvFNqPM+9MG9lS70slTJG3qih
3aH0DBQIqNgeUgd/QC8djA3OKC1shaQLXnErqmtVXarvPDprJKIrgxfAQoA2KRZeTFLCFdCQ2J6E
KCd2Ic+CDzYctI4UHJABTYDFpTKjA6jwKbhlvjAr1FXs4gvq3qIgyS79Jt4Q89JzTGoofbPDJPYj
Lg8R19Glz8+t4OBuKdEqQ2VBTwk8tVwhBoNJU9onRy9/P4aCfL2P6HqpCpuYarzwgD+6U3LYHgMr
ZCBC3Mr3RQoy5weKETtMh9zSF0r0+7HfeHZ0yb3A+tRim1M9hUxL6/BFYPjDtRSIA/PZ0y8PyCPr
jDO3a931u0jkeSPrGkI74Scue8MtYUN8fQttGULDBoRJFVichxGkFMXhyR/vZJGm3F/C9dr/eH+A
SvFsT3yHJHXhBZ7+PPOwE8DCpYNtzs3wE3Np0D/QozDR2dh6DySdTd/7uNj6ddt0rcDA9TIixE9j
HrHytFHdXZfOgqJD0eLpUNHxBBET5ta7AWOb+vrTKwwfR8huHcP9EYPCo/3MD01joDcvxq3a4At6
QBug5FkKvmPQN99y22w09Kt+iQcghHMNyJpyanYcA0y4BhQrvnn9rDwVLCOEYo1KIhBdPlfWfGeH
Zx553q/7Dvftnq6Z4NMq+r4c7OP0AeU7v5w6RC1wQPr7tJ+K7E3xWOeeWiyv/pBefDydP1XzSrgS
VrHVPGCpAHLjk+t8NkI4RQ8CriWSOGcH/0kfDdFWjzmDs9IDYs8RYChiBEC4STQAlrVK9hYcTHiL
qivZbVBW0TzOed6C5gp8A5O3kPtV1ITHiIXMHfIVO2T5gWG5wxgtHAMFXVbfu0CTpmeFXO5msLeV
A90Sp3CscTSjgLUOF/wWROM0aqjKjMXqtPPPbin/T8GarI7CjGhyqfHzGGFsXrPRpD43YiWU7i9t
pstngclJD4YKoyVL9FfVoQNwqrC8rjWUdp8K0XcPYEurIxAwhpBFbq+lSZMzzcLS0LEr9nJHDEtM
IwD7lruh3+dremkTM96P8ujcVldvMfhCTtj0f7MGU+gkmJIa40QW7WAAG90DarJ+S1dLgbmMIy6/
OLmSiu8/LJ82zd3dv456OqmsgOwJVj/8jYTZHt4p/x5RZZWg8WIJnhQlTXA+oZvKmuA7mQE6ynj1
ghwM7YdO3bCjhWTivp4+8r7Vo5XENwvRZqxCyL/8J3Ylz7hSjlf6IxGc2/svMldyC08XykJiptgY
X3C/mK4NPIKljsZHajfe61bnbiYxwuZ0BXIn/FbWWMXnukrWc95yrArJ+V7O/r25N1kbbPDelbGn
5lMhO6REKUt5sHDIDsXoQX9+Rtx8Ocdr82SMFFV16FG6eVYBx7nVFlHJzhd+sheUzLUI+VUMufsy
4zKpuQulBimem3sE8x5qpJhtiiXPwuLysSEViaeeCyi2j4g+Vup81cKZmD/z8dYPgdNBPu3qXSKU
zOYPCEZO3DyjL4XLoBYJs8PR6lZXaNRVCgRLsY9al0uvKGGzJ9n1MPXBOcOvg/9QWn/786gIurf9
jXMOOss/X/yDu0xvs2mowrzOWXXukDSPgC6oIYBrZREAhIVWhmioNKdqQgneD3A0i8Xx7Y2CVTxQ
d5jvrlYLEPWpwwLiYG7rwybu847mhEZ3bLEYu9wClrSudFkHebf91O6t2qRiqXDzb9kxjULrMr2S
Nm6MJR3LHmTiQhZNQqCuzhpKEBuHgA1Q2MyNq54oKehLParWlIrS78u/AGL3ojtYLGTWKWoO5ht3
a15lzvQu6drmhvSBps7tsf/CuNLPF24scz07E025ep+uoeSjAGDwhbbXw/pMVUZHgcSMYoeKajwV
XNGJfp9WFpdbiLHykZ3SxwFOqH5kLO5x/gcLJ/FGmTt1UMVsp8UMuFuAANn7zCRJgY4BXR3grPhO
/AJkPWAQLOeB/TyWL+yM4++zMUU35LGkBKLzXqNzE2pgKRqaQwTjh/sCQMV9o/cMtmb21X5y5YzO
vYA4P0570J1BAd1DoqVmGOd7EkUahmAsIlndQYGIncJRHpmJjtbr4f1dDY51xRHfXE+sdwxusuWl
C877qBeJP+wDvhbxZP4RgLGY/v2/CAuFlORYkThfX5dqtUrwLuTLr+B8ILjN3LeIYU7+wTwz0xUr
liarJuARGwWajCGa6O4Rl2qw8x4O0iwBcebyEJBG7KeKr7rUrU9zQCq0zSXoW/H0tlyO7jlBPtWw
Wkd0nbTklKQ8r26/joRNUxx5leNYuf7L3F3nQIjDF9mqgeMzq/tm/JMUu2EDdDqhVGnSDThpPzOv
BvRTDPSC7ANRIGro9jU8ohr7SPDlU8hRn65kef71BobEmxrbrBQEjAVo+FqUH9PHxkQ9t3cvssW2
aa6Kcx6ge8a0mhhfzCnxYSr9AGykmx9svAVeSiv7iKCgvh2TeXXLXmvk3GC9yRfvnJk5dh9GkH1Q
SDlcRo4VUVwwyeWcrNDHvDn4/lly4x2X2IhJj90u06MC+jbJLyWO2dJOtor8I+7uUooDwO2/C46L
WvYgNMlg1k8DH/t2fvISiSwE/W4XdVYtUBvudELGuzlaNsS6rMvFLBG1qFuc3UajD2nbRbIAEQBD
BQuGikX8nfsNGZWjaU2wGcn2m/7l8yOMVkGQXDV4xZuEcNKYRXE1+WisrE6qrQBuNOKV7bmI6YyD
kah2U0OQyIH006HobwvEtBKxtZScTRUia21jYl34j3qcXIN67SC0KCBtcNBr97S739cDe0lQOgJO
K9x0TfOvHWYSRb9vWzlfgQJDykCDNyql0vyd52uZmbKfjC3dUTmeWU7tnZ0qDQafZijS9zHlwbNs
K9ab1gkBaTWAUeEn70zWVPcYx58zXSauFYKmv/7yQH6jK43757ebbwsc8huR8ywa6M8fgv6wItLe
KpbtXQU8VRsIaLtp+vG4eCTeSb+Vm5kADu+WmPSLhzW2sQAaC/J7S5c2ysQ3tsQ8yVGFQJSNaVUy
lQx6hrO6njwKsDtbz+uiVByvjf/6PbyA/p9Algp4FPnNgSO/MAW/r2vjtR+k3LyIcc+FXvOdDqi2
LcuLLT/AhLdlht/FL2y7vCJittiY6A8Lf5ykuxaKnX3i0/xpI27LKjyF8NaGQ83Bw8P8EDDWCsvi
09OJbG+wNMkk2Qt8dtDMr9xcirUmR5e3m4orXcEYSxzX2Q0GkGp/mXAaUdVaFbWviBkVNKgQr4iL
0BW2XDbRsHY+gXKe9tJAiciMe3iBwbY2D9AZiG6sKmsCmPNlnvCnAIQDSY3WGzg3JWarbJMKw/N6
7Ud3aODGmOEyX2s/7zGsZVq64e2gGcv9r1xK/e6t0z91e98C+LTFj40wBZxDAQKzLCes7ykBNVWx
yzVyRfKbxtkNEB9AeXDRjjC5c1yWRJ7FRA5yMn0KeeVogzSO6WxAi1mHMbiT/fBfi+NF2H3EUEdT
H6LrWz7hP9E1sGsx/AKfvCqL9/9aVZZPtdvksKxrm6CnmVm8XGqnA6mhoeVK4MJRukB4JDXltfb/
0UjJB4zKomqLuZZWkDhzPDgKXmpd0EPtPCePDw2POfTwT9rEa72MWy7qVvQnWtNqQPt1ZIW32a6a
2YFmfxQiWEIDZeYcr0/JefnpgylxuQziXiIUde+WsQM+zoQK54dVokUZ6+RpUzAFf1HUvwNE0wIe
cHYBwgg3Drd5p01rU2JvZU6VegO23/hBUiu7dnFLzOb1Tid91b+Gqt5iclQ6B0/k92MX4c9iro31
IbquXCncg6oSbK8I+64QyabPsNlEsgh2uuYPkfSzTN9rsC6KeAC72CUTQkzbUDq5aP9iMgeAzMXK
JpKxyByY+1P5SLNelAOIb/Uk/IvckbqwIY2MckTGPfPeilxkkkEOLTn2d3vq5n/m70SeHvcOVqtj
pZG0ZG0O86zvcr6onTaHXYoEAwssi9STzt1x9VVFK/UZQJiiF2ej/fAsSr2XafCVC8yHwQtwRJd3
4N49rUjrXFnQehUiiBJqk6xur2R0+nAyCuStNjBgBSndTO7hgwlpiYS+D/4hA6qdRGBUTLvy3+aL
2Rd8u0rbRZv5oNfBguphEFskZH9M/EYzUfI+VAOGZxgX89XBnnmmMQe4ZL/puck++xMmQGvX2cbY
by/6A6e0aT+GjzVBA77u6ALIW88mwma1HwWFOjn4TfDhT8tTCjaszRHRCJxKjMIfdC85gVEAxUJV
KFvmuzyN5Rgn/f/mA3AT5iBYBDYDnxc+8ai2aQ62hHms+jxG/i0sLSfOR9azyV7zYLL9plO9fRQQ
03vb+yZ8CdAzrhKDtdVgQ8UxNiSrFTl2ZOKVY36qM7fNNzVCXXhxLiMAS0ZZusodNPu5krvdaKkJ
8dIP6xf6HXeL+B8Bmjs2MdqiHmDDxDzW6q3KoH65PAc6fukWR1o2Q+JWdeIRXIMJNAs+sG3YWqPB
Uf3v8xRoDXmkAl1ZaZPl0fh2+zGGvMk1bATK3GSBJGNDbAe1LZO+QJYN7pbeLiTap6wMpU8l+cX6
XbdEvCzwKVRdCSc+Oe9iIpkM466mRHfPgja/I2HGT5CD5AcHIEqI2LBz4zIM6ZFi/yGe+2qGREmt
y2DEG58wYbMBBP58/NOzfa4XGNdHSU+GlTg9Lxj2jkNcjRqeU1cNk7BgehJQ5ZY5WWZwfTwWUFX6
TMaEXBLV0pHmKb68MFVKOPWSKCLykSp3/66Fx++blvaTDBVIrET8FbC5FAv2QJOOXpCZ7z7uEJE1
55+qhlh8G3MZ3jm2ISvWq79NDxy7AWVuUFtRktuqETdx9XzfDpc3uKt7bJDqaDyxDf8fUHtiDuph
zFd1WYYV2+VVFWtV0rOVSpR2wN9zvokzh4rI1c7TTInG8ZwJ2z4m+WEXCcOXB6N5YnO48tnVqPA5
Tr8RYaTKlvFvFReGsAs7ixELPeQzqCoMLJ5WIZP4jrVyQ6hpWDm84UfCS7+I4uEEMZgR0ISw6Zp0
AuFWO86iupI6jo3h6Ejy8lQ6DjZhwOGdtAH64zdTHmfz8jjZu7LGTnhnKuyUcLY0hlNDqH2bM24l
U658lFB/mOjvI9P2BQccAWQTIA1DJB1WWMP6A1aioaG753FX2wFLfy5+q3aefPzCyZjauueAzW9S
kF8Ks092Jkmw8DXjkYY9NKRdRzFfMv1mqNguHXUmLVA5OlEXDPQWzf6kliOo9ed2HSPcEq4XdHQG
dvQZieK2wNMhQf9iTxEG8aveBy9w34rXuiwWwt0VJUloKcO31AKkp7kHTZJAHhmD5s7sY7o9vE0+
DIHQ6rTXYhrWUP7Rsquk7AVAbzxc1IHd0Xk4evNTQJvSLuHlmWjLkPnew2oWLzY49g8lXz3sUfyk
LhCYsDUQUDWkuZQ/CW46TDbnoC2e0HpuriJqQd+wlZ6yA6v6QoK8+SDXK2AZJVNVH0rjRpekD0+2
Deitv3G2lpUqY/o3Qw5P7XREZRpZK+3Ji+kGvEj+Aafo5uLCSkowZ9YUyrsYvJDi0JWWiUmbyICT
TdtbAPRkp7jEbQeHw+KGi7O0qgdtUEJTTj2Pe9efcuTY95IPvh6K+gL1NOBZpqCZyKuipraC94nV
piOxZlACL4APu7jZKrM7iStRqTy8k0HhjRVjFjJ0cbY3C0um3xLRbQ70B3B3uYWj26DgeeBbi7VS
2b7++Lr1M6GouaEnYloYKpkTU8palLelF1EqSaxAjSW1nO7i562Kyr87TXRnJve8F1puhjMeY0J9
MSGYkNjZx4WFHaPgjOL/CmkMQoR09GO7C8kSzBJuOGKdgaWzfaRKlME/SMrhy3be+XEIBEWSEp9D
gXQOQprag6ehz7SvxKZa425dSZjYq4lslITpXy7BmfIom6Y4z3fSs45vG6iNNAd8E85d86xqbh5I
Z8Cbq0fjwgRAicFYierDhfsB3jM1qsOKDqtU5Hc8hfpg0HJJ6Ic68Bi6uv6J5FL6yFaDMD4TNw4G
k7cj048ly+ULt/2Wvfj9T6nQawAu3kWc7vSXRwAMEbNNBDJ7Ig6tHLsacPG98ljuxP2cIkI+BAKm
M6weBmlMUCAeztI0d5zYiTWbMUdP7JYzdMtIfWkENhLTq7pYp3MW7wfADd2jU/gXyfvzy8Ygt+yh
D/ovyHL7+c6HSTtE4Y6vaQniuruLQ27/vaJJG0nGsLt9dioIYx7HIEuOPCsijI6KX7kN0rYKz03z
q8O+akvWt2cVxGjOfH7nqtOeTmam2p1g3goWX51o7FVeORgGCRPJZVieWbbWUUCSZGU/hsDxeyXy
bsaFuyBWAFPiXF10urbiRgzz7xxDOXM1FwU6i1hzYLKS14V9u1XKKgExc7ARZP9LGz7ecZgXK0ro
XjxU32SaVuktFqBVE4BHPGv+hmsOzZ8JUDJhw3EbR5LmxXDRj9NufMYtuv9ko2gH1aDa+4xP500q
acu5rkAg35WNfXkc/qv9QJxOwOD/kOt/IRBc5CPki6hVtsB2qKxZyCLA986I5wWA7NukQdv/FHHy
UQmO5adMOtsLZm7IIjEA/6o8kw1GhjV1A5sr08u0m4St7yfH4ssYRT3tmym8H4oXZ2KkAzAR9bU5
I5HO5sNw7YnDdEuF+RDkZqIhY6pktmj4Pkw7C18gT/OgEfCt2humXfhSBk9LeywQ1IwiVWwlUDvH
miRcNtxnp4IAwl5e2MhV9YC2caYnk0WTTeDwK7xL8mDBu6TqowvUL7JcmJQOKGKmMfOonXObwJdv
+tnh7PP8vQD4onu4HrimDaSG2J3rpJ0YXwNCsKVugjT5ix/JAr+FOY+YS7pfiTlsIU8J4KPjc6uD
qgVr6Bk+mZZuqiNU82ZdgSb7HEbJYNkBlq58AYrQlDTuYktHDoVCJzBysZfj6FZ3gx/vkITVP8Gf
DM7sGkqEsGQHVAuLvxvw6J3XwvvymQIZo9l1++/Ty49n5NqqcKZWCJSb8/Ol5HD16dYM6DaF+DiO
pBmhPWk3mh1CI1zNDWDOkN00lo2r/mol4JHUCF2QL1kX2SnqjCs2SysCbtdfs5T4xOSskWI0pLL0
1BguS3tFkT5YNSimtFgRuB3kP3fjEs8TY82fiZXRagKLEIDlFjUCfBysEtCE1lIFafbtgyJrmNAx
7czipP3wflTLPAlbEI7unay6LBHrkptCKvkZ0T05oK5A4l+nHT0tYwszSv1OwO8IO0ksSWtlCmIo
lbSj5xR3cCEcIdy90JLw/yc+qsW6i68R6ZhzbMdy3AYU/EHn5G4j7w1zWKpUNwmoikChv5Jcefup
3jzcb7HjImS2IuSfeHUZtjAz9WgYZSXWaAabJBYcZsLBMRYAOR/gwlnMsCUG6za+8B595hfzw/5p
+IFjeMZ5qy8gt8cOG3Z2Fbju8Z4q3i5v5PUFMvniN2XkVimtioP/v/6HU8uAtguU+dHh0pNaRIbk
J99dU55eTWHO3z5LcpAJKUaxj27vDoZbEoJOmmQPp8+wphbN0NymZytJbv69zQVzXB5c4u10EsWR
gqDSL3gBcqwG2dI1gXYm53z3IViOWepw2gPME4cMVLmfvWr86LIGYlKN0V/9KcEzUXwfz4uOjSSC
5w3YSbA/QjiM2Wcwp7bVczCrAxWM8Wz4hUqVLXOBqMn0ZR5fysNmG8a0b1RY6UPji5S6xBPPqyed
23d2Aw9dLzicaXacrDdEEBJeegD62aLV2iO8I5CslGGLlJ9qrqaS0XjByiHCon+NQ/xinkC1a0jH
RYclZwv4rTqmt6C2C2wAszQzne5dHQg34jFLQMMHp9xsRLQqtqfCUtxZIMAPJ/ULiQLkBuhQwefD
CUJxS//nr6sgXn7V+mwZmM1LvJTv7JpTVNYopOLO5PJp/qdlRkB/JwtPZbq/Hjbrmz591xDNFwwS
c1PncQC1HlX70yKwMAuRJmmHgq4cZCcepk4Kw50iQAgOl7mdGxpXfHOvM5/crH4+CZ8+ggzKt1FZ
cHDtbzJag+7nhDQ1HJnJBDDRyU9wgJ34urU1cFTYS2oLFX1aSFbVv3RG/CenVK0MI+G50Ai60gb8
kbo/l9VeN5Br+p/iObU0LmB8UOnGG63g1kehDj4pX7I4qxqf19bI17S0ZurmUx1eGiol5Xer9t1R
RBpaC+Gybt0g+mtS7mmiieyyREjzl9xKdUclP+alMdxr8g8YFF6H5x84M6WzjMov8KqTjYgBp6NA
bT86YzJ8dGEdL3sjeyx/gb4Kw666lRxoNxaVwySfFYqRwvx/bGWiIK0HYp6zJJhLJhcJbAosNCAi
igu0QaOUcYG7UY7C2f959g+nais/Wvg905K5plaC8buy69HZUmFUs7kdk+1LU7U5r25Zo54ZBa99
bFoJyg9Um9eK7KRPk2BUoO4TO+25pcTQhNurEXM18nSeZntHONFmMLuNwoJeYz2VxsSbMSeFFNph
xB0IjRs08eJr54KtyaKmcIvtDgtSvHiD/MbIeTXbJDu8HJdYmgxnmiFSjD6LcZ4/V53NMY8RJ/Gs
4SxCJ6Cu9xfL04+bpwqE7d579B0yjK7PnXXGokiWARjiM14dHZ5iTfUs3YBig/JWIO6ghRiIFoVd
uOi+m0HsYCo/iddYecg8m0RY0zlWHhWHlykTbVfRHUFd++8MVax95xg3RmUgGOdEuu/hIyW3N3Tz
nY9fJMrCymW5ec4SHGQEb8yogaalb++JPFg6soqrQQRToMNyKVwVXfU1Wqoyes/VxMYNGVd/vr7H
pXeA7LG6YZP9vW62y+3QGINagNj2JN0Cnz9vBAwtrGf2CRTRhuxOQvLfkxWhH1wKaC9B0cCp0Eoe
gAdaSEYvJRJyco59ElJHdilHJgniWZIdRszrsfJNGQXJC+3PK2cO+d88/ORboKw3P4wfzjnDKZgF
jdNYuVDXPmpL9JkiVoOWVoCRe6PBFLIh0cHtJi0zkQc8B9J3JhWUIOysokZrqSXH2NUIwClmxl+u
avRvDXE36vQPevHqIC2FBgPK8iLKWryHdIuhHNVywkdXjVIto96ejW/1mnCGTM6I6WzNE2VHG7as
SJ5tQ9zF50mu8U+z0BZiK2vWaubboF4PsMBBJhyQixIXHTqUK0xtiP5oTH7ojqVN33iLTlShn6VT
ZfLTl1PK0eHfZaWVIaemVI416kCL7RKxAsDNdZ3C5S8Y5kB9Z2ocGGXIDV9l2SFVuQB/FTTXOTY1
ZeqCK5PYtC1QtfbvCAwnHJUvTEaFLnj6BkkiIc/GqrhPzPoIkwx8uLDIGnapVHnQ+Fqgq08kI7Bh
xE5xXox3/7vDH1Iu0KPYeZOuLHImdFjCE9CEIYVmPczzoGhmE9OSTNEqYIRuBarXoGvhoqecUdbc
VmX49pO1YrxAQU51PZxvxMQboDKxE3j03QequDR2NXnb/IkUUgxErrYwAjous1fB0noMD6vr2j0I
p4tfQ5MhNtt6ftj1LKNf/S5tZa09OrG6FKkIjPPGeas0QxBwVHh09Z7GZ1XloveMl3BXBgusIhtq
86sMAskGOMROetLkqUOkOxp/IKAlauYYPiquv6bFiGJeEzdTOkHtUpL3bkzn2d32BF1uCJROtxyY
37OJE3pAWpYbtYf5Kj66rj4tWBGymOzMln14B4Ze9UDT6Hb9BoK37ZZqNUItVYpFeFV5ZHlNT2ML
jB+vcch4MlUrq5qN7N/Z3QXaovc2gT2662KjOtuIFGpf6FKmj8WWJxTQ0FGVUOB5qUOzQ18HkRAm
HEMFFa26bi/Ukot4f8F9s0MRIMT33Ou2OJaFVdqUla5bjjcsWtHjx/4dMBT6fGm9x79gp56nCWgG
dXHJ3Qw2lym1jpSWeBodNiwbQe8xfDJSSZWCzTDV+g///Q8EZ1o0EL/ngPlRV+BuOS6W0aUSyeg9
/cRcw/e45XHhWkeaSzdVHLhVLPFsc7l1P94X63jIA4JBBwj6knusn1In4AvZIh1NWpIMxdX/+cjN
lQvc/1NEwJN8gQLCDsZGcZE4F7AdsI1BionI/UY99fJw95QTa4wjN77GVZMr3tjFrQ3jz1s8Qksp
Fn1C6jN3IeYNHwFOjqI/oDM00wfGZkpMBNd0AIoPYSuVzbstAdcLUT9qkxwkmamFhC/IQGd4D7wg
zvD+nxzDKp73Wv577PwQ3ZEWwX5UlVYB/Jjewnx43EYlVEnDOG97kugRAcf955lvppfjc9Af9TL3
9KUykLFJ5rv1r6fdTTlafyWPYkaZnQXI9r3XkwH7BNY4YibIbzQFGgiybDPyJ6v3V8JyWotm0jVZ
dUrkR0XjUx4DWtoxVwb82V7TYxqR9xLqYhSbg/RZfSa7h/m2uy06rcsA76LXOaijy5DW/9EXzSOs
mlps/dlF8XnhezdWb48ycbdLtaslXCKXGDzoixRQgThFsieaciMsLoYMcKEqc3fa0bKXuaYJtO2m
8swsugoeIuyyr4v77JyAFLbQ2aC09kd7yCMO2tQqAz9jRYDXMa4n8Jtp6Rh5ym99HMNzl5PKlueX
68EaRhy+LMjPHHdpT4qj2LmoOF1KtxVfmN3Zky6gE5ws3ylUEMMh6hpIQ7L33HwNcHD3Y2v+/Kou
+I9qhoNWt87ynusCYJvXn4y8TwL8ZwjBsUL2Eu1IU35cTNW8Rwv0BPuWbiw5D/A1zVV37nUBI3Wo
nx7klg4xAay1Yd1lKK7LSH9jPlAjVyyUQy6jfQaXI+Wa0pEL6ZUk0zFAotu3lR+BWDpEizRLj30a
uOMmneyrs9EpM8bNULrhOAZET/1oT5wBx1bkbUEcez5xIvRVPbkQd7vHL4ZMTey4d8HV8m+gZbxy
Tm5x6xKy168ARbCIYO3qw6vo63I1OFqwoZw7V1lxwvRYlNubT2mF5n8DhAhA3j5lbY628zTEhoZL
Ih7O1/0vAvOm+I9wm1gn6Ggtw/zCJidPZDbqykDdELure7zRaF0aeotd7H3y9I34Svl6n2AGAQoo
wWXqog+pp9mdKC9Rn190JPdd864+aC5Na5lH+wVynERuHz7xYCo27mFqoAa17aVtCqByLQnY3v7q
zXzWAmwz4+iOwlNUpCNU8obNcfnqJ4aaQzwP3DwWzyCogyZ2XTQCLUrSCLMwkeT7NxISHWsZ96Uy
YolExqCazaU+yuDef/YSVrAgxN5A+eQ+HgAvjOfj1jE/4bPYQGg34T28aQUUbRlO/YN/Ua8Xeyfn
xPd7x2F0yypbUP2qgEVrmhaT1Qq7EOV9REWIlRsMmbAqvJW5rpXlwH90o3KFMgo9MEq4oqGe7ZnG
V2e2MfNZBG2B3E/sXyd5ajRbO1SeKpjIAyr52SsgPLHSPQKed8q5QZZJiya6e/GVZMc2uot+GkcO
kfPhpBA7huEsIZMnUVlhfUzv8fyH/iadFgY1IA/mqs+iiioCjJaVmi8IVm/Kq4MGBak0Bn8wXgtb
iSg0J3iw/P9AmxCH0UWTz2W3dYMNrJM/8iIGdxSDz8v2RITxPDIO+R5tKj2MGX4mXrqp9vr2lKRm
QSQ9g6ri06kCm1GMkTPWvHHVlb5YB2Fw+G4wTHDrDMQcXfRG2OhGzpuHQGdr8WQU+vgbzkPWz8Si
y8SKSoXlosKu4n5LLKBBo2A4ci1wU/vjjF+08TS3OB76skiBoCxyi3dSNaKL5byEdqTvxyIxYD5E
gOkajXDej6gCJXo3HX0J98IbhMRL1eZhvFXFHaERjXJROBJdtclCQ0+p52pAdlCiembRwDgqY2FI
gn8rIpIkA4xe+mIiedWbiFVaFEtlcXTl/9kvkVx1zDtUXc0FCLT24UHr0cGVbDbUHcxY5OSiKOXL
MOFF1rm/9GRztBFDaQN82QcFhxh2QFd7Qi9qwHA/x8+OfReEO7hvt1RdaC5Rw4CGMN1AwEGG8j7x
VHxCYYczafXTtISAzl6SdUmQhm63qwaSckjhVINRjinOeGNY+YwnOb5ArMQ8jWD8BG2IXjpyyy92
Gw6oYuHIB1EBtU6z8mqt7p8z10yoVgmCpi/td7hso6IegQgYmLTVal8FQ7s5tu69KKIv37LhzHZ2
S7Xx9+gbuVZ4jLZm2yqpMn3HHRZzXeNroxfxntK9cHPhbJ96jfqeaCLUAEvR67oju5Wl3aEpP23f
dhGcBVrBp63Nvq7Bj5l8Sd3a5ICJnO9hi0dJuJkHBUwWrawWFFja6B9b1ZWYV90tkNi1slis9a6x
XzRyzdGhtTv2AxvOhR+UZ23ggCiSFS8Sx1FqFQ8UX4U/cWGuU18xFbU6r950xmQsiCM7PGPFzbkN
WjH6BjsrubysX8CDSOe02GIwQ/JmygtOpNtm4K2PbkBTRW6VqAWUt3DoDyvEdiPOFLpGGvXTfLpp
1wO+4cvRroOcm4Zmt2sEhOOmQuMvcxBmqO1IzXnEsWBPLfCt1cmKgX/3N4RfSU3wdW5l+a3pasAY
GlQPmlIGDed9SmYpaQHBGXigQoDwSirYUDNyLqoFb+pN8LtmYcVQES5zI5ESWg3iAzGJ+qG3mlhe
sq6k/tBq+K+h59Ov6xEX8GVGE9FzaD8j6KafzAcHbt2bk2E/sict3PH5zfOVdR6o2kqcB9ABlqsR
g2rmpGTFoQFpDKwJX1mHoYykv1PtrG4eo5Isp/W/YGMiRiz1tc69O92wPvMEjoozfZf9eF6VHOcF
Xz+PoINMqJvsTq6W/ar265+Y8Z6R+91OivmHI2aZhq8AhnbV9nTS25CMxetFEq0s6OluT0FNwbwS
7fTOk3IYWtu3gjmeRiorxF6AMIWr6RVcRabR6p+mAsgond2A/le68T70GcZuxbATPXyNGGYbdwAd
YBqBfnmJwUcw+vjoPKLumj5f8edd66FgDuZyI2vQ6Lk5ydn4cSKniiU9osjbucmdz3rYFbGvYVoe
hSauTyBuEsXXgE+2ikoHqEP9029vUBIYChO0vL8kGuac0v2uw3LISY45awlcAKT8gDJooA/SSK26
cOsnpQ0Qme+I3Qe970xUrDWvPEYaqxuteMgwJdGUkNuea8aeT/0nDXbiWHFYjgte5CCcFPP25M6k
3JTZZTp/nP0ihhq6FEilC8mYItuz4xKtlgTU6VTjG6k3+qnBOjeDnfnGlzmWxY8gYQj4HzA1hMdJ
Bt5+ERsks05WO7r6QSKMdvHKHQdJt/UkgWk0rYxuitJJIEPiDUYgoo1hEnQnQ70uXywtTUhIK5rk
M7nsuBr+iOXZ5e47S/Mb8M1XMCYTBbIUIcpTAshPYGMJb0EZevFxpWjk5hZnu/bQMbt7eFAMg7jO
aYw5kkeiOpXG2oCka3zNCjqZOwn5OehDiPDeMB4XpKB9aKlzIkYjVpUyAAU4MOe9pryC7CTJ0+D3
Yl9kHIAt9tJRbbPdFc8MDdjwXaDgbiVOIginsXtMbrkU4cNHKEqv3fgpXdt0T5z3IVCSBJIHhwgi
y1jxAjFinDVD6ccyMvmkQ+HPmQz3aWmFqaxGcUAWyDqcgU6PmNJLmspl9owzU+uCPhL0ZjoyHcLL
H6GXmxCKlN4WN/En2OUOJpc6QfDTIEdWT4gYxW2+vwMSAWCzaIaR4D0vvok062D7KExTaYLEI6YS
RPZjcJNpsx93Zjbt7/oR/eM1eyRjNPMtOD3+q7feJ1v4d/g8xt/V8/IBKezBq+TyMK54xG/7vlnn
8HZfQyq5eEa0heMK3Q0jlPVBelPlHwZjCPJxM+xceBSOZ5b3We77iwaXDq7u8NZTpBMZ/Ev560W9
tgzMolt802G3dvALwP3blCxdNQ0LctfK9Qx/J0mF3c082reUtJ394HIL3kCb6/TwjcVWL3OK8ZSa
iu2i9L89hD0bj09j2xRVMJTGnVaBxLuWIrHiE485M+QkulRyKU1EHP29I6TzMpJbF21u/UYTEO9m
wVL4eCcZkzGkIs2vwVxOfqXIwvQMpJLWo+bjgEIrlpbdiPlq38ttuHQDQcUVHFyaBhTOHTsfnR0U
SjgD0Iye8kF+wnntDeHwH0crOTY0kVEXYGIrPzxHUyv3DW2L0+ejYWJcn+9Gdixu5IXLMuADHWyl
kjS6ChZQrFS1Lxy437hfDoA68arVMK3Jo/0BvwF5nOe+Z2OLt+rh71eSsuxc+IEs3quGlCUhx/Oy
2mGYni8zr5wr+Iy2Mk5UfHjNXdgqezb1k+VK+h92B8CFU3gy/QkG5QDAlA7EN2a8rW3FtsW2RZav
gU31WuzCC5OgjQZYbxlKlayblmC/zFG+X3/JvlM00XAcDlfpdelrf+83W20+PnAxXvZsxw+HHNZU
bXaaPvjOZ6/qevaGRGIoiNQbXSys+yoHVyVc82xoixduSdAjkzgWfUVlQMm/KSX6vHziru6dFimH
h+bIj+LTedgjbsXh5lJvVNOMYVKO/UfdHDb/YzVapj91TtQfQMdWW15bCi556tuyQcH7l6xBVRj1
QwswJNkB5gM5FnJVgkkiy9I5dC9TMF2MMBWDweqfJzOYChSYRSqpnrq75t3EooTFM8MssfgNOjh5
F814gidmGu3Cr4tO2LX0XxyzGyZJg9Aj5K1MAb5It6h7oKaSkigePL+UGrfoHIZIiSXrFAjXEDtc
BbmV0HCn7iF74cQFJ3wIqMFyiUDdDLUGqerBJFn1CKKgshTAQlZjvJRFcP6XN9Otk6n7rGg8jpNj
Jdv36w0UL8BqNvLawQf/g+BSA8sF5cNAaIE4wpHyXqVVZEz4PVnwmFxhGQ2/r96Oxn5U3H1iPSom
9wnEO1tXAyPFcBG4rniS/CLA6iClY5gyr4sr6NWzTc6IRA0TFV4OwO7VmgfUhKiM6bsHTNsTMZ2C
/QsMzndJzSDbkKTmMgRNadwCfu1svjXrrpeVvjyE7AFf8v1t6RSuTLI/jR5Jwi0eV1PqSOZOy58P
6ILNLcflkKTvUNqNHG2vMC/jmNlHmhE4GmHyMmx/cHTuLlc2rJg1+h4yn8wwb2p4RbYzGLSAwUvW
5kCsvpLe6rc7xGStdYRaKoeMJ3o9aV5KfZMA/2TFpfhsQjhz2tARyJOHbKIKlH+XZRBVyFsSiI8e
JPbTe/6KN7FOJjstLL0f39KkhHUrtI0sT1xkEFIbwaZAduqOiEb8vk+iRyw01cYChq93oE9jYLGE
Z0wM/NTsvMaUEYCoBeNqbz6YNSiB03g/oSnXb91eYE5Y2cxRXsiLaDoyzN6xR/TR4Sx1TfSzRq+U
9uqX3Rqit7dgaY+nkO/LZ/gAddIAUmnRtIroL5VrzatfSqhAQZ9uzCHtxOfASk2FeDztni364rIf
gWCziW15RFGG2Q0r1w6yVM15I5UM3BjV/ylRtirLiXSXVyRXxtqu5Kl1TAGMa3xlvfM8Q6wXwCUe
lMBjg/xPW/kHSI287BLFPcdPwctvvfKO1nin1zHqgjdo8qXu8YhYObfD/oWXvjav0k/WG9dWuw3S
1Y3CC5sT1XDxP9TItCQhylO/L3GW0Ls5gx+2HPnY0wPpZEADhE4NWbJgQTff2NkP2BMTEKx88FLO
c13JOZrkIJfTytg3d9mc3BEnGQ8qlzbIeKyop2Y1q7jCxzjM1Rq+DWHWfL6r5n4H2kVFzsYhoOkl
pcB06qy1YmEHSJkb/EACT6U+89vmZamM9oO76JN/dHmHRtI8sKNEOKwjKQmiupFIg7+DBsomUeZA
7n8/jUBAqD0bOmmaT/12RXt53UwpRoBLEeMiCUvngK0NlaAgOYkD2VVzf4UAMqkv3nMqr3QbgKfy
pk+eg0cHSmTW/G1uraxF76RtrcoRVACosinKyIjy+gQCcPzt4E36QKT5zMqP5ix84ZjY66NSRBik
/R/XtTqJZF5RvUbb+WeiiCmIr3OljPK916igsYMZ00F+T/dq8cGaInDY6CBh4fsBEAJ2qTjjuLXt
VaFv6JbZCKj9wgLaaLgHC6+px7pv83YeE96TEyaguSMSB86bd1MrTIaoLwzFNRLM3Wdm1iWmoKi3
QYhkbxdSzZSv3DKC4RZ8bC8elBRLwyy3pWAaHilZaFr3XPgUhkH1i4PbJD8nSGI0WaDMspLdhccB
QmywzLTA3Pi0SlpisrNWZTtx0/qjB71DNOQiw4T4vCzOKDwlbIiR6zftiOiA03MqbbZQRakXaSjl
eJr7Z6yfJrwtzAGw7d2dHCZNWXUaFE5vqjxaf6BIt0TFGCKdZNBBLFvWCh/F/28bEfwKBSlIkUYV
hEHb3mnRDsR5rnL+GflbTUCHFfIpxMqOdEEQWjqimXFSdjEVkID3LACYu8tU2uoe0PcKKbonQMzE
qFhs5k5Pw47bocHicMwpbWfPJqk/f6Jrfaf+IsfYU/E1D3RhEGBNMF8mP3ulY9LDWQ+irinpChqf
brZWiO3/D2s24A1AqIZibvjuO2/pU8fM/ssT8xRKNgdJ6ktyCtrw1vjm0gZQdWG5H/UkCwIMQY8G
4BMo8gzwAQbiIWQgC4PDt79v110U/FyyYIr47DnKNgjHo52nzyVMbYiF7Q375To0p+B+IlmYB3p4
fh8iMY1LCRG5xuvdbQ2eWUXx+K+388aaeiIE5RaP7aORgk03sVUq/iFjkpWYBiHw5ZJonyPOVoyx
CR5fOyRUO/2R1z4FWyty7A80nptkDsRJBjeJbJNkDR2bmzyMiOxU//Pc9IiI/n/O+G1ik6qNaN3v
n/MZm7d1iqaXqAitvHTnQfWaUUa5Dy6dG5q5HiTZAI/hQl8KXjcKQ8qzvdnuc6nvh/4JBEyvpgjf
flvo503Ucp2DnN/Rdj8BbrIhckEabDIk6oX+eFUNaLlu7REHRpYTnP7ltd2jhFWLIVnF0vOyyRKe
nUIlRhHN450o4tUH2GIAHYzNRXzCJrwynY7kI//b7PppUCtjdMqw9Mqfvb09PAibTHMZvyBYQB3l
dmihmw1dT3Cd+WuZ2Kvt70GA/N8lksJlFuC1tciioiaWN4OVpZVblno3xAuDLZPbRetdnx1px/zj
gdsFRD0LuCsx/2BSkFiVDooLNp1dSo+Qe9eriZiy3WLCr1BV6h/MpiyFp66cOtR8ChG1OHzN2vuE
3eZP6KDL5PQraapOtU+IMzh+xTsFVGn4HkiAOF0M4ewbFBfSy8GgmtcJnlQSrR9v5mdmBsVMPBvF
6UHjd2YjgjWeAGPXCI0ttSFxZJluWc3EOQeaUm5kUktI1Ypt3l7cpdZRzlLx3tNEYVX9pc1IBDu2
4r4RVREYZppQz3W379/NRoHUmWLMbwoxG5GXYZ0FGvHpEGycPgJ3lduw8w/gBt6cOdS8TNVnWUKJ
sQtyrPTnt9HsVkuQuSRom6hJ8qAsIIkoc45y2mMheRJSrkJ8+9JkhsUJZ9AQzL7gBHTOGm9kH30h
wj88zpBx45URGNvqAbb/0+bFZwwXX72EKuLh9NV3Z7+oPxRvYNduTiLJWznFIxljTbgeARuthxOr
+uTsev/QSJteULQsxkWGL8ScFBe9Jz6aEOvJ4oiLUgaYtQCwnbteR/9pnTRjeJ3eK26Ey0f0JKan
1q83CHzbY+Bia1g5kwvEpkR5zfSAPgKfWxq86XTRfFnP7ZSxeCYK8a+KHCL1z1b8gkCOdtHXBoqE
pdgdQ3xNuilY9Je66dDGKXAqUlmFF3cOURI7xD38CnG5HBoZ9xp1hn2sIjJD48hfULnw6ZAgFiCk
utU4PPloxveUlUnJ8o2DB9SEJjwEMNtjse7mwpHbYlOAXNphkoWwEtGJpHO4Jl5m6e17dtuvKPaJ
QNLfuIms+/Qce6IKUyYSFAdHQjaxjropJWmhlTDhQ638dnW4ZZfhUa/w6D+RAsMbYtxIVxmBQh4D
HmQB/1wTfmtOZZlJO2LdxcInCEGCzf6nNjcP9Q2pbn3GcgR0Bw+2cf8Q31zyAJPEMA6lmv+v6LA0
+0FEOSRSI3IA3zSqoc0JTa+rEYn3eEOxZ7C9ToYppbt3d2uye/4Ls3gsRX9l0og7Y3Gj8cn5MOEO
lJ9zkEkp8aLRD0EgUnz1FJ1TYgbygXhbr7T4gu3vjGR5XdcVcftlv5iD9ZlFQVr8PTNQB68W1N3+
OCOn3XRu84vBzHsuFLgN+e/t6VHPPetwLjRXdZe2nT6hA596CHV+MqmNyS2+n1/LmMRu0hKk+p4w
u3JzctIPspi3Y6jcR3k8PozNlKevq+DRE7LdNqMak+p86uVcgWqVbaood1Na98OmueUH+fzKuP2m
iEkDtQ2e6kUrpR3pRGdPNmHNAnFvF76IDegZ5bB1ebzFodvZp2/FqAxSdoWFAIPzgRN8IYcLLgKt
PDj/hiqYdvzEIgcE3cFuozuRPeMOrtw9IclWoJM7wZa1pdinAoiSatZks9L2k3XzSkCzwcEopPl4
6zD3UupN47fli4sWeGfuYz3I84CUL4yRSl4oODgAJrdiTsRsKmBw5zUBKcY2ovw+W7yEMnj1guKx
/JSJAPFPCdzWG+HxM9s2bcjo5mMeV4OluyKkUT8b5MTGicZLAfWQriHmfxoCkhMqcUd9YKTuIJrX
DXeu5AWC+5zzgLFvrdOdFbo1fagyOj7Hr2zmHSmDZNaZn0uAuKisC8Xd4G7qezVTU2pMhyKiE8Ue
X0gvYILyDyMFaO4NTUHE6eBHgr6QFQcKIJ/8Be2ESa3amJdnTtrIy+rEZxI3xEchq/CBordKUTIA
r/eRvmsInw+THeOwvyux5jWNw2ZR5UEOuc9QD4/o6iGEMSzLUiK1E/R6bGZmW8yyifMSuaKZYxLO
kfORT0V5q8dyX8d3Wnwa23ByAsk2IvcS2BRPhE/OVfrSJ5KabxcfHzrFcNPUo64Agmv/2Qse9bBO
p/8YFH42/ud3cDkCGAlUas9P4pSs14EYssJgjrgdVRz2mpuDHIJzmzoPf5W4NTBf5LJzSnPKmS3c
/yj02pnkmYWfiy6jjYokSJdes0OzNR0nEmVz0QMehTuEVYmxLBooRTlIfezyu1kgu2PuT3j46Ei6
zEorOaydjO7GASHnJ6lUW0RabgQ5S1fjwOuU9et/gjjTdQduvE9KyO4mrC46v+mfFHYS1SnEHLxe
wYFdoqYYEBkcEgdD+whN+VxgWcxxZh0mnZI4jyzD61n4tUNmE7xmQ6OnFI+jvdtgQb5ZH+7dGMwA
4zTiP2WJR4giHv6722lg+BxH9OgQG9ngjBOLImcg8ZZ5FaEBpmlSln+xLTsM7hbOTR9bH1TYK1UJ
pFf8X8SLWvyFZaQRxjHj13gdd2Vmx88CSXYncgxryW6H6h4dzn5FGQmegSiJIw3gR4CINbq8a45o
F6lhwNNOykDoP3f50CcX9ud89EQktynIYV5E67G1RTiUEP7Wlnr0fzSv2Q1erScLiLizKf0ttk3V
s2iYx64BOFTE6hP+OYHCI1toZ8KV2aWEgpXKwZGtPEpB6LCZIGUb/ruBvsKeZDCws+SMhHpPPC2a
k5bJGK7xQFgSoYKY/fNgIpRfLIZed3GbHcQufA0DQnKWuiYgQwm6qhjeDSS0aWmhwtULncwdc43g
t89DYMclgQfp2EhKFpn4SSHwmDkkufxIXJWIOEvA8R7CH9hMO/vFIDyQCrmfS9jRQ3e+OaurWFpX
PGZqjXo0GPz0NrUdY7gGoa2E1PAD/Ipja5xBLXGX1bhM6QgCI+2leiZo0ZkvHupB5m2mOE8d3Zyj
EWwf9Z61ZFaMJcO8yp2uZoxs6xaPnh1/MPp4SIhC2RSqw+yKGrdAxR7hwzUPWsyL41LiOGdQauoh
wnIpVxNGTwjVyyqmuRJrNeg0dKup29sZTJYJPx5kaBxVyCTP8pqavugxog2sPxVa5LyhSZvbvIUG
+2QOrUFTyXmFoX/l3+qBn5m+7qAWo7tGlM9nF+9MaYEFcAwlkCrE/yYviHfxP0pZocHFUIiD6/SX
FQuTnR+XntKlS+g6O0+/p4QeQt4s8v2UTjdXHqN7fRxVb3owIJEvNc8cLPkYTkegUAFctOWNxDmN
WSZoehLXa4buURDZei3FK0RXR+IgJCrbw6EhVdH3FPl24wcnIRzSq50CKnniG9Bx6S5nHTNmr+2b
MpC6rULEH3kjM36qf2HRXLCj3agXyCCunfdELf6jU0/spGxGaAp4XzxH6+00+a5LsnETTtjoLTIB
ZfJyW4CZJlTuypMmb5jkCkIytInlM7IgjRFAFT6bAw60G0xPOZJ1598S1bxBlhcxOXQ1vANDIAXT
heIou9A0auwTR1ivdwP6TzdI7/Ui7l6rUlkrMqmOO+WAq+OBrIagveA4gIZw/pQOT/JYnpgIj/OX
3pOFiFJhPjq5VpCq8YqLZR5pPRCXITjLAs9uxaJpJrvPNzSFUQexlsmmQRd7Br1WYQ3s2bk9T4Yd
jYJXbD2LT837gxmqGV04WaDKV4LGM484ZD/gjfJmDzDbJ+PBB+G768jeH+51lstNNjNzMv1ZPsHb
h6FoJiVjV2TKfahw5gWmsK216xjEzJSlXmGBMpFR9pquPEdIAeO1HrJ4I3hw51WY5u8PI6WoM+no
mUKDaErC71hTO7SWI4xVMcyg8hlUzUAmlAADo03HzkAsC2FAu953uP9pS1CaPkcsTggIMW7VNFHy
Fz+2/wvL/KRLrS0hKE/PizM7nng3NtsLb19nLCWUmyJca9qI091srueihCMdad9RenSvrVxR2JG3
BqSbiKo+UaemMrUDcs5iVshXWiQT/M4HtHz3TS5KAkkKIhtGa+X0qvracdFvRJiYz+7r93mCZZnD
HS37mC2tYYRVShllVpfxgAyxHzjAwugAEpQlEJKvzM8DFZHTcy53Z7cvqmH0Arz3HhN+5K7HYEJU
jfUDO3RVevSQgI40kbL+o+odLqj1QNmrWF5noHuwx7sDl7oTHcIfajIWM2qgmeF94fHWpfTUaESR
wuKBxYSHoDyM2EVkZTHY15q9DLn/VgZvozETkXkKBIur6M2yAGHGwejtHPpb/2PI/UeqkY2dktF0
dSzwgdwEQMJjsAtx/d8NCBtpKLT/oWg8SHDDgM8eSFkzdimYzQae1hu40XZJ3cQ67IHGt69Ai2iF
/vbXDUoiJqMaLwrdR9UpTd1z4ZPZBj1NVeDlkOopLcwYNfLkCRVt23LrpIKlfR0fMlh8Wwi7CcEg
0D0l4H9KrhQQUiBG5E3xVgJEQXI/vriGVK1GH2uEAJ+wCSJ4IIOrIWQ0bc/JGK5ZgkJFJJQHOwQt
fqHJQfQxRxJgl0U46OxhGu7HLjAKmxayuoEsmDY43q/NyxjacQyk/QH0t4L2XXfnbml+LgIcsymt
LjHM+QZsRMV8vZlF6RyE2k7vakw5+GB2PDSV811w/YoYIoWd6a1pF5BeAgU+WUvhJC2zTKqkJEAe
TCWBbMlXDv8thR6Vo0ZEXHe7iDV1apc0fqv+w/2ISg9iwolj5PBC3WZOz8Fjyo+xqbRWlt38C2uk
y1JdukHmEPzIeRQV9jKdhd6adE5AbZemeDVjAupj4B5RIq7diZp9DIdxHTAC6P8VkyY6gAeZIoa5
nEuI7trf2sNiFIEjYsfGph3FM0dcYa2ATMnA8VWYQF6iZ5qAmhKgjRW9qgEHWkBHbo+qN4D2qaaR
wuvhRWSmFvuUdQMdZn3oVXzAvLjbV04kn+eCWOsbR9KLsBtH5m4sLk2188jydyZij5t9geXC2oSE
+uTXao6N04Cw8K0Fg2Oxepd+T14nB95EbqNXbgwklmuXsZVy3/F0Hzm2ON7O3Idb9rKzyMOwjFPh
9Gc+HgRLpb1w/6+TbWdQr5i6LbLaRFBMkqtfH+bV9LYJrfFvSJR2iqY+o5NyBvU8e388OdSwaPZq
8Ii1avg6aRzFKMBZVwQfzEiDTxks1jf6R5Gwv1o2YnQdb6k6GEqKzRVgNLfdFknNNK/cs6mGDfDn
UnBkGZ0EY7SgX6aw3uiPlxF5ozY2F8HHbXLFGuiD0YV9KeoAyV/9+aWlR5+mPY93vcneceXewn6H
IBZXawqTObC6//RnKtJoHmX7yU9a540vm9qm+66syrHhAQzDhujxiwmslBlVezB/ha81lHVGA5o2
eOMspzRAU/GatbB2y+unVYW3lVngSj8yZtKrQOFGdt/I/1XWXw0TYgrqEtIFaJeS72QNvLSgSCbP
6ivi5EZ69W8xPTGHil4rSrN8tQcgJkOEFuiJ3RnLng857UAJYahjEdZ6oyZhuQSukpMIVeEG74lW
4A+hGgmu70nqpuJKHrzO9YySgWYQG6jHNx0k0T0SA6UX/Z5cI9QLdOMDnzLI8MS5PnYPBUVoDmex
cXC1u7oV5qAjbTudv+ys4vio1SKpi084XaAW7JiQftqsEKkoHv6YMVTZCHaRK+oW5M0MxpzpgBUm
U/lrGmpSOdwafdW+uKn/wQ1n5KRzxIyTZ+ggxVoXab4s03EvXzyyo4Ej4wYoIRdcbqS/eji+iWSY
kn7pK6iaLOjHSgjNnN5RnEqQyl4GpEOUON0rhQlyWtHA2cexcZOPoLBoYWToTv8KiCO5THKxlFZy
At+FBoUhTPV2AP4KOQaMCZwJD+6zphkdijVbm8qwfeeG4CZSWW+HMm4VHjHwsmeUvhZC91ahUljL
megPWdIvRwu6bVEOF8GgRVWVLssb7vK6+gwN1Wjg0CYAWNeCBlc8xBLXYsLVWbFnoMIxRCXC2LXk
lxqxp2i3rt0IurcYchFaXO7+4stZk8H0/dCSVTaAU3XT4VDwt9HhiTs3ZnreyKrAkEEKXW2DrR81
evrdVJpgJNncfeZ+BR7vIyeLQqk4Pos35634SNuJ+NNT/0OyYUzpZOseLhyfJ7eEgq9Xepfg0xTv
9Qfe9o8XiuYw2+C8TlI67Vg2AZ+RXtrkQmg0Pu16zz51wfhESNJfyTR1ATcRlntKd1Hb+T481Rgk
AyoGEGlM11h94MyY++xriYsUKA+j19k2xDH1wNo0U9ldzyDLQuWSwdgjuSzEKTUF+nOWCL9O9Oc0
l9yWZkw4WNT4ln6ugTnM8tFRdVNLnTOhOrclAmdsNaYCTuZyjXJ64NsEkixlD3S2aKA/mWbA63Md
sNJifX1BhcF4QOZHS8gFmxvgdITCWZb5Z+KvqNziqlBbziP240PKs6fmiXU0TjaAtqG2g6LZ6rdE
uAYTZEV9ZRqnoDkatH8onMCEonTkHE0rhcdUcee2uT31Ui2pd4LhvAS1CWoQIvO+ooSdHX9sqf7n
ICM1cr4ejsakLXQRruc1qSfcXWB1fUuZl2d4mgXC37iyMPk9sgRdop+RDUEjQtOgA8Ur+7lU1MOB
+b3zC/narPWpuGrRLKoJZ1820yG0tb0hcLzvCSNw4yMdRgVSELFJS4XTCpUwYi7Gz0/N3n1ztjRy
l2VWk2nthDcDGvvoVdlcHdw4wWSrpIo19Nop6Cl+KTXMK7IFjhgBAUnQiCOl6dBtprDwyMr+Li7i
eEk1ZaesXPeygIJNejnXBl5xUnpDyU34WIjvx/No6X337wmglJ4mri51Kf4pRTZXMZoDHTAtGtNO
/GyTB1a3BeB93CqYUx8MWl8Nf/7Mrp5dwpzMnN8VbutxW0KVWtkMiYDdBP0tIheSyfUCsaavlrJA
XX6/A30GX7R2ve+E66ZINqNvbA7tHKTAOzDFdlN7tq57T9Hh2IBO6VzfNUKgBRv8SFDJ3A6d2jAH
t79+vRF4geqiTooYnB/E3dn7ccmvEd+3BoU8Ziz8W9B4GFzwPar9JXFST9tYiy3F19JKIYfpXrMJ
dNiVSEDdpWPI9xOcvZP7AV0Yg9sEeW2RtTVKHi4hABPL/evQq4M0sIDpmSKZfMnyhOuPxzMfpEki
jMnRxk36LqO6FfhXPxeeMlCGiF/9B5smF/CK78F7nChyVc7jro9gYiwqERZVGopubS8yBFWaEEZP
tiJkB72rUYbTeB18niJvwN6r+SYa4jGo5an4Vu0EwUZwaNGtpHG3IEHZcQ8URBqvL02G7b29LTOd
a6X6nJwvQIVHdiQqmL+SUHzXwKxLjZHJZbjrO4SKksipaf2mKbhV6ynKHVkyPsL8/Fq1QozbFdpJ
noDBadzkbcDsgtB9D3sS5pXG1EFUX09wMvOIj3ks1YmhJmgi7czMeTifFORkOASWtMbRwOP0ckZe
vAVy3gPQlQOg4ftd7CMscB/165Shhd5Et+6McCIwkhbP8xdE8XMBaz9UlUO4eNbF711Al0qc9P4L
OUNyQi4GO1U9ZeD3Xjds0r36Xt6ceqACYegg00TXvgpiR55RmZ0cLokZMfUJ0GW9dN99fFXtflWL
WQv+/nGj4iKAteDbDf2TAEVFyeRLJRAiQKyYr3Ketn4NQmoz+J+KbK5FUI+gRaYQ98WjCctcz6gn
60iYtlqQxXrGkGpB08zPlkJYwhTbXtrgI6Z20dlJiAZYAOKfNqO9TpBOEMyxHDTRBUArDfuU4bAM
OEv26PwsIfJHgEI4cT2p0ivtw3eFgwnJdTOTbTeRwQBajivJLQbrUqOOcAvP/Mz6LzJBgU7vnExr
GEEOPPhTwLDexVfEHDpAYEuAcSAB3bVp2BLVCGwTP9Sl9fNFElRFPpaOQ5R3HwdgBln1G5O3+TqX
/4TLmCg8itnJszUPyMj5dFxdGgIStt+81ufFvLG10jQF/hgzRG0ZGA5s+XKhj/pOwMNirSGGe09y
48HPV4yKUhRXKw1QQ5SyR985YIx2l58XLURn3uLfDextRDUqfZvT53k17mh5W0+kFyWwk2ncQRMX
906gc8Hr7Nla3iEAaL/kHADyzrDX4z7HNGX/hoMO+3/ibX8Bc1HxsjGtj2CWrFTyLuBqyKHbXULZ
nZVnXuvsZhKeLnY2xPqox/akSWONQ9q/jUSEy10NXwzCS8/99Q9Zbup9kvg0X7D2VM4eJNIRxf9K
xM8E0r5pIN34HJ0VKtIk1n7NKebUXhv9sql/dDjI71O95xqS5PlJnRSoSKWMx2+UNN7dUmXtRTXl
UvDSGlELb8McnbwGovbyFK00KX3eVHlv9Pq1yL5DcbgtnRayIW4KVF7emy1bXOx4SR05Ypld+jQi
FZav99ZJhoB236mo/pRWMmttGUvbstXjlsQ7DbDr/vpzySJbW2reBoDqj4+jQNbTikUxmumSdqZ3
0aXM06RCwjjUc6ExXg8v9QucsSUWkpfr1VdpHtu9RhFIunLjhDvQ3ryBBWMZ4WRzOQ+1D43W/dkv
fMNfyCW9ns6c9K6HQvL8W1PhqhT+eOCi0ED1e2I/H4MDJnY+k82oOeksMvNr9JWhVWOAidNnKJS8
Y4fC4+HlVvx5TNCiFpEDciqGvIsCDXYlm+I4NMzyxtcqKKPseQNV2EOk6e6834eDNFizgBCED+5/
AK+UnenPE2XB/GB/sek3WkhqXA61v/MME/Bj7WFN/+kmxTMVBRsSFKxW6G+Pl/iczF8hbOXPT2vT
tPjHx6zL7bYkTFFrYGxKaGR/BrAUNj+01JohXLRy2xOwloa9faJuPuo0rGplFtgALbt4Wr/vny/a
FNSsJwTrrI0lLgUrHaio3XhZVRF0LZVizJaI2cvLvoig/Xd2pdSc5rkBvcET4gYgQ9h8lDn0f6wz
91yTdbSmrO6bVkYVJ1kYSKtxhcFWjTPu6qsLyNGTOGgcahpW2+tEkUCdEjx2DtiWrP3x6DxTMOkM
GQZ4s+qm2B/kjcUF7FlVIqvj/v73j0CJ6d1nV3Pw9QriVfqLtWUWIE232DuyBSsiOWinAMZhQKJG
xZZNVZceTe8ALCbNaQGmQy4G44I//SCqc48jbq5H11+owKQsH9AaUU2PZ6c0rWEwgGviRovOuNjn
1vsbp45CKBab5vohtM6mqM/m0JZB/2kapy/Cczz9o9lesh0iyRBxkSK8eNcFUuYfxRtj1oXmS9jz
xBOtAo6rXJvswqX1hLV9WUxTp+1/U//E7NXT6N1ozQhkAa7gEsivFxEki3IIFeEL3rVcK85qcCHm
H76XkxRIiIYNPcjMDEiRK45BQYGC6Rk10fYMhyZ1o/QG6bVm5zzu0tmAZrOCKZ4p6aMCBBIUbhZN
zIOlpOXaxMYIqTidLv1rFsWHPLSHPMdKzmNQgvRr1IKNKCkSYPeaji4YaiSdacNcQF+hIR5CiR+o
R/ggNcsTqBhhLXfsXDDq31dNSTcZw+1OiQ02Nq4dId+4MZH5rCL+zkErxpJJNBD18y/EIZLexhnu
6lcR2sxG0HMQVy3Jfc5xKvzwU7p0+zHgpF6fvy8DtI94qgtN00tp9UaBOl9N7fN2BTHsxbM+dC9K
YNW18Z3ruPuOXfu5BeqCW6q7SiEFogqi8lFQGveV7z2gvnr2duyOFTkFz6jmCeWuRH3mb1f/VSpT
mx2uFLeZ39l5oPGrsRP5DSvVUC5CeTSRLGFpJJsYMwk99JVhAAqKlVuwA3NoUyTFCL5LiseIvpwz
s/CC2dUK2KpAgfzKChV5JJZ1aQMgTsFbc2fyL1Isg+ELbhBGRUhhkp05BDgVfcsDqLw5/OIStIVO
tVOUuX7P+SHOwWVrcgeBWLFJ21okpxT0gqXz+3iI/AESOmWUR6mnrALJ+qL25trlcUKVCK5WNwzG
ogXs0gXCxa9h3rOllAH4oh5vfLMM9Tpylx5bhmfwlO333BItHEK0rh5usmQUbe8rADiaG9Py733b
scmTDg0t32wx34EcEbgyCNoXakFjBGghgWX1DwCLF5Fipux1JeTWoTR1zRnIGIhh/oExkIgiGJ1n
Ryj/d7QnnIM+N7JlSgcLnbhzWYXE04DdIxy4TA21eDyw0z4TuVQpGNe711WTGLfIHI1s/B15Hl2b
g0ssi9BO+lHzlw9hD3LSbJwjzE3jKYV1kdFtwJBsIz36tzz49+xNHEXd0dShpwHJ/yocDMNpKex3
F0WFdXlAMbqO17lNchY/wy8XVJhwAAVnrJcG471QjScAljvfgyaryzFwQBJzfpvuBmp5HrWbD5de
3N1XxDwhzOpVGLrraj7I4Q9ic0Qo8kU7I5ALzFxKcQJ7XHx3xz2JwfyP4xhGBchXexsDjL/2UazY
ma2J7e+Omdy++BJOmX0Y9ojMI1bY5uzd2HYX0bwvCNyuferLvKlq2ZnXCwldDIZ4FCVBOOlaZ3gR
yia+20o1iCm5jQaBjuI+doAo0okEixzDV7QIWMeYmHPgFroC9f6315+KGnwQ/Mja24NonG703gzR
wg/V7O4Lbfnga/W6JT8cXF3HPme1VBDFlz5qn8z0ynJqWl0RtpH2EPfgxShBUrWBjU/0jEgZRXXC
qido1C3oWRK2ipNML4daRrgQqUHGJfrI3h4tEc6HauswDY78//7F9Fsoizu/uCgqTq1CgcmsnUp0
/bvYsrip+AVWsEY/0PU6/5CV6zNzRBax7m5Hcl8eO3/dGyg+BTx7ijZzhTLuCORmRy0l8wP5+LmO
0Bfs4cu001YtmvXIdBfqGpGE9ohlM3y++/Y7I7o9tBlWddQFvOuRglmWYoOle1c1FZ5dCqqNPoNT
9OtGdNeL4YEg85UEgXpFT1asGkposlQ2Tiwq3msm9hqIHU4sm7zAuaB5GSZowGsmXz+ue7/ao/sa
RMVa3eoR2iDPKl9hLqtC7ITGS6voqXqiu+dMPli6C9AY0RjUUv6IB85Fnk7cqlEFxi758AMABQRs
PODRKANJXKZxESzFKqnRb9v8lVBH0ccRYmFYgYPxHlJGQsBEWw2CeRcgbO8OL0KQnARFZebYgpS9
I7TVM2E4+LSSnBjrc7Crhzu2t9j1foOaf37SJhxYfQFsRCF/a004F8wXnrRoiCVReyR5QDQyQW8Z
0Kzi/0dOdaGXJyM1rtpLvEZ5HInu5o9F5pUcox6Y6DlNTTxlGi3ZIv57+ms1wSCt24KIsC/Ev3PK
ShdGYanhAR020KGkbqRCgEYNV+hk5ZK1tcwIX4EVAkFLTG9iC0Yh3ALz/sjiSXt1fnBDb8ATzDCV
B/kDKJtVWBMebBqKu0+UQvFs0IOlWD0F78Of+v7vsTxiXHNvSzAs2S3t60jFIHwml56oWqIcAJxv
ZoLnugSrPLIccFAsOMGn9oaZ/OqolRf5zN0jvfZErb/hyNugfO4KPlktZiQI8nwhwGdPupVWjZpv
MpJ6shOQeWcxz+osOYeCQQjkLc3AbqWAlh/X4l+i3z0HORVqpyBsmg3L04DlHW3+c5AB4H7tCjka
7FIHuktEVCZed7+6eIcM9fhAapfnX/tc/isP/7LbOBJenqjTqAYjbaMU/zgNVk7of+Cdz/q8/ubd
5UFSao9KbanMNf3oIuOwqGm/6CJY1Ffb7zk7ye+OWtUmAUJ8I9fJ6AAhAWyUEuGIz6iCyagZ0Vih
3Kk8vojLZsIjTLEUItmnwuhIKvoyJhtN3YdMQ7m4LEhfS/e5cEnxdrrWaFFnsB5Hr8pXkimypS2c
bzi/jZmxR+nqGX2v1LtIKreJlIbD0dXGVB6jArKpPnM+MoxPEVe6WnRRChqA+bUwGOjJMPkt2Syn
4TDXbCo1nd/HvxDlMmHn78zre9ix7QTwmb9qz123XFDDAuh9sk4783mAWGXKASpD5gdw5elWPqBf
HKO+ZAbcKQ/NY3m+Eq1hIbk/UsD4wdf2e9/LHvGjtV9yafTyywM3zZ+OZjVGWX8ioccRyVDPg0e/
QDojjxtaAOelP6796hhdXhpKDt4eUZoAqhi3cqtnlGezxBJ/hBpDzpRoq4KyF+0QtjOGFKbm5slE
q7Ltn7aWDKkgTXOJN+7LdqxHvMWiIAoTqpbs+yZsY04TZc0oPw9l4b47C53oFFsVuBaKGZ6B6XFZ
8W7ygt5eCCE4yxJhYVcKjafDrtmBc+y2WMSg/NnmrSyYkMPu5+cJrbYg9w6SGz9ASYVxGdRbw8zb
ck88uZ3nMvFPFaF2i7Zy3X50cBunToEaIBoNTzzebPTU/nWoRs0OTdr0JOREG+rpkCYsAJkkU/Oh
MuiBLHlFQLniUEyoe3wzl2Q6RwpgZL9bNv31QUZjkuCDbGTztwZ1HuBDPmJCrCQL6ipX4tfnmJYD
QIuH15ibydqkOxkHPmjEED2HyLw13THVEhOToWhfdUrGkuEFNJJhYvZrw/2+YlBceelTnkx8LmSf
3yYzhKXfbCdr9If+oscZvGTOBqfXJ0kC5lzCFYFfvTq8gdpdjaYgzut6Cy/YVZgTtQqWl861sgOm
FJ1sTdZxwwblET4Pah/94uLh6WUsMPdjyA6K675sImUtJQogm1HD27DLba88SNcWdXGhWN4CMw69
RNl3R8yJ7JtOVAKXEyteS2H6myOzRg3AUIo9/LosLKOnXTTcbJ63RkiFfMUx5i521Z+iVhKBLEgv
rm/4X6LYMhL+q7lWee26DJNKaKzc17re0TfR1KB/sCepnIkSoRYjyoGQYC6mJwZX4e/q0pwVziLu
JtLcnkvJbAo1OAQyMpsUP9ui0JhaFYiixiLQAi1IktkTsqIGVQ8LJ2FSZv+Nas9q5Yf3rX55FlxR
kIxb06SGi4UvOkCKFqRmqW+dz3qoM5SEm4UrfUTDlJtZyzEAnxb0Y8LBFT8K3sv3ur/HfMEgo9Go
nEHgjvz5wOdszH1/JtqnGBTLZmGBnIlNLbEiszPluLrG2Zdpx91pP773+P53ZvB3A+lwVOXZ85uZ
XlHPTdwLLERo7/HjxycmixRTWJ1VPhSw8JGSI4lsWr+G4P1gdo0xVkKPAXDXAF+UE+x1A0EFE2sx
jTsod4tDxNK+NxB+5xODyq+9601Mqshs3dQLpWGQRhlxCmaBJ/yK9sLyHCOk9RwMxLfJbkXVhoXl
gn7FRkPeEWbb3YQNfJSoMfsYPZEL4CAGjRHl2QVLzKJxeTv3BhlBohEHFnKbCiu8bM6KIOfsbTYK
ZZHsjNL4I+mrT6BCkwi4Pk/0FvJt+0QFuqM41csU4WLfxSgqH03q/UtBt4k8WPuep+YDfujX6w4L
IeRGUvm4oQhYoe8NcVlhy1vMt4EikK+52segY9JPvj7R4vyZNjY8RaQOyNP471jZaJTsQHc2GI/X
OiPoUugzWM84SVN9/XyVqYaGsHDw1g4FD0he8GSTIZUQyGLSZNEjTRMc9uOeIT9XiOY6u8gv7aBF
+KwkKXb838Y85oPWGcu2IPtBniWnktcXRd9BwWuT6bWKmXmzczeRbviWj7XGLEJzryOt97NjLSDK
B5fYYEWYrswIAs/vdqLEASh4ZDudpXfdMbZbGb+GkKaD5KcBptElr0Qjpxf36CkSmG8xn/JnH5xa
/FmXzXnSfFWdHRlWxK0M7/boJYpfcTgNGRwFnm5Opktx1KZZxAqdSHFxh5E7HOvDbBeibVPt4bPv
8xA0iCZcu8jwutBzOVyMdh+uf4jKyzEz/AZofx2XZ63ivrrLiUpEXwU+0LnzLIgPdxBRk11ol925
88YFqYTfE0BNfFefdlnfWZSZ6ZeZPRbW1OOnaK0Achb+dLG4nSrvDGCY2S5JP9Fg3hxM5uyShX0C
rG+CcOLr2dw4ylnDwcn28dFelQQQepF2R5ng1hkfP6bszcNR0sBtyCW7m6baPpsa0goZOpKhK+nF
lzEPtVqINYz1Tk22+sNYIbxlNn1xidU8854KXcdwPwfXGPaA75I44KlM1fkHcPkPouXsWJOESjGt
mZ/9SN5E6SgfP11DGzvws/MqE6o9jVBnZ5XJIlVPs2b/o+u7d2W5MKN5534dxx6FvPdNyKEu9ip2
IiVEeDdukZpDShja+vYydrQcBnoG3oJdzeZOmwhERAR1Xo1kwuwjTWZXQngYNzNkARsJmKYBfwZj
WW7W7jzuM19+Ws7nKodlQFl7g1HeCMMbbs3+Os0Oyn9ctrpULKwq+fqOLmnPYmkaw5rGCOezkW3b
6I6OKTbhMgomKuIKGPhR5Yv9T0Cyr4S6KAmzT4OgWmMpV5nYnRSNPARA695xhRrhUUL9+jzdKdDW
Wj2+45ztXyNeB30uPdy0tLZ8jgHDg6sUsmboA5QtmbSDfgXyUqKP14ibQA8632coEfin8ZiArbDW
t3f4awy7XN4NspuDyWtmFsTA9+hfpLEfxs2Sityyd5HfdtNZziPgvHkIRIOkNwHNhHxqMi0Kcifc
/BUlUAwtAmQ5VKSoy10bjTwsxQhxhboJDoR3mayqrBhZkL6ylHHuEafeDxJ7YGF04Sd2i2a2lCxc
RDXtwDohJORGi4usRUDXPrbq+MYILgpoMZUrLOkZBuWoVjq8RObRiQq2q1Dsce/NPUzLT69I4LCC
rnb0cuEEtZOR79hnj/y2A9e+hqNA+ioK+stly+BEQgwQl3Reh2ZIiyiGfqeahbWOjsR41aq0wKuJ
DCO4hIt8wHzWweTNqVdel9D4qbgQPyS+Vwem9lluRpEG/YMWOAomUbDNRv3vC4PWqvWuoeXXT+9L
NCJowjrLF33/OhiwQQO/3CTEkCTIYSc42sOwfp26gSgLo96ogQ4UZ6kVkO4OR+M+OrP2ujVpO5YC
NJzQRZAoxvszTnj/kgB8Zqs/zrrh7jsKv8FqPttO3rbvfzLCFcI3vByWInZwkfU5AuI8GMH3Y8RL
YomlaxSp5zcxyT5H6SURMJjiW22dWY9qE+6yJjcyG9KEC/39GSYTStVDZ5WJJ926n2Cz7uuzwvN4
vc6h7uHzUbgOIG07oT88iMrpzcrlgJbh3NK603NOxVLARkAXTJNmK+i2QuVfCHx/FabaKbijlWs6
tYOw9mp9XxmJVGsYdW25+0jCAunoSjKYiNhgeMYZbscP3qzlGjtnzDcW5vrfDRJKJFQgukn9Kme9
t/seE57RK0Yyol/jtpbY7apOTTDrALPr/8xWf5ZQJigM9Vtj/6Y689icLdlJbLx0KClN/hKPfZcU
/72s1sPUh+it0yuhGEvGMuGHAOnuKv3pV956cTXENy5dYbwkVLUcQWhncCSTG38C1HHFwZp2/51E
trQcjlDnlE0046TFogGXpETD0+6jvYwPmYy6H6V0+8RwpzpveXK1yg6zDBUsdkWN00fxvSsmBktz
GqQYkrkeJbybt2m9cDHc7IMlepKQBBrN467aDtyBkLzG+xo70/gnAc0dgoceul0/bDEYAuf74KOH
SGVRKxxHW4wN2RCKBKqdeCnQkqTGLzdX6FZgfRr2DOp/+Q21lT4cuzYOmZG+Ei1L32+IlrdCZ7oM
5bz9yziECPtwJl68p7ZPldV/IVyzmrMwacbTzeXQwt3YD4Hp1KLI/8rYrhnDmU4hBT2u5HSz5sLR
NmF2PQmUWbCuc/+FVNrulylJmadS33FTtzN2wGVLDhFdk+4uLu86YCdALDnfhawv1x+gO+/OXvmS
k2I2xtYHlTQ4lEAWPj8Gh3vlxZllfKms8jWYgKKIelF/frjp8QJP7EwtbRK70AZ7c4n2SgIR/SNT
0OeWzz6YEwu6U9RNyaHEDX7koMgdbGcHb9kG/UD4ovOtnpfTgvgabBYp+BzTDkd8o9p1CcdtLtqu
3LXfEnQbCyR6nGmLM1RKH/LWaq1aBdTB/h2RaCUv+/NQ/wh4vsdZHma4BR271THqyugXReSIFKxV
BZ0ZflknnxOGatTh4yU4MoRkXi0y3XUjsURBO+V5p06sZ60J76SLWdkfL0z2PFAZeitKdQtGrnPL
64SwIwaAo5+owv0wnmrk++n5NIOaos/DzIF1b8m1H3VlRcw5KPVMvYe0xHSKQ1qESEf7j5VKfGC5
AKSQ0NnQvX+9ooKDRdNdRtqAhbMr8DemFSa9W9xZ0oR/FktirEr5Cpxypr1eWzUTDPkRlsYc6i0/
Laa0dkR/dsJq87qtedJRUo27OL9tJDIEsB6T8bdVE9mSYLjWIqU+5c5RFgiN25KK/PAuTBVo3/hP
KBnk7LeI+FtXC8ULkiV0sjL76jHrEiiG4PoVYZLp1qr/z8bWzz7ao2MHDVqUyMRk2Rvo5HSxX2Q1
bvp26sEwBBJzSp1Vd70f27ZIUUqGEMHTX6dhDB55E9arWa5J+ymhPNC5eEh1EY664wXVd/03ubpA
KzEg0Md3nMHQOTuL2+8zjkye/JzGsIvzn2nle6QXWeZyPP8OZwsYeU7LkrxEMwETaDK2e6xxAmOi
SwR8h0dnuCP5TEsHQyxI+v6OIDVmcpYi1PdNk0bMp30y5kiOB1fm+4g3T03lZB8p7tnepGm+czAK
pEzUue6CwLjlJy7aFE1dY/XCfs1ZU6B1K19P4ddgP0ubF6OdZgP3RoqrTDzN/Uk+WFEGCRDjIhpV
3bf0IXEZ6i1rrmK0rNu3TtBDpxbPuhMCU8KSpIfUW45JWEfepWvrv0/+VqiRTZOZCIt1GyX/Hgkf
PjWXlJdzCsMRN6JP//th7g5qv/diSCkU+upO96JxS2XmlUCM/aLF52GLJccr/HRid/gzvntyuiTN
bCaFO89a26V+/4974ZUVT0NzBYPRC1zYlHX8VNcMXsG73W0MURVBSEJMpKuLqZSio0L4yJG8BEeE
DmpLqVNoW7j3yvKGodqfhLdtyytA8K1iS1vHSS/n/H9nr8WVixxhPbTuVSMEteVxFbIgCa88MFUS
IR66ZBzif7nIwhspT1g7zXoMjZJPRz5l2KZBryuj2j1owx1hUG+psP6I12fzBWeUeBZtu8YJL66Q
L7tbiBpRAn03J08gLrz3Tj5Swk6Wc4BgmlXNheQfa+UVrHFKI8qxlDmgOnPATZENclYGMffKltfQ
Yzl1C6iOQcEjgfZT0XGM1C4bH4USSdkSN1RhetpDhrMvOiNJXEmTyqge0c94yylwiIYC/xe4UeP1
SkKd/E5kymr9t2ec2jZfBl35DOsh0AFCqSxJWwAoMcGsXtdP40pujXqt1r7XNHLCzlV6WecpY+0x
32HtQABSvYb2egqFlDjx3KBXwrfu5xNooeas4kiGJzVRKJn09UG0IN4A4pr5tFL3ENrGPJ7xUoLW
HI7zio7D2NTeleZTfNJrkF7P9urgXU6P309krAYblRL2fbSdNo/EAyO6Ys5toT8Pd3d3X4OoEe4d
71KR8fjOsaHm1karLUiU7W6c11ikIXE0xQZMjRbsqf72vwUH7aBOGTQNoGjFmcTeCe5dyj2oFb3h
43xBX/486fRlQdFJIQZZPaf8LEatTq3yXOZIiNcLo+fxATwzpP6OCVTobFEQBxuuQ+XU88yF/64d
lnjE3OheH7/g8rsw39PjOvuFa3qmbGm7iyfwU1T/8DXEHiK2izASPzDqACIBkDUMAXlVlndrJqnz
AJtOusRAJDb7wWH8rdis2RLd68hQV4/g+SfP8JYy/Sm0PYCCxhSLKtWxrs5uBXzwGsmauNziK31o
QC1M5RUnmqCrmWZ4kO8C6AboFL70Nhbr6C7DWhnslNK+LmxRrp6SKYXkLYX+Zvu47uWTl1J9NtfL
wRgKrZjeBwWgpG4CzXBsMvO8rB/cK4edHwy17vBYFYCiVfMQwkCd4ppfWD49qwnu3+jo2jtM56hM
cYUk1I4DSYsa8NI+YsKXC2BLWdbLi/9XFZo37RrNZCOPjhFWhX+NGWDAWI3pNSxOL64AJIsGk7ev
7TM3Uv9Tjrrzkuo5WeX2L8Z9RwFcJ7NCDQjD8R8oFJlgSj6r3nDG2iUQIevH3oH23EaCIevhy3R7
wE11783L9jQ4fvzvy1Kuii/N29Tj+brvbHcoVr/s7ySiQI7Z6nPzqw3BGqHtEu60G12Fh0GG7fUI
rjdPwgF648Pmq5OrsPO8yPC6MRkIvFTtewm8pmIq5ZSmQjSW1szX5yxcI5qU2mt4j+ssGZ6ZN5sq
Tt+axmovJgSZyU1AxTMUp9MtPhH/L80TQ12T+8gee10fXmNuFVubLsFP6y7a4PPPZKyST8alEDAO
IToEtypmPqrYLl4y5DRMHCRee+FtPChTHxnczbSwSthJTfVY3oGXzkymqv+3jqJkJvdfZe8mEPME
GaiDJX8lg6i8yooMnOEqzMOSERLsUo/0tNGdaw42jH0m1cseZ5HPv3VhUmfZnesl9LP5AVchLi1Q
lRZ+KojqN6wG8wwXCMLf5WXP2lDxMQ5Ya/B0/PLVVySedhk70V48OJqrLq4/MiH1ZOqy+ToBFKv5
nX1fVmg0Tg62BacVTx5lTkp1Fp5esnsRnkeurJ7VjZ4RaUqw5lO8X1EcoQICWY1M0Svt0u2qznxk
eiTQLA+9KdTJrFldRBeFNMBwIN3KhgCrB8pnqArmJqh3YNd3/9kLfPEkZyh4W8Bpna+mKXXLW7xJ
ZVu9zHC9UEHIaXud7K9Mq2eyvi1X8NvaCN263dGbYtsLVFBxNwpi+f5hiFMGhtygADcVo/I004OA
pHKslbcvo8T1cryZh8jfZ6DQejTxDRppBjNiM5TBczkKyhyPWBql2+oJuEIoDE0lzrDNWRAc1Eff
22QPis4xZhjiv0owz9oVrDvlUAEBtbBOoxinfXXNy7734T6k8ObpvUjWV8H02XpIo/vKMS0vXPn5
ALjreGgVkI0mDEzdDP1jHJsWjeU43nsi1xubaWRX1SHDLOleUKGEm6ptEQBBTT7+20D4nbL65ZEx
IWs3MIIc14TLnwPnZCoCBPiDPmqRsehL2UTzTBRgsTbuoNUtwnyJXVnk4FyZIaNl4QxKLGGFcpL/
egzYPIVya6Hrste82oP0DMIcN9I184IsnX2jklFhc1j0e0fBOCHxWWfaq8zpoBEkp4Ej6U8W6QRd
kjv1BJ9DOdAzy0z2aB871TwMN7tWs0ewVmWyJJz0KvCgE7zdVMl2f6ONRsN6ekla0VxxTpQuHrGy
kvVmrmhJ2P3cPHc9rrXRMSEL+bCJ8Fzsmr4iZVBDKvJl/amK4zzr9a07S5nUN8CDQbN8+DWJk8Pz
iR608li+DcmAQt6WuJ/qpJu0vQYDo5+DB9xJggvhXTiIRz4XG+dTsDdpjgtfh9jETlEvQIqfVDDD
r14FUtfY8uwUb/nSeeAiE+jiaGrhDpYMXIKHc2oJmDe47olPNd+Vg4C2L8pOjKDelgb6IOq92l0s
Jt4NVQzlvYHbV9FPmNR76qeaAT9sULkUugJsUdusaYNdinRf9QgeZReRBUPja1LOApXYNEXUv6XO
nMaTQbE2qoQHFqgF3BtrokVUcbmysCLe/EE7z/V6eQ/843Fephu+cNWL1Q23huvGg4QSU+1tQuAM
4ZDCCAQPQycehXV/jIMv4LDnJMGbvSAyoXQg4uF262CHwAAFWkYGgYJWhMI3ncg54Doyf2tMfcdQ
7hgkfLDfdS3nCZC+U5ulbgqrYflDiy2yodVZlY1602+h+7qG8NZtw/vD4LuDQlge8plQVzBL8sfz
796u1R34HO3lnDdnI0v3NDrT7W8EykEzaUhWvgZ9z00YdsbyuM29+b0Oc0KpukO2uyhAR8KV52cJ
3oRNvmUcb6LsHrnmNok1125YPlelvnq1dZ1Bjghcv6Jq2cZ0xV9sLD1HnH6izJh82m8rg8sN+RpJ
cmv/fC5RSD1fv8QqaMTdCy0yYAx1GAeniIIrTJS/Y5CBpbWi3/zPysxufBy1zfKpu6mCBz3OTI8q
zTZUj8WhenQUKTdoR7LJ/g8CJH4q6xbPLlO++NWtcMyHf5g+JY59HqFEOJhdqpJw2GI0X+11blYU
5Vc2+ZU5LoKtoY7vKZmrmmY9llre2Jr1foeDF3EJsiWcSxi33+yccnRkX+DFDkK5mFkfTaEC+DA5
Au1qdML0Ss+/bCzsvQE+NoO8VkR04xuv9oPm/50vNUsEv5y/1+cRXLq4hdZQyGn6beOg71VAhuTX
hnwlUnUaMaZ4YwcrxVupAjyhwCMZrTz40nUGElhruVweUSFmyX6ohK+VMQSYOUvyFz9/GYlhon5L
OJ727wt5xWg1GezRkR4ATqXSmo06SzqjaMtyRwQICEXrxgF1NGtpwv/tr3goDktMLJ994HL3Vctn
Tzdh7hOEdkZ9utd6ZxfJS4IhzK/pr5ruGMIPpH/6QFPw/Qym1w+28TXkr6AQgQJLtc0vxd1jhr7P
PqKpSTnZU+QcZFLd4M0xLXgmkzXGJXb/6T/S7/XSZyiAWC3Yj0ZwGwHhHxWvRqjE6zxiIXcVHw3E
Mhk6ITXUcIzweFmyQSl9sgoQHkTXLsjI8p1HF9N9Psod3ps3u+jG0P51BX8Tzpf4S2cXilnWLiEC
35vImxhR9UdwwiQTbptsBsCZQrWXeWw4U29VhPRu9xmMH4KT4a6qclCkWR+Eyi09GdWskboCkdAn
+ywhwLxM6XvigAOGVF0V0SoCOZHjv4V60cEJUczaw15PBw2exerYB107e+Ppyj1MurUMeS9kZ0QN
QH5xlcJx+GN8HlKuDSLZMKwnk4tKiyt+b1DIq63G8k8sq3ibo+ODqY4yKtdh+ijYejEAI6FmKTty
u06fU5aTaxaSex5OPSUd8GRzVGfEbgOFI4sMQJztaVdgc9n1yuu6W9VGMBV3c7EepKWrb9v4USqJ
FNEtUwFIR0DtNaKXX0eegL5LCYcMLFD9LTQTnkNCqoCY34yQpxqtpRh+50N7Z+G01ct4Oub8qtx4
2wggoimBudonhVhvLIjwHiB4xbuNF4JEcJJliMoAyNQ1V/24COzv30MdvK3l5ftoT2W7qQls7l/E
hlwz0v4YgjtquxIOdkBBnxC9CKuFV4tzSnQFISz59lG1ov+cHEW5gvz74Qh1bkTNor4ZKIuST5XT
nXTtvc7XcK+FDS/yVKfWSqngf1pTaIKubQkZtL0EdIu4zfT+POOdLzJLRzMUTy792sW/ynOOXaEZ
UsCbCg5pQ1NbTIlIpin8jdOH1Ie4bu25duEekZQVZx/0SobFm5JQZmev0j4lhUkAldcwz2KlchLF
SqjyOaxsrpSkqK3sjAgyLi1H+okenhZMRA/OPlPZ3S1qkrC0R1wpHFwlSb/bfQOYISrnGJahQyK1
TeFQPHxljurHOStMdmgrKUUT+5ELGyK3P5qGvmAseMUQ2HJwBYx5OZFS1iDdpVxvWadsv0NAAJWd
WeT6aJ7bo0FujQWAc0PJBTOB8wXBvQ/uhGLUsqGIPajW1KQQM3XL3Y+NLMaJpHGXPrPkcIkZJIH0
UZNAjhLjat5qj1uEQAl7jWnEL5bQP4Aa7Gn1yltFsqnKDcXZS4sCcUyyvFrT8R2DnJh7JdoOqHyO
PLSjJOXctlEVu7vl4cpKTEXou285WVhJinuAGdHaPj0H/zNGFIEdLoLm+iOLBLAvOi6c70ME9q37
1Od7Mnzsj6HiOVNX+jOKNmAEBUs3BUN/PgMWlhwXbQd3pmnsTUXVQhQ7U0xLJw0eGfLcIJksN9GV
0KKHTnW9INKMaA1nFT+Vh3uZSdCaAluLWhzAHabn0ksSPhKhBLwzOwD/b9foAYGcYqrmGFrmxLl1
FN+L/4il8eHGSP2B68eCdzl86BOGwUwDWQXjZ29YPRoAool94Q3wzC6UT4D4Oetrw0sCjT+MZ7KB
NvO7gnvqx9xPvC6Yh1NjY0gihMAJfJx/2rgEbtTqi5NAHMLZO028+Tvo3efSoAJp/P06KJv2Yi3v
xcvDc1wFv+TWAq0eVfktbU3OpslMW04U4S3xHNU0k/6N9nSVcEICsqm2lyLsRmbLm/GVpMiihiXP
XprHOMFc42XhFwXYfbRYUXMEqm07W3QgL2H8mWghNAJb6Nthm71fbpOQbmjE9zTP/Y44NRe3CnMv
3eMjjqx0biejZ4h3hZw+LfVhedKQtBBKpkmlHRe1wDMHRGuX5/2vKP1Q0FGbWKKtwbxkul5C4/ru
r2sJuNOwPQVaz7RqFTtNIIVyTtioea5xHax8MP3INgG2Hfgg0Lph0wiHzCPNbwWhPZkSYw4OFjfJ
AXSdIttm7Fr0nD7kC6rsML9YlRLpUfTbaetCpio08pa+QEi4DjvYBbDnkw5Ll7CYAZCAegtGkPa0
JBqOAbxcrWWSxmITqaN2ta7RL9kEJT3ZOjnQmoRLD1hvVmM+8Y6Ztnf2eyVyveKSzxDCvZqF8HDK
xTSEyFaYpFTJYNgLqvInVsxI6e9bXdJPx6OLP4x/Gxa8ActbLOquqQsGzoWMGuWUn0VWTVr8JdKm
FmeohPLePF6QVLe6MPsBNMioQKXzyS6pfFv1eTLZ6DsDoZYQWeCHqyObivZrQk1B4F16smQGiAUf
m9VZcRzwODpoqhlKgus5w1nK7gjWtmkUcPJvRQQmFRGvquDpz+uJ6cW9SU+DT9oYKrXvElDc94TI
ZVlH5HBfpUYNUcC0szsyx0krzM6oeqi/6iqO6u2cuGxtWx8GywXfGpezcHGYAXx9w42IepzEecPH
30CL84sMrWnxfRHG9ZOS4oKs1T5pBXHyJDYi81QB0JhBPJhxA2M+9icIxB7dyJbKkOThyw6t2PhN
Hxz4WvS4DbWbzzbxlX6GmmH9Eykg3k0bfeRwQXFmaUACAsGf30JYXWajsktOjavsUhcicnU4psds
tFekYUhTWQTsTl2zV2QkxPF8fnt6t/F+Z1qmstzOy1y67cLfgBp+BzMTGYEILUnKH8kLQEPnRUGr
eHh2x0Pn3tAqWooYoF+90UQiQEltYt0supri4lPmHjTUTllnjFwzBQgr9vHLl3ZTKJTstliL4qnv
u369DbnC1wV0XI+gzLlBeQzqL44Vd9di9hVWssWYTKJEcxgU1Y1V8/udXmSyfsLdbGMHdUNjDXR4
PlOppKFEYOkJw/bT2gy0DdkAPi7C0lGF+jkMYA58cauR7cKSCduEVtUSLHAGunHXrfGJsgtVYdAY
qFMh713uwBX3TekfDytFzzZ73BHwikZOv7SBqfbYByA0/It4fOe4posBTXlWI8gKVxjQp7HYiFKE
gvfmwUns+bSdZoIsSMNKW4JUcuzF6v0bzAgUFa7nIG0vxQheCklxiW7n29dktKBOR3ugoG4pSf29
PG1IdXsgw/Jm0W/iXFE8DMQxQiHgETScsP4RjmucjAn9ZeFbgTszAScuCC54gi5Hhrndnq03o28E
MM3AZ0C0mHgkDAaGO1pz6d4/b97YqXVd0K7x5Yd/yPrENDbRyJkBxEIDjj9r98irOLqe5cML8xbA
Z7nO3/5qHBKH7Aj/5DBks8NfLBsLWbFEDHWlQMhcHjxQhRfb3yta1F3xdHEXI9yoCqQp6PndrIMu
KPcMB6v5GOkvjDZcJnchegp7lBXQ0bihileorkkYV7eXDTh5QTqeaxmcko9RL5nYXRUUkSFYGQr7
JCtSJzLrgz/vc+jaRJqz29ck+dKA91mfzs+0IZ+9EwnFuzHKbVZzYWRb5kLUGgTsCqFbsi3jsHPj
pv2CL5cetOceguqx1bkjw4qQR2ziVtfHjIvrdp/bR4YOHJWQUV7xBzvJ0Qza3tAiNGO+qNBPjRjm
kHPLRtQ2623wNe2qtoBp8pYj/Vk9tyEuSpgnJqZH9VNqg0tGCZtpEDiWWVe6kLnNQvuk/O8HXLfO
DE0Rjep8hBHxENZu7zHylBaD0t3A22wzpbQKybTekYzJ5a1VZqsgQE+g4om/kQYsdW/QsZfWJdmz
HEz6QSQVPAArElO94E5uIc//NI4WLLKH79vdMjY83SO1AVDd7YH1at3RJ8f9vMqC0iHe3JhKWzJx
FKJDlUVz3bNqNXLkQqu+Ki4P9ZqU4iRKoWMj+inbDSfVNqvDPQniV/eQJBR4krmJlStHrkzOzWhQ
SuYaNIEaLfky/aa34WKxDAExhTCr1V0K6fRUyREvu3vLSjH0YMqripqHP7ke9ADvyoi1O5IzIacf
M/PObqsixnUDtWBpI5uPYRd4bk5ib0d8b4F+xlkJPeDgKo51zKMPZtzs5bUedXigeOzb2wpn0/Kz
I6Bhr17b15tgQYT5CxFPztqrwk3Y8IgCZf7bhmNJKyS0zc4kHzsfkUNscp7xw7SL03FCJygLmXzI
XhO7bnTB0n0F+Kf01OC593wMYkRuq+ywSt4tXxmXfU6WGbHYmZGCbWyB71O7Oe2rs2biOXsYKQBV
gNYHgBKMMyKu2WcLuS3gFs1bFchRCsRV2W1Iqgho9KILntvXTpxGnn14BI7eZSdQK24FAcHDo9CZ
IlHOSKau6JHXaE9jLgDAZTN50VbRyeNsaNPYP7d4mFuv4XM40Xjx68SfauWcSrdmON99j3idDzBA
dhJnkxZmt3misiJZEVqT5O+h1iBQxj2IPewZCwfRoSpBuQ0jyduXvLGk3DuA0yNkQ/vFxRv6agWD
afz4wo7bEMLH44Iqd4IXk70lXgEr3/K3AYQTfoG58+uqm8TAliVnade8w5b4/lPSZ3T1EZU/1YPh
blna/Xclut9CQ/JAT32ol7ezS5+sD/A2qNka4rfqLDrj5VLSNX1PpO7RCupCz8oxIDnkJhYMvCmx
RG5y5pzFKruB8lDQhDoEh/cLhGmSmjgs0C75rnBsf1+gHkX8gx0E5qUu8DPfvvCEkel4zAjObSdL
afCXnxqfFVZM/Khv8GnhEcbl/FooVsjDEx/nQh0lPfHCIpTsnFIcOzrda4jkhLWwPb4kdB6uQmrl
zKiliFrmc9w7aRKFBxXU28Ne+OF9/3AoSyaX6LwOupMzfV/kEp8Iv+EaCDF9a8jpQtUCWzy0Q4aU
9NHvZbqHr4WXvXE3/bgDfNav8rcw6b0P1mwpK52djZ2F05BQKXcji1FobLH8gDPOtiRBqu3kHUur
3kCPc4F1Wqkc47C4XZXclNGtC6nxeFzYUh7MWOh0z2PBLC40aS/AuNegkis6/EuFTEHkubJC8EmT
RRs1IXrnMGMoa87KDkfFAA/mmtDAqTYBlquecBNEsFLdeL49mrTvarDomvnnh0A+AjAF7tuoGbS/
k/uDY+v9Tm4bLNiLFZjIUiUOJNWO+3wLRH1kJ3dNZTF7yWlHC/E7ReoqKp9Pxc7MJh1auyE81hrm
MzmGTG2vnLisVuRXPuSyPIXpsMoRT/bqRn3DR+8ecIUsDY0aLWwmQhYHrcb7LNv4x0aGWoXM+/9z
i+fWsw6lC5VKPHlyj54U8reBsyvNT6sXuFRzHn7JvNYBs3ffndt0lSQbVpYBEQKZ8gDSGx1rvGIw
U1QFmTWMxzrHI7BFnbY4YhyYlk1zHW1KWX7cfaOdvSh8m9ESzPWaTbynh/bu6G23oP3ws8bH8fzD
fDSqKgIwxkwmQyONn2CQ/qLHBQO+35i9SGWWg7nYg71tfKtTbONSRNtgBsJZa5Iqx/x5UXR+OjGS
lNk2OALhMSyLqqCUet4o8cglQ+cOvQFFTV3BasbPL9vJtdVKAzPUpxm5mPXMJwxeDTBkIuIO3YnW
LkPUGvPjEqCZdUccPXYD5Xzd8wNBSvD8kXa+XmPtKHHxLRc69TSZiNNBUE2FzDSR0u4xnH4NjTcN
oCiCjkinVW/qn6RiaHBWpahSnEGaMIKVhHNinH+QQ3vLaQ3KnLw/R3gwcyuO+6hB2JTqA0OWr4Kk
V1tAaXyb5PGuEq+rlrdQDyiVyU9xgM/+xwbx3xE3En6Bid4i/6t2VGFqinKtPi/bhSqHKlPTkdkt
vxgtqIQrcAtfzdbuc8jyb6/qJfje2c05EdJ8bgYS7fJdLZbrcyXeqS5GrbxUq//KDy/PI7qcZvk9
SDP/YqFIYydwlRZVS8y2uLXZlLocbnCz/8PSq6Y0fMwkw+Ggk/26qCeavh08fsuWikw5vVHklsrE
P+nb8GnnjbP9QVW30ZP33VW88t4LIHVjVNJi+kNU3MTjYJ8gy2mao6j/8BpyLC61DD7Kzosn2s6p
n84V4tIlAZE6mcGReyJaJ2uNMDLerrJ8FbuD6fH28cm8s5Zeych1PdF4vpRkN4MjNvBrUsXdl3dH
WGsjoYU31Gc1lSn+PLCysuGiXCOWBAJ8dy1PhZkau+5vk5I590JGOva+wgmiuM7HZrIJksbqK3xs
iPwoXmnzwuH5kw9yTtva3CcyCKKNsTZeGCeBfof/KRhXwM6NmHfryOMigwZFE020DzgIxI9Rv3u4
++2s5Zg1pCaZuECzh3jB2KDhBUWTVngF3/ZGU+526YlQ1BEsSgHf7ENn0qiIh0Y7suS5er0NfIf/
ggtz6fjXI+X2MMEXAH7J0d/zvCRFUP7uRwOUtJen4Ymbm9/IzTxNidQEOry0SjTgG0TyWrHAO5/q
zamxFGd02qGfqQ1Qpwi2OiIXtV0DMVSDZJBfNYi9a970rJe9f2xlKWeb+lRTbltl8RTKnQi/krtl
jFgYplWJoZR4L/VI6kNcRpy4nXY7ER+oh4z/kLx2YumKbLF8YOmQIfK0kFfv5EEXDiYROKcH8d2K
kHdl6/GoOxo0bo8st5t4Z1PsFPqIiYpSENG5GBRotW8bSyBmhYp6gk+hI+ubdVidemOkw8PXLpK+
O+eip+T8noJNvzzCytu7Mn4sPVx+O5GvoHzeisSpC9j8uETfFD9ieu8Vr5rFZNjkcIU73tjnhEwc
dX3YtlNg7GbSDf5lGiPfpbvqKuGFWWw1X4QGhJ9RxmrL+X4uPiwVajXj4fu/044tob1HL8a9xK96
5uFzMBAGf9WEubzwAyHVqTvX9ZEUjC4KmW4WIXdod9+IlNBk5h5y7jS3xXAFCRClrSC2n2qXI2zn
vknaMIG0waNUxM2rKGsR12/UN0lgaqsq41n+WsN6LIH+E5Yx1MRz1+32fZOjaDVr0+C8dMDD49pN
e6bgJCMpQCq247c5naOGMSuL7YbDTVopMjx9VI9p2Xz6CS+9wApLpcwh4GR9C0KbKQ6NZitBqL9e
XQ0/LVZG2c8ITJ31aYhPZ05GJ9ld6TZp/GEn6GVMmyNRqyESt/gnet9Ag/Rsk65Z8IxKEiZ7LuNL
TR3FSEG8Cfz+9HDr7CrVilke4VOw3ljaIrElgQunRXWZbAv1S9FA/sW8aU+HWeXQ1UpNMxY3aQ95
9z22G+/VAcLdvbYeFnRZVpStVNrAs9kuFpvoSW7yfNjkSMD0aH+RdA1ipTShQO72iSpZsn6oYIKS
rDaP+L7lZXCd8MG1YquZTX/w65gGtl6y/RCYmtiULBfIzktz3/agDL8pLVh51cMckSFQzlVtYraS
SQUDCw83pfzhEEwBXz55BJ24iZUGTOBcmTY6enLcvPbkk4MstewqFGaiud2wflBRtTFU0I4of4TU
bTzuIJKQf1AupnHBku5Ssoli2hvRypiwfR3QpBseCfxMD2N3CAJH5zuGvIHS/cDfa9vt7NExjx26
A2PQbycF6TZV2jCr13ynNi4lgsueQdhFbmdLQICNw0a+iVioHszkCI9An2CqJGQA68eud5n4Ot3Y
4UjCo8R8mSxIkjMra32yuyC2xFNCSIwxB89xuDwaxo/pISVWURWxVRWDkoTlJg4MXgfcwO0XtwRZ
u1dU71ISBF3NG7QcZ8emJzYTWDapZIv5ODyhNF9gmrMVekTmV9jZXSIWFPjAahKt6L9nafHifiMg
5XOOcNciXD/FShjNslnfDdJzYk1n1GuKpvxI0daHLJaS5n4R07L+iK635h8bu2IJtdmKqIkSa3Jd
GlR8fHsNuoV5L05l8FEsQeyW/VC7J8AYhmpuEWE2V0B56ry6q/8eIhcbpwISQgA0uE8jvFkb34kM
qk7oYWQtFBn8RPmUST8bMIMCNYeMw+VQpnsKs7ZZGPF7AV024i/VVJWG75U4+bSwg4HMMUp1WoMj
KYZfdMzO8TrnohbG2k7T9BfQ4yO5E7D8036dOZE+qBOvn+psSkurrPeMc0ORhPVXA1e6+NdYg66j
F02W709lA4PglRR4gcy15Ce6NjrWr0ChdOQK/iecLAtVYxyRLhiOfrWk89+ZeFCiX9xR2+ga8dz9
k5kIFZ2Aweic5HSpcLVnsYSwyefLJYYZ+IErrTvpbW0hHvZrxDhgnKX4wFT0pwZUzvRXKh7+gI88
64COS0hwrf4e/ppIbj+ihWQc+nIen8W472fSoAZ6/ikVM4+wDhzknA+Hmbag5ZtLIIm2uFkUYP00
abmIgSgUrH8DsQq4XCv0dByzYi86V6o+I6WZInO+UsA3p6Ck78ApsSv+0tNSu8/3/2wMdESf652t
NEKW12PhwY2IenKLskyfD5qb0vGizOZdtWBGUEsjrcfkwRqX4h2P+LCgiQhcYeEPLaQPJMGrdG8d
Y0I7ByujdXZ34E57dwKP0aIeioMpyAbNvH4EFMKlcwUBRQ19UHFvMkw77BrO9gMs4HuKopF9d37Z
/qPahJmvIP71jLBZM/hJfhGJqQphSC0zeDTJ9Ua1rQ3NG0UZPN/yk2q2Lx8zaIJ6a8NtKuyxdoZn
xk6SfDJ1UZ+Iv8zx1+NdcfR3lEAnR+ozHvhfibVgv5xRjg9mqpMaT7wNApR3oWh3CTt8typzOz7g
4fGliQRrW3bPfQDud8b9z0bWZw3f0AqmnEOoDbD1ilF1vpvgq2Go583ZdNkAuG5dSb79XtT2f5Oe
Srd7Ha/HpoDntQL55HrsBhXpjJerKXiyk2f2W5s8EfVK1stCbRGsLzMPjpxN/eo+GyJyCiZ+wYem
i+an3AE7PsLswqT23kteO+3cUDWaNbALlUuKOHkgIR6DDNBdeTSK3hT6vivkY3Mpm2s5cZ1QROfx
LpAwakCMt7oDEjNcUZKSRpp+U44AtT+R4Ld8DF9UfHGNyJ2AmGUbiksAIsQniHXnabRcBLnyf0B5
TfFTPeD9ASpN8bUa8OaTRPNaPRMQ2ozGDSA+eifmUIo+BLuD8P4eN9i7ReHg+9TUx+dxus6C76ij
3HP/9DtrGlQQsdXiwo7CYy2bYF+S45lcu8jhSDQapd6/iZpFXtrNGFA+sk1Df6BRZ2HiBqi6RPKi
kFGEsSlAczcJCms9ohyS74dwOGXc0FFe4IYR50e0dT0TaWHmTvyWJ/hcuaf6ux5qoE/0HFd2J31M
RFAcR75se9xl+h/xPn7qiN/WjnzqeYxNlOVoTTiBYyL14MAHvSgSE46aFlimEfRJdDN0vdpwRhMS
ELs1WxlthBWtnaTeeEZvX9Hkn0mH9/zK4+G8Kjc3wUYqi7O9o9Re6zGoNbhE8qQxfoQUiHjTJ7Iy
dnLHn+u0vggSDRCicSJVS3Ln9L+uJxtwhTMHfwugjcwc/fr4X8o+/c/ui/F9pUPgM81WJ0oUaSVQ
Tc43SGPL7NmDbBLZQ/uGUs7uLYLUqwycFRS868o8jQhT13ilbCRqADLXkqdO7/f0hXSJMeVqGxHV
2H5+6C70Gl0kiyQxcCvAnA7yc27ubsoicuCfO26Fc+y85NzVa+5I1jMVmti374+IiHWmKMWSNFgS
xV1AQRoraB/bIO1f8307tk7/+giuI8EVl5Zbf4MTo4a8KAndRLv7MEjEAw+me9LgJOH+GhgxiAZD
3ZvldJvIoEyIwW2n0DPao2swerwdX7Kn8pBKsCg6dGdcfa09BKuV1o60D6ssJp+l9sEDq2PTvaT8
+Q8P894YVogFA/QuHIRNoQJm/rpA4XkidGrGyq/VlKb+9w5IAo3ducEXgucXkuJ+7nyfOJGG3Rdl
DFiELVuKOVqWX1FDX4VDx75ejl89IXqaKhJwc5mJq9hX4bDu/yGxauDWpbytO76QQhRT45mC+AQj
C/zz1YpFQyuzyjWjLLHxjY8mqjyVxrh97cmr43Ar/cX82brjxQl0qUlWFv0n3q9ulU7O+Swh2wON
6VkxLwblGYYs+UK7+M05uWQw+nQC5iDU8sy+Es6ue4LTUXJoXzyl0hxDW4OepCvYa+ML3RtKOu0i
1/j/oME9OjWRmLpzVn6HDUimasqhYeBLUF05lZLUCkVSVL7TrZW41F7bJpT0OEg56ZImVF3BgQLp
1EwFG8zY1+VD3D7GfNrBA+KUTPC8eK185su+UMEDDuEudFsYj7oMA0RccTaj90ldfI8olbgO9K8f
xXIimnY2jIa+jBbX8ZaKXdPKf81LxI3CsG2f7IuI5aCYJXi4gZ5Du4Ealt+uYpNOTJHmre241GcE
z9pV0UQTSs/kgOHOA8Nq7odZMsrhbVzHCH14uaSxRZFrW9Jzibh2Bzboq3SmGwp1/IbjHBvVZxE7
1cvH6clsaJo+PfR/NO3+C6IfkSCsa4T3Ar1bkOTyhUgcblKG+9N7dAEljnnCu21ScTt1vxNgSr37
x+OmataWJZl6PoNwNeDsGIdJNbXtdtnsbyUv38pv4T0pf94fTSZvomaXfl8X7kqQnKpS0PzhzaIC
tGQkegTvQNPtSXeQ+pgCejoWt7bZx+Elc+OFs6lRSrVQc1qKeLJftX0bypaR8Sh9g1pwZ0waCvOI
mzFzzR7tZq15lCrqxrXzNbwez0RJJm1wYaDea50dPSJU1L7wUTc9FZ3EUNi/uPW1J/TQBYLivYog
K6AqZD5XJKohxPbwL8sAD06XtWn17oOrGeWgTP/pV//V3SElW7tkPBcKCge/ku/lxsnZBnUOBkCC
iJBBcQWSdPfG+Yfi1yxNXMR81RtdELEUbl2en44ucSXH9EtQ80cAFpcIFAfbxOaTVNDPJhU5p3eS
M8E/8H2Rhv2/deTua98DhVu5iuu+kxiWLRvS9ywAscQXV3QsrKWwiYxUkhwAIDFLeXnlUgs2ybjX
4I7JYA+LSIktb4N3FooU/f1OVZ7zvkIHIRzVnYh55yRS48IVvRJCKATrxCSQp81J2q0Q3fPD+cZH
Q7+tqh9Th59xNLb56bsNhrWxd9mEeSim3xIsfk3WHljUtV9tormr+WbBhd614/FIlTPnXXAipCIi
uCBTtMYtM1h+fMaZcUcbFn29b2p0eWZbx7mTV48CtOF0CSbMidyDHTMVWUJd0e8GOq5iTCcWhJAn
gn7c16wfsAPez5YMSPl12Fq95C4lgBCh2BMLoDIm7tNhzIIJy0vcvjBO/8N1O6Wjr8m0SaBnn7Cg
v+P42y2VVQXRchTIF8w3g8+3gUal/6ooPyI50QrOiHlVdtM1N6hD4r2svI3cXWbwh69Gu9/wmB44
9NZ38e97C/s6IpAcLMqvsU55SCXD5v5wi3MS+ZMqFt8eyC0xvXKNfO9pLzkk0VpUpqRf/Zev9pfA
gHFdFDrVwlYHiDKzB2ONf62Z8grwAZ+8hB6di6IuwYXOGsMOuNtaRc26Z4uMdY7O0w28FkgK+M64
TGRKth5m8NsUHGx/zGglzttcunITmdm+CWkzq7M9NsCvxgUFyeb00kRNiGPq0QncBt49u49wgbmp
3YZCfuypT+uvPUYUhPd/ayYHVWh16XpjVm/c8MOpWtmDNYTGi91UGw/S5NhrqVEJqH5XTkbK+s4L
aUu4nQG58QHTHGaEetSjqrJfBtcU5YQA2cr6iS9nDf+F/c2Qkyfrm4A/GKbnsZrU28O5Jl57Du6F
RwLxYzvNobZS6FAWeMRUpF/JRBYVGtYFYHzQtdykXHkdx5L6+thD8iV0mjgC1H39T6TIq99yUSsz
1qyUgwThv4rCBvC59oOtGI2MSegtaohrQ+1eRYp9VU71gjV4I+Fu6mqCkancrYSr3uqb/5NtD0d1
2dpXRa5r6AUSVaPDB1Y0bqoXUSXxONm6ttXvA9N/B2jhmc12aK48MkbgeDxIIAVvfLhsWWCoJXrj
MIPtM2XvxLnVGkU+BXs1WAzLcjPeVh5jTjiqNPgeJPOmEF1W2HCZcppaanrngnU5vGeCOjF834zZ
ky2qhvYqdFvvktUGwap2cAuWnvzbrV3yO2sO5cUTOeS2VUqC9+B8k+9Fo8zuVCzzGL0ZXBUZNP/m
RjUaokahZEFXf9MRgmSfN5ILp+KUSmnfq+u3chUaTQLvZrobP4SwwclQ0/Vvz4evuIlAuVW9B+fe
sagssz+WrVRTNW896gIz+9rMuuBKqeVTRyRyU2SA8pDitMtwgo6nAWeiV1Dsgz+qAjssoArUlGmc
GbB0PcRhrtiM1wzwOmwg4usMRKh9vYXmOe8JWg6cMvJ+Ntyth5y4uUDyC+vfWhWO3HeP414R75EX
frcHK6WwyUVZMBe7dbM4J7geTvKPTTI1iY5d1ulGGjrGGG0RN4xeI/NuVKYvJpG42l0+qT0ikUyo
0tzBtwjAuGCv7mXKdnzWatgyF6E1ElabNE1HF/JMSARboamMLQtb/7TNJ2PC1GQ73h9Fk2FSo22k
dbITX2pGxmtn0T8zTSNZTEtj+HzthpFwLgJ6XCVKryqdVgkluenCyLZGVd/oTWVKZS5IpbakPy/p
7yKPEF4G8gL0xVYAIx/IfzQXVEThDViWNMqYvCReA6ea3uhRXpirZ2+wR09Gctyr0EjVIDUzeLdG
5r1bPFkzP8c6a8YkihD6WvzO5CjVyXQDlX9UnelYSEB1VfjfdQlizupfUZQzeO0ThdCX42vgqIcL
nqoZdlctTKVNiZjrMRePHk1APoD3CSDPXmGnsx02s2x4XoG10fn9SIx+JzxAiyDGddtY3/07GpXh
I1mIoZHpXv1rDpcsCdCge+gTopuqkUlbPaDTDT7z2j0PN2ZCUDmY0HlP+tNUTMD3kAoGIi/wByva
MKgzqgl9J7R/WTkW9FXu9X3ZB/X57IRXOrIRAeyUp+aTA9jwc9hUejhzrbYknR6fXGeVXoygQahk
hKdBU2sfcJCV7nhwn1vUTHtzKsftE6kU0HPn/HH4YN2LQ/ytmjI44BncoMlWGB0/HRhOoef/RHtx
5vHDMfQwXg3ns4HkscGIr5qR1qmkdJhWkMf/faR61x8mO3NbvWAs8RFBQhg1AV2cR5b19e1PI+hu
7vdLYN7vveNu7IxZhhFABVKLQu2XddgvTYmllb5EyVFumtU0zobFgIz9jKnKhe1AMcJXWnzlODr7
lOj2kOwjmdUXvFcqbuQcywex+UDEOVGsvz9+/C8RaFQCNVFa8roiSXoz5CL9U8l+u5HnqIA+B6P1
AGNzJk1y74cdIP7u34XqUUg73KoTZ7p9i6on4hHITZ4xyToKLuw+TuTNOyZ8xATSMO5aov/mijox
CkKFvJg3pCe4avjjkaFpGv261BvVJ75alpWg/DJSpR/5yewoxOldUiDCPnLhTkMSyh7PXng9cB3z
aj7udWmafnU+dz4ZfbkoupPHc31KgZ5siK1UKElbFE1qkWD76CpcF2dH2RBeid4w3/9MbfObRrzV
wML9uzJz8id4LjbL6F5yxrcjC5NaCgJ9/iolBgUUvNFnKQp27HUo99VGpAkCAFKJCF2VLyX1NrXL
lOEqi1+czwdUOpKV0KGQFBRewp+3cNZTtkm5f5TZU2SUQn0eSwWnED/5LNi1t2NG2yoENF/De0Vx
OpxvNvj1w99KN2OssagyTpDxmtlDK6WsXJMpMrgGBQRGtOCE3pt8wA+7dDl3EQtC7xxqTICMu2k1
uczTnG9baUSmBh7hMI/f34WxMDQ9KlyqEnayK+rawegBOeoxu7G16ObPEfEyDWCfeM4MvU8HvC2G
ngPmvA/DOb+tq/pbdztHdwZQPXEe7eDEqUpnIBSLRGFvEp/n+IMIHLJG0/ibUWKzM1WG7zYhzes1
qbzIAxilOOfnVgIQIucGvxwIro27kavN8XRxpiNV/eVEbIcOS1xcq+WT9fY3fy/yPUcwM+A785nK
7bRpGGFlL1XPTq/fGw0Fgfj6e62QhFUtxVCtbaGfGgN8h1fXeIXdUhBP8RJxqln92Bhnl32Je9+A
GGCx2ZQJaFXzLQQG7D2t3bqNz63B3roMm85sf1XxihXf5SzasKXuaYbeljEu9HORfsPiav2Gpq0O
BHlZo7bE/chEmeDE4thlNqHTQ0PwhhrGFfAyqzTUEMs3ZWH/aTZzd8pdW13fZ3JckUE5861HMwOy
FutL7nFXUCG0RkBVPU93bvrb/RnnKmtazQ/aD1xcimu8SfS6soDPy1Z8NsMFFSO2/7RKUzKHCYFd
+V9qaR0N8jEyWzGupo/eKPWOt8ZH+G4n/AfXpyBH4XBprc3LvHFgz3N1Ah/kOKliu+otct87500n
ix/EUyaI8tP5Gj3CVzopCSMg3K8ST2Giv+GU+SI8cGKGbO+IvANoqCGyVMBcOFm2F0WfBqcAdsJq
rHOKXJ1kSpatVut3PLle2Ga7oESLHh35l8s6JE74SHLxZcTS7+UoN6kBelpPTNJhvHytVajT4zrY
w0+t3+N8zjafjFPhl8+6z26wEKkK06luYy5TAD/BZseqyu2BKEFGC0IsV8uJOJ/7jST9WWP7IN9O
m8ZcxerJ9fTmBFhyiY7RYhA1DWpscUr2g/HpZ7UX6e1IVqiO3xBpKq6nhtrwr+WVk/r4713c878K
ZU8zmRZTMXWFlycgFpLjZ9w4E61BHGzwmQldXivDGmwKLQJo7cX1OY9frgrNp8fx8yLyZXTP+orU
B47Q01EYri0g89E8m1/0ElepoVvDMEWYPZSdTT4j1VKlKQmgCFqCcDgSHO8KOSBUjPTmGTAhSlKM
ze7HYeWn6Yt36M6QC2HJQGkz1nMMhjAeVM9gZcPQsQLmwkHKD2y50drZyu9y4akBE9CMRRc6uaox
QoMIjc3ew99e4xQ3Z2Vw4ltEPiKv1e50LphuYrSpgES+GWj2wCZCCY8u6nLBVYI9N+Xvv65sgrXn
VNkqbvqm7tao/ssAvE1egZroyhu75j6bTOiW1WaFefVtF7oeNUBPtnKea2FFRC97Wxd9oPmZXJ5j
Kcn8JBgBIW8G+IFWtMcYvhdg4rnPFM3Myln3tCQ0vfQnZk/0JiuxrMFxxoTGZ29Ecmzaa4iI8h/0
+xhGkHcdJtMGRTVb/EE5LAIDoX29dTkjWcC4YKCCgo/530I0uGEm09xdN8WiLir3uQ2zJjYgQ3pS
H65wHAFMXM6xlgpkjvJwuiVrah73dIurTbnVjqnQcMloqKEJ5X3/5v1/vVkhD4jhgjcDplkVnUbX
7zPU4zGgzB3zxuONzKXzONuZvVF3Fjt8F0HxzHk1OG1+i0K2oRvoVq31L1IhCmxvbzbMjd1+G+DB
Yr8LEaRP68SVaxIm/oi59HOo/1KxDnDgmjnCQ3rsmtz4HCrRCsRUrfdyPky8kkgtjueNwTv+Bu7E
0f891/m/yf4nP17Y/ftrxGcXz6umpcbyvbjUH7dPHyd2dq1aE7hG7qsFMuMafTg+mYwg956t786R
NwwP5CyZpOV5Y7JxIIzJZXaSwrkyPia+uXukIiZI/BEqqqh/hkdHfqLhV2WgSvZd1Qybo9X/xBp9
/19cZuzp2S2CLl6GmIB5s3aq8oR2b6xOmx2yxaDXpNFsSl/5ZWbOLMIh46SniKbDT/dvl3G2IVW+
kk+rxw/uyeBN95smRuIEyYPGi7vHIi4YUPFgxL1CpVIydtWV6JQWk26lIHVcZI8qnafaXRuzqGPb
C0rH81u2KVKb3k/zuNPXua9E+Pq41JrX35farfSugKOrhVigQ70FX11Y5UTUlgrnQadOxjtYbJGc
D9kHpAakRiiUM+mNImGOgAjyXQIrpOb8YLD27ks7xNxUBtVbwv760HKoekR3ahoHx4kKtfK3Irtk
gA+1IciP0bGiPAtlWtH0hmAvR1g7tQrxHK1t9JOnL11TR6hiiTomeLEtQQPTiufqyo7aOwE0gd2Y
PeQEixNT0LVkYjjqo4j011pmMG/RHOdXVWQG0lQFRR2YodkHavyYxiA+1gR8w88ZedtPkS4P1iKy
d09lvNDPQYTolGQlkpyc7LL+SotduI7PaFxlXp+0KH7GeNYCtVEQaQlhtmTOsurxROgwx7d6r/kn
qmvtA+Kn0ANorpcdOWYq4YG6WNEHUtm2P3RFHbQxEEhADiYQiDrpcGavEXGTGv/jUOq7rlzncwQE
FvMRxusHNYp89sDivFKgogzAXo2xj8VjVrQkTuAMpByIhHeNVFhmtbm16zZAf7gYh0qOxiQiKMML
sHc8+9SkPk8H6GvCZABGhOYqv/+4FigzlrXaGCosUs9k+Y6dgp/O/BMdcNA8liNQddJgY5QKNzNV
ghtcByfJK8G4FB9JJVPyT4NI3DVNqfEogxuUKaDYffxr5si+UjKyedYizo5UF3HQMAKyJunox2Fi
rT7ckO5YrUV2/kW/wTEr6mlBMa9+1wr2Kodk/+W570IrqZMV2Xhymj4huW+5F5IKyjYfQDLlCzIx
1EN0AGdhS7pR5bakRpIbYy4HNAvpxh3oX3MlrBbvhHUExLv4QFvfF9WJc19F8NqIqAmBxwY2QWfC
Sun2Y0kEvX8Z/nliVPB+LxGaL0l+CDLyUgAXThlM7jZBcsfT3VKLcGO5uV4AmzvcZxvENKyV46Gx
YeOkg3maXgAvCeeSY8PNWbprsxq25i56VdDQE6qSBzhRSHMODg5OPMGZJp3M7JxwVAc3woP9ubH8
wpfcNvN+K8JD7cyri7LNGaKlJcTQISxpEFbxW2Gch8LXS5O8FgW4Q19lipjWmnQh66Wn8hr6ng+p
ZZJri1xPvEu++m54rqFCGXqkImiWEPTfHro8en7RJhe4tVuSwgdqma9rEP0QXNw2sKo5mg7uSGTl
VJoW/qcozvKxz3yZLChZ8q2lDzlCvdxPDKdnPFeg/gwslKq+Q8AwYPcsfw6TEKpHE8ubVyQ7ed5U
Ni/nE8uJ5+0y7yBp6MUn4Jm69XcerNziHIiRAGVk17QJ5ORnayJl3I6w31bImko8fGi4OilcRAxW
3Lz7z+dULFr9PL3T8QNyfFRAqYv6RCHGPMlyQaLyLQdFq+Utq0y3sje+75Hx8PvHOSLFtyXdIUqz
oiYFZ6hwj/rcsRMlhVXXGj1EmjY4pUnIZUzolYtoWDXPGWPjbtqlpJM3mPZPPxJnh7siZKIRmjbB
Ia5RuGZ0pTBUBYcbZBam4vdXdLCMOFNK1QuER45F2E3ic7wjpqkS7417/vuQaZg6Az4TNNgv6goO
k37TuwMPlOWKLx6LJBU0IFOlmU06Qlzi1Xu11sDXDAV4piREni/dTU/I2s+Yvv50ADdDtWayyUDs
BvkJCHEikliNOdcHpmozJz4jJ+VkWM7Kq/Xni7BbFQJyhn1QnuhsnVNfRhQWAnErBTnqdZBRYBKn
Yu6f0v5n3MiVZ9Bbjz34f/lpeD7XlLW8nsChVJMyZD89KJ7V/As8tFcv/0EtB1bLMMTWdshNVX0u
OmiK1nGvHBP7Aao0fJbc1zrbxrsFfHVybHYjQAh6Gh6q9MCkX3RxgX2HrZNM+Ou945rLUlGRVYON
eZhKSiKQ+1FpQSj8sDVINrU2Ne6gZkgRmvqJ8uQpTipgMgz8c/kNB6ov57/tJEepe0lzePCofSi4
YR7QGjNhyW7dKOe+CfX6yDH+yxRk1nd4AkFyfZmVpXBlKvrPX52e9TQ0dVLmM9dKzwJoR3/MuVtf
rvjGkTLkA+8nwwoXAOGJobAiel8EqaqEKubvBswW82E/eonfblOlLc6ThP516opvHgE4CCtaRCwk
5mHckVATwSntcP6d8CQ+RVfQTdyJSVP9/4V3dZk1KCijuScUfMBtB1OdWQicNBFhld+BtAAD9BEf
i+t2Qwv8Zx53ltNAC7UNiLJnl8x4sKEQsUcYuJdR1Of+4b9y60V9YqeKI6wkU3DiO7LwMvbWhGdx
gAH01CVJMDtbf/JfTF/XE2fbCLcjrrHpwEGxWegm+XHrNp5dcr55itd7msh5bxyQ499BwBiDobl7
D1bBuaq7Hxp/wL54jCt4PxJ4X+8YQ0EGd9SqL9DPMWY76cBRybNnc0PfU4j5rfX0XxQs2HbgJ4LJ
pkpi7+8xgV1sP3cGos2vEzlv+NNDfneYEbYkq/Ibc2SNfhUFKyZrlFIZKuShErLbpvw81MrXVNiA
+yROOZgwcpAOoxHFVlHYYerh+dxV6s7EegWJSBBfUXQcxZZugiJ/dNGii7b92jVNDlVQNpmvuOzq
QHOHRVCbXyEUUJvHa4owuncFwjGNAGvj8obcypWuD9dr9aR1ROmH6Jx9Z9OKcJaIPleZQYqvHF/s
I6WMzlWOS3CXciVOdDvcJrZZqysN97tWb/QgIrfy098XfrqzBpRHAKVJT4yjF7mLRQDgxdVQldl2
cHupydI5MjuVcCH5V2zVMOKnuEQVz3Wr353joa84crMKDPwaTnmf+oWwR5Axh7lX4eR5uUs3kgND
+gYLUg0BOq+ijh/tyvZUamOUmbEc86/M6BwV9HV5wQaBJmJuVdtjOzrXvEMpm/8jFwIY3nqOfXV/
ZGhoQy1CHd+QCS6WM7zMS5/a56ueAMHiH/QJKDG+V3OvMa2tPS0SEndMgvvIyuu1j8SDlfw6u5Gj
61vtkB0svScH3RtROyIsuBCQtxLorXRU9zD7nxJixtntEFeiM3IIdUd0FS8pobB15tApDqDU7UEN
vB/I+Xd6ITAQQ+SoqY2H4Kt4aU+cJIlwrvtxNMmCYIU7Ex7fFKNESoEon/8JXywpfv6MQPdQ1l7R
/9m3aRPHWS+c5CwPFETKE3kh/W4zCbrIRcgOlf7PT3vqFNJRNXVEJrmOXjsGS1ZCOij4roKEwkXJ
iwmnBQZ/B6IH3plOD4r3CJyNYDb4NX4TsAePVv3JvqgQcokgq688TV7pcuhHhkHacs6i9hNV3xLp
QRzvC5eMThgylAIuTJAn/EgGf7N5/AjkVsVpp86ATKm9jzmK/wJ//s3LcPAg47TlPl/VIrP5JPDa
tL8hgoUi1MabPGk4AVteld510iImLJ0M2MYbGuJhfFk8A2frb3oc3XbdqmQyiZ3x/0/0VOTWuf1d
JisAnSA2zpkOf0g0AcyI2f0WWBOZ+J6bplBsfZTu3WtAPTvWQGiqtjdai/OLmE5jwpWHLqxa0V3f
kBwwLzQE41peoL0Q+6GHNhktIZHuyqnQNINBMyrbza/h5w64eX/Z5gFOycTpr9Gd9J1t9fQq4gvU
u1cEx8JjuLlVl+3s46zW5h0myyZ3GPdEcm63a1EDQUHJNA7QJctQ/3bc+b/iaePnnNH4in47bcbc
Q3IXaGtCCskCwT9FZNZbKu02Z3L6vYnv6zQrUVJWgv3Lp/ZlF3fp+cDXZw1kz4BdZz84hyNmxosI
2Jh46MnOW65F9iCpUs9uXm/0g6SLC5kISh+PRBX/6Tz3BlIaOIYH3kOGeXPRAqbyCE33ZS9v+hnZ
62XmZYRleBzb2rhdjIlmi73/nQH0MaJytavCpff5EnqFl6+WjR1U28wIcnBnlY6ArFOczweAty9q
qL9L99Vm2tYo+Q5YecrDgzVgZHkxOhl+qpp9dRvSTisPlf6UAtNMwKDhfeXZNhz56Lgea4vK6ivK
HhXS+r5v/u+PNAbmnDoCyK72q18oeXjNP+Zq9XKkK2dLcaKE0Ivb0r/y7pN1g42WWMkMRPdjd5g6
iZH+S0f7p5WQqQ8EVRoeaNtyZoEQFPJxtu4XIq3VNERz2isBdTJ2q+tgrHBHFV5pSJ9V65UafvyA
fwyQ61cg7rU9z+i8iHOXgXCfkwIfcJQcRwqlDHoVQUOLeAOETBUlQySm08Vc54zrl4KAmguz4lwY
PN5w+1kQeh14xOo5/x6dI0Hgq5LAPBV8r4GeuZp3JPMs0230ctp7SJU9gndpX//AogwVi46wa+Zm
cltazsFWJlYSz44mGevb6f1IXn4+oHee0Aw89mdM1g2wDccfo7x9YqX8yhOz6e+9n7WnSP6+FR36
u1y++89FdaayCElPwS4EhVHDDlZX6TldqgWVHb+mW0TIOJGg9iYZqgr2T5AyKwG2JVjfeG+CtjIu
KKAzrb07wSTgtWHEGF0ptPcy1psWth/z99BTvYUkOh3GhH9y/w8rWDUQikmfOvIihgLoe01zFEBP
OEH12DrcFwgpuZJjerVCBz3vhn4eaa5GnTd85RAxNxQlr3h4SjCjGCG0+svwx0EqV2ZYo3xF0MjF
c1wv5t4LJcQuGb5LGNG+5noUBG9Aa0L1Zm7Lrrs393d81pUoE85sBQoQz8Srw7K0jb3ynjwjONVX
3IRP9ohfA0K6cnZh/h5FFKz0saUCb7LYgzc1mcg+mHZe0AW/I2RnB/6LE+LUw3doFaecQvFb3dw/
D4ifdodzYlUxfrgyG2J0P6lUInMGRdHke3+DPao8CSYc1qmq+71fexjCKMdpNCkXucupwfM6es3b
uTUKOOKR/j/PJ+M+kDzbIgdDi0WlkIEHoM5WVVYO2poZSdRjYCOLO00sCWRUHBTj0/LibXDDIwCK
N3gAhstgDjFxsxXngJ6p9RsZCh7HAYWr9+u/HF3HmrnGwkaZXvdD9tyKqWa9yUebdIQ4XqdWXOVx
jNcY2Tt1EzTF0KcWMGDSNQOTbc6a1R/Jf3qv9h2oBeyv0dCHI0IrU+/NuIgh+E3ndIPBAOx3Ry1i
qvwrDv93Bj5T7ns8bRfraHHuytQ4qchwD9Y9FpoImjUHndlPhkl2XHx/idVbP1alzalNKzWm7FO2
Ig7oYywUgaHBRM8vPWGXiZF8PAcTsbiBMwCqa7q5JExSoV9fTDhMz6CoGUyaPQn+xqiA8tkxAp9o
mXTF+nhyRthD1KD0gQM4PVgXfsja9BvO7YEpNCXlJ9PM4Nl64UAtLpVRXuTerneJ9UT7t1wsNTJV
n4Clt2DdenFvXHeRjpj0Z0ugHLV39uxajZWO2tpgKp8HpdJnxBgVB48PA1tL02lkXE1KNxn96IFD
hbjXqjcOTylULEQVySYc1dCH2hYGYyqHX4aDijTFnqz6/71CTzt4jW0mYIebsn4XjnWIw9uZbuoN
VFvwy3tzwm68AXv4p5vUjASTxrrRIuN06o4tXKb4KI+8JVWrpiDgedBXZaUg9F2gbTJTqq7G59eg
dCgzEoXu1qHbHPKrN/jRsB929AfPlr6nUvK+5EnxvQOn+3rRCtrSTDqtVgA4Dj8W6k8aeVWaD+T/
+B+N7oS0v+9VuSjmgvGcWfRoQV0A0wYeeKVpERsCq/G7qFbdyhNHRxWB/hHjr0JPEgYSJXQJ+od8
+CcwfFLR+019YkDAbiqAI3yGb4f2oRDfaivrOBcdl1H72NG7tqwpiRWUOlIJI4HvGjzM7xWf6pa3
azHTGeSX0s2XlQEtAOIptNlUKfqy6/LHJvsWreaMhjNcww9bCMEby1GU5l6yI1FhOogaLDAYg0Mj
03Rev95SUNLrB19kFkn8CQxr4a7nDXiCrjl9jkIef1+Bt4+aMxg4frLIk4Bzy0WzWEoItF/sHoDt
kqv0nqeQEjvRZcIDs7B1o1OcecebYRNCDBcbF0vktEXIQi7gXyL8BKTJ22DKKT5Tl5Hot0Xa+gcg
4NUKEFpyKwkfAGH5vr1RRyGLSUPoIThbtB5zkDJNP2DXKE8mrKUe7TfsKCYAfb4mda60G9aaqR6D
mK2zCUTPnizqCPU5WM69VoLjyqpXA5KSWYjpY8Oj+lCNQmPH1EOOb0ehQMbyOSXN/VVx/nP5XgpE
/y1vqoF/lc63Zf6+ZUx6bjnHKKtiK5+nkvzTVdvQG90Dxgo5wJ2HExtIJ4befxCxLHlGS1qLaeR7
fpTZzx4IoviFpuq5u2lAmIdzV2iuhodp0Zs10KAERMpI+tC9HfZpxu3RKJVElzBvxfhR8jdYKTY3
psScL9Fx6QifXErzISHgJGDFJ8n3UrKDJAydIYFjiXrq/ZPqZegz9a37UkPFFVOchvTowRYFrWaI
iuEKZqByCnSihHOEz0RNsz1BRVm+caarnt6lJkiAX9wR59YGzXlljsv6DNbBQ0L2nQufAFIVuzPA
mZuPJEmEIAqc1ig6ikKFZbNpj9mB/cyGoVLjk4c6HlqzlXlCVE16k+ec5KqRc+gUBfdHHfRD7aIt
lQLA1bsWp0ncu06ouBzGgEKzBlI55aQ3915X85u+qONx9KwJ8p3YG7JlzJMYE2g9K1niuc8mZiQ+
hHZS8H1DKkCHaBJEIBM9mNGU2oaCozLPPHPVnVf3WXI2q54swux2WrQQztNXOFJWq92XLSEIdquW
PAOpavZb0R8K5U4zXA+qxsJ8PE9AQzEKEip0kxyNwQq1Ny/GOJx9GWvhp+ijW+4s9q0QYyymYUlr
Bypbb63jDGliYHOMI6udlnPQbszsvRTIG4H1cPwD/TXEvz3ph7PkavwalzIOyv8x+Vv5VG6DB3Xn
DH7WUfPYsWO9Q3tNAh9jTIEwdk6C/2B7c9Yu4BJFqm1K/gUhOzSEimsic6sh5X9usb6sPsAKh+yY
wHiv2tgq3/ciFmncOfetVvqMYVppoB4O/NWInbdRKrq2EAvb7b4EAkyNyysVI704Qmwl2oKlcVwv
PXzvmA0r5WNWbzOce1KtraG4Q+sOJy4488PTus6xXtr/Aye6rd0tQ/5IW+xdfl2FGjM0EYNMMM19
uPFJ3piVbhnC/8UwRwziD18GB4LVpLUIHeWQMHqLh8kq1NkkW6/dSYlHSIYvvxVwKHbnXTPjao2/
BYt0cpLigD3qAkoryYnzenePo3wcGpqnYSvUgsxI0EaSvRq2Ng90UZT+MRj05chslkPRFo1Qw6uQ
9hNoVNzCfK98PdrJUjvyeYDw+G30upa1QbMyg6AYgs5bQ+MRKSpXGKBTNKaSy7RqIQ+EVachEta2
aqZPcimPAfM5BNAqgp3hrFfrhtgDlRJVG8agks8PeI5Llb8fli4ptJzkB0PXuH+rjWTNEajngChC
O62xRPMRZJL8FTBDMZ1/z9rsKq7tlWCZk5iRo/xD07Y72pL9s81zJ+CctzXUjz+Y/Wq8Yr+rdESu
1+fHY28qcyOxK6YYwzBz75VohEq+MGomW8KcW357+nXfVtY9dmGMwxddrqKp+GEz3/yPALrjIvIm
N6Fl39pcXCOjhjYjiVfn+U6s5ECv5Wk/dL37T7DVQX5uRi86/SH2TkBVECPAr4D19J6unqmrapEK
NbYj/iJLWloUPPpfKFoHigAm5bRVy/0JId7QNZIJpVR9AFBq4iMpRpfWAeLeP2kEBER2WrHLUeCQ
f1ihZ7fM/9kc2JEr87RMkl3xVhPrGBH/csq1xEXkJE/UdkQRV3w592jpnjulNZpYELfyyMOpD2mi
dnvLGuQafRAsZSvQhaht3sRkDi207fafKIRHmzq0w+p+bKi3tUbvEJO81mVQnfaaNY61vViT4nre
l1+nZSrf3LrOFROBe/O/qPLFjFb37NObQsa0Uai5SobSEp+Guf6dJUuGPOyBVA6HyCuBGiBmdxBc
xXWEravF+r02jX/84JJvZS7smwyXUuedF3KBXlUTX3RPNsHB5dvrf3+5WBT+B7cMKTwF74P0xSSG
n8jd8fKoSO5frvWk7fJgGZjHnWmuyn29hvQYWnMtUGJtKteIOePvvpCzkmcxE1It6MNMZtzSlmSK
+klNP2XtnATn7Wj4hieqfWkh1gDWDNxFKdYalHAl3XQkOH1xxq9WKWmiemnb8G6qNSFavTKXnKKU
LLZc3NbfTfAVgtNjqsfAg26rp6WDZ6NWeRJa5IRIF1MG8wkjGN49Y7PN6FChFdnmwyfzzON6H8HG
RbpYDG3EF0vxKwAj4dNjBssrecHfMQVNJ9LYZPM1DMlzWxvRzEZAwsMwhw+rspAdK44vrRU3GuWR
5sekKkd+E2xqsy0Xh0w2278ANFsfKIdkdz4dQBUC0hp59BfBXfQitnjnTskZmp6GAmgzYiz7lFTi
+wkmLS/k/pxHJGw8cabWFH7Jz8mita/fujlufYpfnpcKPYm7GHioRwXs1g7l7Y9tvB8gkRi3aScN
ULyKYGqrLGlnNEnIM7u2PuQbITCfHHeB00R391Ki8dyVR//KEfktRYOayvq35al17m0pbIvm5xbj
cFg+MJPidojw6nmnsZ/ioCxcI5F4nXy/OxI7f8qSYTCa7AwYL8rmoFQV8M5wIidiF2uGF5LquQsO
JOfHmE2bJsmVsy7Up1bOSGImrOk1dI/hVcEpXphZeocObwZdVmv/hkc4hDAZ8bUOdrEB4u+y2nhq
kt8JqxIQ1I0Or4hIwaGpYUHTvKomaMBM57dO6K1ZZvsdUnsOUyZAZ/7p78OzsiRMD+mypIgZjWDd
XIoZvnsNH4ZtMEob1QV+4S7X0+QOV2QcoM8/lVe2I3Hz8VMqMj1vgNuXj8Qi57JLZNZ2REQDIrNc
NjZUMH4CuAI10fhaiIOQpSB6ypQ7EwHiyChTFy8YHGi8IOUN8/S9YJuJllnkK82UMGbywiu5VhcE
VnHRQqUmC2y4qPsSLVUDFsLGY5quVeIpAQjed8z4trDrDYg4ANGTMl9A0ikeJDTAbE3UwLbJAUyJ
aTJp4lb7KAqhzgcLc60m09lshte+pLIsGngUH4BKVgVasaQzAuhkMZ6I2r7Qmcqb3tVXNbIlEE/M
R5z4iCnJDAUR4GGBizz/idLD98+xapTsDtIUDyCuZMFnWo4lXJz5iCUECm0BVYrE0XjCx54Nu8Xs
pb67/HdU1XC8ajGph7/PiV+xZKrVmKZZ+LXllGau67lrFz5w+MFdDMR4+CKC6C9G1bwJLr9lklqF
rnYj7PsWg+s1aMlJlpHWEu2u3JOMbP+2ePT1m9ZKDe6sOlv/USaxLwEXD+gMBLx2c1qr8J5lO21v
XeJ0mOep9dc1FEEX/XjGme9t6bpP1W1ZNSg3+48VoD39SV4Dvj/UVM7xkjugyOVUGdHse/ch094z
x0N9Rb3paNtBSrQIz8oRvkwrlWJM2xkehuW9a9SUxYP+He5Mlo/AKoIACTkAu4Wjs0ucd/K0kme1
c5mU7Nc3Aus6xKE2xX0Sinb+UkW2PH68o7eePw0Q0+gHp86KVpuoXBbhxLBNXAKYuArRRXXoZOmL
9SsPsv+s40xl9TFsp9JdeuH4VLRNL6D+oZjVBW6EVq/VR9pB/skxlIY6nfVTkmRP5LjLdNNRKQve
ayF/k0aeMe9jFFCL/milOmBxfMaGb0WQ26iSlQLEGzWp7NH0e5gFgnqAxC8A/1/EfEDeq/R+i+9m
3loT1VQn+YVnOWyENy32kOo2WsDjaNr8z97t5lAQyQhhLhWT31ECdvg+ESeAeN5BB7SeALQHBXd0
ufrm42eC67YVAhe92t/MJC6HPxKpefw3EyJohsSqsftApamZb1bYsCq1Prl0C/74+qBh+tHGJM2Y
uMplLupf4C5YGzz3uE0GVdHPY3FJRFzjYVjTQq5e/nMoEqqamWqSfgY9f1H3J0xkQGBGnn/0FXLA
aAFf9f56NorN9M9wRVZ5CYomwMO5EG4UuXLI1/TPV+thZCp1GUFaevnww5cp5Hv7hbvwGHJBgOZg
w8z8ha0lhUzkmZJDBaJdLsmzt6FWbwuH8yvI+e1cRNJDXsW2aEfNk7JjJohStMuzblEDI7cRCgzm
oXkj8B+3Ey8dDzMKuvn0OvOG8sB/5eUGR3cD8HmXb2ipM7GBuwPUZqcsK+1yEZwgzxVzA8o2dw6f
1VMe9gpDBVV1E8F6fUVmahpLwj9mxoQ6qtRluWJw9xPm9c6ksbnZF4xq4AIDBfgdAM4X7bPFg0Gz
OtM5ADyMvZsNGs8VIBuD1J+DfiFx5wa8zBwwMxvngifEfCa7nQ2v7omBP0k/npZFDuoFeSSYC4Ze
DItWNLYYDlTTqe3E1UwFQlxupqikg+JoZ9yyEe0v7SQJVzNWZ2aQNkWj/wCJ+rNJj07zc5FXV8ob
P8zVdfMy4ysMJGLBH6ku6xSNpO//iJyIqtuLfAS9tKhmhMaL/20gzMoLWNzzl2NIbO6yoLQbkJ4w
RGYtkPVy9GPkZylTqHiOD+0g4tnCoACFnhNmic7u+VajKo53eviF2650ANbezb0rkV7dx78PYy2t
iLTgcDofBYyLa/m0ODRpEFYxd6d1aspgtojjeOvSvq2ICrEfGmg400uEAsEOJTjLm3Yiq0aaGxru
2NNhiwCe1J4fyQkUYblr+s7DOl3+QfCoxKKu38C2SOnCVLt8jyIxl2vk2SmiHElcKgn7KCEsXpZ2
QLfo3ddvS1wtxNoMxDSYRgfgvF2Y722up7M8b//abwlgHEU7Xjr9rjHu6ddf9I/0u04q5yzG8ONw
rm/jQgvmSzFXuR0laUdySovc4fDzl3H34BwJ6HeheneZ+LmA8dueMvvrgAzH0uGfa5Xp9P1CAJVV
45tSpNDtFqKNuU0JreH3L77l2+pLssucrU2QLOyzlAtzfq2D3Rmii9DSsz5VvZWX7EZBO+p4l7A3
8mGHRNfzFkqUO0wVsBY0nf7DRH1PhTZdsuNLT88NY7k0nprM6A/YEvUU58dDklaFfPJSmQGUY/qO
lIEJ0r14Ur+hK/yv2J2yWsDFwWVgP3OOW3Ys5SiWyfDRijSEcbpNoO2+DWWWlyh9fyXXMXSebLPC
pjeKiyomCcZA9yHrLEHHwnkOYsGGeW64FRtMfcESRHWysuLdpprOpnJe7zd10QNpCiM5phMFxlzZ
ekoT/Mwmm6oObRmg/zJxSTVvJ0ZlVXbrng+/c1uSx9lRNjr6iXz//AeYDuBNcjEbNqrZ6A45mRZo
ARXlN8JpToNUi05JHov0ogz1ex3PRDDz1VNsVHHsrYERTnA26ZQYwE+2bUM1RAWT4U5meo1TVfcG
OTikKAn7CL6bhpfX+dEkU6LhSxOpwjyf1FsLW+t5ThE6Qu3m7mIOkPZRIDJiblF+7UWc6Yu10d3q
+bBuXOVv9DQfNedM6rBrjq/HhVkikXZ4a/nGxsL22N6IpuygU4rvdMdsR8oG77sFAR4hhf7g0IEz
lVugXLQX8lFHAZ8JYE05TjCkNYUJSfP+fqcvaL4ICpvRimQPQZQgmIKSIxpssd55WtcASVUciO/T
5SQgRQHvB1yzIKOm2nilBQUPDeIaWF+m3DqaF1YNHONq+3gEexIS2FMwpbTztEzfx2VG/tXGjSxS
JhUiaMhMxUZVH0XkfFUR3Mj5IHPjRQMOSDiF53gudryvg6wCt9yjhFp8BbQlz31Rh41kUmSDcAYr
ZoCgMQFxc1omEA3Cc8kushXaFgc+uBoAayMPZLx3nEuDAfJFykYcQ/TparNCCeTPOFAIywvyfXYf
C4ry/oCPISK6aYIrJZsduqDvLzHYInvw7JBlalEnjFZaQOGUfSkmBfvRVMDZjicPJRM54Ov/zBMw
k7j53Xo6Pe5vwQAkMf+kqt4ctBpX+/SXqL6/ycIiK4qK6qc9gQBuhJq7nZMdu8Z3ZWHoNSLlk3MN
gwibPywgJiG4DBqiv2wlLDgNAwmkUMM92d8cU51hroC0PtZYPrml/Bh8x7WSCwfUtSE8hAxAHJJs
CeB1wMRB2YyI7hQk0wBy4hzu8dSHx9WHGlUTtAzqjFWY003bCu2uF5dx9UtSRVXLULahVCNelahb
1jP4yGB826/bpMhm+LYJO0ai+N/r9zgpYDGB4xrDPk7WbQ+fmnbzCwLtJH2IQA9nS8XtoYJBs0R7
aBoDTVtIYBD2s0/0H3kqFTy+/9C2DzToLcofBeh3htDui+OlhFyG8Hi7TWq7atcG1VojIEPwRHDC
33UAZGd/UEn6jOm7PFeHYHXhAy7jUB0daBlvgj+Enr+LnpQOYhEFbooxyEr+iI6mwXJOEYPwQ5iv
NbGlknj8/AvwOMuZQchxkCpSjbU7vb8559haJasR1UM4gnAbv8HbSP7r970iLNNUzt3Jc9dG/sI8
CjYVgLd89bB3JIgVLih9zs14BfKLFqpgimF2os7mVf/6YBy/fajRhnWMuIRcwvt9FwJKY6ja7DTZ
4CFXExo5F0ejS8T+mgM1DQs+WVE8tIOADqDfNz/riKl/ydvXa5k2TcjFR8ZMyc3FT1fgmakck6N2
73MBP943dYu4KNOjvM35FgqM6NG748ooYehCumRc+6jyrNLaM9uMJgJMe956qLhwRlSCJMyOhmdD
NJHEhtRHeMTes4rmoO3vojKf2uDmlkv9uiy0Sj9ONnxxVin9iG4rjRTGomlrsfLc8D5uqxFSCPE3
7yD7EfHEdG1Pe9p4/91MrK1LIbchfPMtR8mwinYBfRCwE0979pHnux16BLTD26yTB6zMPkQ6lWa9
tCYMOEjByT1cd4lhS/tAlmivPklXnOAE0uec0hlrsk/ziLgzNl5A2RPe1IUG7TLIeXRODScXn4iY
y8txgLyk1p25WtesmUtllyvK2g/WB3fXnNbG680hzS3Qr+s9NpUESbFdLCBjBCjFhh1Vtf7us0PQ
8CWxYR8R5TYY6TtEdjtfsUXMNTpXL+Wmr4HFmBn9HXQr+ZvyAApiGHABguGxqJ6yuJ43I5pHFo0W
aVOrEJxD7yzsaGKPtY2KXxz8llETeCiKA+bd3TmSQIRacONmSvqbmnePOTWV1//9aXKIU3A0q7Cn
9jWeJ7GCTaRfz+RTvsydB2xrKPFxfHKghBVNW47u1U92jNg+EFWknFVPZXag2vGsFkHloPnz3HlM
1Ghs2D2zsqYPmw1AxZhKwHSQn8SF3R3l3OGltpt+A6yVHbkkjvhi3eerUL+2e2xRj79z0DuJ8ip5
nBvm2TZN7zEp18b7tTYyUJ3S837HjKkxSyRTOQjGm6+p+GDcCqBLeRIbdhET835uzGZ1ypkrJPqH
bGpOPwRPKyDQacA/x0i+HEE5mvLGFbpIcEPfRizzK7sfsr07RQQ+7vQGSMZZRFjpSIBDuzibhbx2
glO07KkCU57o3id4WRlIdGGW74Wj9b6OyNlU4vEcoPWIJEErcj3h/mo8Do6DGqZBe1fLw3P2iPGr
/dOa6qLmxLBjpGFEzoKGiS7GuPiXbjHWThULUIDmX8uQ+70pUYIn82ibdarC8H116HAXYt4AByEy
v7Td+lbtcRra9p7g28kc8DkXI/3Q6Zc4l+kGl2IjAsCJiOwKxMKRdg0V53aiie32lgWjAyOTEadx
z0xsHKGy1QVUKnDRkLFo9zLtMy6N8hQ6j8miBeS/LOGV98p2bWEF7ZGBELsHHXeARSlRe2C8gVi7
1KxEW0oscbM4mhfDDecO13U+OUNeJyFMGsDjQ9C62fQp9iiWoYYeQd6iqwG2SGK6yIgQ9JqIoB7p
Ysn+vnxYM98hyPxJXfvLpm+UAEjdmX9btOb+5tm8HwmVgW51H7fWXpdj4Kwnq9WaSc01lMd+J1x1
uqwasARwELg2OWo9b7bABILmuobLgxWyJ7WZVn5aYD+6+a+0MhCfDl0VFH/fjYysK2AnPj6EhENb
MlkwKj7Ne1NHh8CtOGlJOe9rEOJjwBjU9WgHWkbovKBhpgWQltPRhOyH9m8ImBAwt+lLl7u1XgEW
fnwyW94kFPTGEpBqaP/yuWCAjHVGy2ys/CcvAMfNdWV58dnN2J3G8Lcf5R+tzsFXaS5CBOPOMgPi
glA0pzBZYsTCV+eDsaaqRadymeSuu+MfiD0RPvvjCN0J9pUAL/aPcVs2yS6r/ENsHSJ+EAaRdjWV
uGH4vAdJ1O6apMgmRuL8anipZHVXvtQmQtz33sWeAVymGYO9wkht93HMqze9DtancgUR53FVL7wV
C2byOyTqmyqFrniGMtxsQy4YBT0pDyb3I1IB+CGhmCM5svylGrr7iJIdfjt7Q1cDZRCKv1WAMj37
iUimNnY0IaqnXXOIgWdD88iwmp+7I5icoGLoYEuD59heYPC9mJ+C9km+BnKoFzmFIeef6GN96XBq
XYTv+LfN9J5DWTb5q390hOeCUzdIqg0cYS77fn5Y2Oi+8BWDlqU4FXVV+9i6pFKDnlz1yHMvjIuX
8skl7m4JoFIZsxhnNN6fwiHvuqzV1ooQzZxNexdzwzJHGKuU0x941nDchxEIRH3U7PSiZseRIhfU
N4T3TVA5EpOnWzh6TUuL6tWTMJ6P9yS2yHe9sCvVMgLm8DN1avPY9N/bz4Y1+Qt7HlmTY7Clx4h6
cKsLKIXAmkH3tUjgTPYXW7U/Dmvc/jrCu+CXaXY9EF0yBJwiPZ8oBf1pJjlEw9wq/eGPvJsh16Jc
TC/z+n4+XqTJmzfvcdGVpnf9uiwj4zZhzxKhsWdWpv0IlL2ATi/LiAXotQBzOWOrYeDkxxZXXv41
ifGZSJLa9+IbnXybfppaX+hvbvcha0PkHjkwsUvm0hX6T1oQffnuiZZAUGeVYjM/XGK8x702mY4Y
dp7b8sa83DPpqDlFrG3spj5qkuhmxtDDDhzxVLPfqA5rZOT4jl96T/3KwPxXsAUlEtyyTmTUJZnV
EXbRd/q/D2YZSDAxooyV4MTcFfNoFpm6o5/ATYb5Kq7bTul+8jDOZh1IG+Q6Jxp8ztnjP1drL+YG
d9zso3/e7AaY7bPSEOULi22/0xfjy49zv6tFVPFK3FMNWEdhsKHBgIBxrVpBm6YQahyf7XukxeIZ
vweGf6CmnIr3JPYqWiiOwfsdcrKOAjvWWUoG8yN7gCZTzYPvk2XEHJpLa+LXxgqRWKVO/eg5LRsJ
v/lixTuqeNO4qvF6EbyVwsFJwveiA39ogwNTno1CRU5mFgZbD8FioYrxHFjmuVEljKHzBqtjSXD+
9nxL2znmy/KTlow0lIueGkzjNqLBSgeFmNuPOJJ2LACOd0v8T/2YFHnPRn0ZGznZEqOt13390irn
5QDWxOKDlBGsYJqNx4Ox1a8DLQwSHRtslaeO+Zwz2qp7v988+YFvbqRT/TUHpYXESit/dg/ZtVzL
3A21extOwb/UKfI880g8J1XwMtHX8wFBTeg5wwevoUf40Nh2wSenmrNFskq6xbuStoOrvx77ymSi
tT4jyq4x8KI+RdU4kfWYsChb3af7d/odXVIlKHlCM7sPRwwIik++ErsExI/Jtb+DRdVJo+Ak6IxY
YZuwJ0ACdTC6jUt8YgkiMBeo/p7yVUT/6kNWjqYMJtJ6McZUy9KPcazJqH33TLLFjfoPEMm97R9O
o4hin69uSj24IjfUgqYGwVm949qEBU0XA137Jf6wkDfiZgLebcjjjG//bbJ00mWlBUIlnIs8mGWS
oAPGzJuBn8PXtvMzWie+BpD4TcEmAUqk2vGZUOlJSNb+KOCiRNToMj4Nue29IeKg7YYsHtntdOKf
/qWqYVagO6Rg0TLBkNcCr1bNXmrrkQ+jB9c7fQB0XXWZsnDNZuLhloipjEIGerQiUgsWsJkfB6C5
kKVQxHdFmhyWh6fA0r+L0uU2hNVec9wshIRA7M8Kj9EJ7R3ckl3o/+opjY9M58hrE6HmlKd1Ctfs
qsGSik/t4E3x0mZouixhKVlIKwcxmk1inXRZTM/qzWZBC/FwNsRebeEaL40oJ2MJMXODa35oAn3m
kpjnPXr+pTIrcTju00L9yndU3oE4OWVKQlaqTPUhshJwkv7dHIzsDmHZ3ybgw1M5Pz7uq0c739HT
euJuo2OmR5EQRqN9OHbwkr7Qctf1YxyfezJ+sDsj9Y8x8nsGrublyH5zcuu/SW0jmhbCyUCP6KsP
F22UmHvRqgsu98DuRs/qNCSev/KzdoFBR1aq6ogLfNAvEwVc4QLSQmWYev7hxjfvVnTArOMQUsJn
oaYsW7ai93pWcGLSekTjRt3CJr6fRrIrlnyrF4wv7XUR2x1OiFwYXey3/FX4fJpW2lMD/M81qjBG
gY/SNAASzJ5ZlZXVBsJI3tZg5ggE17M913QcZzxDZthfyO3iswh0BVsWo7nGMA//dnmb2+zt3xC9
Q7eg2KWz1EF9j4FAhldb+gMj4UaUCU2TmPo/93p6+f7Pegq+Lbjzu+pCdMDL5FoOBxJmHFTUXyEW
bHxKcbgUulbOKTLixAkV3B7x4FaotKBvxIcOd31VMyF4J2sH1aTJD6Ji6RvwoWxV8vIpoCxdZ7EI
HPd6WC1eJFrXrjAksn7hbjyPgmn8AVBtJbJJxnOK1vF0cEFRB91CWk1tiLwnKqokWj3o8bSrmTjy
JvK8plzbbDLdSFhz4mwSqUHZMdnXoPiw9cdSuwqHflkrtYG+Z8xb3RfwGsIodYDArlXSi2yp/VBT
3L/NB1XpzSi52V584uqW57rjAfQuqDAaNjeWZZ3Y2qN2eWe6nPOyJLPfsJzQw3C0jzTlptKfOjLP
hc5WDWfoniQl/UonlFgq7o145pvs9u2bc0PpfgoL5kWhk/ETj3WtjlknALOevMaJFqndKymEf+uZ
UgHtQVkELYZ3fpAZgyCZOhhl7HMefdVh+ikEp3LA4o0Y8L7kKZawO8LTyW1RaVg+ABYhpa20qstC
00gieUBXQ0fhxfzYVcG/XcQwk9MIFCvZBU+UiZOLvWL4RoNarDbWvkL3UAS2iQOJUJcKuHDA7eRP
dLH7umFyGuqxYW4pcq6TFVL00fE+n+upvmPVpMLr7vpYTFALWGG2qeqoeId2Vo5lJMdoXCJhXacZ
snKaop8fcyEVV6/CLBor3iwBEGsNs+E96Xd2NckKM0rsSQH/k1nmennoGzJ5hX2sffT1YsZUDAdz
FllUgmI6q2awEeFeOn3KUYsG2Sp3Bq3KB6NtHmw2FBrCJLxAXz2Ce65WJCPh1ayx14sSJnK0CrZO
IcaV/lcJMhjLaundVCGBQzovgAOMQyLZPslhzjIQlnqCFBcaEkK6Gosjg9WK0+iQseLzpiYS+QMx
99Kg0KZtEvb90pFwx/+cpUm9STHkwgUoJ3hcFwxcH5+XUBLE5eKjo52oLlnTbvuFCd5EW3GRy89t
xkJq5belTgRuYAx//McWGWYQc/w1SXtMia0nCvyP3AO9n/+tz6vrzahf5GqA2w2vIpi6wS+T7LOJ
GVn+0TQDTTn+asoKnrvs05RT6A4qpE2DSD0ECaTZ6mKpDscDHMU5PRUtgv+iycpoQSquw1PuGJj8
6FnIA1kh088vJCzhRh0jbG8pLhDX/vqr5cjdQ/ca6DPci3gPPzzUzJIwoPfkrehDRGWKX1tIgZWR
1b4+PFClZHXeH5fEr7ygVzrBmjdonLanxdeu6b7X7X9ZQUuvpbJcydpiqpLLWrqp2JmRgCCTm1U5
m/OB6DfqEhV3PhBB37R6KBPtX6W3W2NiGnPyBreOig+VNYakJ0HwsZmQxOVpHBdTJuZUT75Ah99e
rKIT/sG98oAcYeXyL88eYba4LwbP3TJ9cocgz7/sRbEsOlwfDi+YQkFOtcaKBPDPoYfIlODl/xmj
C3bi+kQHvlWE787HWii0kpnENv1Tr2/+vhRvyX2q8nRlcr50g8tsXcBydQUaCeeqr1FIMxgesHNK
3pk2vRvcdnmCqHqzD1PzpXTcZSj+L46kRIslEKYkfdoVpgD/8djkuDZyL8it3cOGS1LGofABFcDD
/LTV8C+6+VHs3OawkiHvbUT6z6GCcJ3bIBWbDGQLIDzehWo6mJLOG1pRddnjbwgR4HgRbjeAERnj
uOHxopUbazEA6sD6zbEgNzNX/BZAbi/T/AnnW97yBtDOU1MALu3nSfSkAqBRCTcuzY+tRE9UMDgy
WqIae6mBk+1cUSiOG/2or5kcHNv2Q9175cNNKMYntEht0cZWGe/qNc4eExxt0SvygIIZcRzAbJ/1
aRFtvvnDh79RdwOHyfQ+GmQLTcvnB3A0SyRMJxNZfNbgZz79mGOJsMtZmaK0xHI7VWtKSf1ee0vy
nBfjA5sAbtHR3PEgj31uU8OZzo2BdmkzW3/Wt7nzYztK9gp/EYBZWrRCJhKft5TQMZi2vzeGzG1x
82adiheNWRwvwhyVq895Ivck/ti47hCTiZouK7WcVhw46KCJJQhvAx2GHa5t5qNyRUbex5NPiQnq
djyDZtKwbd66LyO3E3lcdYPVWq7RueevhF5FybDzcqyDg7plKYa5W4eAcC4kyZtDcOq+EIM4Ey0A
G8uOglyNXHWsh/4j+3tMuMLG+a7s6HmU2V9i3gsN2LbVavXzx+x/KM1VQttU47phMW0LySyb97pK
wS805nwIk0WCCOzPN6cg5FT7oZv8s7vidOQqtBRAkKAQbZGsTrpofNTFpQ6DR/MNzxb8woLgyf5x
oWn+jKgaZFcZWAFpLRJyX+zA9QvO0T9oCUR6+eO1zpAa0xLjqgTIM39ivgmR+DbHUsVYJ/Gl3Y/c
fFo4xt6oyRxWfcsMsGFKFDSWLn24A30cSgsOvlz9ojgu4ejQzSTvMU1WQeiImdxFmVMm6ieQFyKe
97pfZyp9orgtQAoAKOWmoQZiRGy1DxBfTDPv4By/3k+vEAAYC9NPlyEb4LXCfS8iFa6Jna3xt65d
5+A/QEMBXzjrh8wmWmcMYwcrEj0b8Z2nPRkMCVqZ5Q5mDGgnDmHafGYsR7pg0Hgnn5Th+R584Dk9
pXFh11XBW2s8NqDslLIEiyBtOpEfYaIs1vV8O8Xf6XxP4e7e9fIyJ+9FGCGeuAlLk9JdF2MtIDhn
JJamoAKqwMy4XSlZFZy3rP4qclNuh2lvrCAK8sFcFT8rHt6n1iR3o/Lf/Mt7cakpMQnDHDRi/sKI
F2Lg6FEDSoOhSZh0IBDTVz2gMegz+Zha3U1xkXqAnqrtSNUXzMxjfryg+IFVc74obVQ7WBNt3q/T
AGCyrLhkEIsf3o6n79HYXKKtwpkxnR7f/j7LN5WD0h2WQuISFGb9TrKx1hfeUDEFACzQDbSx36u+
brPf4Svh/x9WFqCjkLkn0Mcs7goTVVNZhMLvpd3ktglw3+wFqjrMabDhJRNwzbcfNddo654Zaoe+
QWt/ApJ4XxghAiTLII+WI0aAESF6+bSBdjVY/dpM6zNRxnfk+eCLwkfQddsCJaiTHXSijt4M5JMW
X2Q5WnSk56DVHmWFQ+1aIXbB/u7cQbybmCmVzf1PjmdnA8UqVMgVulMLkT/iDP3OB518F6td76xE
hyzwXzsHOu8zJMA1ESaJXseXRs2lxfhrYCafdgMkeAq44kQBGwsom8OuVohzxCRjPXHtluTeBRti
9u9c1tX3OVVRjh/RQc50JH3udeL5V2dUDJgQCqW+/2qPsfZsLyegyeUgAYrrTCWcxlYiPiT3Qn3i
cSxfZniPdr1f9Mdhs/jLg9KcLCdeO2JDSZLZaJ5dwCdzcP7VemOYNSHQIVH4M3Cywjs+NNWrAkRq
oynD3w99SIzD1wnPqBjMMOob+ba0tlo8Y+DyFiiN/BGQcIY0x8z/cLPn5z1rslsN67IsPUSMvBmH
ZIupzeiljJbtUvzId5qV1yagolI0L30DNzIfakIeW7vMWfNgF7qxTiiLR39SEw8sVKTFE6e8PS3h
ghD4H5Nws4k+y/pM2eqiW5+xu+rVxw+rXt8Xq9cUisAM21t66IvXrQty18rqlQa8K/RQ/CocZT5F
A2QQ2UCYQmROWFCT1k6/tjoC8EpjYsbZqtI0i54bhwVlOwnVwEzsdzd4ub/nX1f1intIn3uccRo7
v42A2G0+fPIFVtN790TdF+tcWlDV8H0FarefvaeEgaOUvh5j/5twH4Nm+HoLgoLXC9e5EmeUzQPe
wVJvpEzdbnsgW0d/8Wbr/THcnvQ3eje/Nq2M42Kye5xXS9ZzyDwDtgOnN8a/QgcMi9+dhro+P0+6
ugOeTfg/ahFK2MqBYKD4no9QUS+GP5TDwgseXnqNs2VNXe0YmQ8OC461dHXZ51Y/p90XQH+0D/XH
qTODgwAoLXt3ViwIwZ+1PgOYITlciIhKIW5qmY440NcI1WDNrz+r+hk84Kn5+5vs5WIV8zw1mrGw
R9JzN1KiOtQlkRC1pBvAEHnyPcwOL7tysubDLToFv9U4L5k0VmD7vnHlRMksrQ4ZrtUhN/Yp+jfO
Yj/XsEMPNxqCAl1PYdII4C/xOlqY1boIUAIZ5coJkx527Mv4/T/+148YrUJnNjmEdNNialuZdTCH
C0mwGy2zgYf391bx1v+0qLdS8IpkxXRowbRXTtmIoKclwivPdmXcyG1YDNOHtIew7erwAtCvn7XO
wj6GGUc7cl1pVQUzluTfK9KB9IVT0B6iDaSaGVdn2vnXJ8fr4yr7wvdAYWWtuR5aUHuti3T3/wZP
ij1zt5fXBXblb1tl4qmZ4EHrmUZGCx7CBaE4A5w6g5Y7NgcgDeD6FGyYJVJUBGPsZBEZVxl662+O
rqFAc94vxTVukHE3NLG3aw/rhBx2Cv/NTwtAx8/b3GOrT7WCJGIX/bLCt1dHHpHe4MrtD8KEuCGd
XiGixJUFQLx/UA/mkjJXqQ8CbbkXpwcLLY9ouA5VnGS99Ie8iNxKTB0Ar5kHR9DyM43bF/XSOHV/
fuzNdM4jUkHjtLLBiCPtZEQ3Hso4l80wMV+R3xWgI0frKcJDge8ClPxxk0XkugluVGpjFDJywuqb
0+y/VwJ6viDlT/ezUONdeGlGNXqWqbXN/kf41C5M/LPQWqzDr2rUAY4/hv+dciMBh6agHFkD+KaX
JVFQrQa9erneZ6C1zPKz4kntU5hsM0oy62EvZGduDSiLiQ+oV4QT3oBQmWU0iecZs5Se8NffkB7z
IlKrcgVt0OmtI7dXDrJVWugbhWWRNn15AdoZgfgBcc5IUE2f5ZzQJ6skB6+9BklHaYkNFNKLzgrX
mk5UEOK2fQuQqJGn4cx0hO0bjWCesvi6ET04cZZonJ00DAe5nCVlYIOJECwN2DlA2uLZncobqdLp
0Epubj1Wc2S0xZhAs8yemwbe0SUKASweAFmZD8rKYlN7AAyBx8IC5e84cDsGPpSqhAWGCBNp+XQj
4V1ol4wRdIfFcROBFCPak6Kq/+/TTv7w8iM7VOrjrxg3JCxVd4FPdwwG6zzWbBDL38g7UfnEqbYF
aijJlAP3yDNMrZTC4WO6jVeCTpiytpIeZgMSM0+BuLrpx/EeJkEIms12w2bOF5+XrjzJcxL0XuHp
WIeB6+mwQPqKComdYwJVqhmj3YSdvHKMkD12hd4qBK+ERciqjfwQ8qe9ALTsVTSs7K2I8BCZeCIw
GK4QRc3eKXI79knUm/+Rg4nrMDcYGHkkfKQpCIQGnMoLTCQ1rxRZpgBjk2RCdXfS2FTnZe1LcxJF
dRFqt/XPrIINqvt/7VpIU2J4XwuPnC3sVE9EbReoJA8hHogQRdhB6skAWATJRIJwsAs4ujh9GBsr
LMDuJFA+WkjLThJni5D099soa5yDKqQUfd6yV0IkePk1Uk13iJiaEk+oR2nSqF18Xlla8IrY1T3D
l8PPvkG+mxyi0R3/fMFv+sUel29PlrXTrTOvuwjoIWU1d9eZZ7k748w+BH+cHBXZJlkiuuUboZOq
I4+cVj6mxTiSl1cTZlVMca7VN1UrfYUSOEYjvDkIkQtG8dXzyD5xUIX+e1SUaZclw4/EF6eBjr2h
ws0hnmXttdeDEFXKq7lOO5cOxHZ7XN7twyoXeSkWvm8HrBkDTACZ+2TQOcC+n70PCupIA/3lHeNb
NmCLtmbRfJN+Y+IF6xd8xOGwNwHVA8N/yIseLCZyo6Y49LrtBslKCGakgTqHcq1j9QnPht8Rwk+1
wZxn0ux4dBv9V0jzbladalw2GOKKPgyKuuuQ86xO0Q2QlNh0jnivv5GL6Ju5wlB2ubrqijW5HHl7
GQyVVfBzDE82GvYXexInDznrawCGaRRTMrZcfvzlZ7f3KtGxK8gW14sVwwgw5xqp4MUFvPh9k0ki
jeRdH1s+VCmnOlx2KK4/fi7kVG4Fxg60zT6MKj6/zDla36Ofj4/aMS4/mPo0diHYkLHym3N/3iYW
vDlKy/ZiTN7illx6VSBM4dttJDcyFAkdXhGekrYJqSBUqscwGfbOMBXeojhlTUS/4C6E4257DZB1
IYv7Mw9wc4WDjE5uokb1VmOiRQmiYaZgsv4dM3f+hfvf9ndb+yfC3JZt1ah5ftciUsIgN8IMazPN
2ymNyuA8iugv14Xm8Ry7Ey87wZeluPzBaeoXSYnTmHXJ1m2CXFZHqDjgMAB9Ee8Xv97c+/i+xkue
shv/m88FxTMccDZ8gPdt0elLj2vybZi+QiYw+q6XkR5P73yvmAHYU9QtkQmQemgqu5wakI/XmoaG
2pQBm+PRw9C1o6Yv74GC4yJQODohwaAMRoywLzUhhm2W//d3Er52eR3In/SXSewVqE166ILUS5wW
Kc/Ybvf0bjWVcy3TqGXjaYlEZHuqne4KSn+qiCF5zv1P0ZuViZOtmIv7mrMeIjC+JH+bfTxQT6Ye
xRq8/e3v1XSVmWw/z0b0WNtQfWx/4oty1Z2YyPoQPOIRsOTbAOZr9pEXMbUhDJMaNqetUbkH3laz
bX3eOHsLYbco+ftoa3KavpDPQtHUIQMKh3slyOm6qpV61OAkWD7NuRgoAz5P9Thjk8Yg/wbfatpo
zcygXAIeRYIsc6xQ9s0wnfUzc7+IYaaHywhp0prad94DvFO5jvZK+INPBum4S6QRgnvliFwhJYMg
+Wu9e8vnwbDwtxahB47uCwNnuklDUM+Xw+CymfAD6TS4vId1I2U18gMtF8o9M+XtLwJqHZqn3OhU
JCWXaGxXE5oH/+i/WZhBrYlPw0i3BtaBLdhr2emGoLNRbQU051hw2xM7Kvs1eZjsA2OQFx7aysMc
on2J1FczBJieUhI5kKYpzxi72tYdnUTloni7qqrTvgeiTM1bPJnSpAmipyF9L5W30XyHFZ1Sr1Oh
9bZEsaXlHz7YGcTkJVWwkqHcVk+O+60iBaQ36wI3ZvBoFznXBkhtBrf3ZWhM6jN2Jje7b29JteJ7
Wamm5PQGkKS5welw3XqJHbFTeE9s3n2VALv+mNEkh2toVYLHYk5hvp1c2ZeJu8/BdZ20MJhJeQ8b
xfE5GQ8E+sGULdVZJ9+syMzenUcP1MUMf9jKuYKcA9VE75CldcmM07ur0XRwP/U4kLCsvfmpxkm5
AiXdN6gDvgtChlDZxxeX+4HcmaCzu3tkQy2h9desd+yau/T4cTfq36O538pvpYFadWk/+VGKf71Y
zmb/P/RkzP+/PPUR4TUvTvRXSWY1PLwmxsyVrkoB+sUhKmDzb5jZ8xuqM8WBu3RoFvdK2cAE+wLH
6Id0tQ1nVzVuDphQvzlXT+SheTG8DyFpWDPelqLcXEoN+qQYfEzpSKTlzI5bTiLzJi8wK9bFZWyc
xPifpETaPbHz150VIZqsvc+aBhcURHSsyWNIR67P0+jb303unl0D3qFAV7F2TEl8dOdLwWxs+I5s
8oDCUXj9r3siuccCyjYmJ+LUO6Dlmig9YdML/FjI7XE4EWJYMR5ci057gl2S6yDIUCzeoyjGSObK
3Xrn2Wlw/58zfto4odvSZJ+5godr51khzNaqJUyPvREtxneONzc0pjkoJnL8X+1ziYPlEpwHG5Jf
09bQY4QK/ielHJPJIaWbRyD2IFTrLONsoPPnpbkDZ6Sh5m6dk87y1WVyreSbHPVAGVupVfXdURLh
xf+BIHqSxXh6lyy5Y1Cl5c/GTmnsRBaKoOOtqGBB1qxkjxH7PqXcySJpEWVzGUikybhYrj95q9o7
LzkBMalo2NjCAWmgusyO6fTeh3jwTuJSAxTxjOyCMJISfaklq0BwatOgJKADzXWlcoZPYGzxDAAG
luqQTbNP2R/4nFqxcosuIeKTGwZAZxyda2NuSB5vPPqGn/tM/T5TDS6GxErUe/7xzExy5eupehDd
WETqKS0NU4zs2u9RHlYGo2Ax56KcZ36q4r48FK4acuvh1uKSXYICCDBrTNU6VOFKeDEAs4G1yZIq
6S3EboK0pl9lGnSxLzz6xN9aTMdSG7fGTeYzgle6vcT8kB+ZhZAbD0z/jyrEcdApx4RdMwYJc0F3
dzgNkM95YC0JoSTDcCEqwYR7t1XufWbkOAOr5zc8lAEsoq+ezmToZ1/wmw8RmhYJc09pGLoLESI3
w6OcTerjSe1pkH2STWPo9p23GtTtxYe6kI7wjnbcGRPBlYdYzntI9Ido94dZa6bH245YYKWumKJS
GhB6QunXqdeiFp4hi1f2HsOigTVViTSXkIu6S1Oo8vJuJq1mAe9iFhE6125VmqtwdK8yc732b5tB
gW26DG6JDVQgt0YExAZmneBjUgI7CJF0ckcYqmtOT3eZVS1qlnwDAMnJpgcWUopqMAiXBPX7d17A
hs6lna0zXNWCtfatVY6K8Rlx6fK1Lo8v6lHFxusTMglf8LiaC4K3a5NyNg4OOv2b2Ht4v5DcE3ok
rYKUfcnfhziea+5G8uDipYdEndx9/atXH88GjKuQFzAFRzBVkVWTWyYrmSp/kX6/AN5LDVlUL6d5
Q3/kdrmydjP/7nwajMsTLxoobAn7SxfNOlVshhPFBtT/I7win7E24Y4q7wge43aiHeLwNc/2a4+4
9HLoEAWQ5Q9VZp9WNOqxdoQkaEagvrT+JLQQv3kOiIEeshnEa91qdx5Nszq3wxGvrN6wjyxSbmwo
aeI4In80+Dp+tWInVaAYIRQ1rw9/0Q3SklHhDsgr+iCZCEzAmlPgc4K4hYiGIHi9E91htS4/cmiE
5YU4oDmPHU9kjZDVXmLELy6Vubqo67N1foBnNQ8n0SliT9DoDlN/n1WdehE1s1i7vQLXTj+IrnYe
5h+4iNsWwwGcPXd2yZqpJAtjx4hiwxtJOm2F4Y9CFL1N+8d584z8N3fSHNoW9J9fhyvcH4mt3dx5
Rqx3TSrgqGq1BeLVk8a7pN8ZSXdkjTs0fSovRx8JrMEAwtBi8p/u9W5mFSKsSv8qVLb3Gs31JhFo
TKE48hff+qy7RDBFhIUCtBJyRUGBQF9/TEm7ZHzZUdjCwCqQHiA7UxT1ri8SgARJn4+7NCToBQx5
qEIkqD4swSuDhT8ynmsVkIV8HKmRD/hgMAB8oEx7bQrmp53TibW/vXJUQyTfGc2h4W1x2O4jLU+8
EA9HGCGrSLMSD/rwD5Ny51R6EvWzWuhEHRlRnmyNzkPWPzdwME4d9U6pu6yBXXNp1KWYF7W8+/TS
JZxJuWIg7h1WCmirvmOcMnkaK844h/OTCUH0sp/JWgFTxguG6xnfazYs9KZ4SM3YGoSV5kZJOx0U
vmez+UZujw4JjdxeT0QT6GurdiFshVXq/CyCD7jGJAmbMjFBjgDKDen9Ky+xmUNAW5FzyqnZoOBN
g2L/EL1RBJS9vTaMgQEY/3FZz/4zh577P8sN3LqLANa9+9aw+nrg1x6Dh288+rLl6ErCo/954NDj
wCJoEl9f1mzSJasDCAKUgd1y0W+4i0wqKJw027j33YhYmu5ca50ZFrwAqqDw9+8CrhXiuavZ3tp7
VibxGlUhM2WtrYZVw5AuFzTGPD6M2hXlXQCWxYlwW0KT1/xVYurSen2en/UuxKtFim8k1uON/Ghn
ipaEPAr1gcsbMAioFgxA7yR/St7/HLQMX52MUDgM2uo0gxdy9FHUR2mH8ovxfimv8Y2Mnhi3PE41
FwHCRCTWLh6D7W5Mkb8dNmPnHpjvjEOLZEjcdY4XsQSlUlxRYkSnxtEW0oFCQIUvbZsog6/GKofl
vMHWPBPlcb+iUItCuAqWivFQ9xf1USWZd7WdWLGMnejX3RESkzfCeyPqmnOx82RWFHyC7OEK/N2o
xKbDHDa7/7YxQ54HWFlCnIpxeD8TXgrVnTkE9cx8WAteRmp2tbhqitvWJiSusxcSTECNaQR71aq7
F246yKYWYSAA6RqkMIfLZtp2xywATlFlFpa52lcIfqoo0/OdhLpnWrlZUoTdcaIONhj2nyb7gd/Z
I1MNP7owQnaG4DtOWz4udLIObAKWVqWOpFMg3h3kal9f0QDokms7lpoUXa5hi78zPEgXKZWeF42G
S6w9n2dhFj4T4m0KbsH4wkYtGrbq0/ggQxUbJ8zy54eGkmJMFQnCox2icSsB5Xwaq97xJBoSYsxf
3kYfUcKNZjzoA5jIGTkgR5AopBFc+OkepP2342ZRhM2q+TmH3S8RRA8Wgr2eq/qZfCUiLOR1XsQx
y1vVENjKv9x0CUno4ALBUc8zt0vZt1zzWED589FVfzkdlL/8zUh3m5Ha6Egd4/aOsXZEP26pFHbl
IBBhf0lZhyt312gmPCs/ZhI6o9xoLygxHZRpEdnF/4qEAq/nQkGMfXSQ4Dz059kdHtgfstfqoSlU
um2kE3PWedQp5ENQIMxFm4CGJIaXDZwQtN0wIlbx73L8rkrVWohAwLhJ+l1rM+VncpUy8hoMv1Z3
lXBvH8TGG5gLB1vkbwVCwcnwva2FJEHKGOsfCvagW2xDiNmbfuK1pXsH4mxBQKCyl443/Vh74kzN
sxuKw5CyzO1sqMfiJaxQEOwReNXD0Z98bxG3Osa9tMSLSSWnxjiD9OstKCc0EfpCwdr5aoLGgivV
gTgpIF8OE4xGdwzbmiNZ3iL2By8/kL/O/sbeBdRTVa1gMC8nbgKCkdKos+ZLa7CvuxPqHez2GdYB
HuWlRZjC6OIjYG9P9aOk2vGgX06ULOprb62JwKfQ6SIE32nFSE/sfY7uayCSt2TM5dRbWExDPwJi
3A/JY4p7MxDona5t6Zsd9xMrnKpqU7vTWeI8zRTXC2OJ/f6mz1T08wrzQe/pVcmocodjJYaFsf/2
x/o3+2J+L1B9J4ydMyUyy8zu5/SlYfONJgqMRRLbTfDUORVeISIm8/xJGt98HUu+9xgN7aorPzgX
++W+XxxN6XLBB/0YWnLXY0k1Bt/W27YQQavMxT6XHuQrKK0nFit+TsuVfWjffXP25HD6BtBwaFrE
GCXt8fdX9JpvxO0m57SrLzQVx2jjn+LnNQUuUti302+KGzUVltNHlBVIfOIn7BvjnZuKwV9f3VzT
s0fiAEhag/p0v0iWUdsxLzUTpPkHcyGG2UVypjlb5Ak7eHHOwcHm0iq//3EwcwaofGD6mC8oFzke
IJsgIUpg/OoxEKIQnEha5DGUb64EkAXA0y9yZkBq2vUl62TKW7yOY29gAXvVuVhfcfyXviuNhhkM
4L19otZ0Ihh6H1woZ2fjEidknNdw5DqSU8ZTsZbpe1mgy1v7zUdJDw9fhyA3ElA8H+H1jJvbic8m
T7qkwq85vt29UcnLVJmsGZopQwTbcBdexEwQkhdXlER2qkNFqN7PBIxIHfwRYXstUo8lutoLTJG+
WxbrKYaXn5RIEM0patt2khI59OAVJtnudy1ATbW29lxjAKbTVAEeZRYEVxZvxSVxI/J5Apf0Xxf1
6yDomVjSu/36g90qSj3Ma8Fl3CUDZTs7O/FXK1EtlUouu8pjSQuTPD4zYKA3wql+YiXomxtQQXbi
5vTa+nr4nqMQOEQE+90AqCWpfb1a5KoChIwMcTf8L0IJld9gAulxHD7UEzYOyLJZqNptLHxIq/Wn
0WppHzJ9JK2skTTqzeauEG/KuxPQjreX2xFiDRwS/c/1RuU1HDOYuBdO3sZSZ10rV7W/ygy7wu2F
mP0QOkYi+AvBSt6mEm9aL274I6PQBj548WBfPpu2A79hV3wzSA8tUa21wMT+w8CekOCd0mUcnDzz
KRIA7NFtHzf1DYVprZkXN6UdHA7O090Pr8xsLaFSo0aQDTxS4keXoA7qpu2IfBHguFpAHgY/krsy
uMsy5+3UzCrza1CkQWDtuVMQcTLBK5KTzMmV9K/SSHsfXtOXQ2rDiVvagl/ffEXI6RG5hYIe7dYh
+8Lxgi5MO35M0hxbeYZIczepcmG7/Qb2RksGUMIem7KVo5IFnSPgghF/j2hjszJlttEGbbj1Kuhg
ivN4B51r22FpE0yUv6sbfNMOvFtogeMp+/JEsOfFQ8cTn9+amsWf7dSqedbQmDCAFWT+1I8mQQ9A
s6+qKbTkZAyNmnFkMvz4TmFmNKJZj9aJmF81JHHiaTY3Zr2w6w6f/EIvgpoNCcXa191k1pbgmjec
j9gwI7xIDdC0YTNEHaUGoxppjuJSGaL9/udL68UxcdkPCoaYH0aXgdm3OvGZa4/FZuJjJUrTx3R+
yZu711nuI9Wbb6Q36HPD0DSCh3EmgJxJzFV49T9mPFkOhkleUUJpTawa/6cUy2LhUThgCAmqhH+t
n2zcVK/xeReUsbn2fSsWP9cvCd7uqyYumC2ThaFjiSEdg8WCnJONacX0Xji1AVJAXeMONzruACzU
pPH46lftfYMtRPcm47/pzLh91TeL3/fo+cVRu3l+gsReahVTvJmRIwNtYSq2abFWtYET6yuu8do1
SH1UnIvRTucdDT66KIAau2sIMVkPyHcnaV3OamO+8Nszx7XbDJRk9E5ncHJFqUsEjtzVaosi6SNn
KHWzVTffOWeHTAdoxHVqLMsBX4h2pF7Q19Dev9/CjgHjcCmyI9mqyRAHoAHwKNp17vHS6o4+Orvn
ctPv8gcWXYzB9UANzyJCT8BEgrjvAgYieSQi4wE83xedRuMboAMBU5c0u7hZ48J1qwacNKO/BjAY
hjItQNeCUie7Mhj3F/mqy5F7TEmsIcXxRR0bpfGg+GbL+ZArbyQXXu8FMjDsvIPa+lB6kBzYCAIG
6mvAPLgXR21pkOH1vZVOqQPnQf6C9w+s2GVvJ3oFcwC5vchi/2Q9sWhSxn5vyiXPcUVBguo8aXSR
NYU8Y3SYF/KBkaCAbL44L2yZkSeZqBfdswcAq5ad98dteuz0HWVat4JFTAGPjhFGR3uvQNq2G1qb
ld0wHbjtN7B+xzknelm/GJZI2NB/jOblX8TixcmdgSyCMJ+YCuVlIkfi5PIybuRb9E2SCiYqU/fV
0sxYBczLza4nXd23de0QHIR3hujx3SztdWufCkf50RP6LLxGQMQpHiZ7GWzfZYNVnw91ZeVC5cGY
9JIHzQzasCCg4OFV15uo00bDyo5sr312NhJxRBCh2E5seHvXLRZ1TqYGWFvFOwAHZy8VChZy04bN
zwKXhNyDOV+zjBw2qQcrB2+VYnfPmMgrrMQ0yyyi7J9quIFoEipWpLqcdBKQ33ZKVaridu/Zo0mk
PewybVw4o205ZUssxEOfIDwhm7PrlQD3G3sFX5YkOsRvOU/tu4/Xg04eayBjTVZtN5nYqjcyx+D5
94mK9JCCB51aNh3/4edWNnMFPqxy8MVLdgmrPbuFBa03b5PAc3qXYUDDIPVM+XGI9BM5EdnCxkz+
pzI+EGPHbgh3ghjHOJv9iVzQnztxAGiTDSDtRvzFXwn1cIvTJrCXQHhdxMWJ7ezJ2O1g4jqkb4Ly
6n5ftkzVkLtbb2pNKF9G/YRMDrrp22kR4XWSoz1YbkleGUJIVelQuXgKxdm9lvDgG1n/Uv/DsWFJ
uuEmx9X+XorxX3OZp2yg5cuFIiVnLcWeXmd8PET+WXo2QTpxogtEGmjPsecbT9jd3YC+IhCeXsnw
YisS1NiJjE+1CsMKm8uRC9XyKH1wP8DZvPljdt5wgveDhH10S/SX/cQ2x3NbuAaYya79ghCoCuIB
rmfasB87MrbdZnFZM0H7O7deLGGmUXFPf6njaVlUulBtRVLtuxL1x/BJp0H84g6b/hW8k1tMDZ8b
9c3iSwz4avM4/Ov7qvC5ni79cBtrgkIg0a4OTTzFO3MhaRod4C+zD4PnHQCv2H7n8JeFBQSQMOjy
1B5al31QATEiyHXBLV2Z+H4K+fbWqyqLoeVvSTW69O6Z5U00ZYxjRbhjGvXzqtjuFQj+wf9oJwXq
xL5rZ2BEJHa3gyb99+Qr5JcTeDo0GartX/uMQfGVSZzvlDgXOkmvZQNnGh0rl2tKUPyTkcYjUvX8
YCbGxLbwqvMVR5D9fZcHxaf9V6VI/4V2DHmGigfrgQzw+A7Ip/+ytfjO1mL+XEnLRpcLoxr7IoID
eKMhV5mRjA4UDoxSqsQ+YO+ykOF3XT0t85Cb3CvQdubUTP3Qr10MwAOu8jpEqME0TYD2YtWkKkkf
i4FuxyV58FTu1lYb+lxdBei7F+mcxGvKee1N0GPhMxAIrmGCqQSz1IskqKpO6OgvBMj8EN3p3uVI
EWf9vMdmRmVIqBGRUjBkom5wFKHMO2wUyjyQ7XZRSJcsEchQ2SADWvRVthra8/3glwdmKm06o5xC
ap0SXcccl5ErjveB5GwWSr1WmtOpPUWq+tCMEQCsRSoN/NwoG2bs1x2yQpZz/pa8s39+nGDisrSa
Yy97+M0ut3OeiD6zuwbFFgucCrqmjEVhZ+AEXl6i8YSRQ2XC95hTpkIwh9va0KAxYbczf1VdTYab
oEMJUYGxsb6k9eakQPAQhMgBqTux7wwj3RKX6EWEP9G2VmJjgmLtHA3TuFrHhaZr2LtkhMYMlKX4
UinU/nELIYkCfyE1KD6szzSOMwRaSaXz5WYCi6P/DaTgDxoq00bOV52kWHJUxDFzctmsQmv4eYZS
3xX7eiNWzl9lz6NfEDQ6b5Ujlje3fD9lk4L5skF2fxekzDl6Y54nF+ODGKEu5n+aneEpbX7Ez0yT
8mWTrlsLjc9keLc09lKz3gzlYz+5/8U7CsslKn5azXtyuTP5xwkplkWOqhY53QksSFsoFax/Tmkc
5VBRSMS9mmdliVmEU3/wqe0PyuZp09Wv5F8Gs/OhDmNHAfyZE7DvjRiDbCBkJCzKuAWalIduS3wG
Jynl2aZG4Kp+0fZlcp2+V89Xz8piM1H+ht/T+F8/8rWlsbYB0dLRrxhDZHXfl3XQFljk84bAqs/p
Cx+mfT0Hx9pjbmLXEdhAG4bNvOX5o1EorhzBZUgBbr9m4T3x1yD7RZ1OJN6y+O63cyJ78vYsXKQX
ZP3p+s+/stFzvnQP0/CZbsCcv5Wkubsx5BpzCQnLUStDeirAlCGCpP3BN/cOYyLFR5zEGaUs8TNT
OeDvSyaAtPQHCEQS6gxknbnwtKGgJhOa/u6wMQsxbjraGEfuOoepc8YTR+SaKJIQsVJI+TEMGN6Q
CRIio8AhFtHvP4N5QHbmSedAjTenbKmLcOg3sx63Opz1PpIfQ95KevTHak5igzuW8FeiE+0EvTTV
qTkqUDWBPN0z44UJxFwSDQW6qOCv+Jbj1CsUZQXBrUtiVVN4Xhig21ab2cBTP3qriEJm+evRtTDa
kzcYFHUOnsW/ql0g4gnaOcDgZYXA7susPlOe2SPEyPByXKSKWZsz+6m7jfZ+cClDaBdy/hvlNcFI
gTLzqq/aJPjpC1VWnl7OtsTOlU5qcbnzk87+FEQDTBuwsPFz3z2CdQFFQTjg79Vr4QuOBKrowSNL
pOYcdQua/u5U1JBBK072kaSD70s+P4BxuhDdIC5xF4/1eNWL4tHL/XVePHu6oMM2RpLFEiROyxol
8CZAW0gqY4RejOvL58tf8h+80KgGlfProX3gzNb8XwF4NJ4iL1DmvfIyZo0vUzwiF47z02dxa+uI
rtp2RLsT/GZG3flXbUICJuVpSFiUtG9xIzxwwmvZixjkxQHf/FDF9NkJnEGv2KdIApjbvTDtznVO
j18dY+TbgtAEitmGis3+92OoIvZrV9rDYT2Jt/E4aX05gYs04vCGYxUYNBE9t7aCGfTGlEqRBycm
71mUeqhYfReUoAW6CvkU8+Mt1cdMD755jAuoekaws2Se+HZgmW5R1IwhZdS/5gR9sk1+E+qovGtK
ENxTzCq3gRk65HbwhryfWg04Fj5E2LoGqJkKiLXkpX2kDn8N5R5BCh8F6ApdBawtAFxqTZdNhT5t
vzbcCKgPyH/UypMFBlDHtKmW2Eq+9InM56WuS7JCdeQ89sxkXY5P6CiVZC/7T2IvgQxRTUMwbnLq
iHqihDtA5a0VgEeZ6tszquw9cp5vZPqwCFRdtT3JJQluqRykjSoN8qPWJ2Ozz9FRxvfi1tjkQW43
wKwDD8k21WPbwRnAz7HBKXTCjHtG0svs6yxz8Xm4trUvtMhlCkf6BlzVLGBp2gA7/Ia44VARI6hO
mclRAm9V5N8SJJfSFz2FI/kQAIjXxR+DECh4bDnnl0kfXX26WGrEcywz1w53lL+sMTg/PQRYuSv2
uR9iG9cZBiCgQFkvbWZL7ifVefcfq1UeS8d59LU+djdbFzZf3yC7wkUgBimIf4x5ft+9zq7vXgKu
DHZKwSkoFTVIB6cwYNrdLuzBiY6Kj/ViKelVqcOGpV/gCYazg1e3416CUntK7ERzn/8VXE21Mgqy
ag56YNuScfpAYlmftRW1GZni+CMbwfuQEIxoWPDAQ2Y5Q6FQblGvpvW/IVEq9krk1tFPeoYrhmFf
khUcAzLQeSc7633QKq4ee8j9swB5vkDyhOcKbHgMywX8oSZz2M8M3B4ziyoW9HdcHX59m+s9S4mY
eBYRrLFS5pAkPtX4TlgOrAmjrK7Nu8LY3jJaj9eEzQp0wfPFKEPh00EHBjQZu8S9zATWeVR+aoYL
xkc6O3xnPyA8jdIEY57ittOM1IZV2hjlcsrlU7FvdUNmGaSVqPw9y/y6s7c+0OX1lhFuIN9Ykjwx
1WdabxdcvD2WPjE8xpHK2zruJxKvdl/0dTQNA/0oBH5dI+MVQcK+LJqSxE2hgkOmEiYRWqZEO1qF
4xl4eMmiaP+mOkdCAPdem3R7w++NDxcrhT6I6oTGZ4UHQsJBeTS9UaHDo9ZMZayKL08vezXdZT0Y
3L3Q5O9QaT/WUSqHCyPx48CagZJ4/Q5adlxtnQKouRLxtL4NRxwoJ8gdvXNZsl6zX8TEupZ07IwE
gpoJVo6rDbWlNfEFfwTN1NfldQEFRWaK0dfZ2YB/tY+MgHYd8NIjOUIlT3yfgqTVEeIaPOZ8pHhV
9hWWlF+ayJCmzPLKyQdtUXRwOv5bsQ9f7h2Bai/JWFHQ7RJ93Qx82YUJ3ey40iq3kOuZr+H/kpfX
YJUBC86Dw/A7PLaG+dqMNMnJQfQBGEFwfVTn08OgLembnE9jJ4b0986XHmVgDTQ89e0o7pqtclnQ
wF1hXcoxHrH0paLsBMFSrE/SO2NTOkVuZE20crYaEoHW4U33esPOEQ8W9XWJhypEAwD8jIRnnhhR
BBOUB9ENZtMx2xB4VZYBFHZ9GYMQiN/YBsi7EYTsuVLypAHRntAT1Kwogra7Z54Aw+BNl7SGkEAC
xxTq0LNCep4ym0iCEFb2KqGr7ebAh3WcIoBSHxEGK+dL71L1KhnMjCWzLhyvvsA5PgDt3we3uQfq
u3CUUOYcseQ/6pFwlKwB0fgFf1kWa1v8joO8GeTtcb77tRIcU8/kGq2USiq9GKSCzR93sbvJ20c8
a9ht+5TOgsk5G7meAPj4Qr4xDr4bGMMNnuGJT31OisfCBM9LNs+gDMKyP0eSJHOuclGWzJt3UP9J
mud2UNeh7eX7k/Iyy9itCqy9COPp44alCMLn9LzIgXT7yxPp8uWfjlDY+gaUH1j2idhHxeRcaPq2
BsSctfzLh8GOCC0BZy37GbvR8btFn5pYs4A9V+jBnKsioTLcAMqAWXEntcuEjLAf32YcloH3701r
6S0mfA3VHF38qkEEYQED9e4ZkWIhww5uCMmoWVy66CVXAabWZRX4k4dAEaG1dMfYPHusCLaizd1N
X/HnlhDHktU/SFrIFUe8uhhXAY0j5Wsa3ros0Da9TnPe0etJLJFKhoIFxBrR9/niW/kj9PvgjsZJ
OmNNfe/7KHeKOaBn8P6FRyV+sqxR/bP9mB/8TSzAIDltxm62vopMsEP5owmnX6Lb7jvCezeOg0qF
X1MZMVDrs7kbm82EV398TWGi1H/VdY/KmoL0Md7GrBUOdwQkRu7kIFHXynLwliHgut44u4MkCSha
mCGGjEnYY6/+DXJ8bS0wVNxhfraAWFA56XvVa5/A1osO6xF/B5JV21zIJC65uCqeRWdgj2GIYCyJ
LAh549bY3RWnscGXQn6A9in4gbXGzUt8YeZ/zl7HbGtRBxbGkXPjcbX1UjlDHi4hKNHxTv9FmLQA
k7NEvo3guNXbs+s8wORRIoOEXmoK1whQU2gC4o/5cRdjvFVTiGKKGLEDrjo95BxM0jlA/AERXp2w
5HAWGdLEVw9wCB6XwqYTnTXDKlgLkjijdzx05GvCiUfAMsdrxT15RCu/8bAjMi2eBGFvBH+Dqj3g
EMbh8cKiUczXyRjf/tzv3yfnsLFDFJ9APPyhZgME7mqZboNDkS4T5i5DtFyGzk8lBsQfWzsM2BVr
RW/JSOgYEDQZb5gPQcRPAKV2jLC+7SFQLyAZKyFG0qHc3F7yE2uoM0tNIFwiUGSJQFFVbjYpJDo0
bq/4R5S2b1sASE3eLen9M27NUjjeeXQ380jKj0M70QxHibejdg+pQbOqw5APR8JWWFAYXoQaZnKG
km7F5uY94T6/K5Kj7T/hQ0qpAEB0Z6sXvwfBmlqATq0RgnNbGvgKieqRTkDStiuqyG9O83VnBJ+n
TnseTOyyONH70zJJ7KMx/+dL1YcOzqmhjkjxxns5T0K2DHUFQpIqlWgOO9fR3TcM/QkkuNQyf3hR
MpfKE0Lr/q/PxFOKRh3cyYwndQ2tqmJM4Fs6sAULowPP8sWTZtFt/5bpYj7NIHVD7l/rSrltnBkZ
s9FSBQNIjrRRQ+qkVeFIylr9Gg70Jspe+PiRiljhSn21/u1/RZPwFTLmVGifw2wVhpRXGCjczd0m
JX8ErW2sPnwo+WnuMp+HsFGUZ0INZqSo/OvQEAkETtAZPYNB/IW+E6h3nfixs0b55gDBdiRo/DIQ
GgK3LSJYRNrGfAo60plfXv1q97ud0Ttyb2wvjqsOaccSq9LGdQCH2qP1Idh6r+INvscQpoLwKpqU
A+HwM/ww1qrW0IX7CRoKGlTS0YWmiT2elCQHmyY4lGrcsZEZiV+gZ4fQvZIhWcAihI7rlhBKKc/j
LSivQmsAx6MOqqz8/e3X3+iNwHvXz0T48xHEYOcYu18K5I3AbpFsElh1E0ShkwOXmLy8IdMevl9c
d8xV7POmyevgOoAgXDL5fgNQ9CsbCq1xt2HPqE/ktEGbqZkCBrLRdStazR2HZ9umZFtLcc7tOxVQ
OhfA3GgeV/4cAuvH4HgFI9pyPPNcLxUINPRnEW6zu4Vdp5tZKmJT7gBwix3yt4ihucMXbw4h/Hic
/78cdfbBgKOOair2ASl7MRp1lk9Lew6Ris91X6GFBoynuLxqyXGLykFbL53rpWnpq9N+9kagRqbG
cWeZdVNCwyEKSfX62kAfARVQSIpn6LLGehtg7Cjstsuyhm8AP3n6DhqTRYHHFDtcK4JmfwusvF1f
6TZpQWmmC0Unj5ycyXfXreo4s0hJGTA/S0NrZM8QELB3OETmH6ICLMBlxC59Yff87Q4Oh4wUUCgx
qMOGAjrvMYcx5Sp8mCb9U6LBIK6DewapF2+zxaZargUqw1N49CAexew4RWDGtWaQhZo9IhDRffbo
ctC9O1GtLzLYN0O4RfAFGlE5MrA9MgvDtx2hPi1GCN6r38ilvK7RH8GqzCSkk5DMzq1Kere1cBVj
wKi2AiRfYT1C7dnDtTc+41r7ThgIwEjgdP12VOZv5PVh2RD4G5g/3bJ/WA3tiMuNtgtn0SAhf/K4
ZFIpWMsq0+EKCiq6cNAygr7RVI2urPDD+NJhnuCqX532wrid2hI2OqQDhc2RPOusyQO93DvHeJIZ
a+CXZ4++GXAnRpl3cyccXv4Nd2n3lbHERHl3S87RHieOxXE1YYp7KQb9ORa4EpsMBxnS3YD+32O2
CSG0vizqeiH+cW6ET2+aYF2GHUVTzdmVVWXfwI5k5QYRXf0S+lIfVITZ/WQJZi9rzfgP9c5Yxihx
CwxwnQgz3BEAChkfIdHUOus7DMo39neTO4HVLM0xLACVTh4Z/7ynY2ltRaz52hUlzR/kpduDy/8Y
i5bzVLKpotKyGTz68LgCIZ4qPLHxmErlct4UUsTW7pyAoJxuJtkhieNPUbTSl9nUnXDzcPp3R58E
Xyvm2FdSgbmnsn/oxg1nKAVusc46OFBMy1y99TzsJMU+c1eFSH4U1u1CZR8Ez38Fhq1DdDXV1W3q
DYHVzWjh9YhrN2NqOW0ch5xPyZjUmMfet9+s8FPPYnvkdcsHOn5ryStBNMmOlsNCXCF1VyVN52re
C2cWIM7J/qqfG39JLyQoQDeE6/vnNhgP2CUIQEjG0wG8ot3U++/twXLkF8s+onLfgKouQpVogNm1
21zzRiYeeclZZe8GycO4jesf6K6KycdEZBCDsj0cCylnwiE3HK//3uFJ2u6QHVP6leu5bzJ5qDLr
FAIhGsUrn92Ex729lU9q3D98Zn5M1IUtZlQ5sAhQH1eAvhewp11e5YzOleC1TAWPTvzsj/wDbCil
Ol1YaIFzomnEVchh5amooWmrzOZXneuC6jeeYy3bh5FLFUVx35TIELWbCTmhLld/Iq5VvYeZ3BHK
qZFKpkrtv61xtj/NO8FFbd+1tmaj4OTSMVfCQHMGcy4syGN2uYhdbN2aRAzrTmSPEKRIBU1aGfUt
KBLaJ6KIWCDV11uPRdyzRRgNP4ilA95zxoyWN/BpeAvl9AS9uI0q1FB4E2Zl4rxPWo54AVfqIGin
aZwct2i+6lMgR90/k2YgyLjQjbRt/bLrHKdhkBfYB0YZY2KS+qZ5WGX/8TpYljtpA5kjp7XQIKwO
4RYXh2AxXRBiU37RahAmQ87q2/aSZJrJgdnU7K0kHXxiq4ev2PgEPu2Pl5O710UPYzgtS1iICxwg
Tf8SgcUq5kCbWB5JfhJ3Gr5t6vodUqS+8OmNou6XhU1cdaSoGwi1BPpR2o1Us2cUAwA2fCGuhVgF
+Z/k697UR5ThXyzxrD2AnRyAyL9HZx9H0T3DEJNphMwyN1odAIN9JPavXM9W5DEd1SuPnrbuFSfM
/sR62EtxFG1fj8OXHvpvSTY8o21Sk93FQmh11xw6F9a4ui3eJAN6nprinfFyOxVdqSEAH8n/jN5+
Y5Gsnh5DK/SnxpxGMeqQx8PK4m7/VOTCLAsPV/uaNalPxTH8/SXyAksHbGZ3R8GvAMYAh1N7CTgl
PNC/9FyLasFnwHFFaHAFt79orgUajwKo+ApiAnUgyOC5mbC01R1p3jBoahYL7ymHju7svbUtfYmc
WHnVgg+aL1LWqHY88e6EV27z5XL69+BRli6Z+lQaiiCIhysgwR5AWkDpjtlsQiBh0SGV50xfuZ8L
Wv7yI+ImakreDUbfvJG9OlPWgDw3HYQaIJ6JrjXWIy3odbmMccIXixoy3PtNR+CKIgw/wo5ZKJP3
iG1p6c4mjHbMSUm34AzVjfwxWOCasNnNrXp1fUzhUu7u34WFFa8uNZVnbzXxBnP+5IAeTa/yI7PF
YTl8yKYL7bIlXOQk80u5sgKnp1FfzmFFyW+czgwrofh4nnqmd0hyA7HXxX2zSg6DQBYINDkSVU61
iJ+Si0JSwVCSZzHyO1+sY1Dol5QeqmdFRVzyoqRtiW5qPA+diMTmRzFzd+znOXgQWsIzbR8JQOap
JsSiPyRI1Sy5DMSh5YMem3bLjmeN18X7bjuZ05qlgcKemhU0MEa1k9BwzMOrubgZKT9RtPHbXaXv
6Y1kA63T5M1OgIPtkBYeJcBkYfNCqyLXYko4XaC04xl3tcU439WguIG3WRdflBu3tZb90uuV5kSr
F5xPAbs25pQmOUGpoKtm7fWlOoboJKpPVrL1KVS/6e/zdJKKcrgIugdhMoFLqxab76yB61JmsO3n
Tgkd7ofL5AVSfwU9wfOTudkZ1rD+ffwcs4Oyp4WFctPrE35JfXXxFSN8ySC3mIic7H4rhYNLb41B
mUrA/bTNcDqWH0T7tPMp4omQgmPHgx0Y8bOPghVDpmhq+/XoVBOenCpR2TlNcgMvpmHVxdnULM1Z
qQ8aSdgERzypIKbUYYmRJ7K3yAV7EyETM9XDJu2Jo8maixjcaLZ+Axwf7dVsCFGB4pcI8Z1fvveI
r1bytD68TB4pHLwa+EL2pI+AtUetLCyzhaM7LFx5TkRAY88oc1tVrEAwq0CE1mjFM+Ay+AICu9uG
tDwi0mRlpFNjdNHCBYcZPLiOS3Up+FyCZN2V0FX/SpiAzlz2/ysNGCzS4C5NLvSgek+/y+GqJIED
gdatz/0YCFX+lIUDZrvc4cDwN1/fEStq9MZHf2eaOreBputsElDIG824WjSfeMx0EelQKx6Po7wq
2iGiNfpdYJx2Am5sl8rJEdF/SY17LtT346+bwNFOOAaWX3ejG6ZcLlXnSB5ngWxrz3jaoBB7ibKz
NLrcF8KfU4/ZZrwBi837ycsEWB8kEAc3GoCq0PPmFlT5vChZJBAKF1kDAi5qsZKX4U8qA/4iTpbN
rjVaK5DR6Q4rbwMAZugcP7Z4Ni9UDKIYigqvP1vSjE7HUolkPLdKx4HDgvv1EzquLsu6aYOpPVC3
7K9OS7AFHs3SV+gD6E03mv2OCbs+QLmV4Mv33MoGQMClRxmIQeqmhUSvM+FryEqhCBwCtf4npo99
AE8/7bj+dlqT+pLu05pAz95nBCgc698a96nisGWi1U6WnOn/n7CkMxxcrg7ZtCMVku37iy6/1roq
PfaNDPJhmST6o4CRLrrgQo6pIWTeHPa5/ybv0oZk9yJbqnD/aNz+l+6OcJu2sW6H62NKh3eiHWHJ
PREvkqxouGSBSGBqALK7L4RO3FJoet8zkjBjBNSP62gtizQd6zCmwSqVVtJc5AmAtoDFsSHvknvy
HErob8mvjLSNSQYbqN11QFDUHfUFKYlanWQ2+PWHFAS6dFOOZHA3WuDooCJFgYmkfyXRwq5LTVAD
2pmWwhIm25LfYFiBYdIbY+qEjXCE+BLHo1ovB/5t7LMkHWwgBPNn+9SYMN6xlHgH+zss8Xf+buj0
8Uclmh0D7Idzfgz1Iv2SlTJ48ZEtze4So2FZoqgz7/cC2ZGP1rRspOCs6+we9LnPXxVKYPw68WbA
1YhhmYxP/b4RWJm57HCmK5vXJR10u0kYNzijedMI/445BHzN3GArDb6Ot67hvPc4L2RAa0j50p25
X1ZpvMd2vPLJ2mTxDuAnfojEfFXBE2bWRs+N0DZjLll2LG5wVeGCxm2JF3eXe6GIB4GpGbIfpqsG
EcuXlH89A2fhGISsVp+t0xgJ5h7iFdENe+fG9r0mY19JORdpOoS32TbKvwLEn1hw6c5FH5YD52dp
XchNz2zKiZ1E2WzXzg91YtXkF6tgSTZm3WMkIHtbEgG1ztCD8FtNhkAztD/AooNXJbx55hpILO+I
A2+/GlpzGf8ONACdfd+IuUtm4b0NmdVe++xwXtzmgn7grEYWM7B4tksm8vxIuqF/wp9OC+7ZNCAz
azZ98LeIGrVSFWLqOCFPyJpayTFA+6ObqzZcrzMWstAY+Hf/sJ0Hyu/jnDqCXToX+JMzFjcDwnJU
jNroxyaCDZ7JDv2C+YRxdMhdjUVfldoI0rVrjjYUNhk07glCyOJ/0xPtLFqLuEJSRrM1gGWQ799r
wLKlIfjWaIYwyfSW44B8wD/TZ3YphHVGOQYNsoJsVUv32Gu3KxOIps6pMD0aI1wH55mnvht+QW9A
mblh/gy+hDROiQNkDIq9VPxh1ZZNNv5u/IMNjn/1D/5fLJjxU7kPW+mTldpfMBDGiZdgrNhigjKf
nBoefhbdLdg4yYe4RvEMZLpWnH3l9s8/dtBJVD4JmTszUCRg6K2CqqJAPp1ELcCDRudms5WV0lQx
RmPg5+KAy76WeQLBuqzATceELi4Z2BRszPC/xyaEre2HqZAvMFb0MhXHkObUGuYY8m8t3sTBHTBK
ZPPLwbUnPLG2sZgg4DC1MHiY6glFXbYvwtTntnrlX02EpKjj6UfEw0pKad//04KEX1koqsx9zp5o
4pCkvVQBoqajFA76zXLdsIyWrfWDAn6UElpw1BqQcpQ/mGZbf4MC4qViX4t+Kor3AriFaooUspuN
8rtOv6FxVTwMoYN3f43cWnXvdFtLleHHU86XcOfzjZXwsYV11HAeX6m+BdVw1lKQRglMnejMQz9c
QLotpsgVRhU65tduCRIcf+x0FrB7u6gqYSxVMtfK6QmZ8SqzZTe4YCEstH5axOAXLMUC6ccXDRzr
irVh8NBnLOgQsr3QZB3zvGc+3W56TZ1zStkdu02/hVAmVvjztDTDM9tAz3SuSeo+AcPRrzaLcoV0
iKonp7Rs9yyt1G/zPWP+2EUvZsqQH7wF0NoTuhC2XaEVruigN88icbZbkubud9NN8b9xB+haWu+F
AfEQcYGBLT/pwPAbDSdvaM60zpUZGnw3dFhcW3w5f175F0PAwXdyi3xXPi0vY3OiUQA76nSAPZCi
ebZCElFT3XVxodQXQsE6GZLi/iAqZ3kpNy2kAzKrnz4lUPi1oQdh0V2JhMjC1IyCgqmtduWdCv/M
F8SxGknDpjsZjexFDa8w7R2nqfsbrwVcp3NB7m2OJiq3i0vNZXQPqhMwqsJ7ntNXDSp2iTFxe85r
l//PLJnYVU6Fw+WF+v+R3As/Q2Ht6vmRUokja3+6CzcT43EyE89dkb2KVl++T662Pg3PGB5Y+U1x
x4OtPjf33aeau98blHY9SbxHIWEaxyBuI0/o3GtNbG7JsshMSNjp8RhPbdnRi6PKk6aDhYCLUVOw
CA6+bAjel/0UmjfddCKsqtSvk6Xf5SSMRp5KoRnRke93PBBknWfmniYlzBk1lAilHsanNiIorNw4
c94VxCK+A+AnLkv88sci7SKDdjzhWHSYhHJN8RgiCdKBzxthAdsTRXWEy+NI9qZGU4pxF0qbyAdB
P04jGab/mCRs2NkaO1md485gV/2rgTwMgCxByB4Xg1AJz1Bi7pVF57KGWLRe+bhdaa0XWWITYLIg
4zoue/fMRTxs1U7A2MRF3/mcEHXLBksfpySVHkxMuTa3s1pvih5HkDkPwZ7/qsZbRavIVMjaz4mt
k3UUe/9fGZa9lnJDgV5qPL2p37KdX4++7wmnFVULLeGeivVZamHc+rjcYSZBOmdN1b4jSivlaFoX
Nv8+ELmYYF69fUkFwDGFtix8uDJoYRXnWF6AKLKZ7oqcA44KXQteEg8eYBH3K0r2F+klp5Owi5v/
V1E1DCzuMQp4CdG0ANEluJ4Y7PsR8VqF6N115SvAaRfblLu2KuUxM1jq0BkGsegmYpfcruPrGdvL
FhzZTh1P5uLTfVdsic/RiT/Kg3aem4cKCsHMrPcu2oGE7Z5/QmMMCs310z/CoUpn6g9pzeDHgHh7
2F3tvjx9lSY2jih01xH761atxYw0mY5h6/q2NHpS3MNBKbRosK4UUi8ZTkaW0jkLB8RWjSSZRoyB
ojhKTm/wU/Z8L1Pudq14upb4hdanRy5nq2YmpgzjguM7k4mCEWAMiS6H3YLe/cJA9vwYgQXmpQeR
kZi2M/xJRTbSjKM632IPL21Z5FRLRUvumlWmm0o/rTdP1K6K03aWV6Mq0Tub9EWmVrG7lVAI2AwY
uHuKfOs+T4QKshxS5StLOLAXuLiT+Yyxaj7EDB3ENqWv9Dbl0xM0y7TVC5dlKiJTCWdBZrJ9L0ns
AmwUZiqejIK0DmwWBr3LGLV/ymZy565RAzBabKbNU0kYV3PubUhGthzcHH6iMFvvHakSBOXhD5Qs
Gnh9I61IdaEQsgNyBS05hjMNfUvkzWj9Amxqqh0R5aOjy9KpOdGoJnAenZOB12RwK90dqqwFYsJA
09PwdyFadUoPm/XcRqODT5PjsX75pebJB0GwkMzrrO5ToNuZnZT4uYlhjD7vlOcPhlt6RufkXKA2
2jKHsu3mM2iFFGFjEnI5+Xx5B1oY/zkN/ecE+WdhqC9xzivPJ4q91Do2eg47P7a0Rg+xnwPH5TYj
faQYeIg/EOIolJm1Ib8bdSp8StrGIf4juIkP1JYBAzgcg1nUx3VHO1oJW2rraR8UsP5j/uh1LJ8X
3IzXldE7UGlyFt929gLSivUgrWtu2mHYCHhhhQaQX+RIIc3dpeILAJeNcBFqGnyNjua9S3KhGW3A
a2vt1inIQC2Rk6mF1bLaHM5HJImb55uihixZdGSM3WUKvuqLamIKBiyuXhLJwqwEtR7aWMHDaozM
q9Sey7YQ1/lsUNHG3o7dl/439k1jYJ6G5WLAdACvyDC60TcprrXM+HGw1tCCrAZ5G3r6OwyWYlVR
5+HWRhFvGtt5Oey36WcKE07noEuc8vyKPY1L7VLmMGtiainu7PQk1QFS3+77NMT12Zt43bzBbWwd
3z+3FchXvy0ezxbGi4dbST0/ozBKNNsT/iVck2dSHHizCsbgELEABMtIgFw8SE3JHPnC/qTKHGN6
cZVwHMxTiyf12Z7dnMX+/4MavileJFy2TsaPedCMNw34XWcYHiah7rmIlydiOuWQ1AbjYb9vrBN+
fNVx8qK+6jNPcBDZcb7lukm08z0OV8yDxXB421wrxBlu50/5ov2h4lzXceUvFYOMHlZ+YL5Jkicm
2xbwisLYC+zQWjbZ2k0xQ5sr2427L+7or/Zt4+DNKxqDu+413AmIhoHaPxhdr39ubSIq2bgHfHsN
z/Su0CRWC1T/len8faWzqcq7JNSnYnqJa8RQC3qvZC8Hgl3x4+vIZFQAOPj++OhulrC9+CqUW98X
zGp+tiSse5x7p68hUUewuZG40kapc0j7pbWpFy8gsBAnZ7JFbH/c3K9bnvXbvVmdbkQKQt6/g/4e
YT1tFHDJ73ckkAxCdXPNaLrOlmxlAxZbVk7pJZ1+Y/2GP6jAwOJgE44yQzB6YeDv45I2xJK5MGoF
F4ogM11Uup3HX0cajKwgg3RsG49WedSXbmhI/RUmu7rYypD7e8zZAST5cSWjUW8gPN8fwFySxOgv
s7PkfRw0ijm09t8UVOwZ09t60YhZsQdM+wHVPaU0WcntUL2jTgI9TZdGRXe/k83Mj6DCSyJyi+Tc
7MzreQfISqjsitJSqMDYc42hLBFF+ZM+zuBm0zbwQhqpE9zqxmzb5yM1k7ed84QMf3plqBcySps9
laEskt+o+BrUOIyauGaATyJB+xpxc5aLHgoVKWpd1QHJtlJK3Yva6HFK84Mxr0i1WhyCl0oJ6NZP
Gy69LLJ/kCAaeIg1Rf+bMV6w9wqPAzQeugs2vEO6+6HARz6K+rmWH4+GIcbQqYlI+IgJa2Oeytqm
8pMBlqUUoHSAnEUKgnyZPJm2z7eLm0J6O+DSoTQfPzIUKEdHh2bmDeAXT0aiIYL/Ia87YmB8bTtz
4Q9ZViqejRirmTUFmJoordqdDDZrAqHmXt1NZIbFW88FHEUefl/jwj/HmF3/sTWBVLCI48Nf0aEp
WUZBkm0hngLYJpt6JMJ60ddCQKmOtyRjUPd6BtunkH51u9oaXnS2jMKf/m8fVVRO058e8xCUPggD
WMz9uYZffzxyy4tJfJ87CjUIWInPM9076OhcCvZKO4Uwy/dvLqzTnWNGETke2WGL5QJmaQOXItHc
bSA8vC1pYEDpkbtjU9Ve0X1Kr/svrm+EVCzTTcYCjU2H7EirkTkQUcHD4gMsJ7WI80pDKjeNv+b+
Tk9R9PhaDL3+Ju/GC24u0L69vR8/BNTkdRQujn8Ir6wt1uYRKC1hlxv+z8KnFlI8m+vVuMkM2nIC
8dAyGWjdNf4zcoOXiO9IwXUsIjvlXrlJEgL2OBuoznILaIcy6EBRWLTCqYdZfTigzydWxkUZuFNu
mQV6+llucfFia4KyYseKLgcpat1AEs/H17IQax7GNVwR0z3SHyqmlJX74oEa7g12jJ1FnUYhQ82e
SAvptgIBA/CMU28XfTtvc33dKirdxcMLsAxlZttVQjMyuhh3VzZu7hrSvoUpTPvhVGxOrm6buJY3
60l7FthTTTp7qWSqQo2qq4C/ywDYjXcMbejIwrJ616Nb08v6H7/jiB6sII3D4aIQLr51bFpCpyqS
ZyOFh6bkrJDdzTdYpyGv0uyqE9LVB0zVKFrS3n7TL/upDjMiXLCjuy2ARG1gLZ9UL4vmeKJv9QdK
HHF6EvzQmXb/q1H3/rznGMBHgIG+r36tWtru+n3vnk+8VpTIdxovNk7BrmG1mORJFPyq9uMpvZsf
kisKK4raAXmBD5d7aTtj5fUWRIlu3JTmHZVutSIKZtfyenOpuUq9SkeUEqHYSHDHyQr9iKFgEUB4
KKsMw4Fg/w+uOEGTCgX4cRxtHS1CZ9pMzX/F21IO0uPYuMGIlInqZnQLyW/uoQTJLYFe5TLgjYGf
1rN/qes/CQhIlFeOMlIvrNZMP19wR24hXFV+ueuscXNkg123MNJKbxPi7tO75jQDnI1vXHdayudZ
a4//1cGrtatzreHV2prwuNaRf5pFr4BEBW0HdYJeizB9271EcstK7C4Z85/SzvB1iJC9on9p9gLr
B4LZry2BBX8OhlwE7VFgmuHnt5bdymYwNk+Q8ZYZExrp60RmDCGK+1TOe6Ff6J4LYrfMGoqLrxzf
mLX3CjTwoT1Usj590D8suLi9qvr5yqf5gLwAfR+4cBcUVJw/WLZ6WLlzCpLWjD5uD2N9L5GTdNzA
Ob4T5ryl54H0JnqTeZTTPdY05FH5khiXf9liQZuC4jiZ8VqYBba3U+Pg1esjOokvr77v6kr1A17o
ujlahrD9GUHvFVHWIPqZQHkTJqMtXaLosdl/kGVWcKqsUjLn83JxxZuOxOIFD5yFFm50vMC7RFIY
eWRQXbcAlL/DLNbUlKmGHz1ivMi6t1BWVQMW4E0MRwBqDhRzJPJ6mZM2YISz2yui92+hbdOabDRv
SUE7BjQYUX2jKZEb42n898YfWu/K1Mp/ByTNHL9ex9RrCKjAgO1KaDrCXFnYtlqFgtrM5K+giCFH
IQGRRmq4nYrWo9JGQ1DLp93L895z9mlucB2oEX9H+MYSxFD2rt6TFFNTcSKeUdmpeUAthxq/eiFT
9jKA03e7uwDCdBYM/OYwwaTNWLaGwBF6TPhw5mNaTGPkHpMCMEMJ12ev8pOphRDHXjXqiroHVMbC
zW33iXIQxthkTNbTxCRxIRqjTC2zd9QWfryW/sACH072mw6iY0rXbXNuvnCOIxA8CGM0dP1ps4vN
nfR1BwrDSDKr4uWACOgKeC9O46dI3eVC3C+WxeB1m6pVwBfZu1DrsBfrHDBW1ZxrQgQk/LuCNjei
JVD9+fj9HeQC9d/y8I76T8A0e4O8Y4rnwnazvv/MeP5/Noi0vKe5k93sCfQb0EILgigVuaHFbFTp
S+5lRls1oz1Hv62DeZOcYwBHUUFis7EPf8yG3KQLJyZ0Tnu2mQUsD3U6K8Vr9UxkeakNgELXruye
b6rIjEvXKdibFcXeq2ptdgbFSdT7gRshvIJyg4Dnt3B6GDkPXKIy+eV6h4QRYzPs+TRsc6n1WGax
wi/wMmOxK+1wLt+DYUmgBurIxGEmhXo22Kc+iZa5nzq+cxy+3qW4DMaN4lUCd1ckZtHb+2H2ZgwG
pr0FlH0hByDYyHHWYABeEEo9V+3x48FrEnSGya1NrsOgF7u967IacVGvsW6IQDdSgmv3GHpqeeLX
LoQam3tWzW3QD27Whjix+rTPwYoaRPQRUDcbXa7KaEa9ekU6QfVdEuv8dxHYEs3OdqmF1fMm0ZvR
zJCtsHcOf4fmdc7cbMyfsXiVvZt59F1ZHUCBiObScqwZh69quhgyy+I+2TbEURYMzwwvzRtrshm/
Os0Cuip7KFruoSi3RcVsXkoi8F62YdkPJZchLT5PCDnBkxFwZs4G5qoToaN8SRTlXvo3CTiw57Xl
NNVo0HpKWJKZQ3jW548RHVmSZ8M7Aaflinf+65I9XJQkoZmFND75cAgK16a6GboS14vUjTJVoCan
MYYOScCw88ElDixn4I2BkCTz+L9hN4mhBTQbOs88L1ysazfao12jm9GdytgtRiUw1g7a9p4Za129
TYYP3BuLIzgdXjqzjXM6hpQWQKBx/j0/GiNuHREEPNoB41igA8qd3fuWtUSN7mlmnjYHv1u7rFWs
m2tpBvMjt6aXc/UE4GyOjHKUKKcbPltQZY2wCt6x/bqmB14xCaFczZUBDFBEEQjAlSa7lwmZAkBg
lL2rQ/MhzUL8F2BqdM83qzeK/JsF9P/XOxTwj6WMnrN6WW33M53t+IRZIDhXrJCfWys8rt0Q0PnC
X+HjpGM1Dj4jYQbDg1wg2bcvdsXNQVutU2mZlTgMudViECvawWUBDDDpS8eUoTAZUoEQTAkEZ8rd
l/adtkqacYFgmqiwQxPxSLIxjjQpc2mIwi9toMJXK21wAu9oXVTCOhqrvb6XO7bN62ogxvJVNpOX
Rw2DS2tuY4HGgJEbYq8RSKUukPdySg4Bxwb/o1mfV0wBUVbZEANUQgGm38dN/JcqPvZHQsudqEDg
4sp379Vv9J1C8AAo6frIm21QE0B6XL9/9JDQxanFOi7nY0npoKUwKkWITh06ol2izdUVZbuEipQf
NvoZmsftftNmaTOi44+ZMkht9DBARuixOnYnrhfGNSehSPLHI6eViu7Di0AI7+2DwzTrPl+3UUww
pjLKgfmBcNWW41Q4YRkj66Uvt0LFhf+j8GUlSNCzqbTwnoRG4eCVJIzzZOYT34t0bTYFvQliDJjm
loD5sctYWpn3XSM27WYcxEh9J9lKONpzDlTkq0KXw5syQxU5OLAIoKiGeP4NJoVG1ek+rZssUMhA
4bvNBhT4LWG9Kau/mXa5VoCTCvsljENqWp1zW+5gYeAc0n5V3F5sHWfpHzYrCrsU+r03xcuDC9An
WRZzeZLLk6dKI/LKVCf48M9/Ayt0drBSfyPIbEOxt9mL7Afstj5mi8y/hEam7TmuZMS5hCFxDeNm
NLPUcSnnXIxIdLcf+OHzOTwmPhdqd9P1YxSi8aRhQurVakByBnMeykN7BCmFUANG8utJoeqKNn5V
Ov5hmpnZwFdoTnAyfOuur95Ta3/nQO6vUO0GvUxL1E4o0oef2XsXV1bi5ZLOXP0G/HYDVKSN5cen
wGBM+d6jALgFKGaB31z3yFZRtJcos8ggZ+1/xQkGRV76ZGdPNhcvpeBVZsZBRMtd3OHOH5eooOoG
o3SvUD8o8iZ8zZwq7GLfGzgrXbnTTG3VXyG4tU4xHsao5XJ987b9HNtEYlN7koU8SJzv3KBUGjMv
xEYV6FTFfbAPkvT/pDwIdAonBkmVk4G2a85WoRY4/BC4RViebKRvPauv+YtxCoVA++K//CcNE5xJ
R65pfoaRfYFe0nikD+Lai3KT/e9Ump9jsJPJnF3/mD2oXWyuf3Y7UktQNYVT1EbuDJD+AK3i2Y+o
8k/fOrLJSUvVfhWwcsI6/5lo1Uxy7QqY66Vv9MLTwldcXqZ/ADBf3xPdrr6jv1ObyGt0GXNDD68d
STAqqdEQ2UMfdm6Z3leXd8owxqBqg2YvJgMYpm8yXm1aVU6ziVlYS1X4AA6oI7iGY6reMNrkcV6c
nQDZz2oPqJtBgsZwP4VwICjuSihsLrGYfdvNhR1/Lb4pU2+oSbeBGxe0GjP/pdMaKkGUF5V5/sIt
psEr5JA0znDHRkciDYn7wYNvQarSfvBuZAOioBPl3R3BZ5wL3cXNa37G20xCur8vywkzhN/VesY1
Lj7MGz72b4pqaED+0IPudNKaPK5HR0dhkin1nFBkisqKcfLxKFYGXSZ0AjIgGN1jIC463B0ClVsR
xl/P0qwWwo3yY7Ts5EJRierDZMtaNLIPz7sYwMadw3ugmeFNR9/rJztO8cQ9L8q4hIboRg9QKuoA
w//7kEjanlG2dRJ5kJBvB1lmHjELaqdn+zIdjFiBMtwC5Pgi9RD0Z7OIgH7HtLY3KyYUD9rSxZVm
/A8Fj9aR2/HvPKgCE4LDZL4Qt4Ecp4Sa8iv/3i8SVcpwgLOAEvrd/naJlgh6gqTDBBS4HxMVtETd
mJBLLlcUufMhbrf3dnxwHa+BcmKo/Ip4xsxOub69INqi9I2po6Dww/WfFyXYvDyHLpTJVwaah6zX
mFLDI15x8qFPRa8qLBGVwmgUpDRajVbMbi7WmdQ97Xc0ZPilVZo9XGFLdBDfWRDImwX40Bvv4CT8
b+SxukcgfNgzC4trvqWk6TrK+hREvq5f3JGLGHmxd69cW82qCLN5qxwT/yDhv0r6kD7zHz4PfiYC
ka0hvVdMBtBwJ5XPx1xsEgHQwXb9K5TQM3UD9oojt56zhFuThHZCOUpGcExmX4VDuK34eT5VNWn7
44Kq9PE8A5Sxe5zFhAX43QM9+cM7ds8RsXq2SAjmZbacs2R3CpfjT/yKfTbwrr1Y4UnZBOHEmjwL
xv9eAJQGPfCPsdIyLxb6TQz861TCJ+mwdw7WBc//OgrTF5ovvVPj6YqQHWNmgzUvrvqVA4+3DhjK
zi8xBmoR8N56M84HZyxjqOzG412h4+GHNYFvzA9Ru9o5Q8QA0MMno0PnUX8Asa2KnLGhZW8MTGO2
6tkWGKYkhFAL0S2wKizbOn6eUAu/WG9nClmcP+Q0xzEOTbJiLdP4HaoCh4spYaYHAEM5BAu6xb3q
fnEu5AV2M5fHH5Vn7gQ6GQ7v7I1IjK6uELawp4PJFXKZO1FZc58KrLWPk1lhVU7WWQXqOmAw+IIS
pXTKzB2YLWBFDQaAK2GIm+ASkEt9cv6gerVslSLwCV5TujynglKRm2X7ijWYL/6mNCznHJwM6xur
udqU+A5D72Kb/zvFPY5vVNat/0GrDK7V12lGdoNdpSUqKPztDbOVEea/KhzgiCpThvi1l4lQxVR5
T1y+Z7lvW4Yf622NSGE6b33dSJsD3Nmq9W6egBU9sLrGVgu0Z6WLzDVmbIPZYKXW9p4Nui3JvUY/
4FimI4Wuth4AiWeZM9Wa3K7nJREk9lD5HJQKuFYwyVHNIavvnKSrhSQ+KJijfGUkNnbwRAynAUBp
Wv2B9muVPLcrgNePPPiJl1PRx9Gy54DAi5/GxhyeuvI/p31AkZon/siTvLmPp3oF9azuLJX+ptVd
xkTnnc/Hj4+4jyIbhQatnq2EUU9mlr8HKAHqc0geqxRYKp3BBkKwk7QENoySi0LKonhks5PgGBzs
vkiI4HIwM2d7EgwcE4YsK7eDKzQFfGtfPJcE/A3FTtgD3hkh+ZJdaimgjbK5c6t37xNClePmIAWn
ZpPp2iYJxiRBeM+FNPAuRaqGJiKhFI6FhLtAM85dPgB7BcTa1/gdIyLg0h2d468TjKxX3n1FUrZH
0RqNK1MtnaA8DFM1UBpV9bp7yMw6UgfKV6OW2WduotCWMtSlP6VVpmbVLLakiVHGi5ZFnouBVAEC
HDwVjhXDoAeNqMeQT6hjX3H2Jd8Zqraaj8gCe73acc+lZ1EZGV70oWJKqdpapFpZXGLvluL+hX2x
WsCSKFKKkrfBX/PrUhccPMfZTJnzJjdoERoroZUX37CbBHxHKfsaTu5RlKI7uTyuLrDzCnhOn5D0
hm9W3Nvzdz6YxYgwmsh34/SHbJNpM9/7DD7Y1x/Pa6uTg+EnuaKL1+7lP98Ds0Tm+cOMvxM28L0S
SKWm4CwZP0qMzoP4m21p3YyFRAEnItWUQ0Pd7pZ8C0KyAZ9aK4xqIN0AnqS4IPva2Dp3De/Wj5up
Yfk0/qGmcd3obcSvFdmP7nLdD6h0o4dqYMT3RDZipn/cIjS8g3B2hnKXy0KTstsK2mJ/6/d2DPyf
g4Yu1TusEjJdDQDQAM20PAP1CG+u0svig6/hsHgrq3DDXInhgU8B11pJj/Qs4oQ+awpQZswzd1Gh
zSUyT24w288Vz3piElZDfFJRO2onNhZ6SaObPIlO3o2DDYZEp0IK1WrZyiAVENE3jrLVvo7j5VPl
6yfLXe8KXWK205q1kiWyPNWhG141wb6aQlf3McsJtywAjYoNlA1mr2U2h0P7utuiAHqm7HpkXX6q
UZvusI2KTrma1Zv3+hOXLejmIW8Wp1r8yE9WZGDn/9GutodHQbOGZfWq/ciU0K4Hac81mIIJTRTL
dICLaeZxCCjsH+HejHNFj9TdyHwsR49mE3vSE7P+/KFhfk3A/ZqpGe3L0MHsc07AWSM6G5Ae0ALm
3GvbBoii5WGJj8RXrN1UK2FSM3HPi9xpf3ZOeQMx25L+dl+gxEZU9eqW6hWYoPO0PGTIKMNDpBWA
4b6Wua28C5Emxxbl8LTG5PjLDgjQrZo3mcGzqRBIi4osd21pZHR2kj7oDYOHL73a6UwGxTStO/ph
TNZXdccdnBzrQNQhOo4/MBpqbxLFGWYWMAwYeIVPHGzzyI4pYQ5RgT2tPtSjP+/PrHIIUxrAY3s/
Nzb3uxo08aNr5VVlAQbJ0iCX2fJ1IpqBwznvttcGrwu9pEWdIG+GPiJjsnm+vx+HhPk0wlld5vUZ
T+IXlWKkUc5f2zk/m06JrFBHLz9mvaHfcw9DtROlGOew3hCQSDCSZCVCfZrg8xAsMFS/jYaI+n7T
MP06o3o8ZPvHkRjFCT99Tj8lNWP/6m3IF497rCZQb29PyeKLzshAVY/490cAQpa5kEaHDZM14uHy
LVB9lDmCoLwzLaEapzjE1iX9OXbEjoDRD9iskCCERGTkYj4KdMS+IXjGlLOyCA8vnrcRjCPAPkEd
TDD0DpGd/v9tPKVDnDORMuI2uvRYpp+lbXWXM9miPdElzlqkzLKtztSTk46eQ2oWHP5gT4oDJBJv
Qe0ffZfPJ9OJdL+8ornySwVwDgPliFCk9BF3luH7SojS961f2tAalTI+TJuRdfbonomC7Y9WfNgP
niVnbDczON4/1jC6WhJpqCBM++aF70IszWOqwJaHsWYC9TI2+xgzEhAQK4h4V7HY4kufuPxUtAS0
uTDAoQ+sgqnhhALC+eTRuy6wrH3dWFsvhOtMDwissGTqv+TiGwx9i9c3UiFmNmUaWQGenzPbs0wA
TcnEwnGYnCivAp7JJMi3yKTzUus633jQWVXobqCQm6r2QV5BYG/nsoxmWiAtVnCpQlwxeS8XA5e9
1W3wjQRef5hKGRxLeapgTIWL6bYxXd4EL75X7scsMibhES9yykReQ2zj9EWUvoEC3pK/tJXymmvg
RoTdIoG70Ig0ESDDrIMvd3QiGa8aoR41tTsIcApfmXlGTIFyZ1rH1XKjO1cV9HIV3U6E/wBKFhI7
GcDKSvkOxsPOTazEUlgoMMf9pxg6PT+9LLr38RzuoS0tLANFRg7qwAs/Z0OiUXDntVzjXrEJI3Tx
G4xp4W85smB3g1yHDw4fP7PBydndG3anfvr9rvdOmDlGZyde8pkad11ndUYq4BpXDOvCe/q2Agr2
9eMngGevtSRqx8zFw9+6gahRPyIQklX4Q/amGlmgmjR5ShfTSKIhFmng7+eMB3EHKlP/JZw9h/rn
U1zMYKkIMepuEwEvhLhy/T/wc+TNOnEcVut82ZSgCqSUiv5EFxWjv7zj0mZJvhO+qvK1YcnwjLJK
5L+jC4vqewTw08R+sIOMVKALI7n/Vxd+z59HgXEC6ITHoK90vQ50zWXJV8BPkFQpMbADnEOm3Jp9
oReIS21hel/QvjBbEEzPCpMJs8BBiaj9OeeyKF2I4wG4llcWJ8n/R8HDNntoO9QZX3UxmscsL92z
qaZjg8EH0tLll2pF9SHgXuMgN+hYthfOqNw9Br9EMn7r0KFGGJDSGaUsCTDBUTxnwD3c+A51tQzu
+fheNpuxooLJuAxJd2s/RTajreNlWZvOVJyCWEfEOHauTyQHy3BUR6DldvhjgodclrIL7AIDDLJu
n7vQqMui6wy5GZxGfjuSGsDSQR/3t5Vmq9NWoJ66Puw0K6e0mXrucbjtxcl5qsCZKvvaX8upaTXG
eqlgHR0RtCeNhYkcoUEqqTKKrdu7vl1crEO8nlRNmZoP9YiSuYmpe+0BLZLLRnlot623N5lmXDN1
lRjDR2JH54oJO/fZotoi5tEzf3xNTkysK/C4bn69la3ugVS9E6aMdTH5nhj0v8uhrnUodzfB30dW
1GnDOvdSH0EKM3fCns5vTBYK362kAV0KYRnmIy5jz44vJTm/11wGUIV1v3R/Oh9EGnYsmqYqU8T6
9pBnkuZ04ef2JYDc3XiV4XzDXggVyDPScy9EU+YVdKB3Y1mEhegvA4nhLQFxDlKekXq+74l0XjNA
b5S4ZxNVfe/3jktumVjIcdiGPXtoqjTv2jx8UbdWfBxNoNfZIeqvmJNChB1JG4QN/gYdXVmLbKJD
sNUp9F67R42m7uWmk3AZ16jutlcZsw66k4MOVCJLumga4m9LrYyYr7PovZMyVG3qBdFMjq/SxiHy
eoZjdseCowylRKbJiTlUvAgrPpaWEZnvUfNwRG0iN9TDWDeewr/Wmz9MuqH0WUXMuFOTF7J8ass7
ym52HmrYdn13+CTc1124yBLMG6WH/0rpHBdtnsbEYRmiWRuP26nphXiY1g8FgskilhAdnUQEv6PN
/rvU/Ya90QmuE6EsCbaXPWNev4VEryxmDzOvtG0B0O+yy+OIp3/GqMI76uATwXMhWlFq8XKtSWDn
8sMbjadmMA9V9JeLYoF0CswEP9Gog2yVVmDf5686Gf74fvsuFYmpFgTycKftKJrgeRfgEAJqPFI6
Pca/Zwho2MoEy83PKOhwwh6708pOv5d91ySoSZIrHuhkCt+hv7idL4dPRcSRLJtz39l7t+cCOXxt
I3bdmd5uSnN86yuMdz8pfykFiZUdYQd1y6ENpsctwIby4IX9QDfurSuWxBWGkmDMWfErJYiifC5m
jPixn00SHHfHH5t23zRwC1Uq/J9e8aKj0gm77C9sM4/DF+G5xLk5xScJT1lMHT14U8oXWD/dEcu8
2AW+XZVEHq/ZYThcgPEhJAL/VO7aIuuDXsuGB4MD2T5DZ26eTfPvMk6By1a7aeTCL1Jd+w3Mympz
SjL436mFOMeuB+G0I36BqXulSC837hxoZAuBw8JoqtnOTqGJCaIsbVyHZ2GsOlDg6JbZ6y1QSY1V
mddKedjW+b/BqwCkSlgUHbVvi1+7PU4x3HZy++uM8Eq+vAI2Qmbz7D0yiMuKW5M3ptSHDoyeN23t
U3DvPCtsm4ZjJ6z7Nwd5rEFYrE3SOfn0s8H+2DFKdeMLZgQJvxm3C/2oIi42K52fiLr1NcPa9OhC
PQkjo88hI5BKUVWTBWYAEJaQAZvndySgbxqlmthtMSOz2DMJHUfrAKax7FJTZ/xrnM57N+ZpB+T0
Kbnr3sC6/p2zNpKNMWibuHNJsWAb7eL8P7kSXiXvdJQ1eJ+e6+GDD+qWbl3/CJvSCEw7exkaa+Sc
f3kjodhyC9JNIRvk7Qm06L2M+kBdYwoJ/qhxA9dsv+dlcxyF7vbconNv0kr0hfpyBfY7hRGJewUB
fNjC4fQ63bA3UJ4tisukqB0MxtY/BpHLSIaXdEw6Yx4E743RI+SBcRg81khOa6TJCdx7r1NVnNE4
TjqniMEhIaTQAepTqogGna0HMbtNuEUtt+hm12ysXzzE+OTmy7Tbfvv/RgHOYvcWbZgKLX8y4j3i
CYcgxB/0Z7RTa82J8uTkC88jGD6Ps2U3caYlW9HD9hb37yU7bw+GsW52yj1cTnEBbn+V/KkJe1hD
cynCZSK5eY2DGy7uJVsz/cexiZ8gwmLbBxtthJS97TwhBIWEbEal0W1SWSW69kMKWe9JIy+7feva
EILsz1XcHrp6uMr1oUcXFKpJC9Ue9k+M4jnAGDwkhpghu+JqvgoEIf6fVifEssLHb+1qXPxE6QmX
pvoY04njjqJpMRNslImxYzG2VULMUbx312/LA0M1GYbwPLkxAO2NoQOcmLjOlFt60HdVN2WGPPrZ
VqHh8rKlbLXXVK/BKMYKWlu6K+CvuslM1bKU30feQkB3pzjJ3M4SKQEJhJE3YCr+qx2yJnonljTH
cCtYdnXd12QEHZCzDX7GvLh9RKGUaQAjUgc/CXt+i/6b2wbIqabgmwXlemDsrmyMYvpL1tomcizf
PwxRDkmtTmiaxRlTAQ6DybJfWrdVl5016KcXX7Lf//ejWbZGV2oXDkqAlCgXg7YM32HTuhyZ1Eiv
M8svbWV60lBEc9AFXvA+ctXRnSrH55CSAvyzaCuEycKwtFdYeh8JHf6wr+i3uPEboXhSW1gtIbux
UjP+Y0oeCi0bVp2vIX8mV6kcSjIa43clGZfhpU5gZkTrlxBJBRdnIQk8DJJQNS4r2DjZtyPby47I
vxE8sAM54FKcY9qFBm+x7WzLoWhqPkG1rs3AhyiJcOSbvJSf2+YhBIo/uY13Ur+R5p5v3tpK1zVy
IIheaJztt6SpDlGZKn5M2pLiJw3x2Ah+HaqLYA0fMqYKUdp8SypD4M32x9okMTNXqTvaxGdAfi1i
/h05XS1XrOTgnlhfG0ZcZg6cxEqZYNR3qx/r9uu3FKusGwohNl+7YHjgOsF5mYcwzlm+7nZ2SvjG
tcdDWtxDUaifXW2h11WFSUT/+GMSETrp3sYPRIGCB4gLmtKRM2XyNFcmqDMLKAmYGDMEQ1gW8nxm
96Am10O0w77+0wgkqVgGtvV3i0214R0HX5/00LBQDHECFNhbSm4BjcfNj2fClEUg2oxYQYunpFrR
mURYsZDzw7raX8T1+JCIR1kldAQcKm+1ip3IU4PpGvcgMSPZ6hmYoamlZrMKN+uRcNXKFZtTSvQW
v5YkVAp1YMQiIIqllWuxj3B1ZBLeYR8NkiPTeFbF+5hsbnuIJjL8lczg4cXotnyT4SHaHu/oGMA6
7AGgPKiN0CWfLCyDoE8y3KYAoZPZkCC2TNdJseNT5x682d97OncDIG2nFq7BXxRTniNFWPHhKmiN
N6B5LRqkT8mf/wp3Hmt+zQzlDSttAIZCuOZzMgWHeo8/0hBXEuZYLrq66DocnFbQTMzteprT3YGr
39SX4LL6o58daKLM9WYB3ObYXuczRiblpWWmDxLBdr6wEvbsrdDugiBTU5zJHrTopC6grq+mJPrr
cMPXlkD+qVbTzIvXWKEWL5k1p6eilxdD7h3Ltqr5bQ37W9eCx5qtyvKTKJna/LmtZVS37O7FqKp/
r/zV+BXujODa+fD3sHxghGnDUU5xwqcB9z8UxhXoHZFVCJXp9Dg0zS28Nqx8hVDsu/bW5yfVp5se
mNctOeArbiEA0pyM02u64cjxIGLkWFbuPqeBCJIe41gAXr4uG47cCub3tOobkPB/UUikSHJ4jFCb
+bZkBowijFlQGgNEZ/+3kAuf8CkYaWVzmsl8hPK4Ow+yAhjHK6CM9pJ91H7pZkkKC64meYVAhZWa
igKW3r5zd0Wopsn4bOj+IHMY2s1Y/HBsVE7iixFVHieWdVvzoc3fMX/JZIh2x9FEdyAANXQspqeu
eLAsgmrG70vBzb+KTrUlTCuRBZojEWKP45CHO9f5EwMAjlEEANJ+ggQSMQL6PMMJh94WY1xV4aNp
IEKn1M4wCYQ2XWrfGg4BDHaR37bDY4QBEGmm4TUoAmT7XzLXqrXlhMd695SKAHDJpoi2GznU3T/x
prdBlgsdltzOyLnfGfTYP4bA6U8xNLE8FT49+k3hh3/QYfNtgOGJ4JVSEqKRK1oxT3Cqpfnhy8va
tlquMcvzWzIT9ucIPSk9khzAa33+nwyNG8qI7rO8+yd0OLw1kzjx2HmCHzd8DZ3G7O7wPvsYY5Kj
HBqhk4dBTA/Tk3uw2djpnk0ThBtUNzld4y6BLRwsMiu7dzhbRITVsDwss3Vg84NCkGWSO/4j8+8f
aBMeOwI7yEoQsytKHs9/Dy9PHSLSalWMC4d3OpIyCTZAlpzocFwu4p4WJIM3yfjTn1O8vwUEcXbE
VtbimISCvSI7b+B3cvZOslQxvCkW6vUtPnTvomwFo8QVdnxsWN035GDli02Y6f8E4+cFKqCCdExR
MTquyp4cW1ddI7Bm2Q9EMxq+pxwjZvpMnZoJ5QXYORTCrgmLfTNiVLaj0MkTcL88vSY9i1u+BFlk
cJrssghHmbjJztQlI7pQJEzNDIrFrUwc7V9aP2KM0+pN9kbENRWQQtM75h3L1qU0nCex2j24KAbE
15Ua/g2n6iwVEzp+CDh6Gd0E6P5LfrM6viu7Hx+l5wYnstGh5Ep+aoHi11xvVRcdLOtz8THPpdiw
WkiQztrkf5EUVy+Gtv3fX+ByzJi9f+2RavZEIVJ+7WKgp6u21NznrQu8JbiD0HPfgQ3Uft2LO4vz
64uS2GXQ11T5uIwwg3WmmnqrtIL6gPYgVZkka0BESZxLF/589DRhHbDIKgZDXhBKMlaV9rln0R7e
QRxpXN4wgs74dVo1GMuNSeEPrhbiZ6iqggoFJ4yFgxwlnaLZ3aBmH6RMZEBq7oLJmEvmhZCpk/2T
soq+TyDrz5l1hYe6Xk0lToYc9MAl8JFkGo0KQsq/r6yx2fAlGKzx2wtB+VfLryovB9AUS5ASrWtU
nkxcknpgxo44ZTSmHAfhw955RIIijb/GBwu1NPKuJwZ/V7I0H+Ve3SG4FNZUMxijUBhQhKrpqGDI
TfqFMjG8EtWtL6IAXXK7C+i8dL5pxXiXWuTVp2MXEYGIAgA55akdNsLkM36u47qWJX50fW162nu3
52xv/Yp05mMWMKyqthLoZXfxSLyf1IE8werJ362XUgFn4xeDj/JXYvkMaEywacQQwMgyGcX3vf/z
R4N4/yotu0yBdUAMYb4jaX0XstpD+az2CrGQrA3H9Fabyc6v3kL7IDm5RoZ0ix8rV1pv4fgDOBRs
PgVpjXjkIEjl0v8irXUq6LxXmJ4r1pURlZqwMamsroCswOKoeHpUreadEwo1XXcq3WtmdT2hlYiw
ml86uOwbjhdtm/z5sN9DSRIM/oNQznDTL+NaAMbsGwUSWhkyffeV2cF/ihAPx8ULU8ChWTk/owS5
FX6AZFClTAzSfeAbJsN1OIDv73qZikXP/2e0fUckiot05DEMB+j+P/hszSRQQHE2M4eNCtwW5bXU
/shNhmw+AVIYiMifSX6Zng5keUGNHprYHjlwfUZ6ZFUvUT+QZ/b3cQiGXiH31//B5WFAq0q/4PeS
C2iTfaajCMpzcm3zSKa/4PZ0yiyq0FPNItfqCSre/bNAENIiAK7JCoOSJp9NWJOc0TwJSOkWMd6o
1dw1urq42c5O5pywq3Mn42GpesRx45XhxL4vUboPVz3VlHFpm3EwgYhI0M0cK/Sph8JVXgRKxuQ9
RcskrSFjpI5BokAy7ilpUWsOjXDImEmj4WVBluEtjiXD3CYG7wgf1xa43wFa+MMnJO/1SYm3pGTo
UMemVT+0oIobq2wsFz4HTxxXOCzrdxaFiecR1meCJR+aMBEEDSD/lhMSgJ2HFylZJ7OFxlIXp+G+
CsG0C/4DGADZ/38CjPjFtrPEYg1Id8t75BG790eTYtUnPbkUlUJpt8x9DrUfNGaYpH8jtzJGKNk7
FGx6Rp3C/BpUF5DkQGkBzswwCWyaOH7MwP3R8weBeZ9sYAcQnOEHXh9JfeiSn6Ulyd6HyQNhmrPg
mwNRyrM8fWCkgBucEay0FYRngGw20dj/usIA8DgL9a3miAIF8/0uFrWxfVds1Z4uQmo8YYWseUEq
PmYz8cfR7OkTzAtbzMOtcHqGyYMw2Cpgc/kFmc3mjKkiRV6BU/INLJbjwa3XOv2QlG3Sg9Bgeuyy
3NUdJqDuxwWvnnwlPJmSULJlvdpRtI5RPEl6ynyikoBM+QjXXUrzqKVgtGvyN7jEyC5JSz89spk9
7yJUypQZHPhXHw1KhpbEr0nPW3LWvmNB+UpUwj+vD0GSS1HvSm078mnMEV4sdydLZ5QuIbahcCKf
bFtay7F9JuEkUZV4ilBpv0sBDtmADxixbIeW+2KPJSAcsI9OOKox3URNgJ40x0k+jg3k1dFzokeu
Zn3aPh6ST4NRYLerxka27FdFavbEd0wlAggWfJ6XZvi8SQZKFYAw0HqVHU3gGwV0Nh82DHnp4mJF
G2HjQbkq8+HpFc3lUf41077Jh/WIhWGXBmHN25HnPIvC24YN/f3oxfmUy5Y7YdjO+aDlb8Hh0lhz
j68vr6eVvSScppIURbs7OxiuRwzMZ/V3C2Fuq/fcKaEaua1W4wXOEEs1jbfrmElS8lXtCoDqIYUp
07p/1hqCTbQB05mMrti+/qL+Ww6Ty5bYN2aVYrIOqvq/avYFf9lp4dRqfOiS3VtSpE7PYUNOMkRk
Jq6pAUg4/VSA7B0SHG1beoRSK9p4CrYa+PbyasCdVjK/zS/Bbqo9D6KA/IWhRlkUvhjFrji8r/lk
17uPFHhYE6B4U1GBDn6bg37xNQ8KNHFmyK1XwLng2vjMNjHMfodgmdMvvRUV4StCpSeqOiZRcc47
3C7HyoemPwB4c9qEWp2Pt6y/HaYxNyuCWBPmdkXrR8kGLzmsQDUEALBjNNtkbU61xxR1im85JbbJ
/uO530Gln6fDs/qlHPDmDhoK4bj0zj8qS5paYMFtm+fOgybpG3L//IYiXZP5aqgNDP5Gk7mEOvsw
pE7utC03rI1JPOigTFUnbyBomBmIEujpjwM6t7C0Cg5GKS71YHL7uKA91KM+LgtVCq+w+ZwNOkdz
ZVLX23/E+UCMSiUNfK79ugn2tTPyUIvHLHzlQDQ1z0LViY1liH+GJXTMFDQ/oHl96q4Pvroyfdr+
4hZ3DTaUDXAhDmZ+weEBZa5Cq8C/ik7F6sbu50TBaYD1FWdlvDHT5iINmIjwjRfjhZrmEM1q4EQ+
H3fIoJWEBuI9WAqdVPjWJrvo5FPaCJCZe6QN8R4xrq0Js12zuCacOPQw6gUmX01ELPqwnb40YcsP
tUAO874BVhkQYp5CyiiHluit1k3DGZyX38GVHNmmTtj14lUB8tRCBF4mmpC0MifDmtVbr6zwt2cH
ogCgggRvmzFmmnu5+W9Rt46XFimj3ytlqPlAfjrOF+zWofbxXq5R+zCFu1RiphNpM2vUJZpDHyjE
dvais+H0BlteDlBB7JXjmGXbD6mz6OJytKjmd4o73neuYwdWtkMSyJ66yzmY/5FD14Ev/HyHZcCH
qkKnjVhOZ6JZxOO8g2w7ZQPZbeZfjLiNvZKDTTx8g8vG69emT6ZK/GFjMpW21Uqe/1OVoewKizA7
1j/IQssBEmGqBV9YGUC2/qGX8fC0zVGR05DKfK5gKQEsh6X+ATdxmcnCxeS9544kGgfHD3GBwYJB
iW7O0G7Hi56NssfrDMyoYSQtkIEE1haZvga93tVdAN4+wW+vFjSXWcNQS4dI6icAMDv3do0A0fsU
GthGEjo8d7O13MVEr00/wzdCQqiukzYiLdz0ejN3FxRm1GgzRDWERPJzaqEMRH5ptS89D8ZKvk/k
DYZKLtuwykKUT4GYGcrQm83gHoxlCuJJYGOdsH7czu1sinNuIEy1GB4T5X9cGNqFqvn35V821B+A
hkOvVLD2tdCyqsFZtFa6IdxT0lkaMRcweegvOIi9VwZMBZozmQFdrjvWx7Z+b8lI/UG9mk7F4871
ERYY59CmSjHYKAfK9d8776I4KluNE5WHPHGvG50FiauxL6kWvOQ3Mb8kqB01F1p+tLkMQKrnN35+
XZHGooJJY2lR6M7z2VI/aGijVoIR6IiodwKzftpXXhupncJRAWLPeX470W9fyPwmK/obN1ktFgnM
KUkW8DCe8nBO84lXuQC81Qd0lUjwxNZ0+TpZvRKTbBq2kEFGGOZYLHdsmqgCQIJG/ppralnRKhXW
7D6dX4DQYekjYVniAaRFS9KxzajhELC55VRTmInEN194QkKQD4XaQrKp2tReneGKr4yOVQr5cRAp
go7dbmTNyeCpXmXBOhlAR/GoCprEiOOlOi6whzcP9Fp3fPt8vO/YeYtsTMIf6n7BoMQPxLcR95Ym
YA6wIt7M/h6TqHFeiP0/tUNmGCMsHG0iDOY2bJaT/AouJsHFNFpyPVcKkVY/I7Otrp/+eGNewL8X
6NBGajZ2rIPuLLnWQTeqCOaw5A81BTN+uDr55xBNoJVKPZNvKmIJsNuZvWtfDge9K4kkXl85esdl
T6ySR+HCZM/woql7lXHLs9MDak7JCSXV8cp3R2kCeGRV4//XpMDfS8Jol1nsXtxGCBYCyoZ25epb
IyzF8mgtWoirHNLZoYBLP+Jcf2bpC+dqmqUicskYhGCN7iKmG4aulL2gQc96BpdBv/XofMuCN99+
X+HfN7n5n9s1/gIQ2eqFx1PJJi3lGAsLRL1xgoI4TdU70tC6rWOLVeDHAetTkFN4qcxuAtDE2+qp
zI+4HdQFUV56O7WVo26kwuWziJ7wJEKiOjWhfjyonF3iCho7L3w0uFxK5gZiVw3SKDFCn1AS+HXD
J82lRc7dH6krldUUrYvzdsbFyf30yXbL9wFV+K7YCbZgM06PAjyoe2wUO0hV81KyM/isv+zUBJq0
Fo/eNYNlfXVbtpeh+C+hYdhpkinyl5Tq7P2qbfsrSL/O8xVSx9V8f6ktFNUrfi/LaPkPV8+m7QQZ
5fl0FFNG/avFb9IYKPIa+AUHBuL8VRRN5hHQw3lKgKaVd9NsAhSdebhmtm9pj9CclJVB4v0WExEa
DZ5Cf1xhji1UgpAPptiYIm7TZHgwZmmt3ZbMVVYFS4pcueyRyWOuNRlep+v/bcAfmqCRGzZFfz/v
0cClvJn7amVBfaBitvapAD4727tGBBnNJ6CmE3Wdq4Ee9SauFaIxvzSnO7bQzsdEfvpJx/V0sHv8
AmYK7QOwtwNdZAmmXsa44lRMhRhM+hta2dJGVSScH4B6JENFmPR1Gj5LnhkL09IX/BHI6cW5f6gv
YFZKgKk8iloMcq1Bt/lii7ycnaGep5TSS9ztYS0YGn6I1QHMOUk5TNIPDymc4ZBC54PWMmzViRad
QARE+n+svEaGBIBWtqDrht0qHYWyn4AJ/QU0lyrx6/Fjj9gLdPqyk/f8ZANLuNcfrDjlLzIO8hj3
tRpV9qjjH9Ffcy3jlQYCOB4OgzQydKN5WRyF6nBvw8AA7RVkjNDzXoPb3YbMviagpjz8h/SyVryg
LYsQH9XwRFD8kbflL7JeGpNkJKLHuRcTDMDAJE7QLOu6YnfMK2Yc7VsHFrR+wI+jH1g5fMO8vXks
YVz6f5jzCmnnvaIJAJD0Q532XsKBXBhy+Yig/EnP0oxfYBpSxmXn8JaYHYvXt03XQl200xNKesyC
97inUY5CqKGf2P+1qnIYoRgv2tunSLIxKBh60T9fHQrTDW/dfIoD5ehInQ68+XZyVGgPt9k1HTcL
yYGsq8AItTziYenXjJc3YP/s+7926Vf8pDaBIOQq1Gsx5xVIyguCzMYjudiLehPT9Aqitqa5QFHh
ZcVEdEvKHAg1zqH6KxkPJtCwkiXQJRtThr81VYHJlBGj97ljBnPB961WgUwSvOqnxsp25qMSpQ7z
fAVsCco3g8icR8QCootAey1TcQRTkSyLBvxX9MGHHgDEhjeDJx0E9rsbqwjoRwgO9d6hdELT3r3w
jG5+pQFqb6u+BoRkZYKNg5VIoeYby3UXO6q7Q59xcx23N1R7jHwJwa0IKOW1rF0ArOKmEW1IpC7+
K5+OAZ4UDMO5D8YrdkSYO6y0aTgjSPntjvA5LXD9wDw4nc3vi9pLr9blqYrndqGjvhldN2LLJPkC
RcFl0nNY8O77QFNLyaaQ6LNWOdiqpSEo3JtPpI2HpYapmIbQW95a8FK9cHIzK8twCveP3IivJPsb
i6TiR5QsvUEC+DMpVDmkjX8uP3AfjxJqgAjsEUvMXRshA0YpoybZpnLa4Nu7adCqcrdWySUhUWzm
B2VI/XNkh07yFU/RJTZmUQWSGzSjultDSR7+/m7qRL7ewaK1SJtgsxgwOgCX22udWRnoTWc6XGR8
BwTRWoF710Jpkyfd+hOUKGV8B9il1EIF09x+t5zUydkvomqrAXWvhU3fh82SMfkSk6HZFHIg7Pl+
vvp728r5e/+2SeIGhSaNIU0MKU2vjTk87exTYTD3g6/xGanactR+Uz8u/jMbg1dLhCFNvHhv3kEE
yM33hMKLu6a9fLN4oEpCcE3JhAmmTD2r+70F+nC7N57zq6qvMcPhzkcvST2RRx1W4UrTGtw5LZ9f
M7TQ2CvyrZgWRV6MU9JzWsVAOQ70nu99mflFhKLC15BRDrJj4qZeFe0qknIqmMfLZslkOlC/3Gun
TH1f/KYqwfJFRpTq9IJwL2fgRuEO0oTb3h9ezFLvHnuxiehTE+4yPOLn0DUx498E+4mluylHmvWy
JA4yOA52q3uA+pYaNFC2HLjSve4DFLOZAJkR5a558HN85BC3iWOjQY2tw1OvhYPqGZnmSdUhEAwa
nio2KJKU+Fmmto/dVa1FVjx3Qc19lPJmooPCcR9JJI2LN+TJGonOSWfJuPDizmUygGypkgXn67zs
Uo9i+s8gOUz1hXkp6YcsUXUsivC0PYO7s01o76/yRl2/TsGPLPAD9hHu7m8Q59CE39GtxDEzUwy5
cijUVJGKkV0DZHN3u+97uByMAvXdvBpfYRWNVgkC9rzDKzIu76PtLc1Y8Zorfrtwr/eEx+UmeUrM
LCoFIe079EESkfZLU9dguTDoni6eUR6vSYahBskqbr0GleWV6LCOuakYgxntNuBv3oUEEQuyQBAc
PeqRel7A7GVnWGCfI7yq5YFssP1QYa8OJW2kAwUXw5ZLk928P4mLEJl9zqjFUAJxXkxC7b5qP+RY
VWKUTH2xSrgMKKcXum80cA2VxxaSZKNd7p6wUttxeMbb/2wPKtXfU3jmjn7peebLRKz0nlalBEse
CGps7tE3K8K5nLNOpaKop/dIS6r6v2MBb+wya++EH9650s1mJw+IASiH/YrudiPlt3Ll8Tu8G+cg
lxZA17wfOOvGqw0ANK++P6Va8v4pQowm+LBLUK3yujNz0IJWeD1oVRZYhW5zwYeob/ZKErCSz8d9
/1ID87tkKQ+rXdGHGsGlWP5A68HUaFjmCI88JanJxgcPMJaDJ2DI4dFjjrbVFZsg/GV9mfUdp3WN
aiT2TOaZiISxfMxVTWmAw6gGAm6AlScv1OY94xOFURSVF8Ci+W53xaKfxAYyTFCZl36Oa3VboFeG
seVflKKZ3sW5p6eHDYgV6T82NEsIb1tK+2XUAmQ1hSuj0hfGXqebbO65Zdyg9CYEy6zNSS1Qqamf
k5cPPttvr65NBcj2z9G6/Sf4Ys7KvPXs7JCt1yYUB3Q+/KaRzlrDVRxPGg6444qoL8fICiyraDMu
VcEcGCEobWoIqXIKzkdxL7fgeMGbXBhHxWqK46KtbkWX8ucwEBG9ECw9gLzY+4g4SbeUgEd1JoTC
uSU+FssUmaHQKV7Twft69QTyWQmYUD9MbvQsxkk7dZKVPOn/BuiFUk3q+iE6Yv8aNRvvMTHt2+hg
ZrPKO48BFW4o8OiKADG1FSf8JrCYip6Zy3fi6UHU7AJRwnX7O/Qla2bj3kZWnwXnElVZs5Tl47Ie
gCPbsHMipmtVbKVPNU8ECftIkJPFdeQphTQNDUwh2/sz3oRyAgxp2MB1zsfxEe6M1GIpWeFrLYy8
NH20i2dDyeTNTB1DIdP96J3TOBqnWc98Ra8Wy+GPjQpnyY91MEYye+vtcuJisIRXvrVAnQDjrAHD
91k59NlLPJEVwMcD6BDeORXLQsfOxhxiJCv4ZLFPUAEC5LX1+14D068gtIFsyGHyRhm5r1Bvfh03
44iaOXJbJtQMNVJKE6tgsvd9HFS8pqyA/uphxtAvJtDUP/MAYM2XvJkMsLNoUoKBonhZ7PAOsFOy
YNQ1RQzVtfzplPEavIHwlZaBER3sKxHHdt2wwsTL+KbLdOYmFjI8NJc9lwM2J/69Ooa1H9mL20Pr
mpTKlqfre5gZLQ7xykAL/OvKxWqPbVJaXnnSs6RuDJB9yCVehfrSo4aHo4l4x7WHLtWr+egwVw0E
GUcWaoxP2YlQy5IsJvTr4xvXGp1jdU8SDiIvgGMCBjKVIIvvgHb5JwhGH7z/g82H3/kY9eF9+RiZ
qkwDgmkQiggkI0soVoHCeltFN2HPIG/XCR2hzGPJH8eI69SymOQcI33vdY8t/GF4Hr0Nze0TDyFf
CHQ7QKIY84FJxFv07gbouBbqHh2dRTSiXhF6zietqEVKWNjHgXv4u47l53WIVqnS7kifQhCCJdW5
hbAYICm7EzoRvAIxihjtVsrJthgg9hvW5rFxi3b3rA0QHb4MtI7jcrxEwaYf07WFbFQ6YGqafkg8
Ibk9HZNza+QtMUH/26Z+3I4iR6UvXrJxjTZ6CoEJi7ni0kHDEjLndauAxRsLieyP7yq9AuhFFq+Z
uF2Ha2eQtXnha4GbUPLZ7umz11CqgAuahShopmlxiOKdC1tU0sj618mFSDtrUO7FaSPbwNR9qPR4
rxAaYnN8MZ5XzOUWpA4owQ07p81Qoh5qUGQxIzlmRmPmiqqfreDGnvuLMtfMa6oXzDUj+jrdOoQi
OJ9xiYwYwheEmISti83Z8muL506Q/doWYX2uwwZWvh17b8Q8yiGSNXtKV8Xe/byISo/Pe5nVk5Vy
fZNmbC/uzRCqFAG7BQcdEq9wTS+DIjlxWrX+pgl9JU+jlHzDN/m8Q3lfuE/qG7E1kf3iBDpWr1g6
dL9YMhqfoiDJjBS+ulowEFvllnPzTvPJLIeNZH5Z7qiLVw+bfB4dkzp0gA2hokGnl9e/EkeJwLC8
yli5Xaj83ZI6zFFMuGFgXUKmCo4Z0avrPmCddmglc3AK8+i1yM9RhQcqzp9z3IG4EVaOAd7ocro8
mMroBoYiO+atioI8vbUTBSorO5f68UnpnDbcPK7rZAeQPCThDZeqFYkGa3GrhuHsICOHfdGSj44D
xo1yJUk99Z7zUG1jaGU40tDTOS82o4VEhxYXiF0n8UMKY0pFufKlc5EDdONfL7kKAxqO1zmq9U2R
1IEB8k8w+h1HbRK8qyI+Cqu1/AfjJ2b373WDb76g6/Y/KX9u+8h1rSocNVjnENjlduqKBs3WU0Kz
YD08Q4CFB4ff05YZuVoPfwgDIZUsL7Kwiz55a8UyuzybvJv2RRmNjb1SJ55fk5q0r0icbERyJPKG
3aso39bpJAL4YMIzvgIMrN1WAhhGJxyLAy4MB8ffGyrr+FrJpppDO1E7PZKWlcXuR/niUsw5mllk
izNxLLzIG9aGpiW2luIz/3SrYliXNPfcrWtMkJ6lRo2jdY+yCc8na9ZHTqQHKnWIa542ab4nwx/7
kwY+GBzaOrUFpp+Ksoj/X3P4LV17UUTXbU4c8wdK+zC6+sIo5MVnU6RrxDL19FcqP1ZXZD6vYfKM
CPxvuBSiNWkDzqpz52X4oCx3LY6776/l85J/aMo/ntONMRYgetUhztylbG9vASL8EEYhIeMwJhVy
AXChXdubi40c1SoLz0W4BCfxJmPsLVXe3U3w4aBTOcEbQeB+ORpvshVX0XHJxmFqAKhcuHmEpSkJ
T71PZgptmgem5j+x9ng+w3Q3902CgqeMWGAGCQblybm7lA1Xhg0gB3GSMh966SsT9YCoTEThOQFN
PAQ4zhLT8ZssM+GZpY65FhmpYFFqgokcJJvXCMFhuGyBeJ2k14VZO8n+QOt4sdPqAacqX8jZPHwx
tLA2Nd0B22CApN/2I2l86WM/mDwIAddZ2GGhvBRLomB176UIjCJ2EgfE0VNDjN3Mp2IIZthhQlhS
oYPgEQJrrsOJE6YbW6Jrjpifz1I9e73Q5ie527w/vVfHr9ebb/aL34zfgi3PjDgcKC0N95ciqn4P
TiIDJGXDSNNnoEV6vUWo5Z9FocfreQ86TDmFKw1beulZP35gfeBYOOEBpDhlFD/3OsajQDE1kb8t
j2fEUXjeYcpS1VMyD9n6aFHh6YB555Y6DRiHTbU7SwupgRXVRtlShOo7Va9retmFTb0XCKJuagGY
EAAY7Mhu/pf/fwxvbdOLROLT65GDMDBSWvFRS2AdpZSkJxE9Nl5zDx1g7hCSIlociXL+oUR7PIEy
4Vzcrk7I0qBXYgXnvbKFvXDUBp+JBzBTEBBxsXdoPMJCNSewCza13UTuA+9UziUIfOnxJ807lwl5
f3nHJKUQdVg5PglgJHaPH5wR09uK0HiGxtcrFG5rvopuGDGik5XV9+WSu/yp7gblgvEc2nrgWy1l
Y9cdJSSQl8HQJIDZiNSO7s8DmsP7nHrsLMVuDxgQ3gmLB2L1wqlag9fv5zCHOrPgh3q2sUQYKv0J
v5no+gXvKbWINHu0t2uaYOlpKSOKJ3GSUk0g0Ey/v0cbQtMpfFyQYLd70IW5ANvqzgbOIte5tA/B
CbV9VNQWysU+M/QTMg9dVmlT9InKvPc2252+jdjr89oxh2Xm3toveosuFEhE5UzlLhGR05eURGpT
zcdMri2EPkbLzu3F5VFr6TO/VJPbvznlTmHeFup6KCKDxO9lkCvztblUzk/SPGlqZyL5QlcyRjiC
f1SfvmAmkdeOOZaKpgAG9kGveruoEIAT5BTak3Tpy/dDQ3c9hrdvGupCQzHPnHZyROYOmhUe0AmR
6fncfKh9VnjN4urcY/DTo9C+I4+3uEOrtNJOd0u9bWSOSrUBtrY0dGBZp1DxKgnsEocYvA8jTyhp
JelK9KteYcQ8V5e0CpxXlpG+PcdfAoCzG5pWyudBdOl2AdvW227p1q+tiYsDZPhcvNPvdujjVCjc
osrk8Q5cJgn2Ik1GhAs2o6YqRPfLd5tGC84E5X0DoGwJzXcQ9JqoGim2taM9HA6zUn1QX1ZUmV7V
SqNCbwpjW6EmK82CkdHCD4BTeM4WO+H0k6ro7YouWZxRekuDOTT3ksJdLkcHtF2BGQsYr5vp40J3
/LPIgGCXaaElPI6MXhbzEb02OC3YolrME5b1a2ZuLm3VF3/cIzoGpmoTEHr6a/muDIgAC1YQu/6t
IQSMIATD9AO1dPNS+SfqlReerR3SZpcOMJhF1x4ZRRmWKJ+qdYljc5NaX/P4ohcrlDLmz1UsEs/N
x0DYWr2R/9/Av2F6UzbcrKBUbuSqZViQkBhErixuHeLNTLVdm6P+NwqLpd9FUDuAemqsW6exbdDl
5fBoXpsxBQRCnh7bY0v8QGXvOpRATMW9mdPpz7anwzGZJEAulQI1HliEfxbMYOXsjqmTFigEzHoN
AlQb0/aUJNYgxqUR/m7LSPZPh6jJIBzsJ4flVoRWiGSvMJjDqdN8926If11a02km97CvxkxDvJA+
4Hfs5XhYYv4e0/BJ3sr8zQUUxzIlRKMmjkoR4BRvomHAs8ioDqD/YDBN06EdFKbaQmqUgnXWPVUB
SAEwXYFsmA2ybQgVgnXMIu/fam8arWbirOhKzhBf5W5WKHcuwAe/sOL3M1uyg5e5cYYjc+K+CJZ/
krPImZgKA4Ktqbd0Q2pj3ZCLQ5boaYDTtUlooZQI8nJg1mr1LyoZO4hdqCwihvwHS4Y5KhaI8h3f
F0n0V76yWwfFTBBUCp73Nm5QCTpEh05rDUalbnzsD+sdmVjIQl00uqEYnaGhMweR01s6jZ40ONJx
ByrcYu0O55dAvGNsGj0pYvfh/VrG1gR5qJD8iZ08tnPdfd12koMOefPNO7haG98K2qpMkBsMdL6r
Yk4b+nXndQRat5Ra46W1Itm8CgpsUWSsNwtVlbwPnoz8LmXUKTQDaJCh548HU+A6ZLxlpAhnscr/
eDBQF4jj+JJP0EZNL02FhPmULxr6quihxnEGhCcyxdoQR7+6F+5XacvbCK4lSqnCKmExG+GMJr1o
s41NxDM4t+PRJVoEeLzlxinkSz94FyTu3v6l2XTH/tCp+pLYaD1Xgvzvh4nGwhuab1Q7sFkqavxA
bPBZL9JbCV2FsOz8M682UlNqyZqL7DlB9QcI2CHGvtRK773/+KRSjF6as+6yakAMwL0GoDlkHK5b
+n35eEdm4pwnV1wKS4ZqVUL0z6icsKRFrstrOQoLOlt2CoxL1KBlfoXFBaqFIK8E2KXReTVFaSk+
pwRMO3iW0DfTnp8JwIaggkLZ7H56cXzevLeqZrpoeRS6/5DzpAjIyQWksT+ZW2r9a5h47z+7Y5El
gvrdNCYDZTs5+kwqTVuKvX8DE+JmuGHjwFrOoc/K/x8Y7Ps802Q4XtWX6TbXYL8c1JE1+dnfwddV
LHhQJFgMaA3inWEaAM2qVmajRyoV2ntrpooa7fKvQsuT4XvVvxFuY4zZaPnWth0o9TNbC6Xvuc1n
Oj24nBm9D9k6SmLN+YLa+wur0p0J94v3zZLf0HBFtYEbpUe4dp34paNwircR+LVNxSzACqoCJgyH
sVvNVRgRIW2CINr/A0CgPgordbfh6coHlax1Vanxwuh4Wg0TrVXn4YOEIap5vV9nIwA+amdMMjKF
OZ187AtgSlp4BiFWqf7dOzZsxiSDdC3yKuv7Pen508+wJzIs6kVqMu2bRLiV/4s0qSr8Kpx9P7+7
x0laMJMi8YcIPBQ9SOfLTgH+uv2AAc4Zv3aVHLkFSGZanWftx1zxMRM11paVFoTJnqzefJKmoPI0
OVXSnfcP29K1mhUk64ytGBrNToOhjl5yyAlKe6geEzk8jpn2ifPIGv9a9nVjiGNozqiCl2g+gFdV
de4VnEKNNVI/PzuGApcYnLgAbOZjGBpZWmpxcHQAEduWcTm5dqpF8/W39UMWE3cgl0WZJZ9CV3LD
OMxSV74fx1CRk41I0Hjvjpq9KsoFx8GcS7oPHjyrBBzCZdvzZSohpjBHjYbzFr04tmlY39HM3pZj
uMQHWPAYVlWsP7luQvsf9Wt2ze5Nh7KLsxaViTQuXxHXckV28ZifyshXkKAYEQqsjoaxNJhvICdG
eyGDxbRXcdeqL0JQlt0vtflJfOU4UYcqFJwAdOybSaEGmSHr5YvDSnyLK8XtAJrsyvhgsf4fB7J0
Pg5t2ejeJv/dRkEHrlRegf1xvfMfly56fMSKWIspTJq4ma0gQE4nEswEYYwX9vGBlid0MLmtphRp
1sQVyeN9TWQMD18MNug2XVkuzMrO3+O8p9MImiFxVhU72BQ03OFobUhGzr21BOCcAhML6Q20sWmt
ftHrqmScegWRAhj8iWxp02SwPM6MMXgSxhqpvm87Q9kwlJG/rhwC+nSz7sfZzQklhJijgxL0gG10
MmNXRmOtxD0WipoqVk3K/HqzjrmO08mGnnkRquSUrCJWXi0W+RXN/QhgXOF72ZkBZ8oJP03Ow56H
DdbfgC/ysMtUo7dL+3FB3Dg+KFC6EbEEe233UdcyF1BPeTg3en8j1RcTyjUbi1V3kBxlDjypo8pa
5sIMHdqiL2O6Jb2Ay0H6C6x9hyGp+uwkYA9sxJ3Gkozev11XbZDzFqkbI1u75FCmHq7edG1gAwDD
Jl2gXHys7zHilj70VwyrB2vlLUmv121f5woSdAgdknamSi4jQ+TwcSXJSF54ZqWukRtkS2E/yi1p
OTjrMjEO2tgsEnjQV44r9GCxqX8QGk2YPMSC5VtGYCrjZKFjLUQHserlY+jAXlR7kxYZKcVGS7Tf
3ukrjkj2GTDZG7M1UNJXsEUum+C5mEYZ8aT87OSHGC4z6FA2irljDxqfGiXOUYwoenvhX058hzL6
m2xSnchc3kkaG0lvGC3OpKgdQRkeZhmb3DYijxRm+QncCWQCnr/r7qimGEnsRNjIj/NZSMurasei
iQ/qcpWKJRhUZ5A3bgJjjrfYluNk+IFQ0r0LfFH9yeKBei4GdmkQyyUMMMvu3VFf/u44BNVllEy6
QPYTBQlZoKq55st42AqoGvWUipPpfOd811hhLSM5Fbp0cH8yVsNUnJWOKN9U+cb9HRG6YKGk32V/
NSxzpYLsYetmCey9WK0JfqggiSfFJZG6kSEnTL7wwkm3TB177XLFEsy1qv35+SwxWszJyJ42XM4D
pqkZbpoAmJ2lp5M+LdbTW4A3UsvRvDVX+mhmpl5J+WMXTAhZsjQYf0JZ0PCpHZr1G0PIy+SiZBCi
HUWdRN/CLC2Q0hWXfeMBpkvTZlA5zNOrz+mBTR1qm9n0keSwP/teOKjepq1k93WlY7vX5fBpsPe+
lzPe1qEOQPMrITIdfdRtAZp5ZgDryIlcA/rL309Fq67fI7I6dvP7+ROjGF+qv/8jqFsPtr9PNPC7
V3X1iFV0QZm9VFbfSnWGe0XMpfklCgMlqSatyZIUcOYf3S7NYDJEWrtMdcLiZgli+PcsBr0Y4Egz
DqpVoh+xlFg0PamKJCZjU1Dy7F0uDMraH6GT1VMNo9poSx8aXUyFHlq/VDCxKZ8IEv90yhoMr1sZ
K5llS2fLCyezB1VpgqqAfxAOLiChRH7yjNdHmurq059bytD1iajz5/dpwojJDK5j2vx4Ynyw65Gu
CFqv3ql8XPaR7f81CCibED4h3Gnqb6hwbNo/FkVPx0ESGPm9X1y46kFzIa7qatILTQlwpOnmIGEl
VRNnFWOTEfSqr7UdGstiWS/vAwWOyAzu3fr45n734SvoYxee65A52gSRdIEqPUsJGh1NW/FKNt2w
eXizjwadVddh1mxxehH7EcxIwXmKy8DY9G+S7MFU65L/L10zfMMFLIDXMwEDPb50oauUKWQfXc7F
tZC6gY3yQSxv6w66QMVEsIfHl+mfxSOW5NC9WtVV/4MNjOZi6ViOqSTtcNc996+b1psU2DzZ+zzN
RpG0OMUjiHzUlr1kNa5KmWjZII1SpjNnd2LMUPa4YaHDh1la6RBUq6pm8loUP1R6zbFHIBilHpd4
9c+Jd9jUXUT+rC+7pE2ycOkJFtnb6Ceq9TgL7gH2YienjsxNfzv8nKVEbXgJsy1mdSQ/hm25628d
79//fzZQ2St9H9SKZm6XxxALLntb6lIARjb9h7ishFhkKgSU8ttBp9M7G6q0JRG7Xqp81KRYfit7
m8WEdQ3fb5oPHAtrtDVufuvdTuNKBzJ40a0ci8mgKu0r+hyWXDV/DQxqHB3p7pzkQG0BCqQYLumQ
rF3ReZfWGqgo00e6ysvmidATaMhIjyX9FbuYDX113KsMHLfqWmRycNdHd9cArDKrnremDfTViA9w
CB3bR24JTyydvGw/kXpTlk0gLAoxeko8kB6AuDpxrWZy5fJUCO/DQCzGPAO7idOlc68XWtTZ1Gbs
7kj/kkvsCDVsCrEqV8Md6rci0vNYlH10iVQPKCjzb6yqO1qbdTSjJCzIOkjrP/7lMIL1Ty2x+KWQ
RdjEqYKYHVUKVFb9kp0taKOzBouT6TlKUylyL+9Kzzx2i9ScTC/ATX4GyXaPztLDZJ8081IE3CpT
Xv1N6gXNecfVH4Cii94Td3Z2f0fkhE8+064OuAB2S9j7Os6Q6v00AiotajqJiIGgGapS8PUijCz/
LDVTgipJ3AlGd6Uqf1h0GaO29RJfSHdXGDsjeBPMOvW9ikk7a1rB8iJ/6yG68YZRKKi/sEpowe2L
s5S3mhCGZsZsoC1gsBG/d3Gx34wD96sRvhfAuICtAsyTjVHhCpl9kAVw+L+e+P6V44h6EvXoUd7z
LXZLz9NgqgVcRx2SgpsLMUmTohHNKQ0y190hTQTrSgkMiP+RGWzlyZ6iwPXmTRfVKXVaV5MEd0CW
SEAXtIVqdojGqTKNXpXFFcAmLyuvGI+mJiKHvYcTmraMXNGFiHOnTY5+kHDtxjpAlEDIqHO8Aq6T
gfWjtllMBc62GVOAX+jGn0DTfS+KtzW4mIfisi8DGCJ0f4mN5HCPXW09cguoVXvUpmMTrKwt4diV
uP0M3BjDsI4e4fbeWdWROeYcuyCGNMqzkVXjl/9AQyIUcatyK+gdUhFoO6qUIoKeZzHJuHJM2rDv
GHRzg5Nb2LGIe3YIkxpYG35nY6PVp/kFDTvniqGBvalrYgpA7Zrn5jkNLSjELm9KseLTcMTRGAuL
Km/l57wRDxz2ijDT2qN/c/zJzkT5tOyFOzWFy36Hr8I5JL4sarDAXusQb7a8EgAIjPKr4TUplmKv
SKTf4f7oimkVCTU2CAj1KBzalC0UTKEH22qKtSVSlQPjAh3CF5V8gdpgZXhwirNmEs4AJp9CP2ys
eqWa6VCAca4pC/J8yLIxgy8alXHJ4mej1DPfrKCd1p6sbso5WPi5FqHqk+gviIFA/NWncMwjVq8q
uwGt9qdgBeAyQFmECC8wMsrvBv5Y9K+C/zd4Zoi059TyYOSXu/arVxI7gi8LkgaNoZete5Uye32I
PRUNy4Mw44oODNm54K4cyM8S44n12YC62ObITUjll75RJ8xx0WeV6DrccK38JHt0cHOAeHraK7/a
jdEkhm2kGK6MKh8+YnNV88LXFh3YPGPvrM95nBvTM4zEImRw2Nz9kjKQGEKUNz5dY6JEf3uqkNF7
MEboljm2gr87H3inKTQJJOXMJ4RP9kwKyHFSyU6I73P8OhIcx07M82Gg8dMMwYr7ZdkHiPvGi1Jv
SDi/66KD/Tl8W0QWaWdtv4wWmnFAhScFcdk1OeK9XZELhnpMYeIoR7cli8GgcNyvJXFvrnRzYrhm
pg7qTTx3PFPFU6GcpY0fYHtYbN0xr22QRq5651Z2YKosVb2AhChlowo+zQc0lOYxIfbCe+bAhoTD
38DU1X11/M3BbgC2qlbnb/77tsz+W5onv868LlqSP3px9ILIqOdPd3IcMl2o+BAs19ITkGnJUt5X
5fDU/S5FTGm/es6764lj4AvoGsfNWou8+ATh8a2myKvmRcEzczg7wO6rxnLET4ABLqu6usq3cykW
lAhn+0hgdh6edUJl4aA8Tzt249Dfwj3tJFY3p4iRvyo5lWxJzvEqL7UT/k51AagNnj5tDgtPOyuF
jyWpSW9NJQwyOFTC5I0pAhBI7Se6JVRlTFhMumi4y9Wo6Fhf3yLX41OBqi97edNbopPeIrKOdWg4
zrlfZIuIATkkYYUxUk62mP20LFGGqbeSO64+iCrpzH3pqqiDM3fJKmXxx714Df30TS7gZ/BWLUVQ
250VLx2Iq8g/HtDKUi0HYdRm4LjwWq9PvIk1/mG6nX9LdQW/7IHm9n1yBrBHDV4IQewBz9vvPGiF
O1ti1lrmsBQOtbMyKKEUFoQ67tkYDCdP+yNfhKfmktW2fI7QdN1qJ5r08ivEBnm49nuQjWYo/XKx
apiYbmW0gVqSxhFQ0tiPpYd1b+Cj1lcFQRfZ03E+jGBYgM0Rsj7dIHlIijBfinESfZM8lhk61pDs
9Bpn1f6IXWAALZqIsX9UjDO6m0xVX+YKf3w5lHC4OjYqiNlAgWqM8mWPN98/Kn9KdbiI+CRdlyLS
fGJBtH8r+IVxsfNV3tvlv9DCNe96Av91LUu/BQl3L4PEY1pGFDc1H0VED6+90+UFVFH6I05lTFwL
yETg8IKyolXU6tkQlQKzJbaMc+UqMLMRFmcU10mqsTtfcPp/FKH0ncLHIg8ma9Js+1qzvPHSkTCM
Y6F3SWPmhHtJvUD8l2uxonl2lcYqUg8AwTX928Kq5ds5iWqqVGuoqHSAro6fsLxqOcC3z03T9sSo
Yh/oR1L78Tm62sPnVE/CodeErGO6UDAKq5J3D2hK6pZgfsmr+PJpQTv5l9ZgKfqM9wt5rbBFMG30
/0+bzepn0DkRR07SdqBMhVNOGIkzeZ7rOaFBkxBYkcY8d10hfqhZx3i2rAbtqdw9dQgW9nbbK030
oQ7bZ8mFlEly6JOeeGxwNCppEx5qB/jRR10C6I76Z7iGeq4hsuToG4xxpAQkxshtlXolCPf65t/j
/vNhGRu5YAv1lcfz8ITiY7M7Jwi9dMki6b0KSaOFygV723w5I5Tm7jAdVoFku1mRi/eUFGdKPx99
k/1JTVlMapSYlm8iG+8LW5rygHmp06hQI+YzXp8S46SYBsfESIdKT2P+E2aS97f7RWs81qSq5ar6
m/ruYl7WNSwSApZvtYJWnbOAyEWCGmQjZ1l2JiHkZwQSx9n+NpyeEEj22DXnpw5WS228AKZi/EIJ
plwMdzKRxCOn5atKOfu2Ep+8HZtvkcQLcADk5HEwHzZp/gJqim9rRiCc2feWrc2JaPZO49xuxU4+
H8Ymhe259VNkk3Fcg0B0H2eCixMpGR2zD5kqva8BaQQyxB/00jtM8wxgmga67p+Oj+3mEzYJgmMm
T/xGWqLywwx+gyZKbbETlMIAjcxz3gEO4Q8vNAknSagi4VugbKyD696ggF868xo9FKQ62c/ELoKZ
VqbYr1O4FyqHLfa+Ng0mI9Nqi6Pl9TOlqlhY/ld7f8YA/UOI9I1wbR+7Oocls3CfnNidhqzpn06y
mmlTvjM8A4vLUtl7Ci8Im3MsIpbo2aP587RqYma+ZCnRdWGlfHr3E+3pZoXJ8SUNRIRUQ/rU7Qt1
+7GTTam15jET9ZDETnT+aVimIesed9yaa9DaUY+dtno5fhYrdxVn9yttmszb2YP8B8Fn/mPlNvfU
YU/Ga7K2URZ+DS0vmVlnod0yRmhcQ0Cp2YQ7NUrJoGw/pxAEKKoHKMlGYjf6PKlxIATHiWvYFXDL
Bl/dAAAzb1a2mHWb3S4pNbYoiXwvNUhC5OJByiRKnJ0njk5FQJLbjZ2k25MVgGi6d1JpByxrH+lF
zZPH3SkY/qaxFqM6wTcfMndu110KR6pGboAUJi5au0gAkLuVHS7+oHdplB3Wggx/AGKD/MX+Caps
T8veMxX5DHSoOI+zUMuzpjiOR8EQod5P7nqriu1Y998r3swgPLWAuEWRBvOEoUetdhKM7seCljvh
feme+Ov8bqCsCl4orYE3gYBdolEcaqKPDLtZWClsTztDZh58dqmzkj3eoZlA1rUyh/CuyKT0DkpC
KaoDZtiwF2zeKXuYRqadyr+othdH41AWmzYkZTaNtbpJj+gBmSie+fJVhFUOepeN34BUstxjZhwc
fSPJGqzWfMC2K7+WODn/r1NKOZp2RWeDNvdAejV95fC9sM17YSD7B0bEKMdQ7gFyAIw1RnBZP5I2
xr6b60W9/KlG75EKq4s0LRsz/0ZxcjeKGRQhZt1pvHEml1ppvHuujYdG2ExlhwuUY6XGd+KZcWiv
WGmRdceY6hdDejIRHsLzo1A04HOKAhJOTakKwKjvPU9hZJcceCyC2xlt7hhI+kZgtf7RE4b1W9tg
tF2o7hsGGc7xZjdLU1bviVOSXAba7Je3ZRluvL9+H3qtfgviIEjkEA29zu6L+XgxGCWUPBL/gFYN
0YQmA12zpgj69QlVbmd8gFf1d74ZY1rxzJn5cQYKb4V0DPLrLuJinHlbl7IM2Nzww/gmQQAgVBDO
013V4mXMYvdXjx/B8Apgh2AUM1T6V8loYnC0a6auFSC/sochtHgpt/Fhf/C5PxfktfXXksepr6c/
ptP0QlIQ9tSY+DFMvZ60f/KiD0ilZJzrqdQ1hmAsz/InCUcOhDS2Uc3sPGNPLP87ZPE6EeVLHo6/
zWh+5LpIr86DkqoHgwW3H/hxyRjV7iVJ1Q1DLpQxggNOPDEMwiTVWxhvbRn8YmEd+gYdwygET1fg
/VN5zixHhsvjjOigjW5thitj7LplzDPTt2ZQCnzgsNGBGjkBG00+sy0MA7AKKrYhL52F89TNEQmk
eh8ztKGkDc7ZH3/D7RsvvhK63TOAOf+TrvQciV/a11t5ILvmEXBBZgDDmwQ9fJ6hlsAg2h4xVgoQ
kfqCeN+CIqNZ0av44WKc3bPz6UHf8VL5HQRkCaebcviRlTtFrxlfq6oj3h68h7ejqWHzqw5E0DD6
Ej1W63SibMFmQWBfX8uPqc4FDT7I01f3K3eHmP9BHlUHIKlnus7T4JZrU1cTaSnVhZWpywo4Di1J
OWbrhfvNL9hUDsbJ4xvC+0cBYPZ5GMTFnyK2nv0Mw4Nfb6s0KoImahOYvXjIrI02iMGwmsduRJYG
VOiNTnrhiT4mCf1vwHOnFse+pSRwGlhVIh+4QQXccfprn7/OWv3A4z7Qack/719709tIPXIQx73o
pIwJRV5Db9SpV1hrXee+a5Irmfq4RD/+GLYe9DwmQMwNZPjOurQDAQdiwyO9fXpTSS0kYVDxiw/x
o73uj00sU1FV7XNIkjBBLB3Tl7EInbcLPK7wXxOULckT10C9DVhm8cXrrYMn0mDlxRhhYmSi+lIQ
2DwzCES5oelrvyo8p/3NGDHnGfLCXqUZKvqx4bzgnxh9UdfwZoazSMheiJUDzNiiieANQ4cyJoDM
1YUq9pHy8AW+sb0nqSpA5o+ezKcPA4F+aSKvb3c2RVlX9yQhnAjNmaFYRp3sJA2thiRk3e7bidx5
kqtc6L+lLMXRFHBHBk940pqdmxvQkx/Qu7qV9CFZM5dnHKS/iHZyZFfUKMHd7i78EVqQiG2FlMM+
xNO0RXlQeMsFEGEdv4f/CkBkT5OUqCRDk70frUpcEv2M/0hrodFhge437DEezkQED7NSaBKI7Wpm
YHt2A1J/VFC9e4iuzTp6uwmhy8MwVlR8qslohedLsXqPsaf/7+4A5xBWoI9c3CfCnsf2frkQq1rp
NXoR3lopNzXNZHFSfex2r5/tRy1QSa92le5MkmhIr6ET0z6tJOVJvAghRnhRgDONKBXEoYlPoPBd
UzCR3xgrAqN3QLJlJwvBXJv1xcHh2OyfxJgx4KY/zhB+7kORN/KbylxSLXzxVDsRftDQAmuBNWdf
JQHD/Q79TK310UgfE9uf5yfP+aR97xZ1kRFq+Ex2lZStR8hDqqSs59Uka1AzacWrSexs4Lvdj9jz
4i2il8Zf/7YCN8jyg0LjGWPkhkgRTTfPi8vke9+JKx7zJL9+KwZFKQJNqCeP0WClD75Kd7+3t0Dj
hAX/tC6/mPJUG//b46/BQZ6jyOsL7a2BMGv+JkrpTPNdwsZlakm72d3sdt5K4jO7JniMNbf0nZID
mjXuSiSfsm6pBMzFjTM0I1n7qYGKjNPAfcJcjRFzKKUhAPIPLALNEw0yUbMHsSXaTD/TPoqo1vVp
eA7vkT4eG+FfzLYObAaJnqCE0BeatfC0Tfyb/+CAeSWT0tztzVphXhdCxpUTl0pDDKAaV6iw8zC3
X1aC9Dlq10WpY4xao0/iwn9MGZIccN4iSByh+Rk1VQCDOs7WH3DJ5iXpzK2fvAFSGY7PokE1F/Ls
pMUNmWamw4BcVBv+t5Axva0RzripQRJP7Q8J5ovdqbFYTwzAvBetNPu30O8pYxky0qqwZKiVCCRW
gWF7LKcr71zgjvCDUFBhslpzpRt6WqINZGbcDck1pJvZeKuJ7SOITF9GmkVyEsmmHTX8dfTaPiXB
hJ4O6/0sktBA/+KO/OriJLUfjnbM54iC1xAfdywf2Q5bFpRe8LhrmabMZ3c4rdwlKGtuReQT2s6i
Mqyb72F9iGFdFziFVp27rvQ1sNjI8f9MtTzhZadISB/i2p2FoJb41aa4FXr113bqlrSzOwvGquQY
1iTZQV9jFFkItJMRFDKEDk8XDOZz/H8XdmxCpvL50SBdpTenUCE+BXAMOUVX7/YXuYcxyNFtfmqA
1GqeeJkJa3OwL3Q5VoH2AHN74EqovOY1FZs9pwUvm2WXMOXeJoEShoUXIn/a3IB7IfPXbMDByw7v
HR0YdHuW52Mtjgdm9NW3C/Mx/3X2x0OnpxaHf5xAylUbIJjWDuJg851UXXPY2FT0rST9qsktO1YH
4BPIEqYmkEmXgNWX8sX66CbB85p/ucbVlZDGLyr0aUwa8HdTphPoAPzzQtzJCG/6/4OWdSXmVgwu
J/WtjNyPauoIf9BnnezVlN+7hglVweebtcpLgDYT+guvGWR8wS12A+GZy3mCbg2x7xkAWSX6zKP7
pQgaekqqlOw6PiX2AP1+bgRtThcsyHheubEZClZfg3g5ToHL4inrWa8zBG3RHwMWVREu6lNTVOfh
d++lKpnhaMcRl1wCZ4q5u0Ni5TcYBKUhJqJ3IKND9kzZyE+KY92yqAD0WtGRdJn/E7GgTFQpr4mM
xnpVg5RdnKinko0GusonMhvcAjaUnLNGEJYCe7gdqq/81/yxrcg8fYaZGveC0GrBn74SRMw2AtSq
lm4Oov5jI8TtpyWh/y6HjbfQKvVksgGL44UcT1VWfcm88i4EJjV16Y75GqUf6OIROkQhPuTMN7E4
RwjDgRFp1kzYKyp5f/cdY4TnoXgxU4OqytzkWNfhFPsxPxB7SghNEzd07KXI1FoicK1/z/J4DNra
xZg/S4dk99sq87VasScA19SmYp16P4mXkWjHkIb/kH1p6QpeSOxr5yODjSsO6558tX5IEzZNY43D
2KdrZr7bbMqGG2bp22oWagrqPyV+Y8y20HVBSBiviMfwHPqGlf2qFNNriYk1pxeoI6rhyC7gGifm
g3m9QOiC/z00harATAG9tEp7IIdildK9xjLnsrCLKXmgNkuZeXseDU8fEVZtWpqinH9W5mV1TjI1
l8z9m7km3QzNjSGI7gpbRqcDqcpgmLsF3CHBIhVaJ3pf52ZzkaESAJoceCxkLQKRcwpRToxPGl/r
8CyeRELIZ25MmM+jTZ4Clip79s7LuEADkAR9jopjKSO335duP6D80X+RIOQ8YRI2FMHgYfQWivzq
LkWFlPzDgcv7mkqS00KdI8RPjli1wv2WQE1vwFjKlVi6NqWZt+N+IoZv+Qwg9Q+pLZAMeWKDcCLZ
OlXA4gDU+vC60bkobb5PbV3THlOVmDB+xdxqW/Kt3hrDIThj87HtmwD58wKDACEnZqoRnVTUMz6a
zKI72BMgGFO99kpp7UWArvQShm+SzMlXY8oZ1hwA7c0gDul39LCZFCGUiTQzHrTdamDYvbFPqsrX
tZVAxE0SjBdqxIET+KS2xI+nZ8mH6jca2NW2pWxsWoPLn2KLBVn6QsNsAPZUjRlnAualEHTEZSSD
ypGDrx4H6ZbCReW6c+huJN60roDGyYLCWLM0Gca3ceIVmlL9oxQCdvCx3y8jZ7UFM9UnzvH2OLnd
Bq0iBhFdeEr02DtTm0n3vmmY+/8mSKyr8QF/GLf5kjvPTGFGsdpj2UBarkCGFcrdaS7+ZSKgHg2D
rBCRT3ZESkX2Iq0v7CvOuLAZHeNiAEeOxy9RK5oeadCo53wXc8nRid1OpP4PpGbOhOw0Xc8LqzMY
cgq6Pud7OLYTC9QQWPLw57yOgxRYtu4QRJ8BA+UwUmQNSBmjaUrlkwZwMFrEBWo+icYxoziJhHWV
CBjKJw/FqyQ2uyh2Ghy8ellMvuDCXrXu+TJV68h90Kr32x1Quy7y2QX2I2XFkqoILbdTyn1tYPJ2
oC9j/OBLO8I/u6Nm6YRUkkiuSK14DMYeYmp6cPMsHXSKD2tzEodXaN0obZ4EQRg92jet7R8LgE4K
3RsFXMdLQGzw5fS23geYQ1LSc7hJYyQOY0CZTriEQI3DPENeM6Jc1+PJmLkCtBdEBe+1vwJX+2RQ
qQgzsxqfLTqEMkGyityai2VzkMuoZXcp5Hnu2Qe+ESVRRtw6pzaFLvW61aEsxablN+QudDxTS2HA
zI0vFWx10aQTizHgN7JXADh88D2UetgdXI5bWGVakZCkCmW0lVjV9eNUjdQbEGd+/lQ/ctFA7OBV
Wb/oqEkkWFt/hprWDKioful51z6BFH1TKIJ7KkITXRfepFi6i9DfdnR9qT6/bxf8SxBamlowclBQ
h5DtTEfuSJC8DN7V3DsDEMmBs9FtfhPZ8op/QlmQz2gpWHJMPn1V775YXX7w51OmgLunLe/lIGdt
SObsmTTFiFwTlLyKN3vbvwkGVwwg5sa4B1xypxK+/WzIq8i90cBu7UAsMGHByFjimGoldxwMbwiT
dejASfXnUEkYr4ofklSiu9Dl5Kp9tkL7p4Vmd1NfGFK6bPeYYIB8vA5rMH9OJWdXiaWi870gcTnh
hKHJfNNjErG7JYL4AEJDDTrFaSvol4Ey+NL3XvNb/DPlVOUQd4mxT2J5qRUmT8Wv7x8w5Wpltwz3
90sszwz7VcXKakbeTcLyT4/xy3acPFwYqvySdK7D5lmWwcbiO6c/tRUi3MCWNXcensdrv+3BRh1/
Fs9GD+AfwRo9cfX15+FUFG9uSMn4qUoJsGNsrlHTGyzM2drRNMu72LHjnCLjuyr7IElSk0UXPcQI
Wi4HIA4NlVLpMAw2bIQMrtwLcNW/iWAYN2AYHNElC717gZ9XL6nVzEa81uHUJ/KpvLQ5vXmrIZgD
c1scsIMjXYKhbEQhbnHPcvVYDCHslipW1sYl3tkYObd0cCJZ0+DfzRhPVMPvGD5H7rxL2nqIoPH6
yOhxs727rLNTOHCSnNYakhs/1zZvd6eWV1QQVQ39azqa/YyB/8nCGTk/kkXCRWNty7ouPu8N1ytW
YjEvU6sphtoG3uAVJb19fcPrsK26DQuEQ+N91JAfOusQiIOTSPmwlavx6reo9AM0L5nXBnypEEWd
DKRxFp35pfQZJRU/tS4EyDN+oiApqW5Pz0rbeQnDdZ/v4pUbiFt4jsjrt/znpaifmIXGVgpf3can
kwqJ4M78YBv3nNw3rtsVMjO/2zyMzClzX/UZBCw3g7mewss4+Gf9Nx8GG1bUCe52b5O0z5Y4GT8J
JbcRxCTjhmRMhLOCH+8R4ArBNtjKK48nzD0p+yn+GjkshaFdKHwXQuwSUE5u/ak6AXuBcRpcXyy+
8ZkFBT0L7WJsPbcoFlgLLVCCOydhpQPHBCMqKim/2maLpNLxc+SIiynK7R6IPh63gj++74WtcRuT
58kzvSxRChrLTYgqiApZLa65tJmBglfVuj8VMXF5QQoYJT+nuQgHQ3S1klgMUwYAJBsBHmyai26e
QhmGf5EGlck/xziw+Va1B64y7cUw8Cn9ZiDugwFQ8WbfsYwixP8bxnE0SIvRMr4lqBhHjzx9AuF/
Y2XGNBS3t4rzSWaoavzNAFZo5Ir305c3QF+oHhGXR33u1pneSR/TAD7nIsVBrxdQ6nA1LgwLS6CO
BFrTc2XSk58IRc3VN9AD2qO0dcQgaj38Aq7/w9bfopkfQqx0RTmnPYKFAYIn7fhmWCwUKxp3ZKEX
CZP7FPD0ucD7Jls2d93ZZRO/BIM6FXewp9ai95pTB1cPnYIjHKMhi1EiMYaA45E/cpUniNS5zVvp
GUDUmyHOMaCxV6U0nZMZgm9MqSWiQuatR2HhBIyiJoxAQr2XSCBs6aVofjTcXX6s/4SCQOO9JBPw
8ckzo3KvpvfixDIVPB51evKRbOeImryPQFwtVNNkvlJ2stiaF+o3ayBQHjnTT15uim2/Z/7b0O8T
wXBK548/xncwxqXX0IPNZyLMb/S4E2INXffQ9Op6CV6ln9RjHxYMBthW0k/2I9LDyQcSOMDIr/MF
434gRgwadtfWZ/I1lmLregYuCIxj4AuhD6fHxCC1+wfqKTjCX+7mlIWZ6BDamAhCN0UTWXbhl8dM
vvNdeEogBmVuUy3CES38X2POiJxyv1EUl6mYbMCBADGRVbezRe9ClQVAXteZB8nYk1PFk3NYNBWQ
h7+CYm8SqCr4UhRTcnAbGkUbMF5CXK6L7tPqFI9p2vL068/bvhLF3Zlxqm+I1wgoUleKLXtsJdTg
MO/Q2xZ6dK4Mthk9NhqPXuLFfFtBx9VGzI76kx/omsSn8RZTO/Hv3K/JMTb5gtOnnfXd3ZcZfrzi
I6WuyyZujnoZ9wEkEp1u6iWtxXDChWrkpb95olZqs0HxWYTxKZHOyRKCgFVxZnD/6pBDZPZUcz0G
MpqhtzEXV61TnpWmCBPu2tymy2giQbJJb8tYm7hFqrHDaZ6UTfh9U7jI2scBwwE+kHoYBg0o267f
OLOxeroiAN0p6uC4Pyznew/NPAeI7sfnOuVcs4uDzxGvjAL3cj1o99IRIG5misMPX5Fy1wIF+O3C
gOi7J619nKxDO4qO0LRNtksJx1glK/YkTWmbxMHZzEraZk+8fuCy6acBIJaDV7ofLHCcyuVDPJgv
vjS8CaHwe1Y50t9KWUH5pPQbg2JucU2bzYElwch+1TPd1WBSOcsVAo5BMkLj2AQmtPcWf7GhDqnz
1X+P0viPJ1IoYbDZzwNkKW5XxDKWEQPTmpXlHbvNg5ivkVWlAkk4/vHiWx6WHvRvDW9IGaxj8rBa
sfQWggL59I7pw0qxp0JFHgR0w+YxgAkZCdYezMBaRtMSd4X4OkT8gi8g23tsKz1GwYL1d4VHPIjg
WRr1dEiWo7WUGQThA2KyZwYV+Dpzc2fIYl5QfZYzsF87mfFTIROlReOV7klTn5hzYrka9uoFXavw
hcFhbHt3ipSER7eobgNIZ5l3POMLEobjDT8aFulV2Q/0wh5z6xcmrpl1BXRnoz59OThYEApOMxGq
PiBBna1l4FksJ8GA+xiS7jkqVINJYjmuIpfPqmlMdtLRT89Q+0g6z6f11RNz3d+MtmS8+8GdoOJ+
z/yd64gWIQcbi/h0qs/0czmoUZXu125CHEi1fnbMN7Qu9P3jTYgmsFxE0yv3zFUcq49Tui0KU1lt
0v8t3/WrSO+BSzkK/ye5dT74iki/rfqZed+6kkjB5ah2dIMgsLLuIMZ+ndszI0HARmnrZ1D9xmwK
/humJzhy5Zpm25kGh3LN59to2WJOXLFDHRUUa/iCmD07LPlF0FOd+emH2PEGMLlyN2ce6fvKwSf+
5E9U5yXDa398aDVkl6lnQf/nPJqHHWyHMo21lxOTvfIEf+1jBuRO0ORlXdedF1XBJcmDePK22sj2
5jFA6gw3X9xWiC90ChGofxGiRvCr5SyCe2uWTKWTwcFDBDDCaDMWuM7U8QHTMWOfMxDT89fjyyFQ
BI4NFmJo02eGbIJoItmwLROURzEy4fm7aPM5968P2dmM6KlyJee/uafCGyJ1r8Uu4n1xYU3ZSKfr
QgaEflgkRL5yGQMXdJKOWY87CDcrtb89j3qRKwUeeLKjUpy/xHZmpIxTGindVjeCU6UZjVjVGqWY
hCAbPw/DYWKnWDG+YQjORx+IeDoXCVlqdocFOf39wB2zl931PIoiK4SJsZM6CK0i6TF+WX+QNfGM
wQjdVTZncvssM9tVH/t59Xo8cDHYJwZvRJnMtjrIV6SbvKNVLhGju+1KwSM/BtFLJ+ijamCEMw9f
93E8bwDK0tjicO4UpztcqTlGd2D3Q7BGR3np4GlhPPf7hJ8/eYGRbcMHawCq42oNL7dJ8k4xaVOI
Q6BAA+/0yo43QW8n4x+pfWEpyqYLXV4BcXmNuJjD1I2jI16VKT3dr3bRThOcdrvQPHWzflQnEn78
3aL6tXIeYnaqyh3GIVZ4wo4UQIXoczedEQtWpXxqXJpibfm/V2h6vqzI8PzuGxI579Tr+PlboI5C
CN3YEnxSbtX5xkvA7vaaV4gijPhAHvgIERuzSMWIFJ9x0y/NwxhsWChx9xgIbbioKDSJo+udBPzd
HVxq7zZjj2KW6OQVySiItrO8MQZMASHiV6CLbM59WaBeigMlDML87oF4Y1BAq5EtRyFHiMuXE/V1
xBsC2TWSnB0Do4RY5WTw6KYCTMBRJznkCfxgDPRev9aciNtZSY5A5AbWjiac25rRK5uUzJcy8NrJ
mKH9uMhpuyZ3nFf4NTOwLdCz3qZq6qsJcRZ/5KMQp9XKOATxqWKcHyXWNbhimrddCvGCEW3nvf33
P+ciEW9SdyajnKfMa0cDBBoeySEeU/8XEVZ0y6XLWjHKr6lIzQenK2UamdCasijWpzxsEY6Zsd30
zWb32sFIQ2bCYvb3Mzr5/m8xpdpCTSWEei3bM+VULHxOCFjVAodh0Dev1k4weNzTnQb6lssiOcEH
u061gZkmexpW+5lXB+UmGqI2f1NbAJZAis26+xFbgLFneooMdlNa2a+ij+5xqbRk30VzFNkUJJgG
e9uS6n+jS93eMDwM4oCr76HwSuxa3FzTjZ/QrwSxEnhrRCvdc3v2FUnxuvp2oE3HP3Ni+jjpred9
5zOYdaw+Ct+L2K9gpCsQ/iSO/mtyz8SLFA+lYidEEjqUzfARVS1IUjdyLtOKE8SZSNKsZAJU7dIu
PA5yrX9D+GVLbp/RoTzuTSZc6ROA0Ded0BWK/ijtlNqKRqQ8JrUUP4yNTrdxURNodMnps47SajWT
zTU6qirlCTP7dTHZD+UQg9ZUg9TBh+NddvMpodqqS2zi8TgkwJ1lUkIYsT7iNTHKwXuzeEwyuzAy
epdY70rktA/XMjwMShqNTPqblvR01F7BG34waY8W4fvoSVl9S9wJtUeWKxOsUIvwsoaQrWDFThMp
aZf3of4rQrjvcC/y6lENQmsorkuNgXTCfZwCsOA9ASC1+P98DDJn10jD8MbbBluUnh9kcaO2xosa
YbKansnW8Is9qDeIxkvGTYd0frfXsUK4VTK9qDMDF9TCKWW8pp7re/UuKcvVP8MKVMbnbmRjr7WH
aly1Fmqq28BSeYdF5HQb1b6V6xevoqA4cnJHHI0eXRVIUWr0qum4nT4dqYkSAlHrN4mybXK9gboK
zWCgCLmlLtKiUlf8zRiykqy8J+AKdJcoWjk1J5HLi7802crU9KtNv4LggW2p/w+Tf9S0X9fqTIee
tlD63aSMc5KolTqQ5pgX0RfqFul9DhpmNezUeA2QNAau/tC+GEz+dwSVyVHwnres4FFgzxtyXzhx
qUsYYae2nb8bndiNJ1rjJZ/AMYg0NdQ4npAHw2bhtzJAdfDU6xa54/7EYWI3W/RtrutjQV5xos0P
uT7dED9cf+U4jel71n8N8F9b6XIVtHRSd73A/wkroQ/p/pfKKV+xay31cGAJml1sGUHfK0e2zQzT
gdum+vqDyI3TEZdbXTtd5MWFS6Gr1TU3G7GSsB91QAaqAvh0Gi+pe08y2bx0gWtuQ+bYjrogN4xt
8XWQwowsvqzE1Dr67dNWIhJOPjR3b2ml7yneUSplPVf69U6GAf711qGzqCRVW6feX35ynALCmXOR
c50XgKbp+p904W6xTxuni2GlzENGD+wWAHL1edgX3Dwv2HR8Yzdq/47VMj6ccoKN4jPuuboDLFva
QZslzso7vxke7xnsw9nXXI2b5s8V1hbk6bbYh+IETUMEWYjPDjK01vWtNLG+fMOpNdOcHbUdMSNe
tKBLBXWy48bRe9qlDMJLc1zmNxkc1vK0tShMEN0Ex7s4GMCtQNOY4ggkXKU8gGxAXVEHEpEcZM3l
Hxdt59lPG40+BhvtgXNmjevVcnOy9McFrmij5ml/kdDvXD5fEKck3cvWJKzP1eejkn/VGWULyFCs
AtoitiyJPDdKGWymNe/u/wBXD5K8b+N6OalIDbxnrPSA+u4nhddnSLMBj59gFcZagiAG2GYNWGSI
BSAw+2M4H9M6MlXqqU35PR8/QnK4LDRQCDbJDA08Thw00YCMZus0oSqPBVrgaGiyACg7sbPQ6mQb
yQHkrz+LA3f7Jtx5YLK0oxwD3EIvXtJ9OJg8scFsDQDHGvPAYohVUgs53G4zwS4wZ90p8x+k9FmK
g2NKDFfVGuhU5QtXG+EcachlLlRqkz5rDKaPxGJLz9PSmx/SqOO+TbgG62z/3UK4wWAod1s9bk9G
fExotAX3kS2Ddc+aIASUH323W7h24Qs026Xp8RiQTq+3GgQCvPTz8RVXhlWYjLWTujf8IAnidDz6
UzZVaIYoamNu3bNeWPI+GTfKG6T+BgF0VX/TzjyWastG7Un1ifKmHieD+a+qqzzgPKjeVQoDplRX
V53+KpvBn/PI9e4HMjMxxl30C1Zd4T+abTFiDHb7cYb6wIZFfrUwZGRKF0TuVg7JUvdGU8EEtuMr
O3rTSQBg1Pyk+RBrru1+FUA5SFF3G55iaHGfYEVjYlzXW6I6pSH0I2mCUyxw3WxChml8mIMTXd9w
lJQodqsoK9xRyK1u29T5sD96lzFYHWw8zJAos4EoCqeWpuuZwhEP/V2pRjvmKHDg4QbQ+o/UvsW7
iZWnJ77KGrmV/YlhhsLV4GoaEXn9/kG3oAywHGynbBmHthQG3DuCrUNOlxwwP7dop8c6qTKFJryM
O6/hi2h993nPQtEXQ9uvsfRuXuPcIH9KhW5h5FiY3fa7gkLHgB3vOxZe84WzUASh6ZRGUkwOPnqT
cu8D4R1JkDErONMdRlXL590cdNglj3V+nquEoAZkLA6RpXp+87OCdglDis2HYzvmFRBzMaFJ53pW
bkGvK+nVKrGbHRni3dJXDSObGhVY+ks6wsnWinKg/oDZm0JkxQGIxmu2gq3eSm4zGAmbyJc9yI/v
QxjeCyOlqMpZGzRsMfPquswkCWYl11UdiEPHnoeN/U4n2aXctb1wcVqPO281S4cSVC3JL8ymjPpl
EDIl71sMWxI7GsX70ylHuiPWJ0gz35eAhKy+SJ+YXhvk0koEGBT5WsPxuUSvxakThTBV6cd35L4h
pwYeDKoRtM2yLS0i4OeQ4MoJupC8QoMiR2B0+rrfpyqAnmgXTLTnsutWmd+SDgRWCBxqNYsDSz16
Yk39YOq33vwdjbQ8YRiLftfJ45DLu4YHDx730vP9ZMzjcb0EPz2fDdR3K6/9VPrASWnuFbDbaXa/
eCiy+hbFtsEIgFFS6KLMNzVcB1LNQ7E2vtzLa1JjHdFDxjiCcrSc8ADkMR+v02GERPsv2/zxqARx
ArU1bmzriCaJRn+Ydu3s+1orqPn50c6ZMBZl0zHUOjMp8bN+E4CoClxLxMWB7NzgF8qX0w53p8Jv
8zwy2UZ8tv0pczb0Fr5kWCpCp48Hds4Ma9fmON58DuZweqqv3oqcoy4uUmjHKBKMbbvvvm1shrNL
x96l+kpKl9LfisQ8NGx5P3KdMHoc/QXjZ2ojAAhc18kEP+/0FxaLIELiJgv8xfPtOtvV24Cw0grr
iUnkMjEEi5Ua/IW42wjvdRNN9wWHGpncmQbMFwZZMfKWH6JPA1HlXVksg9+9r5TYXyLLUDqPEycU
PYVEUAfvw9IYam3VimxMaI3bmh/+JJDED56yRY3ov9w2mAwJl8ZIze9EjISdK7tHiaIrv9k25reb
bcB1wputQ9E71eaJ1zEbBacaEsfgdtB8XTA4IAT+VutoiwJcc0MVgOqvrnynx6b3SX2KRRbQPaqw
qabGxVxn45mQvvTfJ0ATJqsngpODW1xRecXeGxKX2FDP26x9CdNrEi9P6872Gzss9tPdWuTZOTv3
gTNwZV22BMaiO4D3NZUhrGYtaHOq5rJkflahqljJHOcHg52hp4tmb2QpSjAtqQlc1LmLZuvDdsbm
69fDJPzXuuTFShzeR4xjhcUvdv+eOn3FLhGHStuq/Mk8xtdx0C12caOaPy3vlofo/BGgJt1TgFEy
+zECne0L4DFkoNryXKuiIe2ZAsj16ODYo8x2UbBYo/hYdN7H1n24f7znsSCHEqcPNf4Mqzmg+VlS
yCuulZ6kjHy/DCJZh1gWbF3CIPmQZjtVFXM/siplf1C1mFh4OowybrLFSMXMj5RPcGilo5w9F4yd
0I+qZimJvdF5fLvUPuijqkkPfGT82uhe3nFsREFJR61yQMrr2WhtfcEyfbKWA54URMu1Oul5l1+M
L0kOe2B4Gce36rAagVubgn1LwRc/+9KeyDnaWvaokz5ScTHo8VkVoOw1dubTWA3oBJSkLY/RDIG3
KI5+XM8la+L/2NB3kikkztmUVBsdaAMQHcEvgqcU7GeH48ZIi1Fo4PpB5+Asa38ISV5UawMF+A5K
vN8WWHqmfYIGocNl3UdT1wEPLEw48vA0Dh+qETqY2j/LNKj9z1Nq9EoG9fxid1rrq68iCM8yHxvt
81UR0aEGJoVZNGQA2lCE/LY8e+ALMFx0RZvSVCmTs1yz4xU2ojxS5LAhUE6PMkxl9CSFHHUxZUTz
9SpmTj36XRwg5/40o/haQ7zaBGLuo5OOXjAxMjduJOzjVJFBeNvgk7xTXYbr/1tTSUKL732dNWP2
SRQQEXZLtEpNR+I3ortjlHL2v6IV2ZLsIsZ8HmCHyc0BM69LvrSL6L7eoh6m2iYp6Fa0fDUQ6J4u
OFTrI0wHmfT7rZm6s/IhcnaKHwFeGJTsieghiYK3jGvfVdmWk4ReXsIrSMRROz7tf5QOdxFsL4Az
tdXwnDaCDpqAVV17GhJYPAKCZ5XmEFe48+y+FTcOERY8Lm4/NPzGw2rimqrB60zH/jlL82ffIRKz
+tij34VK8MA6Tua6pcXS2mRcFrECuzLRNX7lyrUms3RY8md6KPE054BUsI5nmDhVYd7Nz1Xx+JrW
jJcguufmqJdw4FFRiP1J6cJWhrMybCsMVaFkYBKPdu/eS2BYspZG5jt340ue8DP+xQ2JW+Jwdmtt
SV8VsZ1diLLqd7r7sBQgv27SbYTcal3f95+6cM1aXAP6MNlMNURdJvj8mHxraTAMTPaVqCU64KaW
KQUdqiCk6WREUVti0RXX84aiurzhxxmzrfI5PhYLHf8KTmDUMlNwSup2WTRLMyMIpd4ndGRUFXNq
HnY1AXtgRvFStBKhKUWg4tNVVeOU7lvT6T0ebcoIvJRc6XnrRH0HQqLxA1CpQoU6SYbpIk9iAWJK
CLlGsGUJZF367GIL0sHESU1XO0ouR6LOj+l8by4uUgn/mbDLsqNHcfY42RGvfj7KcrxvMvff0oKN
LirGVEa1x8iqvgKZu0H9122A/UU0PUVafZG73yrS0c0ZHpp4MymAcup+E0KXCrncq4MdIHFDcfdl
FM+PzopCJ8ZbjZj6YOc956u3armHbVqvmJUILqhxMtlkZLCcpQwN/EH3XH29oA3iQHyiejcGJ5l5
jYTYTA7wIWPbu6OWZVd8IWz4hsGqDUlvMMtfmrtmCxlEnoioBhU0sCBUnm8Vz7Or48FLhrgl2jiI
PFx5bs0bsPnlNuE/4tfGMBJsi6M/3KEKVdbXjtyrj/jXTEZGGwi3OXWqWH+QibRIsdJOvNjdApVK
cf5ubimrSYbM/LqVU5GdiufTN3Bna222Wp82MBcmFbKQE6oatwZSbymoDhZz0WSvFprRPFyFMXUk
/spO7NF+szqBuYM289ucygayUXdM4V2tuJ4QuiKPHrMesztvp6tapvoe9wE4BUlamiR9D6TFaDOD
1CCnezJxY3qg/yBK8EMPn7imSTtoHq/wrR+ftL70pOI/3rAXxgLEG1c4ADMeqxPTzE7q1YK1osBe
8whTsV6coyOHj6dQgv/rby51f2ZAoHJD4fpg3XYLm74wIzBVOR4GGVSgXtNkbgDZVZJxNC4PyS9d
gCZq5X6bHlyd5BMWQUvxUHeTkG92FbNdZKxcPxdC3CkJOO8IdguQUJoGpW7lBIOBzDWf3zPcarVD
2YOWCKyC9WyDewiw51JHrQXCwgw/r761Nm95ZDLrEgSNIm+pFAC5wlbmW8WxR37fccDTgDaE9c1J
b6rdV/AHWm2QoKMWlADTvnxa4LxYqQ4og24xB58+pMBOeuAvZeqmqo4u3ZGwrjAJm6asOyFDtYJW
6H30egBdXeRQVdL+KlVpCmcs92idNS+UWis0rIj2s16gibeHN6orH+dtcnZICPcAA2lYJnNLzLEd
XwLIVXf6BLJsoLI5g+whUFEz5PTQouNDEWu/IGg0rib2zlv3Z7GqjkhBe1sAweuMLt+NKsnUx8Jj
4wFD49ajBahqj0ykfc+r+KP1bhIdgnCoYJIAPxF94rBemVWOvJR4dPmQre/YcGToEpCdu/E0Slj1
SDctENHBAwGUTgpyc89jLzzTaVjiTwnRCbPNktyH607nL5sX1ASWeZcWaDW7pGDBMJio4/g2KH3M
gUSR9SLpqIRI1NASlFdLDMhdEPxUYVvRI/uOou+KXjK8+IO+76jwpYhD+bxTT/oWEbnDQRWR5GPB
3SzgiddvJSmej0/u1OCWSBzb2p0ErVT7DXi67MJMSZvXT/48gdXLG8DJNo94dymroNaJl6NpvSxJ
UtazskmrlFmsFdxf/GH+IvnFSI5OpCX841mvXU+Fz4D9pvGCFqIg5kgmwfXFGlpuWGXjvaz4J+LC
FzCYL2xp9crY8OaWHAt5wwKGtpZmOhRVCfMo6LOQZxv32NJ//zAnBpJeyIHkrB126azPy3U5Gd5h
aWPqNALHt5WIK3v76kVdrNprMzTxcVpEWB1O3VR1JBCLNfLVcvF2ZZwnwe+kydl3mwP5cXwuuSKG
ZSup1gQQnhdbdFDe6fBbZ5AUY4WmIkVBDQCVDFGFxrkNFRHa+v2zS1qBMBDar+hXTRMYV/jKstfb
YMgPchhpGJr6QHICxvh04P3Ms/SDWSFhDdQM6U+iAOBrfeL8M8e0U1XnZdtrtRbHZ8ymVB/Rq6RK
R3cfy8lMJpklTJhmG2Raw8cjszqpXCbKBtvXDXnWRGL2obZh2/1Vopz8R1hKxzHc+fFnKjpY7mZU
JlhG7ph0CggrYelyohK8HFpzJaHLnxqCEWZ3nAdeG1T3p5q/x0wRAM4uWaONHcHwIb2gbwG/6Yhu
4/T3ebYeNpokR+P7oxvjRkehR/jnCcGbDlRFY/KdZO2T3byakIbS7d00Uw1pItmoyJVM8q74KXHd
1a6PwbUreGvPxybO3c4EA5CLs/wQJ5Q5dEO75gF2In0vunVdbg6q8tGY010URPO2sh3S5CJLfNNb
JXGLrV9yFji055mjJ7XlAyTrQz2ZesULE1WBIwjJyzzrw4q1O6LTSC/ThKuvIjm0kstU8qQbAvxR
a7UNrUBY83+aXiZe1LE6PChQl1KhDhyHAg1w1/0EbZEKccM/ecEqNllC6hb+O8tQcCKhNs/sdNk2
pu8fclMqhxBMokuryb4PsLbuVk2BKP0eUeIlmED/L9fGw2R8Op+hNGa1DGKuNpoG0r3IeSZZWmBm
HltW2WcswOuMrQXInBsO743ePc7xWO6tTFTYuaABtLDMIOj0GG4/rv1M2LuGmktva3C/ItPPgj+4
Ovrj5GBsJa2pJPbSjZz8cDNq6mtaEP63raRUJbI5yN7iTnpjVEgPYiEYFbw121EPUxFekCf40Exb
VstToufk3nELGtFvOlxCSctd8R5U8WI53kbX/hFWTWrJobQyFPQbQhb0Js8h0JwB1nBNa+MP+wu7
B7YJvxlM5yIH2x1tL8PbshXHrb21yal7HnZXCPaY1wLNO1BQutNU0grT2qb/xZ59ZP8ZNC/nDgZs
ZxWSXhkIXl58iCibKX+OYgwrFupiry81rfw+gocbmKTUNTGQmPX/Zm7cDyITuJjCTyV5+DFaPpNO
XOPrMuZuuGO9TY9at/J9FBm2e1ShAN+Gkl3jVkwpTlPMFYLad4EEn1DCboKEKU8chc3SUovrtZvL
yQpgrDI6SzmfSarOsHRAx9oi5iMh8THhNYa74o194YYOjqOZsxjabHOaFqsUuqEVUuugsKlgEjof
3vB8bzmHCbwx9IrPb+8cSlNg/Iv2JMVSr0o465/CN8yM4CV5SDalrO2OuYLfTk4U5KPgWIQ8fobD
1B4josmaluj8FTsB6w0CrdhHPYTW9mZK1CQQrrG05E+tpldyawKdrLy1vwOA0M8OJMpMZqj7H2PT
cL/VJFiLFhXsBCEC+V2XUcJLoE7Ue4kDVYJYOsGlJg3ADw89XxUODy4YynoibzR8k4oyaxIFCq2H
7Qe84VRdYkEMJapCTMAOkK5txlePWU6pMg6Ilpf43WH+D6tk8VErQpjx9nIx0hSb4XEc2ZkJ7FtD
wZw7/TMgusPG94QyPpnvUP1g8j1quV7umCSA4/jgHRGnc134/MXl15Y6VOnrmtcgPIGnKJ5dtNSz
o+aYQuA3s3YqyROouXodByBC/b62otdqbv8QppQrNNJPDv4/mRi6Hm+E6HXprhAaChmqoxmCLsnG
VBTY/GvKYrkx81B/hPGx5L0vqU9A5iggQ+IEXbs1sWWR9SDnPf4UrPRAGzhdu8FOGhIa4k6KIsCP
4CbBg+Hqto3Xm4DM1DVlLKiyyhnstJA820byzGKJGq094yy3XEcz/QQVF2jRMHJtz//MFaeZ7KGp
Wa7TqfRmmc5+kgAhlZ+pGsBva622yJyQwUa7nfGbjWZNHIAszW6UkZ4rf3RdRu7jAFCxJjPsGn0e
zW4ENUxUwqNlJm7v03E0Upr2PO1fmnPIoIJHdGQrFnOB+/nak5Jy3rlAOrMxMMiTwX4csqH6M52S
vYhxjx8jMs47K2Rpai/GxzieKs87SudP7p532xmZTGktrH+fK9bKFsHqCA3jqwyXUtQpVIMv0uv3
9z7UlXk6kxe1O6NUjVlf98ji6QLyxsZW6Ud+hRzHqb+hGKvO8XaD0RSwttKd2oLUPeL4dCychhqg
DKGdD4DR4uwIX4jC9CWXHbXH5mM+yoBP/kkcqmYvTxlA9Yrbf//C8NnfQCZGxoQk2CdvBklV+mCz
XyPLcvY37VWl1CJtJEa/5dAzKZVQ/UK4phVhbaQDIp6QqlZDKBG92CFw8N/ynWSCKPDgqOt5NPNw
vEy9NBFS/dsOGj+Hld7aMPcPNiRsqG4RhEjqmTDtp6SkSwl1XLQ4q1QBstnBlv+etvJ+JgGu9xG3
01OIbhk7ttNh4t/iruAllTQcwqjwVm4KWxzgeIWVjAqUDIF00gJsk+ccnoVZxmWf+UlZd+PYei8u
iJa4yP9pSff/We9JqbmWbHkpLoKhjQUxTIxhB1MhsCtLMOb9yHLizRpWEK5MUlgyowD8qXHmt+LM
G/0m5wOHoWqLJh3sxfMjCRYpEdYX8EAnF4hPXv8n+2RQZddQV90hx4vrz37cbwuB3Opovur5tE1r
Kbjp6OblpQ7TnHHYVi2h4zIfoifcb083d/WDAWmrDMep5GAFphafUf7XXsZMv33PSWazda4xrQP3
WXN00z2PTF75fiweNJeeno/Jnj8tfo6aJXRMdF13pF4gBoibhW2bD0wC2IvnGwfBbQ4/98Ucs/nk
LUtG9gjQcc4Ji3ZZizbg1XTP7AwU7Emrn5a0QtETeU3eN6emA0ly0rAOBR0cSO9s0MVpPGYrUBYn
wFvvAMTqQFRdhye13YNSoL1myNUiIz+qEu5VyxHUZdFlUOFmwIWI6a2lokYcQNNPC561zAsJXxvH
+KD5jyfIS3hdU9o30NE712evlei/pHj9eH1NMUhAb8vhmKi48n1aV8To4DC2H6NMdDwgvPNGg+hV
+XCM30ObZz/Jb1DWn4QM+mAMhkK845mFxcHN0YjFuLRdE5OXPZ8k157rOOo9L9VqoVHDG5zKoe2k
DphwNKIWlrPsv81eczJs/qmv/qIxMhfrBByf0ucgrhK5XW0qjEHL2UtE3VfXCjzrMVTI7mXVyrTM
dSgEFafDVC1xQGSvEcT80W/io6OoHpMgfleSJ1D+SVM+bfHCtstdpu6k6WbzIfgNEbMWTIpSqbvg
/cU7DR2ZdIG3nztn5FiCSpyAn1LHYPe+mj/mHPcafs/rHjEz5qWB/+cjvuiaeiaf1A/GuMcP8He4
S6jyQdRi7xuZ7Nw88Po6Uo1t+Qw9rKr52nNeXq/ZMiCv1bRC2yTtK3czWS4dgBs2YJnCZmXtoSrE
PM2NGgL8L/a3ckbxsEL8kp+9wB1AMUVhy7VxV8lDhJsB2D8+9o4UN6iNp0REAwy5d4ToBSg4kjP4
/X0h6niRdmGiiUpx5iMaFs7u0+Nb+d/EV+7RLRuILgJtT42u9pXQgiiDM5hDCSg5RUmIDZTnQ0NT
vXe6fHF8VLKOGd5Hg0AkqFpr6lo70JZuJ7NzNv/pEEM16ILWRx/iA2pcxiL10BJTSBJsb9mmMWzo
vlN4d+35mVB3eX2hYoJzr0X8HbeBmPClY57SyovyR3PvnL6raTwz1MprW+ozDax0NvRH4jUmkRh/
j1WhKOTQITCHe86dZeiamyictWq0Qpn4qTYcGiSwITnw7RCG2H7oPvZKtjBmS5/8mB2++DsZjDfu
zJBGji9LSKHKmGYOeGu7Fz+pXe5jb4wCOUgn3Mqi5okL2FjTSOPgTocS8F1Nc+DqZmRVDz3Jh4Q1
xZN2K1BQu1maV6IDL5I9Z8wyMp+amppJ/9nAArvYYZL1kDzkshI/e0vExbtlevYWIUvow6J/iRTa
elAP8zNLBnu2bgFb3TG3EzcXfI442GmUY9ZxrnAqx3eRPr0/N4+SuUDRjzDQz3oixx9BFqfIi9vL
7gsY+MVpqLzZdgr7McvafcyFSNypcg/VrSrDMxSyoNIINbPcK1hJVPcUK31S2dbKrBZWLMS3fGqd
qFEFWNnlfj1RuDTV4mvEHCeFuehD7EhVOYyafXs7eUWsA+lsoFziZ7WfEHowvmaSlWioqED+nUhk
8YyXyVPo7VGNsOrJ1xEI0ja8qJrAUcZxF8QlwjwfXFHuhkUD+XtdVVMmFd44+t8QJqtutZW7Smn3
iiX1y37vYVb45C1HIYC/gcJCb7DHNEIzL0cTagH3KvrN0GEkH9H7j/CcWPEoX3KqSJ+E9E10f9DY
qxEWMHJTAw2wpW7bwPHt/rO6cyX9SvqA/p6ebqxQJ33lu+KIkor1ZDrh7TCrl2LkI5ggjf//lyUP
x9ugHKqjl9j4P4eNB7kHRh7Ns+g0B/t7tTEGbN3knFYw4qi2zdABWYlAp2FbDMp9f3rqXB4AoaAV
SCOCes6H54/5HD+KXaVJsAgppYrrUvAUN3YBTX45Zd8kANDwn12DnFf6pk/VQeeVeZA3jl2e7Fki
4QIaGGlHhonLbGBeOXGLRJqq6C6PDjcin2Yh7tpU7z97dqpINdUaVcc2QxI/sojFtm/niFi60Cep
GyPim8ll5azpqYb1mPpRjNdOvCMcpmr5xLrUjF6ToPw1uy+HCdtAtlVof51ISwlvpQdv1nFpbS3h
Wim7fh1eNGXuyE8gJ0tQrDNkpEEoyFCazvar9anxAUUCcU49jNUhgKsHIJTHzT6J0cZMfARHxSMd
qHRMMgxFx1uBGnQmHIodW4Wn0i564wmIQq62G2hPpWTA2kxDjKXAKxEDATUHZ9a2jgNR+Y5Lfq8X
PGBMX3R/U1anOmPP+EWEUSVxvoFZhqjSMBYoCQhMT+aJVLWxra8RqzBTCvdM1QyR4VTlWu97gfPi
6sRMa8XEG8bfKPG5xmQeIU4LQN7zufk4xWs2C0P83jmUXeodPeVd7mxPunn2j6miil9IcokRdoD4
2gkULM70YwUC6S44qn+B76zraL6XTHhn2LzYbmNIcwZVguO/dXtEwERz9HMXME0FAZMgw1Y9HMW5
0nexF581vxASrKgOtVJn08TOO45IxJ8PdCyLV5arM33HlC1EYEh69JxPQhY3uAs9Fx4Iq3TWsaaM
s1cDN3vMuEn7EKb9UDHpq78IDu+Zm7zQjYzFhtFn+PlwDkOgE8IfTIQnE5zIZKXEtuXr+dqA67/r
cJZo/i85ZXWSO40oIqzmMYlXvH5il9ZmmWxPS37ws61yy1SiP3uqDGOgOGgaYRhqMR7t6QZ7jj4G
2u1ajJwcIk9qseIZqxlIgQXt7mNO6eaAIXn8NYl5dY6RnpmS8qRdBf2O82mCGIs5GkRLr4jgifaN
jjIbRcEV8YStezuiWcW8oTvv9Raj003BpIINA+yDmVvjZcYCcWFYeZVC+TuQXM1jfZpX5FI0NJWK
LKYmg5OhrSwcNPdKr43ZDhHX6zEMDEGqpVrNJCWYTW964hEFvcgR1XSfEdBth5lHp6zdbDTzqSzG
8U91ToHVS0EtClmmMGUutPp42UHggyT1YXRJjGNZUhuCF37FifgiU7/G1MTNN24vnaeGnTpFwRfV
RW5CKYRPKUypDCvh1vPkK5770VO/fGqPrTzF9zqkX3FookRQ2arKUaTacbB18I4qvwbyDb3mNwdo
FwBtO5TJ72IkmHOfYHdUGc95QjtWahTBUdXMcU8dtr/2UIC39qdcUcGY6eZ1rPJJO/TXlaw40V04
tCD0jxUnqPQ46nb0qPPPCuia7CSKDH+hZ8P/2/SDDG1IbxNiiGgMfSqEybHtOSRE5pm4yyOlzp3X
RouIQepLWz0QqKm4pSbVAIX3lEbUTBjYQ2S0eeKtPyn6tgv7HquNHHAfnu/E2/+NHAUFIrR0P8Xe
ieRMiRFnDMAgilUDXoxcgldKNZnso3BJDMUnAiy3A5o/Zvz5dYYBNCE4zhN67vlALuoS2RufcWxb
idEFD4dI9VrMIdyHMU/ytTFTBGMIOYo2/mZnXHXlDUQqGZk13c1uGwDq3afktMXD0S4Jg7KqMnPV
g6TNI0cf75U6Fno9UEmTIfo3G1cnGdmWIpd7M+pX9YsuCn8JdhQNVLftJ9/n40VNPDSZaB7AEnx+
T/evT66X2tKAYwVSRZBonQ48DVGcqlOQAhwbrW5P2hIBKkvoXQs6rj93M8zsEO6t2giRJ9jw0EkI
W1uH+kBNbC3Po6gwQphjLpjOUYpFY9ryLEdcRLHeJY+orkIy8gi64EguOE7rbliVCQuzkEDTHMBG
6sMkqLo/GFSsVeFQxvrHdyXVJE0WeYyITFbwlepBNuiAklqKd/NUEBUoa92YnoKQkLC88omdvItV
wWDNkWwK8ot2Vb92gyaFijzsw7WqinQWT/SOaO9o7BTEEE9NVAYGdDMdXMI6G4eX0CBTL2IRyS50
xQHs0p5mcsoqjSTJNdYl3NdwU0VJC5DCP/9FGazpvSErubOtJVKqA/cATyKNoOqv2UrSXHY9Rls3
nZk21s0L602FZJJgzH1vWXO5H27y4M95CuBmdzosSHbwaUefNJnu/lYdDi/VHTLIrGliT7vh3wZ9
6tSeE7HiTVoqHvX2Ay11hf8vgt9LmTCyu/7rrH9nIoAHKvQ5x0NY36D5KNsV6fbaKH3YoJu2bWmt
s37usJsYAhVHwoJXf7e1dhG8HhCzbJIi39dQrXacHLbqWnxqwA67pxZIdsLYARdZKRWk4A3i2BJQ
QhTec9xAN2QMHg7mhQhwdR4BgqtDYenLWLAhGCCorRr7KGt51TwEVM86hrsybll6usx4QZJO8QVV
NyqX4BWzRUN84Dfp6Sc7txSI3QdrCbr9wuF8XOUzLzVfvAluSGykk0ecZ37kSPmiGWCny4jw3vuc
g61mMlHUMNcsFsCa0/Mba6tX2JgMEyYeGH7NcRxxpjg5h/6j1Rp3R2sjbAOvxohBTCbTUKOZjAWe
k2VlCjRM5apuzhAcX33gb7rg1EB/Axtm7zl03tGYzb4GsrmMH6lPCrFPKYUwbiDQNVG6vBusFatp
EUds/Ij1AM/9WM332wyk7myJAmvjqpfGh/wyryf4j5/p/qy2hQuUdzs6N0aUiiqv9cprKvbiSWkZ
QK7fqd8YtrrxPu2EfkTUheLvkNtzDNnM2pBEdUG3EJA2QSkpDRuIj+VfGGq8N7LbYmJsl87DHd+n
LO3VFYP7/09KJ57A1TvA4mqz02JuPQR9mn5y+wppVac1lZKC183EIkUvg7kyihRSeLpet/3X+WoY
28DVXUawH2cfUtvgWzxUSBc/I5PL3Eu09gT36/AnBpGHnm/OS2nTxPuc6Z+ytYzxdpfWJPlIxoK1
OCMIFHyjENl7r0Besgn7GDkyJVOMmqW7p+udzUSIo8+QEb8l/v4bXYB8sLWPi6TSlZF2cGxYVb1O
xbwzzHej7iXycIMgJZNVXdNnxn6YxNwuX3zxgJpnndNBB3qbFa+nWQjb3yugI4+o+ofWbGfVrJ1r
OX7/5E7/3ktG5h9xa1CP6lNjROIw24GdPXiuDaM0VN7xLy0kmWmZleLstJYqqzUo1w89dIR9MN5A
mpMXkCjtnDiJlP9bJMSleb8ofYXrH5bPqfFPIVlOy3SGPdhwjG7O4hpO5Yti51OzHCZE13zRBEQE
s9a5SvaVzgAUDn/nQcmfgi3DYtFPkBjU77WcECUoGCUWv7rtPoHcIPkyT7Zb0po7LkFTGwD9gF8O
IN7kE7tLr/UXmgg9nJTrCGSsyx+6T0UEDbB5wN3gqpyrRm8nFg589A+1U/58p7xr8kFKumWWLTO8
izmAmlOVr2xdsFGvG46dLLjRZPVYBG/T42+ChhmzdOC6l8fag+OcNt7P/mYJw4ADYVVNDHBORBd+
PDxtfMKzpOxlh6Vgd5Ufjn5yQJLf5EroEBR1YbQh/B8viKNe8WOm61eKBjiaoytgTh7UDXY1JD5l
u+Tty0LYl8U8ahNiXleHssmm68NzolpcC5QTICSNCUelDNuRi4I1NrMT7aJKTRrOzReQ0nLJuPD7
YXP4JYNAgdhStCo/pjGblmC2zahxQ2Qg+SfbjsMXd28WhnUgEoQY7oZPMbHWB5Y37ZbFGJlXwnMe
9DpUuLT4a/wpaHQIy1Bg6Mwps6fpbNYsraN28WUAiTuhr0wJaxNumZBwQg7eC6Ikj/67AKTklGQb
Avt+BC30PLZbPyZMJMSlxiLAlJHGkjpJC3ApcZaDYvqIg0Vi7Zrs3diOPwBVtM4TZ7+ytu0E7Qog
XftiYTOeNUzfe12x55cTQIw9TL0GQz72gqTTo3bcuq4okiFxRo87j9LzYBT7Z/aGY0ELBPd+2rRa
/kIQyBCOCW789hfcNvLDn77cDy41+Fj2HcbBRaBITsxSp7863ASRt7K49/R8gJnCKox7cyznxYkP
R/LClPz2B+sSeJPX1HlR0mj7bo/JFRSOsbwD28lGT5ybUOJ+tXpq8wFTe4xtoRZ4MRYDy8mP2KJs
UDB1zUDHq4bS5Ays2fa2XrQ2Mqj9GAHZDgTEMI4s0w4eaMqQwT+Cmj6ZkIny3/j0eNXlKYs0cq2O
zq8b1vWew5Twp9baCkP3Wc+ehqar+Do5TwKL8qwZ4e0WzQLGHzq8pgrD/BpGX62DFuv995Gll64w
RhPmF+p1xykC6mwvXS8eVc7i+vIZiHrWxMvwpgcdYLMOsAcDWeOueO7hk9JXIoLAx+g7hMrV3Qo7
+FyTn7mxbqN0tYGyATYrCktHLceC8A2JNYf353b19Mu+wM3VKpZ/pd7wHemhxriz1sHx2K9C9MrQ
EYfTFKUlkrcenF3/jzYeviMFnZeY18RgOQ6PlTg7JWcN81TKsn3KAaxRFafkNC8ZZIsH4tVKjppk
+Em/msnfifMPXcVqo+VW7uYXutQh2rpWS9S5ecuTRymjc4H9a92Ogsqsi4Dwp8kwf6OzdIrVDRfs
czDG3fLJzCL/ajk9yAhlrAdlPq1cVxk5WnKYFAVogE29z9LuCjmBJGAxUag5M1QUNbQ/uDrVh6Nm
pUijSyAlCrQe/jKbHa0NlcZNZ6sUkOYGa37MDtKeZqA5rob7U8IJGNR3qXQIj88LT8Ny4i4fpU9U
Y/N8nxm2cOrOpJyWdQ9v7cHiiyKwX0yHxHThUqutXTR2Ca7ZBMCFRtnsPkzAHEgmh0J9WKhRz8t2
Q2jDipftLFCoJjwPRDLxHP+dF2vo/KUtvUiHUwZ7oLb0iq+pFDqcTWGg8+QLkohbLMisruyrcNt9
BasyTC5PJPyIFaheXIoOI++pNBTmB7Qk7C/9/CkOGVAl2narvNOZnPJm9ysQojgnJUpCF8h31XI1
rUFjuttZqJxh8hPF7mHkpY72xVLQoTO2+Sxa6tVYdxdoxvETZlDNdnOrxRVTaWHguOwv/V410rtH
CI4xyMsYGu034WTKklpJgjw1VJb4TLXyJlKyuhVKW1z4UqChIYowxJMZqRd8UjioBKrIg1P+NSqS
8bh9SZTT5pxH76nTr/vAlREp19FQbW9HrXbtzjK/npqzm/dOSNeeqqhv8wOW/juZ9zG+hkORUq5a
mt3KK4ZyAp2LCt7wtqlNoXDDjw4jS7XbxNo0vU9ymf8UoCsHT5PXjTPKnvC1zOzKvIIiE87BBcW7
So+MJuSfsl21bk9j0Am3keaC+JJGW+2Bd5xIPbiJgQGS6rM4jbpzSULHKn4XDJ8we27zd0u1vVT9
YuaXffvtvq5yHAD91SVIrleYGyIr6zxtrSPeJTF66/trSUHEELpdBM5lqRKu/H+7qBi8fBlvzTPa
1s7Bwv2u9USfsXPKrvRQAxSQKwxwpKSk8IS4L5zMdKjMv2l6k7yGTrANA00wEzbuVPZ0OQV6kx5v
sfy5C3qd6lA32OzSeYFCnPrR04HtgHpceLUMhTLZLljLMj7qfdhJMY0VaINygepMSEc9oVHWwouz
ZNKkV/eFZ31lOpGRYdh5dZ5hKHlx1wU0gluaaxYpSCgBrv1ZZzK8cGaQLuCatEvE3S7jlac6iDEq
HoJG2oF4+Ncr2kXY41Loxor8Oi3bOzZYoP+uaZXbEyOIdKhfkavkRs5ANuWraX2qY7gzzDXPEPtR
L7+6BFRbWkK10SAdcxKiTvjR7Q64IBshrgEg9lY0UdeM/nML8Uk68nd07rpm2Whzeq4w/db8IeKX
GrzR9Pf5i6InlwlwH0U+S/mH39OgK5fxABhCN9jkg0aCPTiDErV5txIYcNEtNk3M6IVXB19czzpx
YqA0OgrjLHAsqkASTqVjRcMJ1QSW6qztx49K1iPo1zjJf29EqKQWoSBO+zRyP5883UEbINafn1iU
vaaUe16f/7NH84GKFrWFvsKRZxQs7Z7ykSOFahA2aviREdthmaKbHrIgzwJIscrz9AExxt3IkUkr
7MyePse+jaxPVAxVK5gK1Dv7Oo4KrD10sevOCFbpavK3tjLGwhq+q9BcOywVKlfip5HxyFA8JlDZ
d/Q73twghLQSlJxoaOKP7j/vLK9CqqjpB9Cbqi4uswSFNQ9cT7Bfr6t8TIPiZfadDGkiZP59Uvy+
AMPGBL77wYzJdedxjhxmNZuZMVF8mVOFuCP06G9xbS5OdhPzDxyfRlBy4WTP5zmHNAMSIVuPZ2Lt
0XXRJcfghj9b64Vl+Q8X7nFXrhWPVdXFkRzH7o+HwFeUGXioojiQEmJOl9c/INgBrDgqv531MWBO
tb8mjlrZ+Xo0GXZz8uK0WO0A4g1yIOe8YVULdGFl/3uJaeNcLwcjhUrezkF0u9KVauvGQmRp6LPS
POJRovNdcf0b3SGCp8hVb9ND/VO9UtI+bCGAPEIKZCZUPuO10EdwLgROHg+RtBEnCer3YsDUNWNL
ariqBJHqUsi/smY6hM3x/1s7AMeA8Q5uLbw5RgHjymj1kcd/25QFvK56A2zm9e7hx66imvFm4b/W
ttSZRPM/tgxBQeS5UJTRpX6VwYrNwdjHJ2DzRlAY3yDIQK15Z/u7lecEsVSHXQOQWXfbKNrkI5Rb
wXE2XoojkoBlNcBd74u22bVRMoKbnZRgMSZH7jGXdsr1+xZRYiKvwmhLk1H5AvHiD7bb4xP0VV0v
uS7uHODpQXwfZYQnz5rPd6sdT8iAINP8WsC7QSZzceYMBHVHmFgAX5+qcG1gD4CPnRpNyqAr+Huj
rvhIs6wu8pMn2PWMMx8E6zaPK9nKBD0JehcPzNrVwerEtAGPMi/4QepvHYnURXEGgKCPP+JeCGTp
jGKnJ9hk4ENqfhnG9EthwsbuDrn2MSAh/S1OGkRyvtlCMTU3iLdYFSJ7fz84qrrTAiQzKQRmomfK
UJhaPIHNUkJgTtWrUyu46bZwDzzKnWH8H5zPKS93wPuw82dr3eldjIjGsFWCAEj9nB12Je7MAKhk
KIprwaays4dQDQQ1/kgmYmc6Ie/sRLGFvpy74npH1SMJ6LLP77cgEPuGl8CTNC0fpC7umXFC5YEn
EeCGsMbAGW+Z+5oVh3acLzakz4rFP/wB25N4m8B7zGb7fuCEkITRGz1KfI9Is65Q8liZeTPkIoAS
/2PkzRNtqhxo+NCXQqoWNLrF9j5kOLaLKy03xwz5gqyfNbmoiQLelWaqk86gA64XWrA57OnnAcib
8vDjI+gX973k1DJELdZKZx3Lsfo2KoMygDmaEjRrkkZFsEWxyF7niyfVt/FimzKDvZ3eLZwsQnrH
5u5tjCeKd/CNbiSEPU6P8KlVDQTyuLp7f6PVEnMZiSWLqQ7vJIMOk16tx1nTNWBoRme+nYiCmc/a
UbiWDHsbRClbT84WgryEDGLaSf2+zIM3eKcy7hfGkTTzW7vUD0G3dAxbLyPuW0poa9+lfycvreAq
vfvvAcoD7C3jg1AbH+B20qnscuSeEox48eHR0TqArFprSz/l/8mfmqEbpNX5/xLFhY+a9MhyZlP5
AaEAQvNcxJ47igzDLWFVxeFgBgxOAz/ablN6viv6J+XXgVO5QDCeV2qEHeja/mrynJKDnAJjz7VC
b0v8Yx0h881bZ5XNYrdgo7zIIEZHBYfevUxnUno5sOASgyeLArkAEe50dArayizEO2Mz0JFeW8qr
Nxih9xAfFIqlLT4sw/mRkcPmVGGQmdM5VYSEV/M8gH1kFS0Mwx1Js/JQuno6GQ+hQ+WrmhCz3dCC
Aj+2w5mhLTlCjX/5Ezo87qLVghJrUHBDrHYvw04Ti5KMFuTm+X0PSOtQSYfotulrWXL3erMNz+qd
ohXpWBAqbRPbGUxhNgF26OSmJw9dpV011q3ig/WlW93c5uAobLlar4ibZQXKWiqxDIqJfVlZB1hz
F5CY7OxvJOvYGdWX01yGNjWyigqvbWw1PAR745PWG2DgTDV+sI7SAZFkEJvobmN4Y9F6ic9nAoXf
WoMoQgQq1LCToqJiEcbkwYkXlzdgVVHHl84tSirPkHrt3QwluDG36QFllq4zfT6beNxA6B8LwdVo
cgDegJUynhqL99XDRKEvChKSjL3xlCEM0is/wO5a+K1n29hpKucGp2mqP+pSESPLt3PaqJrF9kQ5
v1vYSpJkTMeP1bhlY+mdd/oPG3hcTcCJrECbMgs4kDxEDHwgM/9xa4Uq0UdXx0vf0v/MncNHwLSN
Gy+o/uCD/5159A3yWJjKS/hgMSNYe12RzkCEcGv6Eqti6dRkh1+kpTVNSMuBwfORuM5IbKa0HL+H
8LiGjdMYlN041TTwmdIODp4MVNDy6G9VdDLODxAlddKavo7gOj0w7Yr9rbV8BhA78D40DYTa9tv5
Ab38yetOdQ/43hi6TpLU5Q/WDdlwPU6lFRpOylGRjLMk0YmbVPfCrOjnUjb7E4dD1t2qFI6lLUts
BZa1ioNEfcJqvb8a7d4BrVfqawpGws6efDhae7jX0fXVRGA2dOFZLzlYElGDZtoavlPrHiT2aQsU
FVr2suq9uFuR4LSTsUqlPiMTQcwYFMM1uxhMHnbzIu4P0iwtWlUr7zsmay1b7WMZsC2qkN3R06mW
LiimpDWPfvCIDkDvxTwRQJfRjCSQSyOzyXbaL1HDIlSgf1y6yamt721tj8yqSCcid0Dj4W5BioKk
LxvOSUQL0Kd+Xz0D9iNSpx97/JBGL2myg3mgi4mbailgKGsFz0dVo8lRiGrHgQ3NeMUA0XLEJcX1
DLPcH3x6MphwYtOiI+cVqNtv+AM+ZCNM3Yr8Ks4ftG75QQB+z5QY5QmkQM+4LdNoUKwt5Z9HstWn
HYEKl6u/wssKb1N/ssTT70mauC1AYHQ23FbmX5fGx0LRLsesR4mF28TgbF6ILfywN6NO16XRpCJr
WCAzvPoLDgICQr9f/4mUuZn+vm942zd3ksMRvEgmSePlM9dYMwGY+hYgd1ZvxxjpmaZSUPIW3lpb
vNpD5A9cJlcD9t8/Q4MQpOnuOVosZjPY9uNYCqTiUU0oeTPEeuELAEEnoO32J8dS3eBKkABQF/l8
rgsuxpOCB/Dwje4M++e44CBxM66I8WCg56RZd+VgY9hnVZ68WdcRiRQhOzltuSy2wYTTj9qqjg/z
IlegdIKxkbaY22gAC/WlX8Uh9nb/64byxJN13Ojd3o3lPd7hDlm3QDDNzdUJLZE1GlPi0kSrjZeo
mnyDzevOBDxokn+AzlQpQC5lIUabDZEM7PkWKD2CYpXHUPKUBr9PcDE+9X7CSzAV0zRPRYaWEn7w
+8maoezlwQ1IJV3mAWtRoLJNEm3msXL7ToSfVu1Lm0WFLt+EDeIhNZ67egQFjIps0OumNiNbBsEY
pZRic0aoxEp/n01cFvMV9pva2t/kxb0pQYZY7bpmEMocYFnMGblCRpuUyg5MqRmZyvXqRcpo6C46
2T0VpiXT5diEAtyq86xEbEenBBJocdSawwX8Z0mw/vyh0zW4O1dnvCzjz2gM7frvhegqEhY9wc6R
0hjo0A9+Do8aGW5ZByPmQtHOLU6VPJnTNGQlR9YU1J8+Xl5PVrUO7ughRClGhAKxsciVdi3ZySTX
X9l/Efoyc2o6BCYUHsBvOrIjhBhcnRPKk4uAEk6zfISIjpjWPfyjMtsCXVbQZg308dDl24Aa5r6e
TP/v3V6+tvF5mMakTtAHco/rPlqb9V10Nn5OSmLyYydXfgzXDSSLZf0pVh7YKFG0r+t8anLj0rh1
2CM4rY4dDKK/rlog9xjSV69pUnIm4XCAM0rhSBio5tuQpBtd+hmLYCDnD8VXMesH4kDaVIDGHYET
3OVvfZYYelmew1WZqPpUDC9pLcKvhvZOUI0ssVv2THVJK0Zp4pj0khxKbbpV83qH/8HHN/QHSTm7
H2nBsJckV1qv8bpvhQOF79qXefVxffx2nvTvDjS+kCquEcXSMayVcdw/dWT3oWollqsmjVdoqwIB
tg6v2Zkjdu9rc7r2PH5Xa3kEmZuc8beaJPFfPzxnlFZaBMjNiQkM9ITh++4wKx8RvNFrmlIFHNKu
AGDbIwsycUNL8PZFQY4TIWypnx2uVQ/HuoAxG2YYo/uHIysRYCUTjpjCE3InLRu7DcqeWXGslmHB
6lmyRGdtlXn5TX5ochUmuQsMGvkwAnaP3dAktMs0w8vDJkCZ30GJj08Zo14Vwz5INfSSWTYlqEq0
LOd/r5cmgTQl9Sz6tuX7rLrTmi4CuSlAMizcw8QPGrcHqLeOKg/E4E+iWAD1cwZLEuQW12tEkIgB
elAsua9m9O9ZE2birzhOUUyRh0ihuEKci4+8RpY5meeZs3Wo7NjPInUF8gTFmd2y8AmvbWPpGIUK
qvPWeXzjRY4IW2B1KHyytnKvh1YMZLwlQG0AIJ9Cq1S8AcUiJrcdIuHdJO1vdpte8YMxHj97WER5
kLCtZRSXh+mHf3uAGnf04RSUfGagpsYKSBcX0V6vWxdUPjWY4jDAMlwDO8iz8EYRkScahFIJNOan
PYwgJlU+0wCs22MhK6XCZbNk1UF1s8n8N2X/dus0Xfaz+I75nYF95SgujluV1rwiFMPsC6ym5/KL
CpzkStmwOJLykWZ5TA6+yCLWEMKGWe1Dq0r84SR9/p1WCCXKu0D8MBirducZ0f7IV9HR2MBblwJ0
Qimxrh9xaFb6msxRIZkvReiXo7mqNu7y48oinpvfjR29NSxl2O8XJ/OcNzQRrr8eIoZcJmRQGzDd
ZWjWwpKD8H/9wsKPPBuB57pUk77i91hMJ4Nkj/RgqTKkgypxg6MGQ03bFYcz3zEfCGdaEd+Unr9E
Ak1wbqoMqlO2N/VQPW24B2nYqGYeGKbW6fqHbg1SQFK2bYyipn1YxIPJU+MBpUPQwaKFGEqde+l0
tz3y5klxJ+cx3rQLCoGfxDYOZwiqwWhiYdAS3l5OFOlyChicVkI+iv6S46hBHtowrANQqZanZsCj
P6jGU1a/nibPjZ5H4ZU0wp/K998h+qddTSHaqg7MCuRPueaxEAnkyYT3CjpmuWsPa4jqtFJKi98j
4pXASVJ64N9D/M8hErEFMjtlwJt+J5IulMvmiLG9rV/mhLgNU90HtINtoIjgNpd4V8zsgvmlfOkf
iNVpJkmlIdXOH4UWEmWE5O84L2LzzsE8ceJY5tXkOiyVdTt8/NIn2ahHWoLCBbz0lBBdVsbWJtD6
2nLwxVQ3jnwr8RECbt54gpxvCmVgbvQE3kmmE7yYkvfqnaKkS+l3Gt6VoAfcYLiICxAasjW6apIW
oecO7FuUrkM88vvZa1P/r+O35OliOs6TDQ72QICn4cvHkJkOfOiIvGigw4vteyaY8BW3jF6ftDfI
cu9WyhlCE360cVImcqwv5eiCXxoaHeSJdKhJrOhavVsjropo3g7Pqx9NA7GP1Wwx6CSeDBP0w9XK
Kqnk7vh+LowYeEna1RkLgJdsZjL3tim6+xqJQhEpzeknhcRrLweWLtifSUige0zee8BVumm4Apzu
6MDyeaAxrKVOYwlYOTPz2W6CiMgPIoYsOp6erf8IQtbDBTeOLl0t1GqwnrMU5PWAoiUvT0VEJ2v9
SPHMm4KUZo7+/7sUBSDseqs+vmY99FcOIdDvvRH9bZhH10Iv3LhYmEPRqL78VJYIbbLxO8bOmS9h
YymPqHX/eFun2bxsr5bfjvtb0Dqh6FoJUh98B3rGVD7zV9hsxo1eo5BLW+BOQyipQg6s8YP6wrSx
uvjQEcpEiWXurLwz2q6pD6aSC5lVdBZ4verO39Qj6Wfb6hn0DXmtF3mwRTD1/STaPLuC9/7Avf5X
BmTGjVaY+i80b7pbrK/3yxhMDARkF3pPdncJx779KNUonv71O6WDpCIzMufNEL3GFsht+A3E4rql
k+Q72Ghx5Nabt2OhejUsLuNngl+lZ5Gve182/3oPbSo+SpCUxgdBl/cP8eA7wiPi/88AAU6ZBhv9
yxqeIx3npH1ytu2HChzkU6kdl1Yb8egkA7InTpMQtBVasOm3yFjjIrKhrC1xIg4v3qNA22f/CWk5
x4J3m9IQGhOnARkIO7a/zD3eRPepBZobBb4PPn1oZotc8db7u8ICXAk1J0aziZ3c/YxXOjpsv+6j
7Heov6aapL2JCYFiMklTFj7OF28kJz1BrpoXNvgQG4Gs7SzJcbYHEbcs7VjKnTtVjK/d242vsH7M
BWZvHJKn6e/xB6cwpqveJDZAyihxC+vjlWm/Qq/8YkKRr/I+ISeOdH6GV2QXjuX11wgNijhJUR4t
/hefWsM7fNaq9TR3gd+VnYRPu9Dcs8Yc+3An1b7PyVEAYlw2nRfC/sYUW/O3Y0k85dURM3S+6z1W
WN2/jZlC+oCwF95b32Q4t3Rn+v3k7Icf+gNTMxGEOuBCjeWvvASLkqaW5mizkA6aqJKVVV+4NR1n
Tf1Dt+kgEDaJT73fJgaTK6k/YV9KzFKQLEe8iSgYWvwbMJqr3lUwidr5UKgv+hac3Jsgdf2LQt56
N5eXApS6kMLeXhI/TAaBtswVzoYCi9c3KGvHvp/9XmjEe0Wv6QqzcFqjJfJGrL5r2qDMRAqWMVT8
EBtvR2CtAjLOisBjFdORjQwUhgQgbop/SVoF7Z6kl6HGM+SEtIHaFu04tfZuxES8UkZ5V5MB62ZJ
zhow8tGH3yPFCa9tOEy220DktLVajBlVutxgQnieZ+M7t8Uw5G6J3hWtEButvntT+sh5WQGc+9mG
egM58Zo/SKKQ1C0enwOtSgMwYZGt6JJ0sA6Hyi0IAuBGtS0ur20ZCnDziAewwml39xetS0l56MEC
JuARqdStGwMV2U9cOfmh2ouE008u6xUU7Ak64ZfDJsLt6JAVaXt+wxqY2xZ7QhqeY6Epo0zCVO2p
duaUXYAugFrAlwK+URryVloIHK9GtPi/K+0GQqnbeHS6VZQ1hS1UpdUMZ3dLmwh3eh0f207zJ6VS
c2f1byicNzjz8RTD6J+GZoS+0N6kp5e0NzgvNe+pnbZQdPZFv1EuQR356BRGiSTmlx6yl30uc7rN
25Qgkt0ZXJSwV/d/twUW7rWuLMf482rMhsdrmYMpf1zXdT6DUeZ3eXsdCyx5FzpfP6eV5AGYewiv
gMv3SoK0cuJTeXs/55jX4xoRhUcxYR6eRUWw+XrVkVFg3rWGUoHfVNKivyHNM4/SQk2M7IH2DST9
mtqD+KoFAFqF+1HFRAf85o6Ll3H1oIqFIxMniaY86vR7Bp4f+hsiKo7CLE7MHQyJnZBh0aoNrrZu
zozxUjkhz0XaYHCy8KhZ9pwNdcg0Uey8id1YmKzkBgyrfHLI5YxAqAHUHaFg+8tLTZhVaCG7g7xt
m5k1RZE14G5xLhSg3SYWOtEfr6UwtH6sKKL9YlidmuMdhp4LxEIRTHzOgUK8DSjZ0x5voJmyw6uJ
WgVYFQVdIhQ/l+y1FK87EUTFqZqnnHH9m+sJhy/Z5Y6A33eCXgPjICLaKN/kS3uFlZCRF4xCQFes
1so0ew81DqYTxfpuVhwA1aPeqXOBBpWCWJzGSU3PBwcntfl8XZhLvnkKYxxIkAfN/wO0DSotBZSA
8FUmxANaq4rFF36idOhbpm9nf2Ul26WlT3s6GMLFGCnM6kDe/mrDxlMnffdxEdG+d3tazP2UyK05
wUPuPdfN8Bpj426PLX8ulf4BDukRXfbYn5T55Cz9tQPhsNP6MQFv5LakDvoSSLsm7WvzTXc/ucRg
fAVRv3uVG2QQm+HkoGAt/9gt1+PTDi9/y9H1siLrrnGo55ShX81hBFp37ThhUH/sj8L67nHFBehw
uDD/Ki0xil0cdtiBIp8qz4xKqGv5oKWDkX/kRjWcpWPgmynQx/WEs7Zwb3FHxwL6ZGX9AkTbK384
KGA/PYYRLFS08DRgX/muaotzaJJrIgibU3IkeAnonRXsKy1Z8cXbNEAVoCmqfSzIhPvmTt8Z48A2
fD2Os/75cBSct/l+fRL8y5/wCug0MEGV0SP0Pc6dcekoE/Eyp1bjwcNTvsfk4yJxvqZXqUE0aREY
3hraYLdvJZ2lrR8JKVtZgQ8SOp1VnpR/Na7y0JOm81R3ZMJfTNiqVrMucoZfCCMgWfXhO4xphGcl
3X2KLqohS1KrGq4jk07Fg+TZYLfiYcCCcjPEIqrns+yJVWxYs7CvjzHsqFk76iPb1QPilo76Gn0m
nco1Kxpv1fYkSbZkx3D6btxw3vT8DpPA1nvypWIItqtJRN2r9aayHwEBFTeTQUF2ywspe+QWMX7r
8mGGabizQ/KsENCPydzRRPZoLJ54lvVHeYvrSlXL4oK5EfMwz99Ra3kKb/atDbQojhCikqv9TaGC
M/cS4FqTmRJic5RXcqSL8cxKD2PBPtRLSIBPWtESlbn0D1AxbXeH9XpgzcQT+IN2/ZVJqphC9DEk
F/ADPFL4hm1lct8o2EukBwYrLh6pl8n81UV6ZWo4u335V+Xmy4rvpPgYhh2CpvB9ALQze0JicmoB
gCQyA9MolPY45AYK99yoRN6kRSm4ER/pweA28m9UP81p6pSq6tU4cIVueEIJ1atM0m0uvSjkxXKd
benx8ZCFntkfD/9l5ebt3swoVdHc6WlCc/bvOBWpoczNVSJxoxTApQLnxGoBMW8GJVbBGrF/7zUn
PAn2g24U7N4X/nnyQsHvG4thethFrjJCz1bjeLWLzwt3mJfYwD+BAylyF942ZFlUkvq49pZzhpBu
oZPABFKb3BY92QW4iViWfeo0S2wot6QTsBAJDSncbgoFb+PTIPIVg23yJskjNGl/5ZSUqb0k93iU
SsJEUgG8ejhZVzOIuLvaOkvsC7ixma0r8Q9dxoskFoYTYPQH+Roozce/HUxdGuz0k3dVta7Y0d8o
goAbHm0fweuP8GQp/cW09btf7PWW2CoDXolpoZs+vUYdETiwwcVzkkabAnCISQSEQ+3+DxhJBi4u
IByXm7Mv/DbIi8OSdIu7DhhpD0k4QuASA7k/TVNT+er7x/ZW4MRGaeL/yNwFeSO2/zdlAbY1u64+
DoxDC/4EL/mr5oquDhubTjgqjMimPIZO9mW2tljGQTmmtoJMqx1pnQZV9yi3Oh2M7rOvVQkH3Tbo
vOYyu/l/AupMrduYxXmpGGlI3aLxzRONuY66rrFgjh6G2rjOYpnfRwet9dJnQrw3rqYQ5TNHrI1e
jkGiOWEUI+pk/d7G7FzlM7szjKRaO0zAqKiuW3BrkjupiHyU/Ge3AXTe3DRnMFsSrG4Z3XLbF51Q
J/zfYwiGX47ZAF7smjLgAGGLKuNxXGza6wsduTpQyvs9VevYnmB5ZT4TJiZvqrVTh0k6/HY4Ieuc
zOeOlmdPHfS7Iiw9EbWN08SD/bmpRJLRPC0Lt8/S41TVql2687Yo1/iIx1VS78op9wFkls9dg72V
xwJhc1YY46BkY4aQeVOB6QmNW+IXH4QQvyUS/F3WPpbEC51qepjW53hkaOoIdHxcWXoG9gOOPLsT
ABGqqB+idhbdbmcYBaMpEha6PaMXW9Y/7BFqlL8To3TcfN3hqIT2/lucldgO47TX7bO1IMk1oKVz
dWa5NKJ7BG4wcrbJS67AJY0cgFtI3+Khrv3tOsz5FHiz75YMItemOk5gDjVjz5sJjOpWCoUIld9M
cN1u6VJzkck2X6L3gC3Ri8RRn2phiVg60IdMVeVd+iP4nrlPltlQlFn2kNjuy0DyPY5BIfrtlixs
qXC7Ph7OEhJ6XbeAJKSaJzychc9Cj+PwhgOhlLIzMTDJ5V8D0IC+O+fGHFJHGyKcJbNcl6MAn4m3
IQH1YOO5JXCtmQGWENiY8QjejO1IO+1L3xbYlvDSVlrwyaZCsQcb2dkuHGqRVuBCV9GNlp9U2wAI
rNLifGF3PcIbTVHXB9hWJ3BRMcpSt3alb64zPsktpxDDH+ysLAjaxm5OI0KEjDOWGIR0CbLMZGie
4UxY+nUNyclR26LOTA7fmOtVdEZY0X430/gfS54Gxtfo/fmjiwTK0Yd2ytDqh5hbxRCKmEJPiw0a
YSzh1LDWnbb0CgjQmugOKoaX2MAXpY9U4kmazcGMC490KUc7MnmTsM0Y7StwOyAxc8mWL6nOuPTm
zRM7LZNUCB1a1CelUgegNlESOirmTMwQKXZF/LEEuAO4BHpURulixe7P8KNqxpcD7LCmd+kYVAvW
jjQ9Ioxtx3IatSjZ3TuTp/sQvXG3vpE7aaPEbRjsUel1yFL7mUCaCiWpPrcVTdGqUYnZtVAMEsg1
HXXWc1Gz+V7+KpXz2Ai2XC3x+TlT1nZ51uTMwJlui5Ua9DKx//jisc/unTaKzXqt7MA8rX1Ys+Mv
sxR++aHKl96RT5rAnRl1+sUXmZoA/q2HNy2EiBypkLoYrSdsR5vkZMDtTou8VpSlwcvcavzCY9/n
mYOxSzonosrfFOTaZ+Jkbmo++KhzxOJvKz7SaodnlOHU084SAiOzpxHdsLKPsAGAZ6NZUwvPu+rb
vgk6NIYmZPMFs85h8n+vgu7tuEXTsYiVVoZZfG/4V0oPw6rNiG2e//tzWc/xwucY4DVTuf55cVNJ
sjND5pRcFNxxZc5JHiU6dGWywk/MoId3tQrP7qWJFtEkQmKNcor5OnAXXzYLmyABLquDChDj+RTg
6zDmznazD4KFMwZr+W7EdXWtmUUQd23zRwzwQ1/AQmMnNOaDY0rEKAWiV+Pa+5BXPdUaXFcF+KMx
UrQpiAT9c/4zFT3rIZBfuLKD3oGCtKyTCsM+YVjMo8MBvHbH6I+1TIH0Xh7jZp7VIXmvppP+UZ1p
O7Ah0g2VYUl4QA2ZM9uLv3feOzwjso0ChZTBEAUbUeSxowRWmnPKFJ/46Fvap8U/Whz3J2jMs8Ul
NnWFhOcEEeOviNgWOsNwXwh7ZDi2kiYGN8xXBtaGh4KP+yibiOFNUv2Q9n5qRqur4n9edJzNbfJA
GHzXZNVMgevI92mN1V0Z3y+uQyC2gE01tufiXBNhDEgYAp/GOZUQuJhEU2ln2e22JGf/hOrqp2dw
QOIyaJFSbi/E9xQ6tmXBFrOPMY6W/uLS93TgisDIvtOttma5xdfj1nXm6EzDimG/+bQGf4kyOikm
7N3scUp94PQKLSgfH0i2heRYwDc9RYPkKL3jWmsgEgt/a41zqO+pIvYd1p6S0EpVW/+gjxvcreir
PnNBMssXXUadXxnMyS4H8RQnqFx0IIri6WLbZN2RUiYuk/dGu9MN6plJN+Efjozmlrs3ZPaNBt1N
gVEoPt7KmVcUD2fgGY39WN17LwLJ/9TIFm/kCm4dOL+u6X/wMN0yse0AsgJB44Pl16zeKtZQ//t0
XhiyFCBxxI2JmkfvyaCHL+Zh3H6/pVENAiR2gvdiKr2rGCQChjR5IYOUnbPutHk7/1JlPlwBF8YV
gFeK8j/xR6ku64oHfSkd+kBQlyp4eR3tPxdB9pPkJmZbXb+LaAGTh9u6Eh23QYHgcr1yzcYmK9Vi
LDEkbIbE4HYB5Cag+ZVYmyFhGPQgQMhaKSLyhbzff0Bn/1zxNbchqOcghoVG+kdlzWtSVcmnPzpv
F0aJhzsZFNl98kurVTeN7Pu6PANQeDlqQ7rxCFz88Z9f3qBKPGlv6J8FBmQIUpW25NmVbmkzKayu
bCKwspvTYxl+J/mbHGQKufCCcO18UoWA0ulpG/lsBbWt54IfqH/4HIGa1I+uaf5MA9ERGqv8LfUM
mTCq7Wd46I3MlsrR3Ajn/QwEF8MB4R6QAjJp0niYSzLJaAY7SmvPoj2ZgMUA3dVYUR8BwVf4V7CQ
5GK7g5XGSNpJfm2KvLeopzmcfIWOjxjlizNYbgFb4XrCsRliLPO+etY3Z4CoXs0lIsK2HO3qKTT4
cqaZmWED9JrWjGrP9yhegEimcr6iWuJhr3qiGq1FuEpQ+2VHDhvI8wPS4igoGYL7K1DzhQmZcaBB
vHyZgLmD/9usx816x9mUSDyX7aNnKsnXUhzjzIZnpQqe3VWwZajykgnD5ZrW9qM/XgmsVtFG37kf
73PftQd9w8lTO/9yCuOOXE+JlgCUcZAmjm+XfJeA+pINC8JWETKJoXqJkueAeVdq7vQ9EpkDPYKm
hbJA5cpCn8HS9zPiamBP/ZjUMCEpXLQ6EsP8eVa+aHyEn+pt0NCqfNJQhrq7L8dvOas6TVPTDaUu
NbeiCGsBrVb4UAQ0Q4cvmm0gowjnhGdU4l0ilc0wv+uBE0G1vHlgGvhelQ91eCiZzSVWlYkP4pp3
vE8nvv0qQLye7haL/lVUB8q/jxemTon9rSqtnI09ikUcpyJfiDXUWQCilVLiZd6fCa+OYUiZGtHG
d5NH45sAecXFXTKUtAbno3VI1z5bj5/i5WsK1f3zx7QoTc/FCvxsb8Q5rULY+hQq3Fq/F2aEKNlV
/X6NxHaEIFNNdfwcMCT2kQkkvW6aYHHiA/x7gMw0X4QMa/WhoeAXtB9oBEsM1J96Ac4GMGNxX2IB
o7CaUsnnjB/aQWe1gaPaCdoSk0RIK2BlzV6af899pOCVyega3FQPLakzFvQDLpNdpPjXQUYnu/dU
q430d7UQm3HrpFEjMNcV5Ikc6jdrSm7jd9X7LkPQIbh1rCfWKeJ/ZLk2JhRSF4JEv9skK6NPte1C
rWrYbejsEEQmB0PH88hFdU4jhOvk171Y029KHxRFc3BIKG6G5dKMZpTZa2zCwaK4gXh8Fv/CZVWY
VVSu2cZ+x/tmqIYOcPL5E7siymngGUQjrH/1GzoLlwBe8xs/NSYH8VaTmI49jtwssb2QxDIy6wpl
yolTliAjCDeOUWVSXcJQ4HWFJwciVXwjCf+0dk/Dc+P483MYGvtSX4c/hQouRgGkmhVNpyWJRQIq
KbcqBBGRTPZRvbbevxbbIIsu4btYi+SmMquvShaEl+s7In5bAwh3bv6Nb1Ll4Y86dBwCgekC2zTw
mq7tmC1Fu4jCHqYVLBCEYH1BovOdjDfuPbtyaQuH4TVuYEijuryxZMp9stsLRli6OiFO4EKTVv5J
1UARUhjH8LHCQ6cP6SdvZTvpb4FJUZSuGxx4rww9+e4EfDZiZk6n/iJYU3U1iAil+Ysggb+XXEF+
FsNqopYMDRoSklnvUvVsVNnLNK/3VRgbTyrv0acWMILULTlVqU8Znui6w579vNEAqRt/MOoJCJvD
0lJebX95WCCAlJU3zoCP8kga6rPwrAslL3Yl0D4KfLEnd2XZIsQV/xJSIY7m1FA62DViABuLSVDu
26v32t58CrYWqyuvp8rTubNGTF8Yj+sIMN1St2888YHV6PiFAJae0qRASD2r84RAqiM1JEE+HWtd
KiD6tm4u1pzcAZh3DMNcv7u2iUkjIcVCqOl5DAjllYwsGAfBhowPzqL2b4mIxHRcM2KzNVJXIwSX
MXennFEohxUv6YWCZFHNCpS+ZAS7DK4BL/Sxn/VmmjOeuxoVnozAEN9uvVT3eY/2qvix6q2F+rSY
+tkC5whwC4YLz3IL1+mb1pkKPkOlwp9vRiMTy9Lh5TxTXffmbSrs6RJSFJ1KdQgbQjyYRL/rd2ga
0WeQLWskrIrryk1vYKXzKXW1oE0nlJ/Mdwpvs9Zq85aQ8yp6McKeMQnEEthX8PuvHy6xaVnW310v
CPeflNBnx1tGteqmsuJwRFciDUU4id0+TBQBgDRBoQWD2KxMZ0v0JEvYTpzW54ivfleJCuztYGIl
W3FWM2Q52ptj2spfWIYkf8Z7wwLO1O1xsKPGtXj++66u9oknL4oUG9sRJUlZ5MaiShN1tMiWM4nI
eejCjaqJJOrj9TF9jThYlUTcLTyVPt7Vc1t04HRjh51OwZsa+LnbbHi/wtyZYXaS+pxbLGrq+S8L
uui81jzH8KbSdool8N78hQDmjsm+oHC4PeHT1NGL7l4gi8x17qov0wRT18o6sVlyHyLWmGrOQy19
bk1WBLNIGfoZouPbBHI8l0duXAD8zrptvbdzPY2QwjWqp8NRoLtyuemmsfC40N0UeroxQSJUHFoh
SD01b2/gJ1r0NXoI3u8d8lDns0uhKlmJFOmar47L87eyzxEdM06sva3Y+8myxmq2CCQuG8q2SxlI
TKqfxJMQOM7LAz64sW3WBsqt29cgaq4VTsAbDGSBpFVnq7mEoBBTYrCulyVrR8CyhK9XsvG00gtX
TmFgL1LGd+BERlRVjmhaegLliwZnCREeVJztwSHKGw5H5wnr4dXfZKt4t/Ffvl3u15fECNyAWh2f
dBqg8ARVOkq+TCEuMF9t0P/U1v/nVDgjDU3NVnaWoKbKj9MslJm0u70rRwJhw/9JU2/VCQn39cZT
pRN9EmtpY20A1mUIz9jYDM9KBKIidD5ohtrywERkGCISHpIktTGrPXcV6p2SnEja5sTID4/JB//a
7sBMgy5o1Notf2aPLaQlgDOqvB4GOFotxvQy1DzyPL8sZyXzyyVO+9EuHerV6HjlhMhNhVQPtrAB
8JPRDIR/RV+Nkz+vl+G2hC4kc2SfnZGXvY2886MSzumXiUi6GoPbQoMnLschPoMvgdyL+eoDYzp4
Sm/b4RT3AzPW1YxL4buG0+biqUF0HnrnriFRa814r0BjbU2ZMew2Oan1cAUdcBaEuR7elwZ7gdgl
+N9KeQOaPHsbckUJwhzPC8lAf2mV+/GA0KBj0a5kVlM/gfOQFw3YJjvbTU6WBVEulT87Evc8YgXg
Ec5CdldXB/UISzeDjmadVYzGTleqsVh/fdZFpjXxbHcuecqw/rSAtC1zAXiS36E04g5tMW2ujdsO
izFldx9rtAjpkYrgaOE/m2nTyL1GcWrNphR3NsdxPrOR7b0U/JTIyLYfeZbv/DnccX3CA185woY/
yrAv8GFcGodADXNsgbABAKOQJ0eyO6qjXxngNSkUczF2iafaRq3xDZHGHkENU5bDm99kVv1xT9mx
SpDfW5MAqcAtZd6+AK7+RXULxRbZrww6rgUL7Le0/9WP7p8fpgoWFEzIWHNTesiuiN/DWcXqPraD
Gfqq+THEevqhCTOKRhoLMSTD8CYbcgf+SIJpWLAyrw42NkorlKq3vu5VPkY6//2YCTvrOC6v70uR
Znvt+mEynDb+GSbX1xYQpHJLBnYBwO84b2lUJyePDuvs/9EDQdXl8FJP7C5iUjq807DtOPtA7q/W
AoJn2vl9cxegaiDX0W8+useONuP376J2wESMfJ52DepYOEIExdL1aX5kcNSQ8sHQzc5fxVrUJHZW
Jm5fkhbyn//DhdeVA7k1p4WfP5uqR/faDpjwz78MGi6sVsKOLIxZ9wCWaGbnTyqxlwY6a3/h04NI
K+wHjb090b/7PeCiTuWQhb20WoXjfP9V8kjo/ZB4tdHvOxdSUp9/0G1Dewf1JigCRww06PfTSESK
i0ovmxBc7EhfJKUJSl/ES6xH/jyOUKzTtYcoB/yfUqVhQjoV+LzmcLip8v3f4OW1pTkds52ujTLi
s0QFA/HxCYe1+3y5eCu36M8NnaRCj0yy5Odohlz0YuTzwvh0/IbGWDzouUcZ1bxjlcVdStqGo0+E
Eprki4JwIC6TRRPaFXYB3sjiyQaHaetug0iW6DEpXH0qQPN1CPJUyQycaLDjEyQiu3yYxSx7Eg7F
9kQOngAEU7OhUFcF3UAgJdMNhizxD91AqYNgHltJbjYAv8WT80f7RSA+VZ+khPQyw90BmxoFR8/x
+UYvSvZQ2qfDDvJ0J5mI0Ev+S9jxrQJIIynfxiBgvqzp+gF2KPdBrdlPlNJNhaLqNgBdaTt03o42
MQkPf1oVI5YLPXWQQ0PBYozQ6wRKWhR6wKqrFM1hpWVNJ+uMdIRPxyIb2hvmQBaZRbWJ7XAWPaqx
YDSKa5neKf29GrlzE4I0BNL+GK25YJv1KDAhtUzVuawHjcebus7rxwpVMAFZvn7lrDFBuEoIeSWM
c0aFN6ntoAzOHN69O5USmNDrob8QUAtUd5dsNxqDg1zo1dAkw93iVPZkjUkXN02qwuw9jkalL3Bp
+xfc6wzldFxJBJi6iXd6sxsoYYgCSkMFUP+6NMb1mgmDxDCp8vyu5LcwoqzyNDsVnYf8V7t6fjs6
LKiZzDDs7u16M41qamfg3F6xq/f1nXhyIEe7iTsyQMmrFzt32cWYf6GJe7MCp2lukCVfNblKMdY9
4FyDmWhnIMET26QWBq8FTmO5hMT7c7qTEBrZVAhi/NV2YlGAG3xcFuvfP4jZPofMdxyERs1u1b0L
pN5jHFthMMEqcoqKolRXVMw5tPapjakvaJTmsgLBGzlDM98X9jQzr6TrN7dpEqey6vS+JkZs9KEh
MJYdRstxAhPNfs4HVYLZW0DMqxh05URE3ZFQBm9Q/anjEG/KGK+5iOyjcAFZKQQk/StaH/3+g/E9
08XEWKP+VQqv4eEJC6IF8BPnV2Y5m9IXEZjHH8kLNhLmOD3d6QmHgpydwKFHO89jMwnvp5+d+wX7
TwFrfiNUr/QZQ7a52qpdSySOJ8y06ugfI7ijDIGhVPehdDSBXu62ZV524/TXGCgd+e/Zp9bYASIx
JUShoPPJ92XXsZNUtXQWVPuEpzaZuDgDun+bbNSgcIxZ5YJfgc7pohRL3e8AWfzcpxOe6t48xyV3
MIHr8TsBnqysYtQmbxvvrnUuLK3EZdwEBNi3Q9EAbXnFHxahjkU7dICJ4VigROaxxiTfCrTUNAg2
E4fy0Joyb3/TUuJwjE4VqZwKekEQfrP6ELAm/b86jxBrKOKaYmoQe3i0XPXv1BGCHd070vSC9BEz
Dg/+9XxHFALpTfa0mUu8YZAnsPOX6SRw+iRGw1JBiqVpTufm8vFrg9hlERj9C4QmhWF1zwI8FdUM
yo8Xaz3319sjovhkJ5GNq7niPAo1+/3H8iWSEiCiMii1LUX97fJJYyXWvERBWdQhpRYy9CahUHca
K+KbM15CU+NsTEmIKt/myR3FYG0uPkW04EuPAue79HmPeJCO5SHX7r6hJBSck7bawkFKx6vQU4Ir
J1zVZecLxR4v+MtlkDg5Ruribd0IoPIe+MiQRq1japS2TlqTu39/FG/ND3rYui+inNLDIVC9DHm/
8YuJsnD/EkNDD75JVanNxLKpitAZhyOGg3Hc8Xi+dTKYYOkoNqp58uU3neYE4bXZC2hyvWq2BUce
xoqfs53Kt5K0aUmr9BF0fBhdgTavrI+D/OtIaSAHGc1kSTqPfqTdG/kjjzW12z9rvL/CNzYJqxJz
yauMfXN85OplkbwSJOH0CgVYndqT4iMKT6LioWbgUyljp3zHy7FunM45U4YUgIC1qdC1FINnpHTr
O5wF74z//YjTjOn8FzfHuyblIilLleQrI59ANqbjHGvetqh1YR/DoJQ6NouUbu95o4x1NRwLvd/6
HftPPvi7MpN8hFWoPldAjVyBclN21Yr4LH0ImyH1Q0ZR3GivR6HJXwURrB4DSwaHk1bnc8tMZiAa
5o3MlUnoBfMrdMdw9/RXVdVu2YAjUarSu5RUT/M2pSbHqDrU3G+cL8MU4U1gCF52Tu+4Fj+G2LgA
XB0JCmcogXaHa8HOmIQaEej5Px6uIv4e/L+HjL1iKhKm9IoC68uBrWVOaWOnNYpFasL+l3GORXvt
3ZVVYe39xJSTXMx+TwslGhceuueT/Qd6sYRImx0mI2babwSObs2OpywzgVs7AxDVHofPD1DtKzSR
pR4uH09mAYvb6Q6bu5YUfqCrkA4pS+ACNBVrUl3KD2UMWOMTydKQqhmH9Bn+bScuedZurBJY4g2b
1KhprNQPEt+5LZWrOOTQxU8X4LiB7t0gIUQAkM0xNpaokfF/aHFT41f4OyXZzi9MLj8PSxcJ9w2J
VqOZCUgQaJkBgStalyUqXCPqcqDpWxeTOCF1wCs9FR8a0Vsh4v0FDZzXGKBPbOGZz/wRUTYB0HbP
evu7pHY1r7IJ3O1K60amhP2ftYG58i7HDeZjYAMHr8j55AWKqfJXWElqgl/GxHmcd/SAs+fuYTyh
ZShHn2asVxddao9a2fKjdMwurtT9EUZdN9VyIuSHE/NIm63Lh6gFK1YL7BdtJv4e3k/vZT5byM9s
MrfxbsCmJwPmbFz6pLtRltS1dIQSZ+QOpmq0bhPPi5OEbaV3bnM9Nl+TLlacniOUJtCjiIJMAPPc
k7dFCmXZhfv347KD1xV3NJnHzWVtW2thqCJJaRy4Nj/tDLACiTW+HIuhpDo86XSLG5G1PCNFTIMx
ucCVCyxFe8n5zKX/btzRbmWTznGu4ilHHgWEajj077fdfRKECYJ+3I2648M9pi+uUtFJkCc1PZ3o
xluUzx1TCYt/+fYgGOvY+P4nsRTesO+hAohGgax0nkS7M5L+114HDf9gVygTFfyA26CXpVeESrk+
96qT9kEZlkfmoeO9eAsMwXFMBOzcp04oIpY1EKAVVF+b7sILOKKUMXBJhvUNop6AvIcj34l4hnMn
ULLYlf4EF3qTXyjl6Sf5up11x6PDhGMsEtXY+l0gkn7Szv6dunhMNVWUczBa3AxAed2PqpS0st4c
0rgGhYVQddfno3XDdfJaANqobp9LOJcNWTI7uFkR0ZVWV5I8DarSxS1G8bnMTpcqpH0fT873wIOd
VzfrDD3L7Pyc/F4UH+BLV+gvtujSI3B+A0kZY2gt8hNr2tGyPzOp6m6IJIVr+gyfHCDAbIhUbLSU
JV95mRJE9PejFCOFkCBPwyWIk5Mg1xcvUoSlG9EV0YGPTer2hrRTi5u0HDC4wEI9Rhl/mQRvbh9b
Ae8QR+0p+aozFdakBqf7xZZIdm9wM0qUS8A1dhJUxjPdNF5vXKJnh7giEjUDB4a3GBTdYEsiWoOP
kr8VBXEEZxHx4XXpN/w4YDzTQyEyj0cniqRSMfpG2Dli6nJki7ZQgOqRacIN3W4GQpWn60xuZ7cF
4D+60v1dfmKSauQvw5W/E+e39lEGXeuHc5UJ1MQibmdAn2KrX/Bc/xgt+4oFrjp3bdTSv6CG8qJS
vxCZVFZm1Y9TUFVQkh3eQxBDlaKhvhtzJ5axPzMCN+tACKPRo6f+T6zoILjeiMmgw7iLKkJhg6GA
eNhmsi5GR6cyfPugepYTuX5cIp45XjXpjByG8Clw1jo/YL3jpfWtLtVwJmot1W71bFWqsUs8k7ab
LWqcJujrOBfhKjriqmXSDwcnT+K/atUCW283Pij+Pf98IM6VNybxCV7DmlDraHflqqhedV3nD+f0
olZGWef+CijQ302Egvc6IoYLamexoX/6bGr3t+xapT+emgt4mY8pXn52vR125tfNpHfgGzpeyy56
nlX9Bbv2QD3O4GfUMSmxz2vniC55UDyfC892Xvm0mOKIM/ZXhUZjOD+a2SHlM9A9O+1P93ybGi5k
KeZ0AmsAY1DfeVFtZhuWhFmvW3v8VnV3Vmbzq9YAO1lTGM6PKdlv13UBJoMyIlQY6zkh4tl4XD63
1WTgMaMzHlDyhSqGIvo52bVzSWAlznGtu/VM8SSYSo0u9KZeUpPBLT3U9JLfSUduxwO8BxeDgaqv
CK+fjNnf4IiqKWIlrO2L/jfA3VtPKg/XsFGvuVHDISjoQyMjpyFJg+f032DHYpfWOETIyiK5r0rA
/bIrlp2qMrHFFOBb9fDxWZIeQhqcTdJeYkqkuobDcTVjKTEMUEjDJX1CzkffHBzAuztqVZnTm7V+
bAqaNne79xMmM9mfT0Jj+LNjexTtuh77Yt/PuPZuziDxlAp/GrrF3nEGKsn17Zh7zczMBgiMaRI4
7/DfjJ9iZDdJOmzXJXBYCGTXqZ4yMeyvtPb2/R+iuY93vl62MrDINznBBcfTbWZGkT9OaZOlNaFg
7w+L1PHTSc9iy9nVto9gdR+HpARlKJdICTgTJoflj0LkSr/Hz7i4tvlyKvIku6DypcyNb0I5GQmO
P14023bCt1D/8M05rtU6hzA3+IQFnDYueC5QohCQ6hf9Xc7fwTs/TS1yHskaZuizaB+oQE5CyF+a
15LbmSIBwTJHEXol5h3gA5jmWJeFvureUxHi/W0XvwnTUNrbwaQt9tjAGtg14ebgbguPf0wkWAeY
KVt5OC4JLuJLbLrTSrGB+VAxWQEi7sHWs0RWJDzNPeuwjCZ/UQ36fg/8s/dZE3A7uO/kkyJM9GDY
nybtajJf7TXW3/2Fy9+Znlf0z/Id1/bMZH1ITsRrd5q9EqpQ6X7im0rPvHkwy4GL3zqeAHw9SHkr
1Q3X9DhbuCz+OIPSlZuJQZcH+L0NGnDrlbY5Agvrh3oePsi+hFyz1WUM9lGiPGJjA0hfUHnP0Vmu
j1UQmVePSIBME3Din+Y03iSQyjpDk1HQ2HqFQFMepplOU8H0DEP0q/rQ0W5TVCqleiNRPzCDMhvH
fVP6E15rRtm/kRPf2GfymfADj2snp78uhseO9EbI4YAxSbBj8VqdAFo8L6Y71FPbPkR1yvfhQpI1
fHvgjrudCB92IRo99LxLgLz4DsSBKwX/e/2qlQBC2TJWUzNNY3dxEsADTM4kqdvkwXcoRio3z6i/
uO7cjNoiD7gW36VylfaCqTNNrD79xLU38Zaz7Pr6iHjblDl3AIxH3SB3CgMy9RdK++NrrzXMTr96
2u+MjFBrGuzxBqPdV2jYmEatDQJFkxWYDOYA1rSezbw8CAv8JQSYkpKsXrdoeP4gx6ekBXGzJ9Co
lwsIyxKr5IQgich3DU6oTdtvHdPh/D/0Lu1Da8Jyp+M+v+6TGjzqIt3tcEBCs3PMsvtaSn7apY6A
bg2VQBAj3w218d6qJZ7mXN4ZIqbcUkElCqHPdBB9cUkbUEJ/mt9A1SXbsQHPOy1pwdN4v8nQsL5H
871wXp2vz8pQKBCYL/ymWuAQr0QsYyp/C9B8oaEgKWY1Cptov+vbE8OYuiJz2r+sIX4W85ymKOjU
TW88jcuNFLYyT48d/+T6f/bUHenU26HYqT5IVLVWr9deJD+6aZZWNhlHF1f+0RU62j9mSo3QmiqL
hmS8FuuzZfSycbDMrMvFQIbzco1sJ+1wEGgCDVy4kCJqDk+arPKOUjR2vz36UVbo2lB9PKIxQO4G
b54LIYYO+SflgKLeEHtAJvaFnCtmsL6EL/v0k+tB6kYI9V8JbHTH4CXF1TPStWyPeaoxfltJvkrF
k6UTs/G1J2zEG8GVjr6RQid9DJLXJivyt2aD7WESFSErZtT4CQ3ZLx24uMNI+iQ/tXVxTiw0o8+k
+OunvoyuTGi9qBk786s8Vn8YmTFxyDg+lCSAVmWqxtlJmJ3TGBH/ua7KmBDLFal2tI6SC5dMgDwz
lv5pzVkfYTIiu07BhtDychqO6iZAfi9ACAeSU/OYM2FMDJhxTLTZib/F2MgnNfCC7LtQ79bkirfh
Wsl/s4pM7NEYzqMi8wM5UgBxc9JO8MREOukuI/tkPwosGjqrGTNMw3YEqdH5BbYhgpjW+wcPwn4W
en+eUv3Td1aVf46W4pjsOZ03CkAy/+3LMMC5xf79Ekz6yipXXt16TuSM79vCLZFXZi6QZLG24+CN
oikQijRP7VPmVWWBuhbJ8X2kEORP67PLaDdbPAybuzVD/k4k13Bwbc4AwyGH0hj87u9vMATNOFye
A1LSvODCkI68/4IIrJljNvIemesmnmkNf16S0oIYDLYZzTHYLxJtjje71y8ieseUFX/o+15PIeYi
QgeRJ3tWCjun0DoHpGRM2dvtdyJfbSaDJry92sLC23o+z2zo4QpUZOf88TPWPTiOFOOETJZvu03g
+9I/kYa9wMbhjt2z1nmV3grNXD3sr08rjqZekJaWJyOd5vtDlsJM6USg42ZMcv+WoxPusOXAsEyB
JTWQt1Lk3eX5ahqSTqnY/WgZVANljeGSBqRWy7DVG6bN/mQwGwEEP3S5WYSDVDxHZzt2Im5TKvdR
hswpIrOUAlGWEHWdmJ7y0gOhYK/Rj5OdaJed4onVRd8ThmGMxVquRyn6WpOdvRaitM0kazz85SES
EifKlq0n4dhZv3LxTVvVLykie4Rnr8m+5CEYJ062Ti+Bz5PqW8P7UWa3YZR/jvG5kfSb8E1eJZAP
KQ+G8M16Cy7qL1Fl8Fiir0Y6OSlf5LbXRsJDjK8S5L4rYVyIMv8OJdc5pJQTj+5eatAetbUtthGw
hdXf5W95kvs6AUMC3+V2n/a2/+IdW0L1Qma7nvv+TCYvV+UN5ZooeWulJajNvlh25AgTd74S6kpL
msQmykEX/gzL+BGl/+qR5UzCSMmj91scVHHK3KxljImGfDO7rDnxkn32DSTn/7ClwvrznREU5hPT
AZWeljcoVlkfpwuvEyt+EqSYYSYclyXDseYFWXxhtLPdlPo/eTm7qRfVTLHvbRTGpf3hIYPNZo46
MLOSV1pvT7EQc8shEGw85R+vksynL3ezhk8SkkmsJLWDMhUiPlbkOnyYFtp9xGMnlj8UeVjlrZS5
zLX98ig0z4VTi//Bai44H6jPZjKR7Mq4c4InYcQLpuPAcEG3NV7uyX9RVFubheNr/S8Baf1DBYi+
KdXYPj/wX6jJT511kAI00AmnRP2rz5in//kmZdl2IW9Ca9Ax/x3jMn8pGptHoOYDMcVei8YCvqK0
6BuZwFa76RjJM1n7z2YOUXsfxTLExKwHwYsakoJXpI8/tZU9QYtyLZMCmXgvTKTh1tNicUJeJZCY
E4IykzGAyli9QxamWmQnwkEqapxEUH8JpAmMg4ePz5c1jjvxT1rTB+jGyWpUPS3MZNnTpCUIfzVt
Xb1/IY/lnQcfB6c3agOhCQVCOuPY+WZoxwd7J0g61k+ccvv9WIv14oZalFACOOYnA8wVK5AX2vQF
yOsGbQo5agLCH42fgEnRvdCSPh/cjK4iLOemE+W/5M2uihinAyxPSqRe4Z6Ji1M57ex+kbWE59NR
VsO7EMewUdfIW07kyQSSnUQpDpGdcuUZqJBMeBiEEOQ5ceJRINOUBg5noYgIvKa+xooziE7wdrZ4
ODr5xLwt/nsftmvOwVrZpYmLl1T9Rj27ARaYw8SH3x/gEtvJGbQPSObUFOD+rhE8oQvnQAywPgZC
P+SDVAxPo+EKk0HWXcxi+5NUKya3Nm8TMFqXT1QLvcc/zKvZ7Xl/L+HfBqkv8QCLhE5WIs64VkJr
V/Ayp4ahmV4DzvqjxNq3HlGm0glF7VgWINXJn5fShL6aljEtD1L9lwpYxmcdzRDHajxcXneghQZg
XOY8vwJt8a+zZMpb/RKQl1E9QRoFjR3/AXhjikHqRZSFOnTFno2V1D8j94Ff2koBwLQ7eUh1oNy0
9n+mUADI7tDx3njOGUi7fhcuyMLFIZt19xfVourbHL22DlTqb2bJj/TI/kA7rb4iSMR0FMwBx8SR
NwdJk/TKgWAHx9L4OBEMHdDgMOa4CTc1hBnZFEVji028EJDorlhOxZPnUnyJedXamovlKDGO2BL6
ovcqADbYKNW0/Grp2CK9Yp7vEfbX/A8fwo4SboZPF1gCYd+IwEsFaEBkkIIJz/7gbbTt7c6UOsS7
qPlqFr+pW3dR45tc5NryF8s6PppO+rVPQsA0g92nc6GmL7BZTQxBMNXMERVaZsh8dnDw8z9uZKf6
DpNWgxyTCfOkYSXB2MuAA85AignXFuAY55B4kjrVLQneq8wQnw3FoqznFsC7PSTHN9kt+z0z1sJf
N1IwN7/FqWVwV86Hg+nMNXJi+c1gKFj3iFQLjv3kWbEYs71jmWyS4Yy9ErFVfL39ll/1VBLBtJyZ
+pAVK2RVcdqYe0RxGpoqE+MYrBLgCRALchDTejhoRbsd3+3sj/T8x3EvrO8SKTbYaJhWb99ZVsDX
HJ/cPSi/mVwFh2FnXKEw0Ocx2xuJokZTbG+Z5UbTIq6ZDMG8nDwR0PEk3+VQdQnzK2nzILFRGEVM
jJKgx/iPKD62ytCQU02YrQJGFFNty7PkXUtvYJDHd6Mz8e8K4MQBU08BW+2oi1CIcuo1jxBxT0jT
eUfnSuQuuuedMLN6ZFbK+HjBDjUBL6lVlW5ZsDv3UOqQAuvBvAqp94EA/Aox+VC9R4mic3JVwyE2
qsQwodFNQXdK669nwwXNOTu5c1xJiJ6TXwQV9a7ToFTH5rb0TDmxpe/gHC8mzzyE4JrhZOPRccQy
j/jJgKHnrN6nnxwwR3l3iN6j4GzZVVZSF4TuFpVbFFc/SQ8LO3C0PZMDcOuMxYaBytZLGbwRfDry
t13cqPCvq3ZpsLmIYXTsbRWRtbqsdaV5UaoRAosV2EQNcfTVkG/M2XUWxd/4qoxGuGrIOCSOB+pI
SId7xbIFD9JsPmG/mb07/+vNqSliczpkpjxjxwKupp0vGktzV0/MhpXDv0JzwWJDdE8PKegy8G+T
7IHtfIQOMaIkONEjCj02P7/3VwejknPl+kCHNyPsaKfTzOanNF7yrq8wOeoNtMFp9ypq/X22iz0o
dTucpws1LG+rTwe3ET1DW5iLmeTqvFKYH5S4f66oAqQ+nZa7H9YldNW+DNPwY9D9a8+PZrrY07/a
4VF7ZOZFIq/WqoaiVXGxvknlmVFXHGm8pwk4O7s0RRv2Ye//sp2WQZfdOLzDigwnDvN0nXyFzMTv
CsSujbHCqBjioZGv5u+y6OkULRFP3L+oubb2F9arJoEj9P/es4RvsTAoDM2tbTVjI+6i8Zzggt++
Ae0erOkKrXmBkMWr3b754r3eR9y4rl98OnGOx0eHqJ2sKWYMhoC5eAmuhFTYFPFq6/QkLqftzoVH
pGOtIotwSC+cJVuAf3vYz7b0pogeWMSnJkF/u2pNvVBYEHuPt3Y7MjFTuP8FrVGhcjOQqZBiHv4l
ooXUALFJrIyuSOuAHv1HCWFmAmNjefY7Ksja2gBt7f20mscLYzf+FoPfEUkPYN+PVhipH/Kq/hir
mnXmi3Ern2bPbDwPGvaI2a44xNZDJ0Fnnc50ZLPejlmI3A43aMCxxRN1FPbhTHgWDj3b78AyxVIz
0WympqhUmONzeZAFjTTDeHLbU/uDPI/1CZkXmJViHWtTEB0lJICjcZ0+tLm67T5KX7MHKwxFp7Mx
LP0YOIJNA94vu+ZG/wTDDMNJSTHw5ILbzrgP+6bAqacQlFGnRdbNFo9T0zet0nxzhdoKBRPFyaeb
lb/eLfkeT0G2pNMMjaRaqtTWau5t3506zk2L9/Yn2vavNFVRYwLHNcJstX+pSGnpJy4wdZZK/gDA
yxENycnH/PDbWEfs3qZhr1oxY8ITM09W52s8W9+ZP2crG5Dc8LUwm68eRoF7Zzbk6Ku6xl/LXIMZ
+e/nFm5QkNScSfvKE9YbdGXx+/yIW+FDBNljMh7g3+F0jxlMwTq8DX6qCb3gUf22MafdqF8v/sGo
Y9+tjxDpqxvjMGM6IwkAGCwR9aP9cWN2op2NKXYab8TOvZ3CQ1+4aZBBLLQKYvG3KZSTUDu2wzWn
O7c1+V2z/PgRxA8IlRsmYpsZbQMxlOA4lqzAGHdaU4FKGcvUDaIIHec+Hcx5vegMblebKG2/B/zS
oqTCe77P0/1UNVHmmWxITI/INzk/0Dfwrv3iMRlSpjwtHtWrPsXYUGadadhvlWA45h5mIGLgKdQ4
iMz7NI5ELWei3XVigDiaQGVTGHPKVtPVSYLsSx0/+Ojl6944hmxITKbT+CFUwOwo57FhVeQidzrp
m49ph0Qmi0+H+YgwXB44mSOHPXp7qJcpac9nAx2QlJ5QSJC32q4V1cOmdu/sVGDs+ZajF5IWSHxD
yxnRn3lZyInldFKUJcjGUVBm2ayWf/AtlKtWyIA42RJcY8HAtceUrnP0GzaEpcxe9FIrV7uGcaNp
MxcFMEh2gb1lBA3+cy5cIIxBrcSp2CL/qDYi57tRJ3ACfAAH2q4BdubGDzl1wY/3aTbrKkaKxJDv
Oiw2NY+PwGZp23PDCwYgsA3uv7oazC3UFP59YrNh86j8xvAZb3drKeGj464ZTgbUw0fIvHPk6irp
a5NFws1LJO/LwHE/H/qBSaNjBWxKv/rwtasN6vK7wqy2gCvZxI/6fZgStqRCsJaJGRrIFrSGiDyy
wJElSXeS5/B0uIM1+N8acjf+XHCAHRDyuIkwzWhMu2Nzgi1PN7M6m67KTMPgdlBYtMIOaR9K33IF
cx+aktoJ8hNTeWdgHa7tPz6uY6FRlGUsbbpNugqjHQs1Vo1S893K3t3F04sQFmWCy7ZugRs4sTCz
w4y+RhA+5c6MXtlO/qHQ+utFyzrNhfxyBfkhA3Bx63zu83rYvjoOA+XzJ0UXjll3F22lhT4G6gLr
cPINsyoESgsrLaTmyg+ItqVSxsCVglOEv51rN9bOm50ybRroBCcrpSWC3bQ9EkMoN2YHn9+1rnz/
8SDRmlUMaFgQjpCW9ImCqBnC8DgnXddQEysFk1Gjcd3AYGXEDRg5+HcgV8hN5V96WX+jidXKcw5i
/XC+eyCzFOMVISa0hwJzKWchUbST0Zz8KMWxS2hkpF/atCxzx1ZDfSMVhvzhzeU7Z2w9j5m5x3yF
BAx0TRHFFxlgm9SW1fHTL7Aoim2JsQYQhPUBXfuYOOeQCjJ5gJdjpvvPB6OC4KM+9hNm6hpPjz6h
Ev9DvPgeqKZn76ovRWnCm9kJS4+vC00e3mh5C6WpWY4xUzG/OBIVMnOCIWs+yQYeypf+xmVvGXnj
gfA/MEcqiwYIRJZy7lZMOCQMK95nJGpGdEdqi0ICkNjmP9tlsbns4mP2u4Vr/NmeWeBO+IChZcnX
7XK7RcKXOVW7m1vmVtnXSzWP9iJ+lM35bwNUfmOVeHRowsm2Zmeb5szmuhbU9SpnQWPY/JP/wk28
Xeo3HsDo9kiUaLOUx6YweVxX44tzI3aC68IVVKoVpETH6nIKqBncsYfL53tq3A4Gy4jIfHjn231A
imWTeH/N5fg6pKmuJ14TYp0rGOrn10Uo3ws9WZAnqe00Z83Dl04SNcsCjfVuV/UFlouT5dmGWK0H
MRQpMebR2WHSDaMcLMWiP4j7pY6qqHqL2Ao4VIH2+IEFhVdJnV4w4PofPDZIf2qF6IY8FgSns4jt
nqOiAjWlloOLhYY/ws2b0UdReIPymXbw93vQgPOjI60LdyLI4E4ZBa2bsCio5mXDIifseTMzylKv
GStfgkn/cXB29Xy/2WcjFH3RThOsHv45OYQakIXQtnTHLKMhUWX8tp4U4w+1uPBbgmaDJd/DdeZy
he/hLt8Pcy2FEBjS346tk3GKI9cdRWp09QqT3pLye9zRHMua24/RQKnLff6QwckpEB6/upIALYxd
xYVLz3l9Y0X4NIDN6eTi6yb5YHZQAR2PsFLKJt3rdXx0z5X9KNhhNR4xWqemvI9dgJ00T7Ey/A45
bL2rFk41r6aI5fEl4QOqXcFYh/PQcST3OMkqMa+VENh/4Q8WWvGXcHCVLV5iVDeTrzWXWnjqhPrl
l+wDJ3Xteeb/rXNJuBNn//2mzd7WWBZQC+NuScBvn1iwQQ7ibuT/7Y19y7nFVlbpdc0o7RmxDT7v
VBqgiZHlHpH1rrTo6ACuTV9TqI9JOMTIKE0oOt5XHReR4CXYeU/oJt2awP3D1sjZAQPW6n+mPteY
4QJjpctt5+WOyWXb440VAL7XylMtajBE9W3vE7IFSNWXXrjjvvfhlmJ16fjXL/vqiw31D5pgz0TF
2k8rKvDK0fUElddQVXp5fiht8o7GgDKa5mztCv+kWTge3rUpUTaOH9JaEaqeXQR2U1XGQI2XJ+Lh
qSrhnu/WpAQugFsS6L+wo0gxVcaFXOYnEvY6tgQeJ9qf9a3x1VoCdca9YuBO9tB4AxvisssAi52a
PF+0pJ9o1CQG9NUGaD8wP61qfBbsAEEk9DeXw8qSeJDHmg7DEJCRQ7GlISu0TEoQTQoA5FNVGggJ
IdDSxWRUYpv8PFftjtnHIMyr4Xpq0C0NzRkZhPPGz4+lzI2WBzO9yW8vF/YYjo33mtyd+EmiS3MF
pn7C4kpc8Q+gY//RNwxB74vKBnx6L7Amkhzd6vzMCeidnYooBH0He2OdZhY4hBG8uDtCBEsgpfS8
tSfWz05rYbZrsSZ1LU16+kbr5ZEBZKl9sIcaMpcMwGazFUPt49JJQdFAVjFfeu6S9KwdSrC48nkT
rHAGkwhmklyi0UibJx4DeZecXaipYria6BXIM5NDeipLgn5A+XYPxgb+OQ9PplKF2tx5YgUyy9ah
pZQh9Pp1RIqQOjWABW4FyDH9eA37I85kv6Vx1vzgIr5/TJAzX8MpyImsrkHZInIm0RJF60h2II/j
9hoXWFcGdZHv7G+0Khkx3jBx8sC4G+YzF7ViCW5G/NyyMScOCb92yg7OPqUBmpmrAtGZV+t1SE52
rwXU7/pbjp6oyPGu0QDJAeqUdzMbxpAZoahV4KG0rollS7XVTisLODzN2q1DI6iKJA44Y+nnPoDV
v7Zd0p7QzkdPl8x4Tp0P7tFNse7H5bBQeY72bOFKsQCUwmFFNqSv52mUUBZndcodgWsakEoJC8YO
PtRJs50s5k3/tv1Tqu94jXg2jeeaVmcjlxsXouO26rPLTv1Q9PDHiLEgBjRn04iRNDeK2sJr7yrK
VvSRpGaRLY6i5WQ6eK+UqEqI+IuR2m8FSvxjntwBXjS7mRXmjOu0KxBBqtMkeelzpQzSCEL8yEa/
9bxkD1m4j4QMAcr/1f1FgIk1bQHguQiO0wM1rXpeth+MHRZblyTcoLg6iCg2dVbNngtXfyW81szl
xrXxfCnI6hngM3wLx/BPv/sUrhj19BpUHAk+2/bQaluZh6daZzOI3RvnQHaKuh4ehYNq1vbK7jgJ
1Ul0BI5JSPicoAsGGovRjnCpR44cFkAhGdazXQn3KlduHw+a2F9QQgCwESL8xkKnLeYPzcQeMqh2
Ih0747QGXFMstGCWIsbSSE9op/16NT+8/Hzk0v0o7rHTExNnfjLOBJ73Rsp6j7RXpN84TmlyQP63
HDlXJvcwsew/iJRATAnXtwJHQCepvdf6ffx5IvxL1bXuaUGEY+FTFyCiAv+vFRH2Rc2wOfkEKTXP
OMWxEnMAWipej82RtFZguO8UTZ3Km+t8e9Hcjgruejyg1/4nUsTBSx1PL4ump4REDhqiAoTnbfUM
XKstyuy5M4pZlb9+sf+jYmHEXq2zO2eEPhwU1HFb+OlhKbU+0yFOkPZpHncjr3aRjuz7ckKz7q3t
mgoLA5rwJna/+i22hrShbpXe26yHh3jmaXXdTL3faMINgXV3yljcF/YhNuIYg+lWoBHGcBplSmR4
ehb4P5URFLDN79iL1eg+moB7D1ZZArymNWuV27+oS+NaqR4QtI3BGzQt8glKsOE4jvYxUjkmozn1
7hINNKjSfhrEfC+YktuqHRXhISmDE+87teoI43fhelZlXlrzqZyPZYVUDlh7GxppthPB/9aQB+p6
6XS81HGUUlhL6Pr74zA1ijC2/xIgIxXnPmoH20aJKI6OiWQHIWvOV0PoFC9HAL6w0UsLf1odo4qZ
SNMb+aKsdzHUAoS1vz3uiKM5R2OB2g9Pexu5lqTSliQYgChcTPK1dbMTpAAOo7fTaOYFbd/njlJ9
tyTYY6cGAxFBNj4XP0D5deRasvZDRSukmip4rl98IvoqbaQ7pySJ1Iwbl8lfwGAEOwblF7CVO1Pn
kjV+NdXZFyEuVh/lQieaC15ED6Q/1CZ9QHNktgW7gb7GRjyRppZgKEkdxZj9vreqSY2j3LkI8/sV
doeRzMRhsNvfeIKHCGGo4wpD+aS+T7JO+P+0QgUxUzryoyjeGV3e3hrLDznvyJPgcrNnbjW5ApJk
DDX9wZZfBIiLLmSNh2a/vQbtyzGc9ognV1OQqGHC1g7osF/XATsGt+ect7zUkeXjB9f9UfdtQqjr
RDWq5xGMk7pF+EQuFuATwV4o6+K29l3+j8vzMLu0ocbBqgVH61wFcJEm4uqN6zPWhIQhxMq0CsEC
zf/dD/sjp4Rgjqr29ru+P5+UKLFWKIDudNjNxOvF/upo0bJOTS3A7bUURw9EDAW3UP55/LLkWdA2
Ww59un6ai0bJ4G4bzMWXNZhyLXMIWq5khQ8oeufODuaElINMhkk8Rr6MctEq4M8oK1mwF1r2QAUJ
KGnE71ZI+P0p+Brg+2Guezje4jKaH3EpoW4xldozBzSmT7G7No/5VDKFpI+UYIR0QMY4Niz9nJwJ
vRXUe7i9NWb1556ag8DWPvB5iUHnglspytI6qX7x8O2+HMV69nd7YmCTlmGYITi678H6tk6842El
prl99emnZ+u5eDXYcDFTb915Z5TO1D0kfYK0rZiHfubYOUEMiURhvuJb62Sub74ggQOV3OS+5WH/
oytFwacEv3xIHkwxsKIjR7xT5YUAoOGjF/Scjl4FvoSxPd1dv6fsXALyaeFDF3j3Jm5Dkj10onki
n2ilP9Y0vwXIKnGcKBwteRuKAITw6pDBAwr+dM+iNBnT5CnE6QJAF55xhaxTYhojY2JMOD4SXsPo
Dro5XbqdaGxm3Hdg8jdrlWpUcx+/PdfoEus78bvWgDzORVP/tmDaDYjp+vCHtCxrE5ecSUdjGS4s
5DoNXT1ZC13H6cBHN0yOIxkHuIwKoTVT3X4as3UayPOgq3hC8iEXRPWOv13YbUXYkjtPaiMIDzkN
duBOSoZys/HLaIIc8YSn2V/S7ZVclnce0Fmx/zbho9DFGhPpD+xSspKqSVudH+TO7SgeawAYPGkn
VpX6uxH1SAM8v6Iy/2NKgb3EEVhSUircJSyxJSkNxnKLAAYQ/QMy/xUeswJHJWRqyzdob0Hy+3ab
dN3RTNConc7sM73/GWetIGKfa7xD+BqIwHC3Hh441Z7h/oVWSMLReRtDTryd50ErNlEDCo87qXgi
Xc1JiPlj0h0vBziN8e+JBuGnVa5/i1RcvD3eeflS6mlNph6lxDw/t9iEqBjo7V5I9xcAZEQiEM0J
neoPDQRq59FghiM0cJKwVSXo4c6TD+OqgVTKxNiseQbVVTTAR9s6gOsGjr/rHpheTKlSfs7VHp9z
aVeGXq9gQGlOwGIf4mbOx1k/KCPxjrjDO49htTKT8K5u/zfL5XTOQA18qHzOLXFFdv6rJ7uF5+y4
6l4zJNHnzIBVD/t3FS9jAl7pAoadwDvQshYd5+B5F2Y8sBRe+AEnt9yLLrq5OTFghVVCjPDW/ywF
7x1IJ9v5RgZj0ycwbbXsRHU8VWPQ6HOBZdLOq438GqClPGJxtE5gh2NvYOoVzC14OhV2YKFV4txv
pmP4Bmlkx0YBkT6QD4bhDCYU66ENq1r0vAy53NTxxXzDvUIJ0PBbxUwHz77WzPV0S7R+M/d9w8YZ
ZeW/lvcqYf4oYcNzlbOJTT0+frA2OS6eiFIO2XuHTsSOeuUbRxVMULIkBrcWU+byMqCwC3orLie3
bOKvqbV4qnawBiwYW2T0OzMwgCp0AsJLd0CWCux187v8lzbDk9wWDz6AGu257On6qwPk89OTQOo9
kC9yCGo0fddA2mr0BQJmwWJIuZfBUyPyEqVhZYOdzcmBPm7EWPeFhNxuvzP2J48iio5BijzuBuXo
04AwPnLzSpHEIpoOE5QKVv8lgJTA+BPSQiPEhqp9fArXgExJ98j0cHe/r2DnMMJlUEldtI8Jku+R
S+A3G8NWFC+lbx00RsjPhLXdFrmwxbT7nLGEUDtG59kPNo3Ki20PrvKgh1or7LcOnPuyx1YLEAAk
kma9yEqPVebUTmVlK9EJ3soiJQFftKchyD8BhcT42NsNpULsXzuRAUJbaBtmwedFjBbhb2rGURBW
KLSFUTvmB2abLKMSZ3iduSMQfKa8NcHdKDslf8v9BMUtPDLpRXFn7CMBmmSBMGHgTJR5DZ00pJlP
Z+HOpwbTVxxABg57swulYjh58WMvOfscODTbcjCc9fseu0/cbWmzfW6TtLKc/aUH/3RUWVsLE4sn
SL8dJSw03eCfErfcjLR0mqQSdEMQSalfkehk6f8471HML+m+5blgxjNLzXY5oZd/VRZ9GEfTs72e
jb2iPf3BHJSDhGOqxA6y0qlXOaHM9t3NomJiK6rOFe9D0Xlq0K/IYmKm9Y5HhWEGLkAUDU0M6XaX
Nr+kzsyGWNreUkI35o7q2un536YRUG9cJ2uSUwjQsdqCbTeAHTUHVycFAb8B0lTQk3oeCHegSRQz
WyxXaFG1bK7QjAIibvNzxySEu6gPezpEWJqFGpme9MlEDLMayFJBCrSftSXDnyrSVwD2EmN6RL0N
bVhUebaB8uBHZ6LSFFld2x96bc/5/RpnYJRVyk81KMgd4LHqnJZ1T7zSAXSLFmU/gYcmptB35BKj
tEjNwhTPUvCm116uvudNDDP62t0r/wM4lVM6gsoKdNRwVU1hDgG2cjM2CUp9+ph739OCqzVqSD7z
iEiRiA5NpUmd3D/kH/e+BOs0Awtr4B80HdmSFo62tRdz41/d2LikR/ei1sXkKeDgmu1tR5tqRasW
Zm1oQQ0U0oUuYAQQ39JxVPhplVUOQqTIy81bIixr5jYtAS9hXLpVm0/7jLQ/LvIrnRBz7iDf9Gbq
4fV1EIVx70Vj16gDXM0BYJUwWn7tvmpqLtmQpJvME3ij8Xtvz5jTgNDMPwk7XSlrElfz2OpKDX56
e1CH1gg/VoUVPdqminhezhviSsWEHlWX0CR/uX/+sxe7n3r9ePkP0RtJMNw1w8UgrjWIXmLF/ab6
NaKeH8keTk5KjTjZSitifFh2bD6Ttly0D5B+4CEtEPtJcd6XmNchHTNchsTd4Ou8YIDWs7b2RtdP
XWBOaGlhlIC8Gu2UtdiZ0zE7BUc03oRjJPQvMxCUzQ5k0MFj/wNNbWf8yzU/uOTmt3myRbnwNIGK
IbABgjj7+OeyYF/OiHtKkaI4W5anTP0BxpXV6iJqY6ANC3oEmxuwZ4hTKINVAy1S7zvLIthsK5eB
X3tJBsZC1L0+V5Vm7lr7CLQHYK7t4ngn/AM60HGNBkm9r6zU6rmj0Lq6foM3mQzRKwRCWF8jxXqH
vzggXblQ8J2RsBtV4xr++f5JfwDgrbajFrd39Lwo+zJNZyb2+cR3wBkvgBCOgIdCiqF+iuRImSn3
k10FF/0jgGCgtGJ1QJxTu3trbP2bMFUm/LvFhR+ak6ijFiDRDTaKfohT3iCzBpr3kgp1Cg+1kj69
mi93DUZ7yz1SbLNfFkjlwENY2qch7rwDICCmu1W7GFjPa1Eq6HAyp1Oik/B8lsm3b4HrYFe0OPGg
yrFz/j4ub5sFTTV+U1mfMnMzVbpNbV4gCFACMBPT+S7LjR2gfcr19HTwvD/aHNq0VxgWnMId4iRt
LYMAoDUzV5FJFWnWMS4+WdwC5to8Z9kIBiLyyJpSFTo24rSyZkxBnKQBcuKVbhL8p8BpIuiV38oD
igY381Si/nS2eNSAHMNPVBHM5BwRgdK9b/cbyLiVKR3ZFf6ZD+3dyjsbRTs/zBu+cno/LvKEiU5N
l3P5L6Do1Tm5NU6q0Nip3XSQ2dlrsZAU/rIyVc/sL/ybPd4xZs63XK4PepXm37204uJl6DKXR+6B
c/pkdQBA2eFiwH7c4sd5vGTLp0vrW40AzQ9K7HKxtHFa/9vzxodF9UfAAak00AoFI3pysGw26aqQ
TIXwVQcB26rgEcRbiAd+fghMEwH2fcXaUZDgfeeTtch9NNLH1H7t1NnPz7Wvlpam4g67LJMHgZMk
3pDSJvdLXTN08zWHtiEb6ZGJa+pIdGAS7UazY0cx4M2VkX6moDPgWV6RCh2rHq0KkGkzy9deeJsB
Gc+1xOBLvQEb5HAdNFmU8tnIvXpiQ2efT31Rq8U+WRhhQCE9WDpduUtRUGf/MC84q61TbncxkjI1
oKAd+oT+DS4owLO+ZjAZgOL9oV+kbQ5UAgpdfGWTelPjQO1GOKhxtFQggUdnmaMM0HkPuRol3azF
uHuzTVIwdrOr4XlvqzUjiaZnv6sIqDZ2ZzRmvYCCWu2lIJjrUYt06oT4uZfzquCaDfIA1ASIeFkR
HUOQBGUsDJNTFVQ8f3Saoi80aUtJTccvHV9r4rBMPjfemfWyps+SzZ+MCTrg7M7M/uGJirbzyN8S
WqcCU1GFM/y4koZWQ7HPaOgV9nH9ddDxPe7SL0yxWpKpuPGSc7220lb9mJnSFLfamxfh1o3AB3At
oB9YVuEPK4j9/z5ZEkxcDCEufauni4eZbBQkU9GWu0V+vEmtFTodoGZ2U+/RsCZ2HZR8ux52NwYe
PxTEZAcLZFaerqlQplSqCCqiUvZqR7J7aiCkhhqyfKWXypCsKvBGiA/nMIAJWhJ2J4fN1tSn/IFJ
yIfffruuBr+gzsiM/Lq/pr6LMh3JhZFqErYNbPacqjzeDbZTLe3GRxZC+6rH8Sj/h6xcyQuvSfi8
ICphASczN/JpYxINKoP0hrGIvkkm5TTWl1HfPgjoOYHJZYGY10LeNqn9lOu948wH3seFstGAUt0l
FHs/+leeL5UnqpeBFxb7SqOK/ZytjfNhckZhTddTDUmZAedQ7Y+UMMbyfKmh1I68Q7BFTiVsjVyY
6jtHDOwaY3OvDezXmnWe9D4OKJqWrvA5ZrlwJIgf6GOtRsZEilyijkPT69XkQiGrSlUUAdNixFvZ
fVph1FjYkIb8BYYQEt0hG71kJBNfOCzSkrx0SYmNGU1iBzR3BZ7WNEibQhZ8tCyGkSgG0mqg3n9G
pk7QIsI/sKRoX2UcCIXL8a1Oc1GfTwXTslXklw7o4ihL1MeyY9cmEY+fAXZM5lAfdzpqF8W6hao9
9pZJKY6PG8dZzgsIw6/tA9gb7ViTpgrXUD5byvm8fTIB09JHeceYpuKmA9encxIh/6hT0ck4sAdu
4fbpQ4o6plArAb/3l+Tul+2xYpKj/w2h4/OWybLMuJtOUfDKS7NRXQZ5jBCbI8/X5mIPDXedDYdX
yAeoasHMAtfnkmksDlE1429mfLrrbMNbQDwxEk+ULsaXyrnUa9vNrbNgDPuU9Ax0FtLGP6M1vKxS
JFq+SKqC0mWJw3NSKCnP38KeHgOC+g0Khqux6ROY4yVO5joYUXG0mMErKaboKxmbfQJcQLjFLCjO
lWS58ahXRSrFNVd0KXl2axohM7QKEvxjpT+dXzMxGD1VjN/cQH+jzrlt3zc0QzqKr7zgox6OTlxz
dzxk9VihD2FN8HrzHkHjzXQ0r7KKeCkanm2OPiR69cIg34CizFBKZqkZbdV3ihgwt3IsR2fr5GQg
pa05Y9gr373HMtliz7+rc4J/NZgTge2NelTjTrhgHgc9RFXCAy6dxaP6TQ7Ae8xHQdeYDYkZtv85
piXEMjNeXNuIgNvTg5V1zqbKfmzQ6KBAr9+7xR7FT8qdVU8nJICBKIZtEdAUxu/21wHFLNQk81P5
O7W9v8Z2gMvxSNiUmIeQbhFSLrUs/5dnEnssdNHGX0nhTBpf06K3kY64oCnK7m8kLPqxUvDueAAL
F2iCm4tprdodEjbG/zud12S/L9f3bH4t+Hogb1bgFXDfV95jqnPttEui+8Hb05/SGQpXJU/vgG9y
XTbcK9JGo8zGlhCkC1vXkLQra9473S2efKSprZfUHcYfo4Yli9s7L2g37XRfDqKCk1XKxrxHfxCR
fBVAsLnor7J0H/GLFVR1hQWGKHKUfIulbZpCQ0uFyHXRi4//4X10coSPVh/x6JsHkez+KS13vMLc
Jd3PQ/GmSJb/G0wd7uf6cyhiFyZRFImqq2atZxfsG9PNQqjkR6MpzTiZVNKyQ6JbruXoKo4vA7FG
SPFni/Cr5zLLK0g/j3YUsHSFpnlDk90aX1U8QEeBuZXN0OycXnB3MbYjDvZOjpCp15h+ngv4GCcn
CT6qZRjssyWHky/DL5cYnFKG3oD/vACu7ji9DhvliNR/zcLMxWjgfZY35ZlDe99b9KFWJzLK9QYf
81o+KXcQY+34/EZsLJn9NxhObL6zmArmQxLUOU7JeeBtvWIt6HcIJpK/bJJ+R17y3xiXxr/SE0PB
S/ZnXWvePlut7CyJbLLimgKEHbQiuMV9VrGnKYplRi/Fi1Bfgx3yoIY8iqg0qWLcvj6qP7rO+lty
keaoo0ctBcSDL+0fkLoYrcibYl5qYj5/8+pXTAVQIrsnxtuV8cQKMDK1VjltBM7O6Q7TyuE21e1g
sV+vHWz/0fO6xi37OsSbZKwuwRCESSWFsEJFKV5ZQ/08zsOByo8Xd07kA1g0+naL44noAL8FDSlT
fhs/IrNYr9uSuebQ3WR8aWPGqvLoShlolEvF/DoRLAH8hDvb0gu9cwxETkOcy8OOfoWg89CH27DE
Wz2jbuIveyU82iX8ECAqxiT8SdwUM2iOyK8RsPiff/5KZQBthRvJePbRb+Xf1vL/VVft5XfkmTtA
RNicZpfk5iOOFND55yATSwsQ9ympdF4zynX9ixhaeUD3vVje3KU5eLv5Ou4FhHf/dCeJDjN8YkNi
XLNbk6/ZcZlzHmMJQO3QdBLd5ma8P62kU4gK1jcgqBnzRjPRuP/kkl6dNuOPUiXLWSte9mys6uMR
Rpp1sslX5LkOsDf6/hvvvF52hcWVPuqPcvfwEXZqi/FYzolBruXvAnWmIAZtsm1Zh6DXACWu74x0
N+Eg22FxP2s/JmUNFL80kYjoJ1mAb6BS8CC/zFSWsCoLzR7rsb3SOoVeC/N+L6PQxAiln91y16gD
5NnkUVcquDha4tmlfpbD1FyOl01lIvVFL45VIgmOyD+A+pSa+kW9WrZkaxSlsLa0ZRS9fyEEcdU9
yPuVj2fV0NbFWEkeJqPwuT1wEaAwSq4nlXrY7jmacz6iiDc+xFBcfA+bTO3GtNW4zp6j/2hVEwbH
oQX8PdHufz30JW3pbZEjosILmhnRyy4hkkGyWv8nKHqiZxP+iK7J4tXptPqZFJD58rwSctxKuUhY
/TK+uOGUBB07qVjg+i8gAlp3TvACTtaRkQjFdPAwp749gwehsBAoKyrueqAsuh5Xi3vClvYKzjDX
pPSMvOK+yTmGRDTaQCERikVVbYLHGpdRIVoJMP9SYEOFxklDBHpJs1wq69K8s5KFpZ0lGM5qNDyo
ySJ56GJ4FbDsnWAoCQbx49qP7EqCUjhjX+56MgoA3d/O+NrvaGTcjqBXur1AyMOtp55j58MXm0yL
stZHvnpbeP0gy0UCIEUP4fx3HuVaqe8f6UlRM5hFMWwUrTskWOV8ZC4Z431Gbi7aF8tTSZ55sDwL
H1yXr/0HXRWs/lX01g+NU/iegonmjIj1+Ux4n7iYG4/zafVn1GQo6x9DyJJD7ggDtN0ui3U324nz
X+QPDRWWOkbHyXsQTKbfZRHOCMbxoM74zxeVTl9OOssc2w46rtiJGsOCG6X0qwFG+7Osomk6kSVJ
PvxRXLsdQnS3wwDjhjP81IDhQ26ZSSULdz0IWIcZH1MK9GTXI6+5HLVCzrJDG49WzftkUMKYBqw5
LVxkK5UQgxPvmdiKLlhepr+cgCU0wZOelNaVEDslSB2fLvXQtEZ2/JLGBbWAPu6CRW+Idayfi57O
2PeMugHMM+I1r57Y+iOxrICCtPaTImX9aPXuhh0kFpAIyx0HcsfKNBNbTaJZ2z+PUp9SCNnoLtMo
OtcifRSBaNmYiFOk3LAOBR6pld5folekWi3xdBZ9qDJJb/hd/BNH4/+liVd1zOliX95mxKTGJLsq
zXie2EdZK2Y+mKnTtgrPxUblCd3rZptnvqBcU4EKKX+4ETiyp1NsCmJ31mce1yeFW4vYLGb6bnY7
hB2Xt//u3OQYsVdFKsrI9rn3+tCvoqd4LMTIT9O1ZTsMRnR3K2Yzp/9VppDUvOrpVthKONxU1HAv
rDgAC9Gx0RL2TamjHv0pWWB+KvSY6UpT14OYzJGfZWJOlRHsICuMJHLVPJblfJGScYzZ6cZRGye6
+CjLGmouiKG7c5Qekcuzy/1iFhi7gPQLs1egrIj0y8HhhOHpMxaeO6k71OwEs1wm/N929PWasiTs
XgYoG6y0cDfePFCYZp/hU5fdMlq7+ZpukbYu4Cfp4zAtga+hHGPumIDjhoy3MlB6IrJa+0LxgjeA
KwEWRQQESf0H1G7QMHKcr9ZB/Qddk7Auc+IiQ+A0NCsG9PtVKVFODJfcOuMeV1FD0LMUfQDShn8I
Hc/lHl/iG3JDFmCsdQq3GGaj97jcDnX43oIm6gbbnuf5hbPH+YtHiYV6l3RuqM78HRl5NnaOAoyI
MtLACtHXyhZc/LU5vC/l9w+kbBkF9QxufHnojzqrZyiIZJsKcMIS0VTl9aJzrxBB96rIQf+c+jqK
/zaoYira+JDb9gPgfBRYkhVV4yAheoERrbfrvQn8uknALLXzvyynLzE6yRq5iCUA5ADeoeS5irJI
ECQt98FrqujPjBddj5OQoqUK2U8H/2tEOcUDO47CmcHN8JM0/DQKl+KZTI8Gb+FROH6xPqYf4PgA
pQsPz3M+mlmOn01wk4vEhXLJhfBuuU21fWA3ARtisflQSzFqa+nLY9CcwCpSQGS8WYu1WqblNpzp
wCz5TO8r6pAlLyUJ5EWf3X2F/Gv9PcyARIC2jslIW1maVU5CkbiuaZ/nbaotdZ5IKyJVHPW09zXO
vRngSzqvScJiJ71sy8Ym9GEiwGqBqC2tEXTKAwOWjpbDnWlQfGWgirjDgeAog+n2IHwyCO8Zbioq
vZqXwFk1r47+ZWWSsQovS/bKjmDm35xy71g3H/9RCzwIvro1e2aFBStQtAAE2mEe5fQlexSQ9WuZ
O+m6d4YDSbiIhE/RjyUHJ5tYC/zgYGkgBHMADjZIg3KdIi+cnP55zLKqrgQLrNyIkj2vkXS4IlSK
h2x9ZKBeEqgm1+GT54GsqhC39Bi4W5P1FjC9Ya5HblvkiaUUrUc7CLzYMLuTnquQKbuM1sBl0kRW
45LyJjxD9FWe3yCATgBVt34Ts3gQvE/gjDNFuldKlu7VCc7b0xzzyNsZqaadlKeJB1f2zvAxBvTI
HxLbeLN9okkZ4Wg4UuwdSmmlT6z6i9zmQiOBftk3L2XqzKrZttEGk+goVcUgzGViQl1JiRh1+Ysc
3icjlS21E2Nj3shwYMC/paUqbMSw/UENyiBeqVSs8zBpvoJirmLMI/pMa/bJZQgN+FrnPhPqrWyh
ZAdz5PlAxEV8gVqfm8ngAPEk4Yhs+Q5AmOwBZAEPER1u7AePPLK4gDvDXSaG8bs6t9a02YNrJWSn
oRsr1mZ7DQ22vm/7oGypTJCyaHK37QLvK2KmEuTZW0EIVWb5zRs65uiOfDFa3W6drmPV+j3Nx04J
z5uuCKCT0ulN/HJdHGRaP0o+OS7XYBcOxcHIxmMeJk4/V9ysBMTzpcx1Nt1qjAnp/9JApBH26CBa
2Mjhds1Zd2GW/D3AXMNfCAtpt8PuA4vviYdmpyOHcDlAexn0a5lDzKiNxSr+AC9/VdlZ+Ew80u+Z
MJvY5O2u7PfA+GVk9eWBvMBNI/WKDxQNN9eSLb318CeiRdiFAChUVWy8tlZvYUy9vlkr3xZuhhFa
hs37tjPKCzGweJRpbVW8SwtUARPcxHU+5jPs/MxBuqOpcW8yU3bwhoHzg6VXC4uCVZGPC6o6HGzc
M0249hBau53pgF447fKj5AYjApgGHJnJ1+7cZNWOFOW7TDquxCp9HLcCEyN1X8LVZ9GZ3obilDP/
FAvGE1nP9YM7OymDllnGUM7eatL22169S1O2XTsVxzApgbqD5K1BaAy2cEGNsHUsAzghvfgnZAc5
uaDzNHcqdHRraY96kbJPlnivnKubWU/TCdsFbBHJSf0uNxQPjxXy8sokXZ+MAkKpWohPAmxoL8Sn
bSNRixVDDgcJ7/EQ2U6Qqd1PImdjlprtHlbENQn7pfppD7OrHK1CnQX+oMZFAHhxsFJhWSR4zkh5
x4i7dAFRPQXF1kXe6Xy266lD8VpV3B/TLFPFbJpXCurjF4Zhq5DYgKQcvg8g1b0sD7Upe24lnwUR
nJx0spv/WHZF7LkZZmTlXeo8pWZkJROUqIN0r2JJL2Z94BRiVFl5IziNlXaEgksBE+RdNihSFwC9
/uMzt/BbvHBzUmjN7YyS8BIi/Z0spaGp8EvTMTzgwd5bUDTAIf72872zZbiIR2dqF5qWnFzpezE0
NcVYN+48KbWlNzR3cyp0nlVfMz5PPFxVW61l+r7f26ntftRbM2uxOzwOudLgCRS4yeMUuSbWqnRX
WtIYeiyafy/vRF63WC1ePRgGvuHNe6rWjiYNEj3U8Wg8duZ5ob3BXwtoKluWi935C9pcJvOhKecG
9l5ShyJe9qZy/8FFIsOfUM8eLktQ2Wgvj0ZQn0bci9JMQpemtQCNLVu5QXJh2djeJvSnV3iIRvdB
/zk45oIa1XcfPV3wqQoD5STxMo0liw/+Kr5Lw7G5wBZVTb2/K6KGBZqHlVQo08g6yQBfuml31+Ib
q3vVbaJ5OWP38koL/hydzDBI7hMwypODytsxmIizsgDkC8nMAowcUqr5Wb1y0ywGuzxVzws9PCm6
rTJR+HxThmsHOZqTRxWcnWN6jDvPTtZEYojwQI3XhLEmOkS9h+tLAtQUk4fd+OtodZe0NxhCCcWL
+cjqe5zrnoMggHSFMDQL8nk2cMHsXQMrQS+AxFKdz6fb/E77pPj8cnJbtkQqqW/6tQ2uasAxZyYg
2FVPxyfpsIlzndLHBySv2V6DG7OTTbCMd3hDKKr6gHAy3SMl6Teye/s54si3UVdeiWjjIS9CKXXh
JhA5qFAfQoSRB+xDi8Rtv0S7sgy/NluwbtjUiP/Byv5qihNcH8oOsppNM4Mgoo2aKv7ASLIYEmkj
+4eE+01uAV4klG5gPPqVYIJb4UfMPNmBU+gf1NZghBTMuqX3vCzqAvF4LnlKw7qgmHb7E96nbZMP
1CivYtc8/DLu6BvZnPCwBEHJTSifYUiiyKStcwVTMRxpqKdMQaukPMJYaloP34XyOXM1x3vO2lrU
WVqIPNQOPOIQSIP14zkTW7qcr/DtlCxSa98SDRrUveJH1aJ8/56KgrUtm8KJoW6LmL+1tkXSD+4L
7nY9LUJbpFRdV5HaYoigqVMqZSEuBf53sd84Jh23uoVqUYGyXuzKT/w9Vaq2h37Z5weUgChgRSUU
jIgtsjC49fRQ89MN9hDph3agou4s/i5oXo28cO3DVnF9GWj+Yyq3mnUDj+3smpYnECeK79v/ldLB
NkYCuD/aWKdbSIluGdApdF4RIYP6axh3tOLQWDivrazqtgCpWNJlJijqzVnbgx6pSJ1EDwaRUO90
KmTMKUiogBWCCmfHhDFRNoJCYmDyVS6p77Ntr621YFBkns92TaAx64t99YfJBITndDmE9vHe6j++
RVf2X/tJb8gFIdn3QP8QWkwTwCUa1p7sitW4VYOFPWBGbtUjyOlGmt98q/wVrFm3ws1xsXDpvCrn
UuortYDrvcMCyILeIvAaCJErA/7uPziJE1U9UgwV8O2mOtuZ8SxSplUWJF4kL2NeL9cxW+MAPN/R
SlAddQVSorI/8ZUv0sUtj0JlovGlvB0+I+DXNR+NvOIuo555gMqR2fVWE206KctQI78dy3QXcqwv
iu3d5TjdA/xLw3qCZv9GXA2L92GLRj7VAA40XvWDmOLxgROwSUIigmlqDL5FtjAEUgnB9eczyHYr
Si392NkP91m8FfTKM696eLVWAju3ZsIn+ws7cAhAK+EyZe7ybLU/P8qjvUyeLUXq3cZaNLjjhDAd
WV4ngZALfetNK0C8R5LxAqMkgP5fZMu0T8auu+HeFwjdrfR3xHps9WcM9B2+d7CfWsMayZY4eOfj
iLZU885v5yDAiNuAL9mxh/SwoAOCeqVXXTjjd3ERKFZWxeE8Ks/LrPzyu2atfPGzRE3jOqnT35EK
EZpWUlypv0rGQvsLRiufY41LHAkMnmvS9aFZVlkpPNN2JlQNDacgvdfBW8HKi6CGprB4jaMnlLby
QFMHqnzyl+OID45XRnRsSCYsCDD+llGi5UOBIFhltUK+Te9LeMAsHyYOHG9bP6+6ynieFMvb4Yh4
WA9/Ch0AF/NTTnc16/O87rvnUVD76oC5NzC4GPE0B6uwFZWj9xJVB5AhmskpFrpv7c04eMt5/Tp8
0ukAIO2CB+Bc0niGjJqmTZLo0vzcocYURFK+0WRJgwW7lFOgSYUoh9tt812wGqEPNEtrskjYubTx
ugDC+1J3ixlPmFMXhfQoODYwEaEmgPwWWi4PiFe5gAsj9Q/DRT272Q50LvgCxhBYLLntvNzBswUT
iixRyge4m+yJt0RDVIZ/13Wg4U7zVhTCj+umowY90UJeFbORgTjEz9HFflnOMshUKE541G8OaU9n
GZ1RECtfe2cgSDyB80gUBiUN+nSsqRXn2BDATnvG9xvUruc/roMI80mQODKsx56XORBbR6sUnIhT
GuSyqPuBZPWS7HuF4SMDnQHfRGTw082jJjZa+GYx2fIwqPpdYhXcBvc88cFaYU6VAWj8tbzjwICj
24NG/WnK6Mnh8vWprNn+LqOBGEySsv/66WkAAF06vk59dUb+wDN0CEcaKV4aIbkQTyWhA0wZ3vuP
mObl0GI927x9W1Wk00hGIC3Jw8TWM/Mnmext9JAT3FtP1PiV1Xo4LAyFEEx9IzuRrV1p/0+p+vz9
0rwKUpDYVWcP4dtzTnbfpC6owaUu64Ci6Rrjsq7ZIQQg/8Ukuvd/Abi6Uzbv0cQXJaW3jkxlUDk+
O4/N7mqEmygQFORW3VIUqG/3cbEGQGvJCpB/fjjkTSaYZ0FAiPElEsz/Z9uPIGYItbIL/U4CGPfL
kTHCCjjNC81DCPMiMHEzSADW6w+MGyptOmaLWAIp0u5aLRp79S0MirYbooRPmQQMRyNwuIg6I1Sg
3ArpqSCd9VRfYiFXLozyVQZSpmWVHAxBrKKob4c4upP081myicFnoMhV5bFWydGsLMK5KHM+FmM6
OjbZPoAZ4kvvloGAdsb9p3ENQxuYowypw9xDpEcq/+XR5uSAWD63Qjgi90c594AuShpDLnRzH4o5
bfEdRb5DhIKG1BQABmJ1rBhg2eNK08Xbbbnwm5LFK+dI/h8Pv5jV4mVyp8zWEpLCiGk7Kz5UAUQz
eElZnaVQ0Dy3Y552jIn1Gsla4jfLGqq0zP7IFt9b0mCHuRrmycIx1HwveKretLSBXOzCwZsoHJn/
bpJoy0L+NkrQ4VP4mA8Kz+WnJc+p5LbrOVfuonDAkaVqxw1iG0xhxZJU4/Pxter5B7EyxX9nmIBT
kur6jeWjvUgrWz8JUU5TzIJrHVUCqTBg0okF99VLaFdpyUtPJgCfLjvM+9MUDfGCjY3JnbngT4kg
s5NmOyIGezLBeBIaNPnPQFA93Z4MmuJk86TW7uisabBm1PR/Q0kNqbgi6thxo+W8+i7TaUm/ziJf
73srMIJ3SZzrHcSqAapehWNhF8NyE28gr1+gXPva4Sx4CkwacBkcbJMpcHFHT3m/ZuAXbDU/aYBW
2zitbLr1hMKyR1AHZCkxqjtq5bcIwbr6njKIEbjDW3Ewa/I4YziiLgwbLeXsgodRXIOIOeHIItiY
X2v7lp9iCNJkmf0HaIJjfnrOi/duvA5qerTH2MzY7L127pBvU3Aq0y2KUo0miRNY6ms7R75fvipt
fviRaMAxswKOb/zsr21fL8lW28/yI9YmJWch1J+c0M19+2jfND+NTwAZRkLSMAz+u8bkem/meFQX
gDbzbWuJxFhWA8OoQfUYB/9QrN3poLa6Qfj60piw1191an96R9EWb3MapJ8+szW6gNLJH0rfnqx1
uVsVXBBbJaMhB+OrLyqJywODiSC+8HxXkUDUyIhPrE/XMgvNpYBo9WXKnDF90K44escHK+8NugN0
gfYso1oGwDj50ODeZiOHagyUDjWafNqrna1iLLmwi1ELhLCnxsmCWV/FkbJIvSnefJEmlAKPh/Pp
2AnNIpR8amsdAZuJ33FowXegm6qaXHenCQWRHlL8rrYPZaxZ0pPQNbmsLBlovZw+b4ZSgUepN+iH
yL3NgXZG5ITThB2XqV0pDVmkAGdAGjjmmilt6FTDGpgpf2FBKumc3wkk11TphaQdaxsd14w4gHXZ
BuLKKzfSctIS+nQYAeqcWNAN3SGMrB3SiZucrWSTGjGwWFWgIKXsK3bpW7Jv1aIJLibmouJvpacE
UU32WCjnmHY3YYLCUKIII1XsflbAknx2KRgoxEHk5FN1Sy80SURQgtQtUpBZv0pdYEOcxNowybVX
9abygtdmuDtUmM9DKsR2XrMSGFi8tUn4rGOa/nJ9BrBSaDGcSQ3XP9xGkHBbXA/Uwevb3XryMzBE
BZpJuikw8Ozu9RqlTJyYOv5pbzd07LjOE9z+o23j8fTJM8QIH2Oh0blUXC7h3mGOLyPro2NQElYD
YmGwzpZhn1TV7vFxhs5dXH+6PAY6qOQUB4AHPLSp9V9ot6FOfsRLxmhWuH77eBErAJBo35/Vjsu9
TGO9llwFVP27wo00+aaQpvAjalgySQFSXc/UeuLVR5/mPN8Q4CwYfHXRvDBhZtcHnL3LMUUmC5dY
8maxDdYwWW8epEN3mI8hP90bxGHDPIZcrEVIoNT4ddWoFYBPbGGrgEuJwhgfsrEOi6I0OmdCnY57
NPdmuPtA34yk060Lp7F3x6KTNv+TZ+x5j2Xew+X2BH6FXmwFwW46GGh1EPuXBLgKA9t+NjlOMYU+
CJ00BQfMKOd1XEWain5Uh+Opb69J1WIMaCOPWAV9uaq3KR/Bu5jaR9l3a6dT9TY7oMxH0fiz2GQN
ySnHe2iIi9iAaxVDk75J+2YqWOnK+pyA24jZcg0cfhgFTig11CkEkM6tZnFitC0LfejvB646sLVr
9qeXbxehVVkZs/Lac+OHAA+Lj1Bi8Q8kDkAt9Tn2ej339QzYxbZAn40g97gFxB8AhMPe24CJajmV
BDrxiolmM06vOomICjOb4zleVeAls9g6L98ER49nNn4BeBWKeRLLQFBATr4irBeMleJR6TmO0Pz1
V7tyMk5VBxWKWrkuYjlch1a8OY0CF86Si8ufdNuAT3dkCZ5JkHNOrMFXDVTLqoykwqgslLeYMH32
XSPaCXLcZEH/IcF0UJFDVAQtjC06U5LrIvoS7mWn8WKHzr5MI0/6p+UdQkTSG3bmxBCTbfZMZiAJ
bhlPYPUnANGqJ5RudeHiM4ihF5IJhz5Ek+OMH3aBNSxQPOWUWB8S37vGf2bt+0v+iEGwNo97dh2j
xSzI/CgjKLVXpY2RZqnVW2qpfUdEakTFiMqZy03QsxGjuWsBCoshTyObYGZSNB/W4Oxvs/7cuMcB
ciPaOyRvh4P44Vl7j489dAxzQDOskWW9pTkK5V7N5+2nvKv83z4hLfVxYNpuQIcxWIF9Zc+9O9E+
pwcHxTlzwCJZNQbgTolA/l9730Q8D6Yg1N2S+27k42uL/sRf5nkh3KEtaE1vX2e6yBHXhSuGHEFS
9valweAtxnmpZHD0PiuwvfvhDnUo3+7Y95nWLKxc77bI97+YS57mJPIcnaNQOEN1aApurHnepnap
M73iZ0cRvvRCdudSk5Kse90uOHb52tKEArqYU6/H457oDpCFjIHRgKvOX4EehS2euK3RXs/ov0Zk
2BUhi1LiVrc7VV4YjFATIJki4v04gZbbbRO0IZMo8eQiJO4YRYEPfTQBcIzWSJhnX/npWWktnXam
hV2IHH7lgmM44GjrHR6EP658TIsuw6NImTIqq0lum0t02S+Sfs7I7OW/W1f5YHUloBOLhL1HgpDd
pHnsNsUxbZTDjBs9t3fiaJn3Sb81y1B6QtKtyTzQfv0ePud5O7w97iCcdlBKrMdqbhSF7NSq2Aqi
TNV2eiImWAqZl74pBeykfwb9cuV5i1mIy/KSHo0L8VSJ8wOumNfAmMHAV1rVNFrvwafthinQzjuD
4HEkMH1HgsIXt7JWYKGY57YUljWWxTq+b4GTsCNzu0RQIj2qp9CP5aB0fRu4E3EFXmWJFC//hkFz
yIj94HhUezZicXRUaZz/VG0/aw95g8WyddHVxcGxMIfTCIuVkryA7GnfxyIO5EbYx5mNcktciA8b
PVKMMN+Hc2HP/SS0yPRdBkENKKS3uj5ufe7m44bV39ROZu8YEatoITiE3PaJu8mUfmkYzOQ4oiHO
o5WqqCzo4QIU45vkfVHCRcnPvnjL1SXvvMpKkqVLBJ/KLVccTWeb/cMhiKkHUVZwZVLjzPyHNdFJ
EaIoiKm2hKJk9uv7Md3K6z7+EDCvLR3odp1dJGNumFTsnhFp4caVxw48ZkkxgnC8dWUchkjb3IiE
8wB6g7dli+Cy52DllVwuSF5foPpyggS/wh/pQiDTGRdzZ0Brs84xg6oq61K6joZ+Vdmr5RhygUo+
pap/Oqe0QonnfvfziSQNXfxDUtRCjH4rjBiOImD9mMGnbswxHX7R5Mi+CnYjIco36JRcY+kVAOCl
OTMH5n+8uTEXzku2JljPU0qlnU9g1RAVqSn57XhPNj1YF7WqX0Ggw1prJk0oKU0RlSA6te/guo6z
/AuSrnvUzcXGggY04Mr7F8S3ZkPdxoflbNRMHwM+uwSZbmoumcda4cjA9ZDUg6swsZr1/UhzEzOT
dAgxmXihMAvcPkoBUIUjw124VflXFO35hTKJB0gHNh+WhDWjEJ//ZDw41EjzIzaqZKjoxsT1av9C
avJw1DnXG7wFAB74TrUwv/x9A5HZLEIyx+3PaDwe9QMkGp7+pmEKpAhtVZxMTq1KKNZP2jJVdNas
PkJj6ukWybP6Epjj/wITQRV3T6s7HaJs/abu1ENspKiaj8OWe/bpwWN7xwbFMboO5CpjvsHVg1ix
M8wLjlPrPUAj77i0twBfGSJZ5ug1ETbPUOHZcYHFjGywcIpIj7t8GGSUxFZ0V3WAjKHltQ7NX7bA
er6LAypdbWW5zhmXp3UC7DfGH/VGxo/zFAYRMNzBnIwhQfPa7AErhogoKHvtqFNVi1EBsFUZ5sru
X4YjWItNbAb2YOfZkz6TGp33N+pt956UeT78o/y0NjNKktlUT0txogpT2xS2GQs9W06yRu1XR7ys
OtnS3SVjdPe2vJsZ27mDPe9+CL9kZO9lRfulVXTYk8X06ByUF6peJeItPGBacQBO4zTU/gNC9w+m
E39VntaZ+vHupJjV7s0xx3wY/3k3aBDETjvAoMYdCa2z59jTX/2qOWuVrHJeNA2LUiNeR4ScCLgL
wCnryc3zJ6mKFStOw7aUr371RbHvCsuAeOECW8vGRuM6ntyfTUeI6qX5XStLWMAlF6z1wONH63rv
2RFlQxw7+Svo3mCjVKnNrq5h2vgckyIdRfz5Yc+pZ94sI+kYK/vbfXsfWxchEZlOoZwRc8VRyN8L
ZFosbOCck+96hC5B0YEjchzLWOpvza/5FLw3SFYqPVbqw1Ox7G8UBOUkwvLp7jOnSBi3SbfO+t7h
PzGgYXkci78Z8lvJKYmMZWGcmK8WtLXrMAcy1MIShky2QMoZWbqp1YayHaLMiP+PMNhsDhHLmVN0
lGFGmI8tkLC7Jbr7SsKEw0KEdUb81eLoXs6zw2xgM3T9DBrn04G1IfHIZNCcfAREG8qEKn3C1Qjc
DZuAXWAHNmL32FMq2sY29KeS4CZ7aDEewEgWW7QcOOFdZA9ntYNyh4sNsWmsIvzXquR74AglhwRJ
50az8/umpjEPFJgVQusL+4pGyfgy+VciNlbKgJ7XwgEXHdd2yqHaIkA33calw4O+trPTjNvQWiDN
javhfeGcsKLCv2DJn5bQTNta4w/9eIk54tDLg3i27tK1iwxvHnLEhv43bcL+cutlMDrwilk83ZSw
T57z1ZaDG79ZYCHF0PQ3veGUY8sjL6AJ6BZSWl33VqTUZy0y1UQYVONQdqz10E/M1RPB/rBgkxMz
TslcWBaAxsUPybPhl+nspvQ9vo78gwBsSWul6r78m9twECIofJ7a5JeoQvK3Wu4cRnwtvpIptl1G
3Nlpa8TuGKrXop4FKTqsh6YGtutH/cgBK4wTJQIGcoF8JuiOx0EwuhCZJgeZAeQBG/Wust3qanyo
pJouJF5ztLtchPSUaBXsBWijC5ucPjXqw8ff0HMRxZIarEEhQAuFOPXtN4F2AEtqXjoGyK7n1XB9
5WXz07/Q+V0kM+mRzGLOdzxnmY9tyoQ/XTWXIimIv44Y9Xgf59P0xnlyiJ+dnvLAIaxCQA9GEKaa
SkDRnuhSqDdkMzQbglWCMCJmzrPixpD9PieQd59Tp3yMmAMlZm4ZRNxddpFIYOkuF6ld01tMeYlT
v0NUQsreGcTa73VP9b7wV4ASSvJFpZf3s6kLHfyqdZ6hs71WKGCPi7yDyXypfc36w6Z+WfJ+bgXZ
wsAlPSrqK8a6LSlxGkRdkWNbVjlplv9raewOlAXad6CA/Zx3CZUCRMbf8rpE6zG3cnPxM3NMTokZ
SaWBVWYXarEOD7pmC4c3SeOdt5HlQQr59mPYWzecUc8J6FAE9M5hJ5nURtni0Tc6bvDw0eaY1j/I
DXZdALkLGt/Bdk81+8njZMgXB61Hyn65YABcXi/COReR1t1lX1hhusK3lx8QEna6q7BK00Zk7Yn2
d44XgToKP1uOKyXrlgsFl8M1SqqDc3hxDXPZfUDLs79K07bgYKX5o99l6kAVQS8ZFQssRyCdhgD1
+ftI4ZZhVjOHdwRvjFQQpYhJ/IMH8YvRRioeKP92FRrWlJuQpnIali+Wd3Cx1e2HVkv7nrMqCZaT
+RVZHfeT4I97wRuCT0SnSjdwR+yyMXvmzpI4OoPoerStzUyEcBcnZqbEW+MOv+Q6QKTwky+gCUsO
e42J4fkpBzwNkcsNxOKdhTUMJUDiOS2u6Go4PkpyrJ3zJ0cxMvndsRyz5/SiYGtJTM92d5maca8V
MWtOfblMS+PsbS/Vukxizal4xSw337xvoRrh398JwugnHy1s88dGbBLiTkOf+k0Bh8gYSiNmFCvh
plQkM+k+CDtjQB78cUzOdNySGm7My8oA/6WshO8dU2hZUMmIAvP+MyK5YTMwtHkjdTWJkdXJBtul
M81GBNA65gmlBiF43GZGJBpFhvo0NM3qk+k8jSqDzZk8+NTK1PjFfEG3nSgVgdeqbLDndocxgmUS
PN+w30tBBF/dNcfTb/i0y2MhByDjxMYSLV3G5kZMd6QpyU67ZzVlkmEmotfO/2PxZ85VpAU1AJut
PmlUd0OugTyL0Rr76iTPicXEi5Y41SLs/Lm3LBdPphiASjcGroMZBEHSyiWXpxWbEZNUUfDPAJMj
xWAhGGklF9LALQcgBmxWDgOfxzwIzAkQaSVMG3G+lQvkwAvqC7/g12roW93u81hP708Ex85QqxRG
Jp38Cjyq09h7IS3VCsk2kJeq3cg7fdH60WgHodddz/Y/WV3huMbQF6x0ubUn9wUfgyfIogilkTjE
0eGL9W8aM8UrJxToam3R7fnJ4ZYoz9zwcsugKLxT33tNRQ/DOQwljPQMMftsMgpR/0fSj93eiiax
zJjPo+vQjDydOTvL0UVfj7iGuHNdN3+46rQHnsXh3WbAzhTW5BODr94jtEk8CwwJbwy8Yui8B7DY
aTKik6VGybI/6mOHXsPI5mUaZapDy94EWdGifR7+NuPctvAcz/EDIqHazyfm1sULjLynqhZdNOWr
HTi2rNJ0YGiX9p35nAXy4e7LBFrrhxGPPCMeALHYIH0QiJL5RYDQz4cjMvbE4wWycnZuvnmgLA8V
JKzNoOnds8853mNLduhCU9F8qM1kEfNT78UkGvXWERjiZtP8uJ6Qm8bftI1nQ7w+9uOzT2m3sSI8
ZO6KzIxuplWlJifpK7FbCPWZZU5EZJer7NFowFOq1dJMbcQ6VSRv1RfjP5J7R0jRzDfN9ZGPO4kV
pxfmX+y8F4X1um60rGHEUmLGAFMl56FPOBBlRc9P1chGkhZyDbjgImkVjRgo1DRBqzCA0iskvWcV
IjS0i1oGD8WGx63gaSPLxT8VGChso1n3HLfeWjfQTDyuOR+6tpfvW9+0/MPVH4H9VilbZr7bUdJe
nbflNfbN9QeH0GF4ULB5Djs/6fl8obshFrMwZ6OHsa1PJXdSUYlwLC/iN8cbebYDrbhEH1EjIzF8
A/upewTWY+p5SL8b89XsiOetpcncbpwRWxmF3hUmqcUrpdus7u6dm3nVOibNM84QZ9myqjTVE3J8
3wRIQnEwsrv9lyLRKj8qJn9FSyu9Ja8x5BL83jUxH4M0ORgopRGZ2vvDo7S4BbSYxiMTEj8pFvqO
jBB8x/2Qx+0fHSmcH4Q0vvecUPNbYxE+YZjZkTYTkL5pAdPBC1odvsaXUdEl00CJVW8jExxoawOD
U4Q97WxgQzbg6FSbP+r3cyoYMpI85n2zVazirF3zTBJGQ2E+pahn8dZcQLUxbYlDZYjtSca0cNgy
w2FjoCYADQTwVEobbQgId1v7aj5r2F/6FAR/c2sjzRRuj15o6+MPB4GzK+1VVGO6s2MZSKdPpHDB
r7vfXDB3Cu6ajVuMC8GLM10Q5apuWIhOU5PBn6ryFWCl0qCTIybHwHEurfFVetawC0y3aUBCDy0H
ovyVk/0q+MLCYjsr0tW3Qf69/pTic/aX4Mg2wFpSMjyZ43vhxc2an6g6Cyd9Z3b+RLoQgpIcp+zU
Vwbe44FUZDgE5s22rJypoRW091oK9E+XL4tLsHzdLFeEUOGS9WE+1jZyQLTn1VPo6+KZS6VUasxm
+5VGT15mRCC9+Juf1z8T5GWXOvTiyd2rWAa/UNHzzO9o5AmfvunQS2pU4pDlEKsYngXcRZt9cn8Z
UkurVnIm+7eAjhpPA3MrLbi19Xr4Vfv3bYfzCtOeNEO5C6cXbAggW1IOx0isrwPpGEM95VgOVH+r
pMBEA1oXWP9X/MGvYlUEkmZ/3s/OtzA2I8V5R4irFaxQU3+Tf46GsfA14tap38Zazo7ZxkVf8ojR
HPkx/irf1mrdo8FxqtbvPzcqcJwpcktfbd+sSAlT5y/iDRV/WQxJ7ipManluAsGlVHLpUDs0XtmL
Yz/DuBMgffqOe30yWw72i5b0ECkFF+RbJ7y/9vqytpWs305touEZL/AiK2UJQNEkEeAoJyu9W9Gc
sgltIsaFEm2+7hlYXn6mK4SFyHFNULUWyQ4owgLoZVzHD0iAwx445ODh3SfVbDB3W7ui6xZ2oI7B
mON7yQbTsMHB4qaRmhnxo2nOCQo4DTL+CmTQGW9eob1qwRf8otlMAyRUl1ctiXEhKsqXuADpVrJa
3i2tPLnqzhv4Jfh709iHXphLYtS1M1D7ff8qkYgLLUhKd0ulLQtcgWbiCYEGrGyzs627aL/A0TO9
etMXtP1362xlxomiH25uHdjrxDkaYGUp94slCStXPEmVpYZItT8Z+11PkDZ7sXTsyLIkheRVAYhe
0ayouYMH2198Ug+ivsbZtetuONvfbON1IVc0SotY8Tbf1AlWdCDuYApFyDnlpqlKLjr4977Q2NWX
RzmsapOw1shzvkpDvFs1XIiLQzJhYHGg0bocY91o/iyloEMu5E93uwJhSwr1blq5+AEAKKDIxPU0
EeqKhlTAKQ4jE+3RKY9MbbFkxZgFsHcVoFKNbwgaTX/84IZMAsachc0zeLYxMZmTZmSXEUpY8JVA
uJ9e8zPcbJV3I5Y06hOfiClu8VMimC/VeGLH4jTrIXdTjMe8L3ndmejkbV+E6VTmnlNw6eUBxIL/
xP311TwmvG8Eh1XJf3DyksfcK4VI72clCW1XjLiaQSc356zqTq9cVw3EorBvkvJAeEw6l9ZiqFPz
pyJ89oCiKaqMI11hlbtnvbkcxQ3s9kPQuI1LhUyhaIGTMhfwU9MwxUhgK+Eqn53mS1ZDJmjlZqNR
ctD5oGZ43fLJ5l5E7Nl6cPvRBLkKuj26r6//pMOJmhuubJ7Wo91ZRJu+5p2YeyoNOA7JuB7fx84l
+w9AiLyByhriEo7kUW3ffl9Jr7IWceRw0m85JevxrLfbEwoChx4S6NsnbMw3Rg8K+SxYGj7il7DW
VOWRdCYcd/RZhml+DEEfTpXXRYZkEmE3arj06DQvX2j08Z9qWUjlJeIlBNA6NNqXUlZZJ25vbABM
ZqwR9xU3QC0yZ/9x/LsN+4uxlPG4d+O25qINHrCfP/tSEbN/9TYdAbCFYyXYmlcCVmA5Nbyl1DBJ
44pTwH0OplXEg6WycJ6Q3zZl0jQSkrhqsLo0flC9k2RWWdhtqN3o3jMvgc0w9LTIsx0otmHzU4vi
meRk5CpIiuIrXiahzEbtqmhTSz6F33eateVncvLxXOY5pwcscck0JkcqR++TdQOIt3gAIiL5hR6k
xIv/kcD6aRu9o6bm8+uFw3KCoH2wOSwbGTeEWbejsVsLgpGoP4CZ/PGlz0NFtFWWNdIX5T15ftSf
lSjJ0OoYYG0OS8XM4U0uH+nUyl6OQbB+7Z+tZ5ToF07yklBqZAFt9NjFXPOFhZQoxiCs0cN7lqtp
bhUO9z+BT1x4RM34RcCcX8pOff2+fJqz2qgrIPrErjyDpH3xh62TNEh6132FSaM+j0Sc+CRTK4UJ
ru7MO2lCNuczxZyUHLbUioXqFfs4eRYRpFqMjMV7Va5U5228Oim0oxMaz9idd9iGHO9IVksQ+Ciy
B9xnc77gX9hpjsOJA7EUucA+JFPJBKoPnCBfpOQg3lGsGk8c7qbqJ5eNq/ibNwpGcqVG0Ay+hTmG
qdHEIb0X/hE/01qoZoMgT8ZFrT7XOBlQCRIw0NHt1pA5hy/Co0/TLZmfDE9Qa4iJR02F8p2eNuPr
7W9am8ijKgZtSMs+Nj48JwpRJdEaQn6fPfGQu2tHm/mgckFlI/58PFbU6AYc1lyrQrBiroxFRzNl
lBkj5EODnkkMSKbABwWYeGFvWakcNr8u06TsrMqrQj5OQchGD62itPKWOPjf2AOxr492c7Voy7uU
o2RjwWMB9MAZGoIWoVfIA2/ogelo7RYf4kvxh5qiHoKTCNU/eF7b9Y0Q6Sro/sNb0/o4flyay1z7
AhXbp2g3OANHSz2JMoIRPUMX0mUrlBZYlnOg7XRR2JK1bQ7ERyB/I1rr/P8tJxvcKEPZSdmUSzzl
02wlvCEm5UDtcVLuYjq66sqc0NBWzKmJP0DJTf4Vu7WqRhdit6HHLO9fzW0EaON2IEIve/ExlWwB
CznWBhY57oiqh9E6EIDcu+E0ppH1slPh6SkwmIP5xPK68jWoSZw1DBbTog14xtPXFbh1aI5eq+SI
mheWvzUeD2Wdn6UaeDRWYj7RbUeQg+iwZR5EPCwE/Jp/cGbOEMvUpx16UaAxmACMhPdFyfs6tqp3
S9Arwp7b+YTon/LFT8c6FL1iAFIsG4ZtBx89W35vSMH/6SeGXz+y1+z25dB9HUjX5fXrdtsPQA4n
+obFDs+asrgjTwkwgp8IjFmX0NLdMB+luzahokdH9wdZYdfm3Mg3+/RZxs34fj5bFOhCStTQGlr+
GdHDCYWFG0KI6hdHWIJR/PfxIJAu4YDPYyQjWJucKAm83SO3h/ryKc5ruulaB/KKGvKe5cZwYgpO
s5lT7+MVBNUNFcrWOIZ/LayrI99tNuCWYyILn95XdNz28d+oUZxNmQVmZ9vSqUnb5HL176/IfGpA
YvJjlB/iB/XDI2qMcbKnsPmAwWG1PVM8hvI+/RY8YGKJJI41U/aqDjHY0/z+rMMd9FZOBVFbqz4n
4wnn+3qK1x3C7V9LxwWPSPTWjJnPhCwB2fjihmrEA811ut+TzpzBhZd+IVybaatTblGkxJf6Losd
R/ndFyNxwFZ60PIvh6l4qyTUoKoYmYhSOblL14ef92fVNHVHJ3F8jBP2rpgjGU4S51lN2jmVEZRy
U6L7yNR2YjjG9+o6Or7UuLEct63Ia/6OIbWGcQ8MCPoPW29lE27BETrqMgNX0MNjRVnwEIYNOmBG
ABUMGClTenuo2o3bLuvyk9tBJsAmuLJ7ojYUWOpU22zusPGBdBHqRIPl7W7rBDEAWmaOhfqw5A1s
jD2EUqeNbbNqFamOdYTCTL0EYKKwc/2ErunY02cJesYkrYuTOTr30nhVnPV5C7KTWdWORZ2rGdNy
WVPQMTR5cFU7noG46G2BahXtZUxD+FQ8cQ7jqN4N8CXXOEtgrBFmxeTgZaSWwe/IafOGligd3pwh
JZxEV4SQJorqHGDvODHt3tpS3TClcKxTUE5LKxNrp2JT3Kx4YiAnGlo9uQYkTWabB0UwV8ugOH6l
ElXC5eO+QhxZ9pSpbdZ7S161avJeLZGP7SNTTw7wHPdH/7apbyPj+NARJm9FyE4mgoaWRC/9IObB
EmPKccYMpqJFy4E46PczKNfKDFc1cDaZd7NMvYLbhf+vfAkln9RSW39QAzoFiNc5vnl1AgbJ19fV
ojA0sJHdrVSx03KANqn4FLPOo9bG3DaeNIr+3/ce/AclbCwx5WaBaLtL6v0SbyLhkjYKHXchXO3/
rycl8/jkRSbat8hwHw40++iK3n/ThUrywCKKmuoqnCE25KlrPsRRBRGnqd/Kw500AOn6tjjLx4Fn
Z5lQX2HmczNoChnyQGMV5WsjogNP7V5A6w09/DU1aN4Of+CcnRvHr0HOGlxGlyjG2QZq+J2IFnwS
t0e9xLLijr+Xd+iVkfuqPjhxB+dvrICBVnOzdOBjGo2gsLusYgzOUT5mbq9mEDHloNUl3L+S2tbh
1hoFVZfT6XxoYt1HoKWQZuq5iBLZgrUn3wsfAS8bs6UhdBOGJ0k845kgaeTbTr9MvolUcrpEGD3C
X90eCqP8uM00zhz0xL6jTdFUjDoYVQ044egkWFnozn0iTo6XdM0jG02mrJ2UxHZaX7gFoKjKlfzp
iLvg1QcMyoKgvBuFfi25gvgslpi7EBtaC/uvTjk23NzJ5Rb3+/CGJxmKs3VmZsLD48srjOwMDzO2
0m4P+kun+a8cLo1u4kRoZVyoZ3a45WFTYjtgOAxmzKeW88UcjE6gWwP67ep7R1e99r5tosicZitH
sXK+f8Fgmqj4W9PIOsBizc/Dwbr5adzKope4T5dOotCyrRuem9fZaTkT/S2dS/+kAFKzQojmYd2j
Qg/GfT7ByLvWRc+hu19iql0VCQBOEfvUP71yvbHpKIMO4GMFDZ2+//bXHV3xYSC/Dog4WvXHYpUn
f/Waw4KbRWEEgvg13NXn1zU+IrRuCc6LoIrVWJpwGsMzobzwDXACdxAQF09EoH2zrctgs8mnT/CX
R9f7dcFEDq9GIwRJ0s63guVCE5VekoYxyWQ8xoaKRhixfSsQcoetIv+PaAW2CMyL0GPxRCS72pTJ
i3ozQ6CHcWPTJA7K0hm7pTZy1GOv1wx7Ru9gap4Bhiy0VHS9y2izl9jVJNQ0R2grJGdNrJkIZ+pz
keIGXbkWMJwu3LNxkQdVUviOmyNc1ovINzXN9dONc75cjfunWX3OsHzLDxrXMJF7kk2/odbgbhOV
TbKiTWIcdSAWS2ndTpt3DmWm0A96YwLOnJn4IsoaCHpartpjPKxQ75adLFFVB2QNl5ujdPOCAVlW
u5fxRpqyZuJSm8VO8xP7NNuNb35bTeaBEjegHbvsDp8IMpnIn7x0bGNCeqAUkiGV1XChQGbkVUXe
vm5KMADy9iPrtnsKQASt1fMR1ATfFtGIu0mn8/iXtd03ZTQgm97O82Z+jhSK5TZviOcxurkCCh8E
mo2oZy6HFQ54xVwEfTwmpIsD0WRNg+UQRpuIr27cko7bX1oqQDBzpaNZg96RsDcv3AZJ7jh61cS/
61JgQhTlCbZL86xNxE1/ZgAQwYorI6LYtDhj8brgs1S+ymXwoJyYY9k1upLBuPFBk71awueRqXtp
aoOCxjLFi669QyHmcNhK0GQnV+OEUlWiD4nMiVSixgBSGHqN+3WAUQL/UPF5HKm94RFMHfMnJWr5
1RpEL5u3W23+NZYBeskRr7ham010KAyXPULaECKKk0yPx+NVb7PH97FhB0nFnD3ttP9kKXuvZL4T
waIBCOq7oYm9BJJHwP/25yHI0s9sEcCiQBvGhqKUe4BB5ERRB9IKLieKG5d5CKAQQCCVB37dnsGB
n6EIYkBK0key1wpS5Njmbx5xsm/tdI+hBbogI52KTXKj3o+36cB7TjFK+S2CQESzaMRzc2keVcvi
FxgWNGVWVkAKJCp3Kv04mEInhrHkHEkwu6W9YceuOc/JBhOpj3TqTRxANYaNz2oVfqsJc/XwfKl1
5aPYDSFtGBNrVTX3979AemPyPFZFaL4BQS7GtbSD2gHhFR4/pm5q2B+LbzlwkeeWlQw6dnlyV7o5
AywF8qsLWPXhnDuNQMwEn/VvRPyjYjXWSax1yXX7rDzKLGXu8g2vxFDhm4aXB4b93Uew9dWnnCM1
McLppFgWDFDYW7nbP3pChsqhGTNncHgko9rDYYeyKO3SKgHriOPi08m/i7mHfK6Wz/XZE3BFrWlY
o6nf4nctDmizJWXuM16FlR6OUsliVMsDsMga3CPQZi8sm1XiskmfVrhcJ3JwFGk3X/zqYvQQeVtG
hBZvBzOkntCZ755f9Cf1A4JcIGSbOttOmd9Ozoni4MBpeSPdNTRNl4zVDhe7nxJ2KZrV/yDltVJh
rt9gV0S9EcuC7GL27rDCizeuUuIZc/x07J96lB80b4SVmIZDWRf9iQDHHNaotcEqCJhi4yvI9ZzZ
GhLuYE4FeME/W/4mhmcvYJC9/a4wJy1NAa5c8vYVamOYIJBq5N846fAsmVbWI+XQYhGIQfDabu/z
GUtUyscNNh/dtJMRxN7FC2oT9cx5RMv3rY3WwBQ2RTvJ0lUli2jUAPc+F08H5hGjUazEvxM6+DPL
pARoXCKLC8w8tFE/zdQM1PBnLUld1nNybWem9V/c5z/SxiiTlTEx7wHZEOv4UCDYILiNUZtanV0e
lp7rbasNRxs4fti122sPvcWxTF70DI4YjKo3Y87LMCenALxEte8nQYIc5ot+12VwpY1uxow3XBhn
ckya1WYCZZ4SWly05VsSf3cYOkHUiCMkAqjmPu42RvhxgqISXl5xf0iORuPAKjsFP5Q0en2sI60c
iiUFq5G+TRVC0RQkvZyjSR0MUQGLTdN+zmhTnjQuiei/l8nAAWGmnAng6ux0BXCZo/Pe5BIoSElb
CaHfc/PDDkd/r+eX/+85aymvKxfvYKiJYNZk+yUKxAJs33izB0J3IHPx6+dVwX2joNunwBdtp0Xe
Dw6DwfshOD4QrFbpnhPVrSXN+IKPP/C2IZhLGfACulKrhz7dknNgn8nUOupgC47c6DUVIy9qruEz
r3gv+2IFS/niGroUr0nwrOybsaz6uVw7pE4sCoK8jPg2fGTkWGuGxAiWUZPwq0PRGH/ASCvVRPhC
0mOJ7XXmE0HCgxlrqWc4QuVFYSUe32BMlCgXgQU+t+3ZZbzL/SVwfeLuYJjOkdyCJSNBE67qfovt
fzj8YVXz9KBvMsMHC8DQz6EIZbSLrzuXs0dcxh91biE0FOtaFA/LcqP9+ne6ADfUypYpw65C882M
Kp3RYWILPZlETbA6tbCFiBVPZo6ZnDwQ8szbtQ6gZ/n66OvcFiTriB1ipBqFEj7b5U6y4BMszhTQ
yzN75G6qlEjWH0XdUDbIoypjfoUlF7x0SeymAwLuLI2AS50KoMgn18y9oP1241UUs4HFH79mBj+r
YVjxLlqH/qwq6XjzyPQcAIcLLsDXXBqC206AwvB543oj0B9pduaKS/r4b1+e2rhpqSK5YAK38vuI
rFoVHqaGP7DlKr5btekJBJPXPZ/e2r2PV8FSDpXjPul6OEqrZw3XLiO0ZMHxoowv2a5Gin/0F8zZ
zxcZ6VC+aXQ11hBPFl8MF4HvIlvjQCJI+sClclqY7Z2hwzvgX+9a/bJkMbGrlnL6Ufdkixd0fMvy
4HIPL64/b7yBZOSFO/qD9GGX5GAb0ARUH7qUylr8Letj8bDUb9x6gfYlSoisOcVTqOwQ/VltjtDB
rmQZ3CgCZ1hmh5340t1q+Wv+7qcka3FyeHKG6Jl3grk3lIL4hq4CN0+xSG4nOtsvUpsV9RgSmCdJ
co2zludIoazDVwv5En3xFegIEDXGsvslOIYQeUvpZ1uTjBlTUN3+zNNAHWEY7QLW2OeHZSFlM9e8
/HGZ6sjR8Jy4IXHJ0ER7xPLz18ahiXwAOdGXWzZ3+E0yRg+QtFNvy63BtPIYBZ1fBPh5tNtvkXXr
2nOvBvTsBqCKgFVpiDlWCa1F7OF48uL2yTCyarYmahDSJQ9YQW69SQR0Qxz4ZkYyoB5AzVgw2cgE
Pcpse7HpryJDcGQ08Uh3ydRMoI2fRjzRhgJcHHqpl2VZ0IQQRM2xPUqFqceP0+YleBOe66PCZ9Vb
n7o0VuPjLmFLuTmCFIacFtOS2GSLAKJXl/RVKC1wPx2Dh/EqnQbuJ+1MDZ9nOB4V7ji1sRCHWYLD
KXF60L5tNuVGsamf9nJ5Mug5h4RIbqVKx5Mxs9GfEcvDwioPk9Y57+6V7WEb8zQB9fd99a0BVurc
zqVm2PoLLuawpP/cteM2RLnvzfKex/utLbv7n1mgcGiEPZ1HXVJayFUPy5NVunHaHNFXxVCK4Jgl
XFedzCfbLj3kkJ2z8L5VNp4vIl9TXKYTpxR3367QkPqxuLFL556vSkfJJ4LtiDcdUF3/ZhaKnda7
siq7l6Umt01B/9pu2+Vlg8e4vmbK7gR611m5b2OqZPpSj4sYyhfDDbeXHIub6zEZvwevYLVyYJpq
7JcGM8LcDptkm8aFrOgOZD9Tnf7C5gJcuct/DTeaA1wi011z3i/QSv5+jN1JH54MQUapT+bwT4h6
5S/Qz4roZ0edSEJs075UeHzDA8nqRGevD6fh45DSQ83goHSs+bV9P7hnjHY+JFY+COezKpwCEkyO
9F1T7dQGJ4sqpZwxchlJhUnELvW68e4vL9CcFB8ZCSAUjn+7KtNin65xCpA6KvGykbt2YehJR/Nk
rClaZCpqvOUHnV6yZMWFZkEyrAlODNpc5y4eiBxHdBnzKY34j4ABYPjeLbbhCHGWXVO7bqV8gcpR
udJq2ARxOK33KocSlmoBBsaKeM5ZLWdkWKcMF8YFPX8RUbo9idaC1AyD5SqNYLIwb9UWgQsQJdH3
p4+AKxjgw+X9MlYYTvfgK+MHuN1oxkxqhCg7MjHcIZn7bZKYrXtGDrE+Y4BXmnKpq36k56MRHi4k
VrGbV7hsts63IusFHewp91R0RNpQg4TcZIQ9Hc60i1hloY2kT2plV8012C8DqgMccttFmN3mvwim
rBEYh5H8D2xJ+SOpT/p8jJ4EvcVe6sTMqMas4Ila7jF0M97paSHr13LGXuVSjoLXByeAdUKRPsv8
Jjiboj5pjVDDHWGX3ghp+faEIXwRHHkGQpDCHqYAaDUAcbIYzxwctTrYJoLLI5quawo5bndRzynw
iuKFTtyMZSJOFGeNL3+tHlmBu3Madm9vUPR6TwyWBKqrNxl/gPgeA9idQdKs8bI0rFRuvgbJB5Yp
FfLOblby71DF2Yw3YOO0cczpYVfGn2QyNs2NzqXODBqcd16K9PdPImAeG3zWuxk02WugPogqD6jV
Ti/B+n1hDEx2vxrY4dnSX1ka7kRYyTtFCaWBcPOOlRGlLDEHvI/ZS+tZC42qt0dq6HwYhSorG4Wh
42i7Pi3ptf4Ki8ScxaICKt0Pr/NuGmSFwin/vkvQItclh1fVoOx+gbSc4mIqGRdmSdzZ9ogQNSaz
LPykwspf7q5Z7vjyI4+b72oRn8fXbjwvq1JJjwE5usTPg/oKIRijFREsGoonL4kI/Cf7z5l256CS
EDzfPGbfMK9V39lBOxttypGSZSzHHxWxnfx98UyYcMyPYT1SZQlcPA+iA6vhZOPuYNi/+JTG+DAQ
iLLD9pgv+e4zdQQcZoX7hw+rcqhqd3/0u7F824ljECwwkofHYGI2nS1oJfiWYDgLeKnAWhfhcROl
2Umk/aTfkFpP5ZaMvDyNm/um7vhkQKDnNUu61nDzEILJ+18iWg9IoUpRPu6H9jD1rtHNk8jUt+4U
yJMWrz9/gqIL6V8mcLxooSmi9ITlPLI2b1jsscSxdCV61yLBLFU3LYBmCHbUfuNyChdATl6jZuUV
Qt4jt234za9rmYFjGHYpa98Cq6OBI7V8F2XYwJibIUNCm15UjTo5erL++0iKcSLURWw1oq263rij
QBjHNEVcgDRQ4/itka/5LGTrsPuUwPRjEd7VVgEceh6nTm6s2ISeF19iFTpf1XNlu7+wdHShEhS6
sLw1VwF33A2tDq+D4WlX7tx+k91ulCvAHh80A1TW8adio4qkddzCBoHzExaVhcYrVPufJV50E0Sx
CqcchA8vDOo0iHL0dnfUyyVI+ovSy9fzWX9P/4V+h9EEtVQa5gubF5T3HIt2O6ZWVPQCFw5Gd9ve
j58OcQqNWxns0cuxrQQaIBECXskVH5h7Z2G+kJHAxjSh9WfR09VU8x8WzUcElI7cz23RWbfatGPb
HaAlCy3rPmYuBwAhWQgwc2mS+Sr72ZZirVn+TUzfFDfFiMNfkLBivcqmyadSz05mritHMXlkxfTC
UMITdKebRrBpConihsrgb/MtfQmLqRfp4ZyEv8Z9qqbFLzc0HBwBl+7pA0/xTcIyCk0A8VDSADOr
IKpZ8pogb482q2ULwXGehWOcFxnI7Gp0M6bNqzoopWngp/Bt/0I0jaMzQrFoPW13EU1GZG8CErj8
Ml8aMuK4Pf1tEkkCuU5bnMViyAYzPE1mplFr97x5iC+V1FaQf/aXMpx4J/+sWHBijGRl3jmKti1s
hkn0qhaKdpfkZUpUrBug5i5yHETT8vUuhQ7vr5HybY9jJMBPXiSFVDxPGcc4bBC0T40nFuoYP9RJ
TQtkmNkI+Y68k0GMzfWBtvIfjSbDclFWsVxrIxyQr+P7S2m8exvEjM+8O98nZp/qaZUxUO0CUfgA
8QhPnydgpZnwnB4pje1rksCqXjXhuSjbuLzikaZX5geF2XS00hQ2mDOepX9bUeRc7lHywxm7ANcg
WgjmXnq8X/meeOA7bMvFYEHFPvhhjixLMDyFogjGkz4ZfbeXpFVdbz5fRsVdCgvB7SnQSHHSFao1
SzeoKP4FWlbOUBv4zG4XyJpSGuUovamwUog3PUA70agLXbO1qn3v4EEC7yHILHJHoxuUCI3Zvtn6
TrCuzzcF46XKIEbEJKxXrtKRRecQsxOfgq+CrCOrtYxlJ88xpyjWSkf80NCiWKBXaEqR6EsHIrq6
kFQ2fsr8n0uvXHw5LypizdX60GTt1VbrjhPN+ZotapTLVEjiv7mSULcIp3trQ0sLKCnJgpPUSDyL
8cXA1KWXz1OdmAkKq4QanzHLakvkyra1RZVgcv9+DQuYjI3ytVqwTO2zA3x81EFjth0ibt2TAxm5
6ZIFyGlV8gEtCp5RDI1ic0RNy4wFuxgcotGITDM1bWM2I2+gXGgRfweh0ivTeE/QLh8hLfgmPbik
GsTa59z3Mvav2eckFy7OiDFpDFeBCJm1Z+zuyiWBp2d8j3t51uY8y1B56+PzG1OwY/ELAUa32EYO
mcc6H2brk9A7FZ8hsat/7Iej9svgxQkirq7gStGcq8ic51rgtzP4d2T24rc8/PwHdEU54OnwdGYx
KBw+vzk3LQWwP95Dqy3nW8EsfvuPU3gYShOF+v88TkUpqdn5FOYy+oIvCJ+542g3+tP/B79pKx9c
UO8xUo8V7XTUgJSf4dZi+sENGK3aiaK4GpDiNdgcaxcLGdIkB56GEl0dt0cUzwVW/c5DzIb55aLJ
kJIJq7YgJa6OtvJbnXLDNHLxffiHVDeCj8O/f8lgmN/KTiU/w9wB/8jrYWBxwqOCY9Pq73uhTtQx
34fUz1x8Q1e9+cdkYMr6QwNqmD//vR8m5KREufnB8/fj+k2uwyi7WIrMnZM6rQxmJbJO1gDLbwzz
89Mx2n9G144PsfVt4fC9sIaVTCbdgGcxllKSXbqh9rl0uNdZ3FIwyXkl2LmrCMgtlc8CzUSocEYP
q+xxSYpPZwFvQv36vSfkdm4zigF7/b6vv/YJbwfy+A8rLxSrxCgYNb2ZImvr12Ts3GmTeW/le6ka
QdWrHueezBhcbpDf3FbbcxyzE0nD7+RrjcVWIuY8+i6qOaWpbLr5YB+7YiDyAeCcHSG9cuBtJrWJ
xPXfguTCrAFlF44/cH9+m7wTbhqfYySIVfMcuXLqWJT/X7nvKIqMARYJN53yunqut9ovBxj/fHh3
1qaHGtLhKaFquugCGttPgFZJkhcms4veK734rnUuNg8ubcLsarHvCkCmh8HNYJXSUmHx6e3e5NrS
Lj0SvLM3YhaaoWdhV86oyafN2K84etAih2IdtH6aopjDpwKBRILpGN4PSVye6bND8FP6zoXAoVGx
QuLgFQncNa9vZ3tDM14hilWUYcO5PJHI/pDl/N9Pw0cOJMv/wfuURWdCpUQMlYxoxi3eJy9R+isV
HmJrTqaLj33+DgRe/pwQex3JujlSdlf3MonvE1yFnjkCCsikSWXGBJJxxJbLbk2apOpB5jXA+RWc
I+Tyt6p6S6p9nCVFkDIH6777DHqH+giVqS4cnj/n2mg1H8CJcnjuXbs++xee73oOscSTdBMvT5KW
CxHzrkyn/IgzcmWA1c2hUR7hOHvBaulCtqriVIWRWmzH9Lo0PBrMK49OOMYnLfiU5mGnklshcSVX
doPzxGL6gvIOlbhLxQ7PH/xtKJm/dZdAeDRQ0zAaUaLknblP0MqL9+KvEpbCx1OtuiBjF1zl1iLD
iFQGvXqCNHsonaWYtG+um6cvQWShc7uHNelzP+cVWRTmz5/FcTis61X8SZf4w6fBCAMCfOcqZ82v
RC0ZNwgE8gIL8N62X9Xm51x100qdP1JFsuoPyV7a6f7ljE5JB97Dwr5IlpUPIt1f/taAkufrpw/A
bzm/xafvHTXzyVapeUCO5hu1wS9Lta/egjR36AGIlUVCnacRkjY6u8HhuJkcyIivPHRRtOb6aTsW
os0AXwHX3ui04UE2OrjEBeLysmCodEB1fVNHsVhChVykXPYJrFv3vQOcM7mvjypDyUlBM5ybpT6X
sJJKKyEMrRn6fhi8msUEzU9EV4OKDNle0juunB1+37OZ9EKDaBklSCOcttIVyOlW178Ckb+6Cx1e
EA+U2778Wa5GsGpTYCvyUMrkCQc1EZzCGvgDex05I1dMGCFior5RkAm/rMhDOhF1hhrq5DMGAC27
LaU71hXgtgJqKl8fCnj1QF4fB4lgsKUNlDzsBPd2tas5O74ghSs/6Vq6W+w+YYiNf3q+rUZ1qvQ1
tuBOS5w5VfwCdZQPpyn269Sp3H69jQYxn464FAnQ32lMug9T7dm2h9w0SECsQdGoIHdXFhq/KtPU
8F74ymnUF11ehdKR8AC4qaIGZv1hul8A3Gy6NpsBZvBzNUpAi9ovbrwb9dydnVx1dDIlS8+0vAGW
FiKovPTa6GtKesN8xN4pSDAZRH1I2vZ+8wUp9k5cXmEcJfCBRA0VXicWzc3SVBLDfigF/XH8yH3M
x8O+sDWnpanoqXTylq0/q4vKr/B9bULrq+5qHujaI60uJY33nNvO/loJ0234EvH6I7RkheY9iOWH
rhqczEJYn29GQw+2N0rJz2dtMY924xcSNffbltT5QfTc8lhYT/sulWXht+y7GkaOrAJyfGWYBbZE
ArWMBr79NC7RiV/5fzPbBPmF8iZSIkxWFXySQqnV5bpHYxb3PVnh/x4o08iCuI7M0lg3OmVWtaWo
LhOyRip5GUa195bAgcViKz1nYoW7oj7buqDvrr00xlaOXD3ScrZev9ZGSK9SF2+cBfa9SXCX7ffV
k108gBNl+6tLFzuJBhun7ft7Z0yzgHLIEAwb/0tqilrZiE9JRMX5d5epCuOe56AjJfI9vwC8oveh
+LxgHMqPYucKlUU+U9EFyWDH6/nh1EIPkxf0SaPReNSOKD9cfJ4DrceqDwkyaMuy8R74nNzMoDzR
v/lVwIQQqrzwIa8tOSZN2pMnhBj0DUhjGlCGG/yzVQbEokB9tArJJLVeAn9UZ/IXspiEbQ4TwfR9
zvDxlbXa4W0T2UzTPyx4z2bL2QBueorPeODEqkpH4vN9yCbgK2IvsAaMmfTtKTcy2SKtCtblqIIM
VlaFztjK2RI7vi4IENa7R/jnq61/RuPr1kWg0/yXAHdvzHj1ANI1WKLcFU4CUyoAIi5GgSF/oaKS
IEpDmhxUpTePbRA5k7q+GGqUqJDs4EZBq0aFg0yFqD/lwWs3NK+uBJesB161aFFWqZQfLyalcHW+
1cbUNmtHqEJgEVKnXXL1k4HtjOl4RMKLyKveJLQwLw+ZbzqXMSTZsDIubv7dMT0sXg86sdcUOgiD
BskU06kaL5BRLsDYLVzbnlv/ZWWUqF8ka26FSYLDzNvWroScnvKuGuLfWFhFdNY4cxUHdQ2UaAh2
Ih7vhEPoTkX9h4xxC90Ne78RyFQlxtvJQ274fHc01LPrM6JqtUcf21G+r25PA5iiDsinoORsCzhA
E5gJ4V/T2giigRSURCA+1KJfW1bEMVLZEjFtp4HT+iqioAUj5fkvGl+3MrsLJ4IpblBmcOLjL/fd
/bwaQ4jOj4YrKnTVDJh8ndKcVqqiW9uQqdYmXOdG0zd8lWxMEQfuJchHdiMTjPVscRlixncbeggq
HvnCwDjOHrWn6AYlcbWgke/nS5vRsKfNhPvQJBTdIR8byEniI0aZlF4MXbcrQtoVWuO7T30tBotV
eDlQBZRwVC1qteLpMNLOXZ93E2Jo4E1UTt4wceem1P8imhNZLmDFSfttM9ILH+ZrdJcvtEJgH7kl
dqz4n/sO/NQGHaTCYL7MF9A6O87BfFSXgdCl3auWhox3cAqC203CZke9erGZ8kvxz77VXcMtHfko
PYVWFjUX3RFH7ZOd6AM6maPR1nIoMNDRE1I94QO5L/bi3khfA7CyVoHHpTYUO+EJwI0hRJdicNwI
wBlYNtHNBpuBZZ4N7VSckjBy/Ya3yZCDPdlApikWLf4yVWiyQMUNnOx1uNHHAatGXmn1RWf4Beb6
WVJAnCnkeJKg5TDAl7CzSu7ZoY8n7AAbEaq9o2rTJAiR9hrd8QIXL4DTPCw/Mf80Pmn4RfaiMBXq
ob46F02WKGw/ULAEYgDUnhxYdptsuHEOomwc4lO7hqr3Jeo7vqx4TiALJIYyrt0KnQb4se/cT+/M
idKPazzZheYhH6xZAuMlvcE/+UQ1aleqv52HzelwsMpjoFSR1yDb79WnQJDdECUdWP+VHdsWux0p
xU+X47o892bNg2Qh2LdcEJ+blrTwCuBuDM1Qft2U/w4dBxHzLRXDXs9hV8G5DA7WM1MprnLkQ5Sq
aOm2wSoSyqM7Ao6Kqa/wAwK234v1WAx5vR+iZ3MjBZIVoO4qp7Ooj2M3ChZGKe/Ie8zhWJJJ0q7G
uCkx7glbBMfYZy7unOUS8wRg27fgiPnabIEMNopunRPEYZs6BcQD8K7PMIJZJ3sQqEIJMRVGmM6Q
5BusVvI4MHpYqrxgAFqRHBBsMbrprxeNJuHT10qgDwAhHq3DYPFTyfwTKZN93jzEzkwoJEEhZWpn
4jsfe0wqbTKBrkOJRwIiwvhBW+Ot1v4WmqZO5s2A83kiEVVY50a4AeTs7A4Pad6vfpWVSP9haDaO
gDQjXFCY+Pn8OYEnUC1lDw6mabozXnld4PMYsfNlfvC9DaaWDQFoTSfi36FTgFJOqf1caVuBnnvG
RW55OO4KlOqVP3z9+mhzIukrTfG7Rx6/tQqTqRY/9h5ZiTe9U8DkvRLd/O504AjGl8Cbfu1H7ipo
ZhqmpU5ufAK2MG6exseE9tuUiBewzoLLGf3zoDgiBbydRXNTI0MsDqkjXybSffG6UQnGKaqr/sji
hLBrRH5zH71ygznNMyc0bPIeFgmaVggVLGNA7KnGVOqR9EdFeEQjwPIym1u0EXkTouXrPizbi/h8
jt4jezYpqBlT6R1lWtH4JRptcB75/BE9qcAgrhAL4BDp+r6pqElC+WsEtxOJtA9ZZp5Fs7L3vlSe
e8xdDX4IBVOL8EDprAA/2Xwf7wvLK394xU4p1wxuIbHKbG9JRChXzY0SL/Nu7KQbYOWKWyJhG3dE
Tt0WSapTHCFXg6F7/6gimozelIqpc5iWH2YfJiua47J+S9AaUqoafdFD8TYwPgbaR4Ljh8odcnw2
FFjKsSGB75Y7t4n76yByTK13vbk4wuOIr4c/Ig7Qd1c0aKamW+0a5vMs9rT3tZzJkfkpMfG9wPvl
KYKngmobGNg9k+wOBnQdT6EcyCg/bqAkHLBpNbdKS+Etocm96ofUPhCXRhSGiq8hNtQlSBUG/glo
baJh64meeUC4/eiwIz91sIQ8Z+YjpeF8mzWoM8pKG6VlQ0oGRFaGY6K1yZe8yhEPPIJTUq2DtJbP
BA0xWu0MXZDOe9tbjL4o8W7rqzsz4WdcE9+cVRSO0ZLmXt61ujq8y3iuW613dOY+D+90+E1DUz25
CUtZ3YHBUfRWgkDx3psawsl1xPhQucpF90Iu6AnjGw7EGlfxRkTuG1SjxRmmDQTri132lL6A7cDm
mfq0MYbB0EMZGSsIUvBRy+F7JKgtjA3UPkLy9oJf2r2dQN+Nq/ZjgX99yatZu4favwP8JpACYqjO
j1GHb94+eDdfN2ihHN+N+YJ+seTbYx6xXt5QbB4SGA9lW2BOAE9SMCnp1qZSl+A2+gGIJKgeqlQw
7BG7UC9/gx4IiIctNx3DAnJC6+UW9jP3wxYOFVVcgUgDTfnIwpdHakUrIxGvqwd1mKMEg8qZ1LS7
E3xojAa6u9YpMRrF9ZGDwTO+F9q7EmxBHr2R0jOITxJZl7ANGRj9gs22EKiiPjwvssIONITl6l6f
C7aI0o4cBAES/hJdL2vvYPlxBkRgA+4Z9r80ELEs5u4gNFYxB/a4Yo9Ngpo85OhSXBGDxda10BNA
3yygSfgZ038JFJtJkyqBhWbZ/H4+BYBDznl0Xm5SYagROPzTNYO3mw/wKD4mgZIhF0LZLezYXInx
HY5TliDevuXMdQi3BQVZkOis89YRiLYYdDbWMJ6U6AAm+KUSEHeKapA01xI5r4wMIhxjm14xRn42
2ZvriFdRbuDrZNZU7QjLOAOQeAI+6wVLZdkjlFfs96uOPP+mTA7kBfKXpoGdN4UapKmnYj8O9u1l
o5FeuMeRjhJ3RgsCeYtcRgovfuS4T2BrwfI4MXqDxjnEu7hIZHuqeYVhaRZEEtGVUeU4cNor+sei
af4ipL+h+4JqxvBQtNVkA64P+FVQvdVZVrvj/DGdL9EGzc2P27ukE7zQdf0/d3fWk9JPi8I/FoZ/
dc3qbnM0Prg0TYYAff9oqMW2DafSugdCIUQNR3yyfPKlFehKmvk5+IZqObKkqgsC+mhtw/Luh39Q
tA6Q/hgU4YPMXgxE/RX7bHBzIt3dF2y6O4qFPVieDC9vw/bqDV+57P2GfwX2lkCjKyxByiuG2pLA
RUhxYUKyKtfIj+nuBunYOqLCUzzB/LXaSiOUNJbOjDXleo7e7l0n4GpXr4p4gN7V708L6LRRY0KH
0c1D1oJca7RCtEMilefdmTJvMbxkGcN51O7TBLibYnqlfdnWEOxMxkBPcAyBJoEKD92mnoyUYxYS
/Qg8h5rD4baP+P3Hbv1MIH6n7x0qn9q3CWSXRgAxFu49xaW1jYznoLbWYw+AHPVJvQI7uXMJGBSu
JOtSfYIi2b5g9uJBzw2BQe7+quBrzPnjul+Kzrka9Ep9Z3HNfTKjjW+5Bof+xlikQ+btW25+uVB9
8hh7SXHzrEKk4D+ps+jIX43oH5cX3UnhV69jjlacbRpLcDl5WHVt/Jj3bGmCZtVtntxTIlY0265G
4dny91m6fWWcHV1RJxBWEjxVfi2XlbSzIp4Wlu+mtKvJB5NQd4DdjsZ9PCLHqfmS1Z4/xLyVJibE
9a764qgENs8t2CzU4ZziHK3QTVoy5QFkRxZipNB7iqHg4kWeOzQ2gSaH2bHE3ulIw0b2a3J4K48+
QRL8uWtpwusz/pQ4Iu2FN1ne50YdUyOo3B8ucjtAXxiQVwwtolBB6JK3TJM69PlB8AxAj+tCjN2b
n74OR0yMq2UsllxLsb4JC3nZ+oxKgRQ/RwEXfgeyTbMxRUrj0tt4SPezkeD7oTOJ6Vyb9IpAW2sU
fqQAlZwSPDCyI4Q3PmhaUYORWoa9kLlG3/ZZfqjqwtxa9Ra/QeZKtAlYlshIpqI2jEfVVnmMoRIV
Pm10Owa7zL6fgjt9MbIh5QPfUbEhpv+es1s37tFn+ZN9jqnTJFNSP5HNCEA8f7ojS+fE7jSyS/We
viyH+hhqx3I1Znet04r+N5XqEOtzLMVPourMBlmdsKFCYJ23TSfhA7c77cJQS6jfqtjbQVGpsqjz
aNl39d9HfkUSoHszOAz1bmdSg1vfjapikmRWmF4C2/BeISi0mVh+uoi6vxvS2KcaDSdAYUJOq2Za
qwCT+mDrLhIl8BYB2wuRiHAY76wi93z2zrxsnzNBdS7+XOQPolOZWThrT9YnkIp/KmljphFACuF4
7343dJ2WwRzNTYjLirZofwm325xRw3eV5ed8IqnFR6L5LTQewRQxXWxOcROwMtHW/NDg+cNDKP43
8/pho2DZwBsFLOyxqTbP56jMVBTUs92uXQ8fzH3D2SKnW5PBFz8jHxmtgTOIppxXucdkdAIPqsgG
itS0+YuH3HPBXBo6RwU3EQZcebWDrkTIAbp1BRiKnxJtUdWu5lwrdN0Yyx20GmIzDmgXWyXJdVmA
Dh/W04BlhzeS0ITcTCMjFbshND60xlEKJK2TRqHWtbvqQkyFGccbstHxTsON2t1KOVgI68T5kumH
8673QxmAE7zMOpU51qOP1yiMG6UCJuWrhktMn7l4GZiLOPqsfLTiHEqFr5JCZPk7f18DDQsXJ8Hu
/VGp77lDhDT1GTAt2iEvmLzBbPRPHyUEHK856gHzwD4gLyZB2KP3WtdhUAYrgdeqwn9EtaIR8qhy
473vN/gUvk5S+N8bYHLFV8/Vrp9fnt1NOYBN336eL1Jqtc/xlQisUa9c6cKnh6Ays4huR1Wr/8od
vj+R9vhmijc5uSxFA+J5lX5tTwi7q4DESAFyCGfzX412HgyguFh6j4UVHFMWvnjiDiwprWiaTJiK
NK8u5XnnETS8JAdLeRDTqnKA4xv8+WDnGz0XMUTdfnYQxBYUg85JfxGBsexZ6g62vQNaJeVvulpR
Uf/B7U40kQSfk5Ryx5tbTuKBG2A6jJR9NZC4NxFyhI8hLIpA70xP3AtVgjNmdsSUNjj5fdp8bjkY
s/0jsVm29UgRgstW6mWrAKijiIyMd0PZFqxiRg4/gtYrWTUtllCnHH+stjBpwHvdceLr43+M14/r
+lWynUjNjVy6l9JnCb1aag4j5FElSXtaeopLO89mxtPfm+hj23A14tPO29NhHdRRbAIksF/o/mki
LJV+j/Vj8uGW+UjN3TkdUV4TN1aw7ogM/lBuzCTu0amtWB2LSBSq3312wUbnxhnHJ+pLqDlagVSd
NyQTZFOPuRootIONP6YiCg1oXo8+oKjD87WHiEQpEWFc/w+S3NSflLQORekuRYtSuqFKEvEfqAY5
cmzDdWc301w8pZX+xpFC57fS9hi1F/v0yxNn4SWaTPmRfBnus3o9QGlNnt3DEz2lfqpm6OXAjm0A
M5J7nk3ouKsz3DhRo6YBcJzDu/P1y4BSeUJAoO3MF9aRoT29Jg2Kzb1ASSg//etwv5DsrSuqzuqm
qiUvVRRPYA0EsPkBukMEv1asgsfprmeLzJcBwp/rPbnbzkvdRuNv9HCtyXaTKvzlCOaDJxJMwu6+
Fui9BituKko0xWPLdDsWZMBpmHHKZDXKjarXF9s1b37qeaFvGUGGAkQaaW1aZjfKy9eB2Wv0uB9x
ekxJAjyXeGFh1me15LSRFCJ8YPEL916Qkbj9Xgox7NYlt0pGu9AgTV4ssMgeJ88lSYPa5hKykRJD
NSxclLKFl4D041tzMossHvtqfdu1F6s4PH36pNYaWwgbJOaWOYJhgr2k6fJkjZRQ0csOz9L2IhtT
eeIMZJHxXjuf6qKt7g+EB37CbHSejHcwh4lURxTV0SNv1CWPLPf3jVwKP01YvBWx8BfHfo83+Obf
SUnzflGJ8UL9kFA5oKb9efK4wVDoicrhgIhHSesFSbh/1fNhmqhWXkTdgh7DuJtKre/vW0s3ZCUM
8ng1mXD5ikcjpwgx8OvA9Oqz/V31/dSxJQ0hyDhudfJ3PxLlvQKl3olEPNSLBNlsBVXEY8H6pKFG
V8k+arH94rTanA0eyNl/h7bfrURm2Sxe7j8borFJMt6Mxw5hzIHCzl+NWEoYkXwbV6MyuYifzYQZ
bxu2RSctXaz0CsgMkul4Zya2tpCr8qfq64ydciPOMJ/zPwhxsdzQYBBebul15OmZmTuF0LiLUiCv
dlosfENX6nKeR0LU+eVCuLEfmzYwgSfzZ4kHLuZdNraZicH2el9cpNSLJjXhx/D3Qr9z29MH1kh/
pA4Vsw0huhMMvvZV+kKWWSAgpCbY0/oNvxGDlNOIZsx8QmgywwApYX5qlTAwR8MisEJ3dLpfHApc
vnU8DPHZTD/4um3A0clIjuh5ktagAdUUAapQCW8YWTPvxGCv1PWkILKmbK4ZN+6tDxlkYtTQyI52
f7D2RT6QSupDBuZ+lkH0y+iy4mTEfTgeqirUMEUjALxgCdMm8SL5/W6NWvXH60EXmL/R0kQBJVKB
l8iF2q3Jhvbk/+gSZwMlpdZ76h+MJVoyW9u3JB4jJUFsUJKnMnyqVzzkL/e3v/TdMQ7mndP00Sbc
xcy9BA4I9iNyfcHiXzWsfeoNecTy4BbOHAblbX1ilinM0Z4Pb9GaN8VykPnOIFUrqFMcexWVhzXL
eMuhygZdgQ4h46jzfpbx4Ug5XY2+SrkzEvDSW/VjgFXHrX2sAmonegUy/AWyw1f5x4kamXClTMvy
eL0Yvj7Wy3OABZ1nK/3brnlwGgQVQ0WX8pZw1yuZszAFCokBnHDnXTD7A4qrsxHMuUmXV5ftGPLh
iL2LkW1zAJdeaf0GeFxZP/hkXVMyEdJCtupA7TgpnERfni+L8Nlcd8kTU/ZLvpNIFUck/lyf6WdS
KhNPocwKF4pkN+EcYiBG9UbBTfGkQ1g+GGZyILsfBqDTro63clH4k11dJE20IxD61IYKc/lW+2tx
0ArlfZwFtz/o3R8mkQvj8JYMHeFvAbiOf9V5uHnrigKxerx7vGckI9c3lcvr3NtNvBSjQbV1iHXE
+yRd2LiqFPhvnf+KRrNEXQqHJvJ+e67mW/LlO2YO9ByDvs0m1D6AbyF49Ew1UuNvsVcA9K5nUK5B
nNxlod+R0L1+c4su6OvpS195Q/S41hjTJtNx1P+Fw6PbhEcvGem2+JU2o5XLPu2N+e5cclKVwFuT
WwIQw4NbBphQ867lcqrgOkZHd94nq4tKMP1SdzgTWR0OcvZWqv3U9ZAHHV5UANnY99+ny2TkF3yY
zAH4nL8N+FS+DOPYCSNWeZ8ALZjG9nNowBjax3CayGkB1T0yi+EP+AKQ+n4B6ckCu+icSqWcwqA2
xWMwKChzzz6Qi3pAesNZpfuKjGyGVJKhGsHsgrPgvrkHBoytvA+C3K13qdHJxwT0VzLwP6OdFixj
ewuKH4MrG8mB3URi7vDOfn6Rm3ZRkuAms0MKpwscfKFHZusEgBxJtI59jTCCsBl/sazIpMJV+PJF
AsOibrFBZOgCg8oFtowhy8whdJW0ATsa8O+GXo6xKt8s56gUgOaXYDj1piOhuX4RAJDnoSGU0+mc
i+95meRDdqc8NA9CGrwPvkaZtRC2vKUYwjYg0eAInJBV4yfpLb+Sb2WZ5i17P2Dcof97zF7yIJu1
XMEFbR8wTpl1HZNtxK2HHipV28heC9EIEO6s3DnlaG8sfTvWHJeUeH8RqBrrskVcn1oC9FNrOrkt
DORUKlOHZ88/F3op1uTqE3py2wnwbK3yuMBVDRlhCm0q3mzpvx0HOMqGOHvGUD0Lowj0qJRXZp8f
Ks76KrVdrITCQZaMz7K9RjsDT74CckMN/gji9seU2siMB09pC4k6nSsfUc95c3vp2WMZXiEofD2Q
dVaXlffhwXtiqj/tloqCIe+k6BNDeo9bCd/gZRETrdFgUSo8/1oL0yKeKXIX3igKBFEs4/x2yhSu
u+fKFpIDCqprRVaEiuxrPDEr3yjN3fEY33YJdlWRdYJWglQBXmOp6UpsC5e5cXQdNCSvpLipfoae
QcPpazmYeSGvpDgRQiu1nEp9V7la6t+xYoZ/emroUIr0zBEdKEejNQy+wi/fJy2DQmSKM1AJoWVY
omWVtMSY0U+xCZtzYL+4jB96PRhb85lfmEBS3mMLCg9v2+gISEsWa5S2XUnhA41S10bMmUkk1S8g
PGfTNw1+gEHOvnamLOs6orQrY8k4Zpy1Q6NkIlEBxseHChK4G2ht4SmyG4bM/imo0lXm8kOB11ef
eqn5KX5YpznqGq5uwJOUxx0rDb4sXVujH08vp4TUljW/96hctcPqyKjZIyKyunMhW71CFw8RpHs+
J712CL1WRfdNuSoDFn+NCPAtyuGgSaQm16J/nK0xoTZmZKTVPF4So4bmha1WTqbHa0Ob3Cn7gyxf
1itW1c3vrKekVPYSQxExAywGEmd9HpcXq/NDvZ9Zkf3ujNZClRerqyfgV5mLb0pBqyZ1CXv7qEm5
2eyfERXRzEBKWpFMdeTAvtgq+/wVIPstLjDpmdNQun8Ejdq6yJWXkNWu9TV1MeroycZxSzRXgwQq
CWJ3K4ZN7koTaKVU08hBXlW2MVkg9ekTR9/n95oD10huUrxhzihGEx7q51GYtk6HBUsrmzqKmMIw
Oy3Ep8KJF6EQ5k/UnDN0kgRWJXYXSd00dLPOyDQ9z0ytugGNy24eDJas1C68DzAaonYx3Oeed5BX
ocfQ4i6Z4VXuWGdjYdTnwSzMQT4Ja6qj8zPpZUhSVC+CENItDFJOXqVhGHb5ffXIFF+AfcTB5ug4
W50C5StPx4/C6de2hNvrc1tdQZb6oKYawKhqjOzkogjD/A7C9yZaeIAhm3PzhStiP21cg/qe79W7
ZNSPUUjnNlVRW7zkBscLw5Lmtsed64bzjvyDEq0KvasWer37/7tZYf6OSZko4rzHZDOCptC0R40v
mMBLXygNDFHN/dot1SLorD0pN/TcqNqwNXH2YLT7DL/Q8hfD3xHifhSHG0Tji+VEXDLHS6GKiaMQ
aXOkwr7HyLEfR6a7hLCheW/9kkKW1OhXF6NUTSIf3XljqcGwabwIW5osqBu0kIAdSeQOCDjBOCpB
5dANjC9F79JOztoQXgce0fZ+XLdxpWgG7GokFNJuP20tB9pH1d9F69pZ6yQNMbl+nAO34LiEq6Zv
m4OLLrlVpsJntgHukzOiauomtY+jANu0MRkhXYMCaNVpaJb4c2d0Wt7rd6930NyEW7K0/KvxAcpr
rIaRbFAcBKtpC8pmZNAEVar1Ed6qJFuW34WxXEbDSH8+UfrqQJZVcNzkfIDwsGQhPpy7ZU9aOqic
wIR6Rbr5fmV1WMnBrMwXUy0jLqu+21HxghlAAbVPJekBjMbHLSb0hy+evZkDfTY2XAgCQ+4Q4kG7
dFWIxYbsDYYDACRw44uY+ElldbtseaT4MqQMIrGeZi7BZf0AnGqX5ukUoKrvIjoMyxljf79CcOS0
Tmmfx5sR3wbTlQvrpVZqxjq5s7Qxo1cBslAj75adZJVEHt/Nj14Qlq038wdcohbfyDOx3Y+U2xJW
dWuxy2rqMainJE1LF+ImMlbnFQiVuPNX8fX3a79cY4vA8OX2xyyx+x9pCMePQx5HB3Vn8OLabO7v
hotYO1uEh23pbhdV7xjAkBUM8wKggJ1g1ymrS+BHNgQWrBoz3go9gIuWBQna0IGsbD4kTiuMIWD0
YVUEi6GF743fDcsyBahOXB8KRpFCpxD/RHhVGC8RMy+chUyyAwyn9VcJJbvaR+c2frDlB5BERxnI
P0exHUMc7qLBzhPeX8qFOTDS/RYh3llPwnrSGJlu9EJbb1AeUjDi/VTW+Y/AGssbvcQW3C4YMYM8
kq1WL+Dt1FYnZ1Qu0ng0kvJ8DWzcq3KZJxCKKV5wZGBMzd5mIyjGmffWIrpDL0/Ep1m+54NzUPDY
/mJc906HU6imn26g28Aw1UZEcIKkl5zhw5AlTDGCsznd80hPs/i9IluxMGHTifRJmEwFULVVMtds
TTBOUMmqKIdxTUJp8uA22kEzvAjH8Foi2vHr1pPgFhzplH/WTuiaiJSB2UgvXeYfxt3DN8HZESz3
TyZqIb8LwjSEBVfrVbwbgThJrN3ycEkoVyytDS90DQmYXIjTACgrrPNQ56nkslZWmAk30k+BCi6N
qB1l3hRhGdy28996yw/u5QF6Q7Jmqg3LFM2JHQq/yfFAB4lTT5YHXwf7qiJwaEkaHGIY9FHFJ9RH
/qwJEhAlJijXQjVjQ4jzc5qva8oTkjBFoMjuTm2ARhXb9IlnMoDFGcgfMN1a1NnauzTfTri4aFBE
Z5kkKhgKY2Nbn1SwWrjPQ7JoFQttlstFqhqy3xF8Lumk1QSGGYIA15ph1LX7wCS5SHy2o6zxdDZa
6NOBvIncJomeC6JsFMPnT2S4G/GHBoiv35kMUhTWLQfWD4YVpFocDMMxBTIjkMy7ljlicGMXerMt
/kR6dCOFEmrMek4f/1M/IhfmbkbzRizHV1ZpzYQLMQDUKwbguESFOSMrUhlRMbLd/GqGd7oJkwSw
8eRfd8DRCO2AzCaZrHst++92aAoWo0W9yHQ7FW1N9vb1s03oDAN0/29uIbcCNegYdn9JgMyrjFRw
dQU+ZSCOgi85jiryL3DOHfRiTVds8B9XSYbuIjtXxajtEibzhFSJkGIMGPc0JWfDE665KorT4an5
UM1OeTt0n0CmHEl6jWlA37HkQldCk8rthZsmMd+8IYodyeQ2SqOmx1W8NbExtmWTx/AsFQHIwv2a
8PD/UfPng7Xs3EEWAKCo+GxhTWvo5q8N1PIZHtXqpm6df8LGPRAQmaHkmATc/rjPYfNqNqk2t6VN
tUH0WmJ7iuGgUVRIf6ylLU6E+fnprX/VdxSGX1C7H9u7AYuR9106XIWVsxC24KZdir6OU/e506YU
+altfNbojDV9uHcWnhy+Z5b21UPQ0V1QO8k0F9EXA2SWd9ZxGV+0kDbVz3K6uCY/8RV+MLX2Fzpx
Z+lEkrigJNO7CUO2EksSuEcLEyM/klksjl2y4Y1OLV/8nucFdXDePzwGFqeagYzdqZ8uQU/iAQTY
csgUrvFUQCzQ6FS8amEGrUac1NpWlv4be+MURGbr7gh88AA4hErb37Xml77gto8iwygnbSD9nLeP
1Ti+EnrWO80KeKgF2iBFIxIgbeptGBmawHzhfJZP0bF8tOVghNsxmqmogNl3p3qQjBI7PKOYkaUc
8r0jn+T4LLwpcfTTjGGWpyJX5SKNT6ndt2x7MGz6TOJOG4o9CMulQp3BqoaiJpGMHGWWFkraO9yH
E80x/pre2R+ItLVyHR/ae9ip1giLpMiLPd90z8xlkM6UHIVxvq7wlmo920l9JlXTv5ZmrEyC/9Pm
Rh9pQ76bKoG2yL/8tWsgz3Qc/D1SLTP3m9PsMr4jJPHrxnWHkSOjCBhWdf1ezsJUl6weJHyyoEuY
aPrUJBrJUM4W6srVLYqpgZLMx1SrsruZfVoOIJKpMu7S2iSMSQG1Tu+8vRMYc0lWFPMelNkZzUkG
4RmEISPYktl/wlqS/9gKp54szpFJJZf701S5/Zc6Z3MQCjzd6yidFgMgLtVcxG4p39I7l1QrMuNp
r5iPYk/ERIPcyQUwBfjNiUANMDq/RGF03sNWPODUhImVp+YGbHQW/nPYvCqMDvwusiz8gFraoBsF
s4hTc3WymZMA4maX/kBn68jWPEtiYPa0uA4cbDTxvkRbj8cddFuZY549kKmZAUorZPAMP3hp6ddo
InKOoUyCp8S0YuBaTZQwStzUkOvlCKKnXvKAcFKH78yCu1f5h2Ler3j8kp/od2dDReEP5nTemxOx
SJP2lhlbt4qL7J4oJl6INyM2mokbziDeRJ8thdo6mltyJu7bl0n0p4GqprrXGuymR4tQh8axjvFX
YaqBBsB9+A+p9a0DFnSYoeqSr4WYoisuLcf5Cg52ditlgOXq2fE5SjU5Zri4KdDsoNvIwTmfUnXs
wZ68RzpU/dyACsOZtRDCYgRwOsqaDvM92cQ5k/9cP2njIuwefFTHgCVc9PNwGLo0mXHfjlh6FMgd
0rAyaN62y2IRznYshUUXLHMa08ttFyKUYeeirPI68+vRYTtrytkw0FaTh0acftGwCtdhugOuo7BY
w2OA5GxSzMChd5euTmIqYfeo4i0mCv+QGC2ymY5zz5Lh+3zhZdJNgx0jhjsaK1XcKzzmG75e8SlG
Y6qjQWzUbzA3mb3En6seAQBdJUEUmYe1sH6li9Jwnh4CsnlwRwzOI1N1sF9sUrGYqXp/3YWQ+okW
mKzIUYmpbtbRjpXFKOUQgCyopdP4+esjj0TN6Z6rv0iQKjEEF7K7eLBLL5tQXRRcjpEgeES9zvwR
49SmxfihD42wBvQs1KJHolz8bb3J/goG1YeGybLZQTkH+2NloXW4yGL7IDyPWm1XaV9h7DtlMQFx
4VFbQJHDCsDh+aRSdbXOkvsCcyRgHQA+fQeRV6S9JZFMDQmv1pnM6rT6/BEe+ycvvtSSNFoYAIF4
vNcKRB5CrltWhtNcpMTLZL62TM6P4nMMTYsgns4sbeSpwqRKI6vGrmhdujHM6SJo83iGY78zXb77
C0uMg21eupOjw2bU6N9YXVW9l72TJZYVyWfTZPwMEVs7WnSBa9jLR6jzZj9riduaNCmzucPNBcaL
lZuSbYNHJ1MofXFkEWDjkShUXRnbTtT9qY3lg1+MSyAJIhmwNDoJ28o4szboq16nrlDO8kpii1W/
1kh7uyS4eToRRHrZEmAHFbko7P1DKeFtqubVPVKsbaPyucaI9iEYm7WZ3XFbjr5a5RYIuCqDOgqg
15yMQ6v0z+ExsvUlyfdr2x0KyuthG2rVvpMsPvYuHvuzkyqTwOa6SF32V64VzDQGm6jbT495Ovo3
Sfe4Mv0WOnAP3+fvRij1EYq+SWqsEHTVzQeSi1iaYDKUobddURYDaabNu2Z1BrO/urlcBnmK/d9D
SXgx0SPv08/icrWgPOnfEeu3huxSBBoFwu1K1QidZinvZ7D8Yc8cLrY7mTcL38z0b6+fn/eva7yd
vR6aUnNi5tWqAbGxHZLPMOA5nzY876CId+G9vpZqfK8Su0kvppYCXr6SfCf5O2/84blmkYMxcIPi
gPEj7Yw8N6oNQjnX0ZihcmEn6qD1AbUlZedSFildrX3OPZwz3vltSkueYItu7Ziz6z1qYF/FPCly
fxv8BOi4DdwSBipAvXnG+ya+c/zQt3KEz8RWd6oU/2t/JNAIWntMU5Jn2f4jnx5FLuii0VgHblhd
D+8dIAbzuKJX7xfVNK0OkZrJ0B7v1SU0ga8OCl6OOcRT+fEvZBD3nOFl5d3piHTCIWhu7ijTRa4K
Mw1pymPJH68Ys9wLDD5+BegQVDnq3Kl77mjG3dGJ4kUwSVUastqQmgqfthY4gWq9/4pDXmdnDbWx
M9NEqCwSEAFLTItLdCBhAl1jR5c1XwhZfLAWuIkxwLnokKhREaaSjv3ZJ8WsAUdX+MWa3vJuaMaR
tt7HrQOuLKiUQt4Gel6cV1GbSggdKJor4kWvi3I2qsItNI5sGK/5ZhmK3AtCWU0wK1pAntEr7fTm
LQ3vk5RypN7AcKiGVC1qdb7GzivtzvafGJgofYTct1gvLJJlz2SHwrQtlua7gnKs8PuCBVOZ9OX/
+UbY3OaU4SSftbEfNxiofoE21zqhciRoYzM64WvB23PW92BnVnD32hlWR9s25Z41U9Kftd68ZPaV
tj2APuB0LPnzl3BmfBre5VFXgFpHpp4QVK8ZZ8EkrGgAvhlQv8DEYYWRwZvadnSf/sbTWGUAyoIV
IHGLCriFNiIr2KZNrN23vBwoPYHGnb8BzFjzzPw4L/sWvigR0Q202pMZWw7RFGqQ2WsAiRVyDJZm
uUX5ZmbF13qOkhfGNLycSamQLiDv9zf12ZjOMhGejmWRdcGQy6gWzt5o3vzRCC3doT3cmTOSUuql
mz6YUz1nTyxmvGhNU5F9ol6aChm7HrU4YF4y5hGfexHvPpVtj9Gw1w3bmLFPlkthgPv5we7ME4YU
eNjCrM5ooilw2ulgPpSqAIXbFsHHk5eGcwKQ5V7bxsfGElxx230XAgIjlYJqS5zRqSKKREECuQgw
RFRGcCvbQ5fnbLbBcz/4mdcQXCOVO4CR5nwxpmYj7B1YVTqJvbcCVm6nqpIZM5iMglfzU+JzuAgf
xnQVM9/qHAdXDmpJlXH0NCW0AkkQQDO+TBxmzXza0JrVaSpmOEqW7l2gNSt+sR0taH9nEUc045p5
bE5Uh1ZGPm3ocRL0bq4BdDLX1v01f3REzE3wt++CzEX0GTfWPlX5UMjozO9Ba/n5QEzwgo6uRFNf
mT9I2grXywVcSWI5Ak2LxX5F94c1Uz4S0cI+Y4Kd+H+loBCMYcaO/t9JVmxcwfx8ruBZgzqUZ3va
tL+EeLsS7PgYjQQ/T9uV+P+65qxxPXXJoU3ypnOfUkZ5Kz0wkbSgm0ri3TiOaET+88D8u/R8JzAY
rH71YMFxWPXWSGjnRIjJ9bvi69iwRW5HkuRvvkg20FNdYDOrf8xSMVBLVjKXM1kH7me3fqtFhZIT
HeB0LotilIqus3HoM6FpCNWoMVQy2udK5W8iFIEjLzCmstJGav6/ktpgNeLju11GoQKF4LmNd7mq
Q/8kZK46sd7ecODKOkoUZLd7ZUDZowrEKYGeCzFc2Dhf3O8XnIsp92qBpGFgMD8BXvGnd3o3nYlM
YBV73Z+8ITje4Tz39pa8tyhwLXS18SdTTAqDytpyxXeBChtBNcfBpBwUQBbuHGtRQ5p+267lsvA2
tRlXFCP+vjmc2AplPKm+9ru6KjrS8c9Dc+yB0KlvHSrUeGx6DpF67ANvyvPGQfQJgac5I5JF3TNA
nEakPbqaLAZRo2+t7JgfCMIvrT3VG7ofnUbLE0TTRfrKO7CM6tQtHKqU1aPlb+BYawmgHdW0Smy3
Jnns9dk1j9Wt/6Nnx4RcVFephvKL7IXCfFnb8TJ0N91i2XrTomkbava3csxC+Xn8p3SEhWAK6kxf
gr2uD7u/s8tEzzwwOASl6I+VQalzpstCSvf23hj/x+XVH345qeiY0k+WHEdAPevRIqYRLg5a2wzM
2AgTbB9BSxkMK/nj+q8sVpzyqJtB6lPp2yFnQVdqCDpQ1jhMciJsHxytsKcM4q0qVBlNnkkJwjYS
qB05P9vW8v142BXCqs+HyJQUaUIpq/UmD/tl2B/JCjU5W2vMsa97YccmEGcqrUBgvptwKhBh1CoK
of9PQ3S5sKX+JO511C66T29c3qjCcaL3tehYokg2tFZkCs6kbBED4zekaePge1VrXrA9dQ05b1FE
67WV/dVDkHP+ML/vb+421viF44tMLng4QGBpWnl5iHqppH9OAP0nDInesAfYyMSrLYM37dwGZD5m
wkCwAHCK5pwaK+40ww9UQDLQZynX7SBhq0CL1IAZqw9C7CwS+zIYN/yom5n4MleJYqgnPGhSEkLG
/KtIQQ2Nq7M5vnaKz0MMpCP6mhAzl0Y73wiRQk7ogtpjPeL9bkIDbdCFpHu0TQCNWW3ebxZep/sW
chEk5XKk06cP3JniNttWFsweFV1x9a1aT145Apq2fmYTi2Mf+G6BVb7Kj5z4j0EW3tEsHLyM/KgR
r8ORHU5BuvjqOGIP1Wb91HnMKCMGEVpMviU4LxJbJQDYo4ONtDygFWlOQ2qM4OoeGq+P+UKoxJCi
76PxeiUfLdDuSn1u9e3mEn9BC9mzz3mrUGsXcNUcFoE7C5+oMa8bo9PBYpnFuiBRtAPtc0ivupRy
B5LA1KRnDp3VL16tt4u0ECd1f0rJmWqYLG6EqDTPhnFvNaIqo/p+WDVFTMIblckr0XUGwu09IG7I
ojcebh54f4CaaiRQwZWVEtVrFlGvaTivzmsDpKy4b7zQbK8qZ/acxqZ9TNjpERlaZc6XolGg5nsE
zKf3qLRV1iYkOqS/eK0Kz6HcXcX3KdE/5zWLdcfheHaBSnUc7qm6UskZ62SSmAitHa9XdqtYatTD
6OhrT69rp3tXNSrsfjA/nmae0kh8KlDkBleCHPSgP1ikt2HVp3Q4ZBPbDcoPFHUggTqtboDVeOMv
paZiT/iazxqGLqlCZuQujxacfHGKM/j1dyoykxEN6cylmMq9DpI+8XY0iG2ebc9SlAY4V8ptP7nM
hqkObJ412DjwpyR21wr25ttUcLTEGjvAZkETNb80Y8UEoLpquox81+IxQIGzr/7b6IVBOHmMZvUC
jiwj3ub4yvsAs/+RNwagiGurA7S1/u+ATAcayEWWzZTW3/Q4Ty6ts0puZXxMQxBr8pRdhgY1KJDl
lqewZxXppMVBTJQ7hW/z0PAVcsMPPLr0dEVYb2A+ZAQGjcY2ZZ/DRsiXvDWZZP2JArG2A+yTzkco
JwjHaHNO2rxWi9SGYIHuJ/PNW6PbqcUcCvFJDSH2twZUls5OTI81jqPtOQ37vhIoJFjhq4Lg/YaQ
aQNg1KAdjr8KHlz/fcAtlCOqsK5I0coLie5Q6FCRkIBmpppgIWTkBAPveTJQb4g/wnbs+zVvq7Kk
l7m/NhbyleNKM0fOXrJ9aIEaGUrTjuB8sEyJHeud5XPjODYxc1EQ/UJ0ewadaJ529AfvS/SuQ4+B
o+P2KuT4F750D2GZ/jGzKJlNTCO20GBGkwJxxwK3chlPQhQukj8IspxyCJsujvC35heXXo626kJf
W5LpOS/K3GtQHXG9IZpgzaRxQ1wH8p3tRRo9XBGgv4FJbX6GGveednyNcJl2/zyG1netsgzk+aKQ
xW5cDjNQkEnyH3SODUUqBnL6gvDW0fLRIK/SO9OiRSETz7iGu8zuhsdB6WNP1BnzJ5OmNYpktQlC
DylYPm2ELhJDzaYDqfjT8aaYHT8nAPrV7KZWmCHnBKm+7gHolXnxldZOgelopNqOyQwYZGohkVjY
GmB15fygLSbrjP4QRZ6CUcRUWVdFeoEO5zSEQyZvea7NsXgbXpZE0hZEz0D/LlkgxbKXwXu5ftoF
usMH+TpXgqKMqyVlfZali//axk2W3rGcjvhPQPwvvZzLyw8cxI1JIU2zEKQiS4rBzuVNQbLYcjUo
wj9GUyyHw2bLxXcnTQ1Un8V8wyMuJ43RX1t73mU33XcbTZaz/Oaej4f9BVirrlADrfEqesUDVess
0OFBV28VuYL27Zpkm49aErJasVDi5aFYyD1l+oLPXasIUsow9tOhrSK7C71rVutnyP6kN7RgE+S6
nYXFGkEs5rh5r5fQGMCUlDCQ+R52EDjD4IOBMUynt9N3gs8O5rENTdwII0OdTaplbFBBBbbNUCXJ
wzRINm3GJmgIVc54dzlE3apqVfEU70li6qNzRXX/wzuYODnP6OTHQ+tMphCapVgMaT7pWMpRfNHp
SP8zDwLBwh6KdqMJUwUUFU4yUnXrOkiWJi87BHkLyfDFw5TxWW6pyQyi0zO8NRBabQMzJEKMISTF
mzt9elr9w3R+8zRP4o0Vm1lFKUp7LprZAg4z72+lSRE0HIKFOor7Bp31hM6j/JrqAdGILfJsNMta
tQN4toIDPFqWn88Y+QaI58q7XjwMsGCptWmbthLswtcQGqEw023Nw+eqq5LSwgh7xNS/svqV+WRz
DehklWjlYFQOMDSL1aOW2ODMvRBi5mYZJJfFCb23FPg39SJ7h+KpQ457DcXhW2WJJLSUSTDfERW3
Fx9cw/v+3AihLfNLEevGFtmb9jAPHizszOnR20K4sIUigQ6Mo8fSnyf0ebl81ltKaIn8HWXbCWwh
v13AzSVUo96H5qnEUnXWJAxBPeh4kF2IlOwLg3iQjhVWt0tGzHZjPkcH8CQ9TpOhOkNBpg8D3g3M
cuef1omvpsXVXM9Fy6qZ4Qy8S6VtBeC3qD03pCI2N8ac/xfYl8Qlx31cJqp23e5eALypwEft8QZ3
HCgtz69H7z05muGGJbb1efPBIXKNcaaqQo6SjzzV1VVu5xFrd/n2E+eZHWLYMMxwI3srKP2JLaKc
RHjo2Jk9+IxG9RP1KXZiMBJx54o5p/kfXoQgv2lSH/pQ9BcGCHgMoZQTuNvhTp7JYh3NdiNHzMnE
W//ePWGx0a9PsVjR5Ybh+CX3bWGruIprV8pVjblR+qishKhk/5mDFSLJJ0EZ5+81v4e9sXdHjAmA
BRRi419rnXaU7EkZp3wGI+lSjuKmJOzuBac0Aes+g754Q+jN0Vh/VHRV82Y+wkj5sv8WqJR+FBxR
cajLgvA0i+z/qdJT+Zj/jGq76rDb70y+rWMJwvzd7j8aGVXj2wGXU6esKGH7yelLkd7sln26FUct
JvDF+8ogPX5Ug4Q2jQ1b8scS4zStqd5cBSkX4HfwuIRkEROK2gaxLtVIq9zy1LAxdamQTiXS54fd
vgTz/cXMzQwmNUqdgexaArDAt/A8dKIvIImfaqAf1EHNiazT5FDoHNN6qHxELI5ViukF9k2u4LdV
c3DuTKC+DQSoqwbIFiltg0WvkB/L0iFCq/M9BCZ3ivkJd+/1wH1rFzLXbsPocpBDANzDURPrt3Iy
wStQPcVwx2QKCUWyXb1PBpfGLBFBcGb149jyIzSi9qYyWnLNP1QPI5kFADtl1hZLcM6AcVp3IpPR
X0ThxV5/dHbB5JTl8rt+Q7IAnqhwOqD02Oy/eZOUvJVc+KUGKQE2uBWdl7OGHMURqBvg+W1xLFR/
zZzY9hJRfk44NNorYkB5bVJkjXlP9ak+SR49nZl9yHabqTFea9I6QXBxLDEIsZRh+MA88SsJWtWR
LA9iq0UWKi31D8J29OQR+eE6ZDBVnHSgHTnTTJ59SowSHdEeRbtYttSuhZGL5gUEAJNQ3fb1udS0
2B3KbYIl/c4vq0zV53W6g99rssk2z2vfHb3lRIRh0ipeqI34KjvNZhJbJmtUNhpelEZnH6xkeceM
IIuFVq70cyLJCQerC0Y3lv/kyLiwJtAKg9jcYc+s2AByzRWuLBUGTlEaULExx1s+ZWntzT4X+iTk
ZMAvEoBBSLKZCWDVnsEZj2+QxmXJbh0ZsONsntNyUksPYfr5x5ZzDkaq5rTlL0XQEMFHm1vRMXp1
LYWztXu3v1s+l+/DmnGojUuOfGYocy1zW9zWRvX9ZkMNEOp4lIY22EMMUsLQdqauPTb4XHDd9JFF
qfeuQK0rBmfB9D9781OtdzzD0HCqT2dLBQk3QLh+VzWOwbJPYnoYDt0NycNlskkZD0XAGXy6Gaym
La/wPrnQdwL/fswuClZIuQiBFlxBKkdbuVL+XCju55H4qxJ9axnag4IPASy49iZ94Atfl+MT/drr
KSFiqj6RjRQ53rSlQ5wCV68M3MKZIrKys9vZxFBwRKthwpXJnuy3nUQuuSJXfmn2HgwrzJIgEmQd
/WvIgOgj89A1Ju9Cekk8GyF62+WYZfMzau8B1K+svDPzhy8JQ7WOsmUxdof6s2sL+4LLBwn44GBU
7Fmr5PE/2tNDeSYfNcCONEshke66hop7r9hf8SGMm5PE4YgsD3Eu9NvY9uPD2djlpCBzGPbrcSU7
Y660X+zuBcDQyA7ngfn01j65Fqbg4W4xWdN6kRfV5TGq+n29yyP5IF7giFtdAyM6j3H9kwcUQZ51
EBcztGCkp0UP+Jy7Jr0OYXJzZTQmIotVl4/x9+BICN3bJsV83cMiMiaxNr9vOiyeNhIXPCEHRzlR
i9W6Phh5N//wv7e8DCEV9A7yXLJh2mtXV0gx4/moTjMkapiYSroN5H9pQ6YDcC+sxywO7hQtfa6N
TuWwGTZw2ZIFEWufhc7Zw1t2/AK2x/SRa+Ufj5N3Dtb5nlRMrEH2cCgOQr1huQVqFiG3ickbLx25
yWLfxM00e0LKgkHiZ/EtLisO5zeqT41Ee/9qwVGjCQBMVQCHvFXsSKoYSyYYwU8/8dEHvUF9F46c
KmwzCw1ZK12TB2vaLWy4tEknaFBQ8sJF0kWOxCQreJpKFEAV6C6vei4Ev2BIy/T3VfQ8f+i4qVBu
8vGWlDLwJvdMNDwbG/tc3RCEvnC+fzL9bKq/L9UdBfwojviE5rlcNoK2g65h1KJKpR0ZuhUyX81H
U/j6t0Mffb/ajzky2jJNdmd62NluhjsN7KanFC2u965hUkv/tH+XBG5kD3Swg3CfjKCdiS3lYcfN
fH8rJyLUzyzIwhlnKFc5BFJBcP9XHbG9nFAv0sTHVoHLj4n3ux/LuNxgPKbvBHIehqP6LgwaIHqC
s8hDa+y/olRBalT4zmGCkmGhGPt3We/5VU6EHMci3A9RTM44BRd2tJDk2mt3uS2cCl7Dmmxje5mm
fJTVhCAJO/BklPE2C/jzRNV4Wmv5qaXtRV0h+FbAeNXJN3oF5NGbfNWeaxO2CN8wHY1UP0M4/Ek0
lKqhOsDqZGyzP9fJIprKT4PhFIEVzZgJrpYgQkxwT+FIPrkk0rI+XtrqdTq6s+4xPoPgD7Q0Ek5x
3iCMRxkqGLqIA+5QxRy+fTIigDlP8XaP/a1XveOkBC9SBBqHQaDdUchLbsmAQu0UjSu9vHvqenyp
uZNYS17CSa6akS1D+6U/ffg0a3gIgMikQOuLX+TugInGmHWKBpCh1eCrfzDHnzx5YYW+eezoV25T
g/Gq1NE7vHE+7mLiB8rV+g89A6ceMvIgShjSQvvmBMwCBUE+dqOjpLwLPNdtFnZLzs7QuPpD7m4r
VcIbfDTnl2916zds+rMAg4qrdMPytVD71HzqILUAdHqu325Yk9dEX7k/kkxWtbiDNo3sCRyatSQR
XbtiD5F4goK6z5uCVc9oS1OCLIG30CKPOYPVFCz28uXHtqv8JGaWKqmuFXSpAfPBaDiqgTBDRVzJ
Zsn1KKWgw1SkYagrLu2s4+3kaEmBTLv2cUZXTUlF2ZIBKh28bAurk6tjBBvy5BWFBzwyIc71z3Ed
WMJHPOq18Lkezig/XZcQkoFGSXJiHMVXP7qp0c2jgr9YE+r4CL2NQ/luwGV/RI4v/FWwSX2zhxe+
PRwEpa82jUw4Phm/QbBIAMZLZEfBtMHu0mDHLewnmAkAYL929rfhZHrsZEKXsVw1aTDwaRnoJKj4
n/7ZyrbKud4z4QNPq0THkJrQ5jqCE4ANBtmlSMr5bd3J09kWjw0Jr/NoGCThdsbIXOFn12wSEFN0
IZX/0tf8HnszSYj98egbLK6v3N4Q9vFQcIAGlPYQbgg20OnKqEHDxeRUw67LXliVY+lZ9CE/almp
yFGh0xuf5e+kCowhPqfxxxlVd7JnWoOOP7CGQTql80Re/M8uw1AiCSzNg4SsHPWqsl0+sxV7srZX
CVWoXpfWipEFrkDYdyu5AY9XtpJmKT1hx/zuaRzZBKNzTc0FfmrelTWJBoZeIYWEC/NUfkHzpNeS
TrGUshT0hB0TmylLgmE39ZizW2d2UBhdqBAagSu08rqMs56RKB/6mcfwmYsYnX4UNlcsg/xyYQKq
EeoY61kJ3QsKthybT/7SQWsmg36MwX5eb4VKK4yA5G2On8yF4cSrNiNlx1BzUbRuAvzCNIpdo9rZ
VadsmqPfhes/Osn4o199p2yrWp6aDufUbsSDmYYyrc3moFB9a7mvq5a3nm8ttuRGX8D1huQImSSX
RqxXuEjQM4ljBcgrgLz+T1s38Z0J/oDu+dFcPjau3/p41IKWhNSBRDtQkDjV4r6MYfwhzgrstYKd
dSvjvnYF3ySQSTzSRDrvvxH1xLyrUPRFczR2AgblPhrujgY9NMgE9XD1J2GHsfXarYqjKYyEPhZk
KgAyCLqag8vVLS4ErNR9Zh3/V8txaBvMTSioRq5Ctms0NPD9Oh8OmYajhtGtUXCZiPKloGwoyG/C
d9P3Zfd6BTCnATJ00Rl6OJyJrIIBumNDr6tZC3yuNWh8KtGh2+Akw3Nyz1IQQCRwIwJnnTx2QM4A
60C2S5gCRFEwVTJZDTrXhLZBPpoqpotMGX5gQfJ3MCs9C4ooMXEGcPZlwwv0CiTXct0Q7DthKnZZ
oTm7hG5uExFMlzSyps24omrucW8M5ADH4CQ8pKgMgLyJugdtR2o5j/bZ3vM+IkSt9dUaLH4adMP5
dmx1rN6TDKSgTVRt8Kr5GXNqDdCw/9YZumAIKzNtWXWfmgDNcmDGSDqrrn4QaYTooV+5cIOa5Kpy
GMqdVZFAfFtXB/ZGXkBfrQYjBwfYtbhMlxPKhkXfDE3m6AmlPOabauJhb41Q1389TWbZnxH9IpMD
DHbk8F1NKevE3fsWVzezSBqB3aJq3qE2a4yqoe9/OqYO/o9SdU6rYklnT4bYo9sOesfG6GtPebt6
LTM7PJVU24zVGv+NPpv5rqqdiYKUBrpJ6/Keg402oDaQElyDntlreURnYAuTMjvuQZP67ObpnlF2
r3H5XsYPdM52/KXOk806H04kWODCxTWb5s/yIlVDOK98rl0qb5gGAffAtuoUT3pO/P1h3ncYrECK
A5GuM5/0UYwLT8Z9xkElbm4LFagCWUp0bUThH721WN6CR/Ip5CkYCdXtMkRDisnoOMSKvU1KMiZm
7HyHELbzgIXZjKFILYvDiQxkGtUyiHtRLCvfc4qmQyOvaqb+kHOJEwmkpckyKklpKZs2sosmDnPk
fci9KX0t/lYd1sEzGGgOaBuwiLi/YQ7rbTXEVMQ+dtKH5G7nnToGKql6WygVum0eo88ovQFWKf7F
0ssEDOmtiPmkM/tUNbk0LacQ5DTDHK7DsehEvaZ8q5I42PQCXEUOokUlYsghpJ6QkOCRH6hdUv0e
lJKeGY0rRPqZljgG6eUsO36IHr2Pc4o5NoXrYM+07hT3gQvUOsXv8TWGEPXu3j/2bxy6v3jnrzZ1
SbB/BSjybWoX3WN/yiyBK3iI4Pr3yfGlfdyWYmnoG2jTxBGWum4T33xaAf5E2c1kAg72O1GwgKsh
DEIm7Q+rU4E/OdPbSZKHysnDjLUooiyskqy7G+Q0z54Bl+HFv08HllmKi8XBM0tAgRy0JuILZTxt
YOEl9JwUqFEjGqlnyXJ7o7uJIv7y7B/wraaxsMoHBJN0+VHVdgOAXN81mGD6eJwU4xUo/0smzPtN
v1NzUy3fY6VxjtFmT6cdxGOZ7nPP5Gt/foKuYluhLyNlZ5L0P1DXoHuBnJ4wc5CwezQXLgNi0EMN
1DvzTehi3xERta0zWEjjvDO4iP1EoJcnHZSlLWq/4N/OjEaw+5XkUO5zaqHQkh5dBw5ZtZHBCHqZ
j6C9hxLsvOh/9PDp1QE9uyt3gplPWlqI3zas5UB8zST0ku1sBrAlgnHYgA1Jg92VD3+jUIxzcDDn
fkK+VWO1sR2dGA44Tcc+CihwWK/DbKN9yfppFa2RO9Mwi37vxHPvqDbllhtwNVEzezBtJU0FIvuX
Byqnd7aiKG5i5xgzOtJriqkYDwS6knV3Tc6pIyD0ZDr7ddSfdwF0PvFarnRhOYwnH4dxH4JuV93Y
dQprirOMD5k7lEDAjZlCCchAulErFS6YZ5t15maSu/LjqDk0fYxdviXxM7/b4e/IMfM9hOGA2cSk
LchCYvZt8GUGS/5PpmX2UxCJTcWA1eNBJY9g5XWrNoihYWZoDjbpm7b2b6ut0cf/E+ApXhOl40QB
x1xwKI0BtFKsch/X/e6IprDOeHSulfFWvhRGgagxdgFezoKNeVAi/Naw4ETzB9aKShbKINsJOiAi
FuAjThNUZ3U/BkzdFMZIBSNFNCMvr5cCJtVcG/iTRVP+QH2ake0kGXbUiDEa7Il0zIQS8Rb0DPUQ
hO+Go50ttq5csvmjSAMI7iFeMl2aLIqw7LHJu+6bAdwsJCeLeZarzNxgG0yVjZrnCWwOjKLrOif/
NrfiShOd3ZdSYzveJixv1rzqeYsZaW0H9A0NM2fsw3LjBQDoSU9UqVzugpn+5JeYg3HWtu9kNyG7
vL0cJwM6piBvJk4GvrvNXGdtoWMkEs2uTXGMY8BJqc98w8yOdZG7Uc+J9V2y68lcIy/ZVKvzKRVQ
XXwbnevbwtIaXg7BsTov+BCmBdsLUXdOA62GcprTZ6YNjY2laKWFDfrysPmdGDfT1uCXtFGQXh9P
UUcHOlN+dcWVl7y9pzNYyLWSVMXTb8BWGmQ+IfWnBZIvW2zuMi8QHh5sHRdthF8BSrNxCHkV9RYz
QlHgyjmN1OYl/KVBLedubXZQ7JCqJhTje/b2ZmaTvH0ReP36XQiPvIzUziK4rOJVU04ORjxt2r4O
mSclxjKM0mw7zTk1xuw2tCAecG0ehKB1BeXMKh/Z3LWft4QVA6kqx8uXpr1dGmzHWmZka7TnFwrw
/z3Qse3UTRjTH0IAOr4eiHo4DHy/n9KwHxYSUzIkTcaZGZ4gXal0LgX21vW5J0/EAN9oXpAuOioY
JFQB+x9kify8qTUGNPmByLbHseLr6EJzQxL2bsrmX9KIwTah7/cFXZhUi5YOeoboxpEvYBEFD3O+
RWWv40ONK2qTZ5lhHpdJ+V7hDSKJdjhX+rRDZDx2oQ20mYJhUNJP9QqwVKzqvxaPCJAk3X31rMgB
/3Xkv58yButOxayOuRUvg78w9/ZNy77Pxd/Iui+9rzIWlwxCgKhrp6J4yvaWTx2/lbQMe6vmsS/A
3+x+K02SFdnIpC+Y0mfCdHrJlKgmdO7Si05XvMR4Tkn2S+eAIrhgbvmuhjvOYCR05dJqxkEvfwaS
gMqlm9m8IMzGvp+56ifJ0pW4KaQnWbzBii+1upXKUlyfJwuGXMPJ8XJpti49HL8RuFcdh0UpXwM9
t6YXfAZv4ohGyx2VaYIU63LlDkQVyIYnANQsG+ZY8VMD/FF987RqCwlYnx8wE0SWTlYpDGiMGoEO
FKHAtT124eaNFsYNvniFCvwXRT/q8snPR39ZVh7EF27mDkp7qty9nIMgfcoNa1QxI3bk+A32/wUF
W7vc4+zNfs3A6aW4Y8P8ga59fO2x33KnWoHNkDFH8s9UEpjabLPPACpx778k4cYTjr4Zna6cHmwG
32RUSR1zmND5uubf3V6OnThqZ6JnT5xUphkQYKUMM0ku7CsURcHWEb6K1P5fKxdZ/vpHKjc+rzG0
ZoCXsHISl5ir7DIQYZtBjPhMA0Y0zb/JSIhQHbO+sW9ASTu93vzm/r88ndokInZx3IMXnLNWIe9/
h02IAv4SxUe0dfzrd7b9dTGbRIV1Fhl4p3FoY+/Q7vZygJPL4hIzzrVFMaumGBQFRPZxiwRVWCLr
dY4AtPjCCC/OERubpilRf7dGv+yY4KMdCrXkMcm6i3OCYVFuGsaf4vU4GGna4EZ+GfgSxrZbxfvt
+OkcKueWCaICmWcd2EetsGcdItDvIY52a6bb24Hg3fms9kcevbD5JDrZ4hHM4p++zrSLc5q3bTOq
LaBOS87O86BZ1EwWQ/rqLUGipC2Cb4C9FlW45dTVjGzB56fw3aDQ9e02WPQh1ZmLDqHx1gs1+TiB
+V+MubMcY951PVvmUq7AHzjH+PHuiO4/aBGuSBOe4Jm+gFELqDl+rAhUML11Ush4C1D82KlCRZho
0pA8Uy7/VKitfK+3tuRRMYY7PsSHxShsitqWEYqv7e+gbBv3qX9DBx0GDiDWWjCo0EbIembqIAZe
xgNy+R88gLMFqxNoCgFuM9bGB/26367BCVosOMNwdBr8ncvmKmNbnjolYhZCbf9z4TItHdqeaGwP
35piKfOeSx9LNI14muM5hcAuZLRUTEv1lf5OcS3IpRiQTg7Ht5JCbZlvugJHuGjOcFk6YPjtRJ/R
DSjMMK9nqaLZhIoDawn+pzBcsnPN8yYnDsnhWi7XnakacY9r9CZBoaQrnai/EhbpB9w9GtVyecKI
0AWnYoynVXWqnCxWENyG3H0JaMswlycc9YcFf+DTkrsR/v7n4MRIwAHAE1ICtdsqO5zAHoXbtxwY
Bks7kmcPCmiRklXN71L6KmLD8ztiRMnkUHKSJ8Hx481Tl+85lPB5pHR+N4AP7OABkP4YWZ6CAfIY
Xr0TAO6rYqeFDy9GwUK35tJ12s6DoefUUJ0jPNKaP39vh+0wgkVOkv1YEagi6wYHbUlgu4ZNRNzc
QbPlvdrEYFCSO4XcLKwgRaa1RaUsoIXPE07j9SpVSgbiuizXC7ofpHHSEM+sovLh2xNAfC3GH2lu
t6vL9ZP8GvPeBytYYkNROv30DFeFdiesb7NQlv6W82zZc8QqAsuVKJ2aa7KPi78We46MCHx6XdHs
8lWgPVoxErrFSTdUOhXeXuulN9gLrobtAD4O4Mv8pVMMLpU8F4r8JRuM5n8KgVanlRfX+YAQltpg
qNEQKwQe+gb/gDuwptj2hhBoJkWSZCKj42E5qBB+4lmgnKCD3r4SKqKYclo4HrgWTVCzC9kElKk0
OH3Jextx11q1WWLQi5RB2ybYYGLb4DV6vIGq4PR3AfSYU9nl4rNQ3s6MwIggbywjp/dJuTYbncIp
vtrfBux1/Ceoox7pP2VWHMcLP0TqeVgk1ELVc3BqjXLdtMvlweTho9bp+a8h8iVFAy2Ho8ue3wAr
He5kzIC/QrbTP6KCb0JPrHLTQLswN5ft4ylaBsUUvHKg8Wl+IMpKvjExw9Wxu9VBLeNStsD4Ezg3
pWD2v+eKohqAPq0AkT1bpv+mPce79CBWCkGgeaxTFnA6uaflFsP+u8z4jju7qjAKIVhjAjH175K/
Sf7WMqzQmfEViZ6a5JkxnbbxXkDIuLnkv+8cJ+jNOVRD/dw3WUaX4jzS6elc30Vf3TWeDkFqwp21
ElH7R2DyC3MIYs/+/X1H0sJiMNUrZU1bBpLVfIlo4a/mcfoDWxE7yXNDGG0keExSpoVS1rAUvhd7
zfgFwe4tKmRsWurCkG1OYgLYngRDNApsrQoCdrSWNtsMeAmjY+IMjPCTXzFbNSVqnQGxEefIlFi9
lFzhzbixrADBuUZXzlRxbYpmcquDKtEvBT3GhoTbY0F0tMXfp9uRPY9w2rHrUvta61BnOEYtU8z7
K+209GNVkXJxvKc+IfwQGHK30EacrgpqtkWp6vgGD+EpNmYcQv0XQilxHmWlkDqF0q0dXtmM9tEz
TDrvlTvoDPge1qTE3sue7q5E00ws9zdHV9R446WZWuSoW/W6AA3wc0xXqNq1X6kzwca69qBhpsa7
xnXulFzom6Jd/50moLcBydoXItpQISLTuFrHV6ESlXV8m4adZSQyQ14KTRoQpqXydP++4ootGpVl
GQrT15YuzgJKM6ejD0G2Cri9fvKbN3OGqspJWDsgV5Xh2WW9jCC4Tg//e02PYyjDCjK/nXEsVTnI
csqxAxP9aQnftQ5xCPNq4o6DHlvZB+irtIBCpjzWSG2FU6Jk6Yvdz8XQNu04NnsSgXs9r3QyfeFl
aKUKoKD81BYrIOyZ65uHwjsH+frK86xRqQyu1q8S/ftWwb2nHfhxOTV2hpWCvTpt44XzQf4ST0As
mHE8Nms6ujOFdkM+vZB/ie5qEo1ZCyQYa92sLrbPOMnIERcw/cR3hdV1pnwArLfggke6vGGS9D/t
vthzdsMXKAwz4NogLyuL3KCWyjp+K2CiabvdAehQb4Au6ENa5Hxc/hR0HD73FNKsReFZMmWzOnhk
S/YD78U0zGEIYeh0qUns3awYxHO5wdoDicA84ekkjncKE0b2yV7OcDjvNsqmLzfASu7YI1APZUDN
DfwU1vjPqzHmWWTwNi9dQl8WzvqJ+fPO3UASkLzP/AJEcJUFoG+wgOub65bV5uvpSNLzsjQRwgW3
LeOtnWYY1pE/bdEbJGcMVHKfEejZyETPp7wFz2P8EBh9qA1hs/zm8V9GxqMORNw88mhaYi8584Ih
CB29SK4Rgqav38s5D0x8ztuRosR1X8bJN4GWPT8MChQeY9pjZzlLm3GHASHe0crBWxtV2PaOFkZk
GiC6tjYECxLaAnjeihGIuAQ/gWRI3C4Jg2CxSnMrG6iWhxIH/G/wN2wk+mzDa42KSou5eZq7eCgQ
N76KkinU8kedS4/68AE+bzGYCXqLgg8gyL9FBfy8u24aCkwfvuNzSsSiY9BXOTkUvHSVX1QcHowh
p1Zs+lxqWQ3aw0df0MZn8FjU1GsCaiSC3/soB0DumtJo4Ql3xu3nzK5SRQlAi+0V1++fezCvcu2e
I6Wadm2bJU5Q7htH2voiH2dkiJ//La9Ja6UwkbyeQv6WL3hXX7oQe/LF5luJKYmp9eh02dZmQDgd
0DNQ9rba52GbsbQa8pozdFu0BRWrXIPNcL30btEkveBYeGaukMvRhY+8mx+TdUxhJ6SbcaubpykV
EQSywl8rcoZJufkzEGIe27aXfLdSe0oHM66azqkfvmB+Pv9fhsbDu5lC596Z0M4V2k8So9FU5/cX
8M1kb/IQgJ+tAnrow4ph7lQushnoxWvuDpHSk8q6ncLnxiwS6CKdXS2z8N6s/fkk4NnYkGj5o7ku
0wGGdfJd1WcaCLijl3PlIh9+AbmNSLenVWcSEKy56pBuWXaKXWesjPbADoGLHDLdUNtXAMDv081A
SFw8XlBEQn/Z2Yr9IEtrd4ewSAFETOzBPahXSaHdDZ9ydqpJufeCAqMd+0sYQlt7rCn5W41QCwq2
Y0q4oyNQg9zssHWoftDVsWSNMey+72FLJAnfJpa7GsqRo5S9HtG8WWhl/3lnl+6hw9e6cj/spTiB
Lf7ruvQiZ7p19etJrnzcuHnfk3ZervLPEZVp+Ke8aSrPgAuxSjzdnqlwC460rUBTtDnI3CKl+2uw
8X9NLVz6UFmGf3jrVG0lC577OGb5KRi/fr7ASgYkbNLxbJ+bGoaB2u28+9x00IUx8oAwkHOuc9vE
oFd2BM8vldu2zUbfoilkZXpRopaGWaWjLuIrzCxj15aajaPLap+DwWgLoJ+f1cEGJtpuk0LTYvjR
EVrv48sX7sheSOpPcc6ZWwLJVIEuSiVCgDDhieleR+hLY0va0O5uvmQsjOyi/Qq1Wb7thwb1tMXp
Yjb5v//xlAx2yaeayBTVMsZMZr4J8B9YlS9Krrna4fsB0aJAtpwKBER+CwY+7MOsIjBMUzH3i1lZ
+4ydq4eAF7valQDpwC6TkNOxftDBawEQShG4Eo0egQeLJm6RSXxw0v47B2vYol2xTVbg8slamYAi
owhCrsSfJZLmnspF/0F//gc/i5OCxxSFI5S5FsTpJiHBD+07HVwR7yXiKnZ+oOLRR6xq91oG1oY7
w8OpPalYlIt9a6dMCBhFsd8PsXqL/VVQbD5ZNat8qW0KyGvdm6Uqojz0GC+xEiAa7AXnJPmijMkw
ocJCFhUfwHeJzGhvYvxB6f4rqGbk+sOMx5CprrHL9kUrBGh61/d/6fnQqTE1zmYv59kEkRY5qY7b
21EzBx1Bzn7g4NVbWPJcH5wnbfL5v8iCnk5tCw/z8cmqO45rg3Sk9HwENYR8i0H8XMXe1mPxRbXA
Y7LEAZ9t0UMAAzK5uCIdFiUFnhj6ehSr6YZKR7mLUnvZdnce47pxkEY5nkozN9qEqva9ZSuFA24r
H6swTMdudNbHYQj2AOU25XqxK4NVl3ROphO+bwgYHEBQWZzpIWayl0LavsYXXs9kdNZsJtSV3pym
5c6aZv+jKSaVPx5VuEmImaG7m85Pzo9BDLARVOKkA5iw5pJyGmOzQ0jvjRXTpmJ5YZpbjFnUhYL1
YqIBDSbHSE3s9lVav/5z9miWEZpT08vlH/sevHVG9Wm08DP95ZBMFeyqRa6Y2Y6R2DLy+XbLqAqq
T9uVHi09H72JP7V1ejNnHo30DsHBYPYVUu1L8IXZDbqxHEsINbOkbNz2DaYA0E4sfuKCvKDfAwdZ
Xt9AwPPi5WiGHDlvhyyB7oyLPWL0NnhErOsqhbGBpA02o8+h/VrN9ThtCcoiZJsq0WT56CUDyZqB
QCGq9a2DVV63B+KfikeCPHzqsLZX0zhwD9EFmYcmSo11vBniR6TJh2SgXW0g9qOhlYp92Cd/esqZ
8F1NxcPm/uMS8S6cNwieUcq35Cwf5TxPAckv73w5YPBIFnbiDToBTF+kMeFiXtn6H0hsY5aEYZ1M
RWEMN7wJLKY93gjciPEZ+bMJrz9IYKHVrkgHEmtnfyafGIqrv4PhllXBjbIcm64TXUzsGbq2IdJu
JQ7lQLiSLNm71RGhlGQbDyD1Eddzvlf3lWXRmsgPDmS0EbBr5sAITu05cKMiDqtdmIAJvGH09s/j
NtCtfmikq6OsnqPkpWmJcCwcPyYdrb6FCErolxVbmi/Sw8aVN2ByzqpoBT8flaX1xMecHiMtYIar
2PlJn41LVKG8GHcDhN7NZ1L/PVWwOCn24ydWm7MMTNQ4mxzTkRlLbpcG2P89fUvXIbeFCrsu+lUA
mGnWt6KQT3LLWVMk4b+ra9lOtF7WQKGqe0yOQGsQR46YRePVqypLAxAFnMJMhp4Kbxdq3jDLOEk4
CzteWFjJ4PJB4NCBFNSSfWDONK2F8o1A7/0jtPmLbhN7y5EVBwWi+LEpsVV3brM04lil6efK8AMK
9mIVOkudQjcfUFpKLV6ISu+oxUbBE/JHBTlNC3icV2hwGdjhu3uZBgxYjVE8N4jz1SvodrF35FTq
gFhh3z2Wi4lyXaJpjvpJ8uMEKmTcmlPSmSEgJkkA60GsS4S3c1BIftCPzItNaO6DcbsQ40wK06t9
3TBdLUfuxkfSaVJUQoiGQkrcDyXmvitYsITJ7UpC0BcZRGIN1dZtfCeRQGZ8R2WiwjevIt1/vcRt
20+xRURBNfjHsyb3q7TSeFvBTzRDo0uXoXfrmQR+v6auyhPBBRxcLNcIvz9DjR724hCnky9nyHZW
RWPZMgzY/sTA0Vb+HYdZn57+zAq1WXm7xQCSU75Ft6i2FxFpoAxBomB7Mt6deJHXnpyHQkibB5Df
50JEe7hNbxmEGQg5SKJiEnB8XSVdnq+Zon1wQHEIUyaw/97zKHeBiKEMm1NN5JuqgLRxC3Y7na9W
1o5p3ns1j3Bv019LEcnZbTpoC8BLPEpx+6uU/nJ7uI/NJ3CuUavL3sVuvR+sxC6US5bZ31QrxbdC
Qev3GELrGOG9kw6cxqxz07NYPc5xEaa2V10Q6E6rUQbT1ez/8tJ35dviXUWkwZa7APVcZQZ4ALTg
8m54wdEFBZjNQ+AvyMyxPRe4SoddKw0tJn56ewqSZBYMUgykIyVAQyy8IBDhTnu8dZpCe0IdumRc
cZWmkYQjk+2cB9u6+aLi2TaiIgphxNQCn9pGnHmd7AbUV47YqNLeVmafXRIiCNcg0BwbclQ/cB4u
N8IyCqxgrsR0te3+7v/o10jeNmcZPHN1DFDMrRSDXJ38aGkD+WdOb2QL/7NpijkRwZ2JLh5/bM1P
e4MtYcP9s3ruNLJ6XY0v6XCNd4FHepN5L4F6xCZMjHemG2oP7uwDpjDmzPVQwu+InktUbaPRzPru
yWlGUnqCuf2PTfqICu5xcXudN/bwfR1rhTh56G6yodfOoS7dubfePzALkwIu449ERMTe1bNXLZ/f
Bk1LbElFnE6XkClFbYh82iToZMNjZ4YoanR9aBCs8TD+qfDIn7HpRaydCS8dphHao+v/gLb0oFeh
n1fMylalJ9oxfZuzjPzijLSSUeYZJ7VzfiYSQSmBv3ruiPz7IVDBSU80zVwk1/A+zHCDb/TVhid2
DEYNzOZ9+5QYCMoXntIs0lx4eH5yJrE1JFIkhC7XbiIFhWJOf9bsp9QB8yhFkFRlaRecusJ8Q13E
mrDcP5QC3GU3pJezFkqbdzVSgdngQlAR7vXk48Ciah80wwQpiw4YSuSOgg7nnn/R9kG91713DNw9
hIJW2L1JwRtlYWXmSQMolDBdHxKZYeYa3DcVz2wIx+SthcknDP/ea2QIDZ98joNoH/bxu3Uj7u8c
9RpThIq14iDL79Bq9IVOtC5yZpct/Mw8PW2zCASpHQ95sJVE/Vmpt05aBeIYafZNGl/P/lf+bkAM
xEmtgHhZQSLVHNFnZYBlP/d4E4p/hbMs4r2zd7LGqsS8RCo/MMWd6ktLfG/rVLcRzO/gQBMhg6yh
SxKjvqkx6AxsWCSpfyw+y1/eFVprWhvFH91nsp3PDvfkv3nhSZ9xLXq2bx3g4D3R9vyz1+h7Ls3B
hI0aIIs41KWmNiigIkOEq72+jxIyqFVQIdEDIXl/EfOQRVlws/+7ZSmxt4nqNkhENLdPon8f+Xsc
pxJNdWybTpiaDAzgGYgH31xDBEybnAN9sSjXP0MswGaSjeAnd9rv7bax5ygZHu29gA5RlwvcF/r/
30vXAB21N0C396ZPvNq4W7MCNd5LhbCk//zpEhD0xANAHldeFryZM47SqbqW0UAvrSqBvwJM3sf2
X/2KwJdCo98aXEEz84oIZQzS539XqWiLey3Luu4Su5hyxjW9jUZXRaRVaKXYN17hWnjBxnuk/NKA
pRSdHzLNP/IbwOW6sNLO+i+06Q1hh57wLba4dyaVTC+ghEAiTQjoXAbdArP819AimVzjkWhxcG1B
+1OAQuMAUTmzBHTRK2S+jE8MJsQHhq4T0ZY1b7rdQUhd4BOQNc+n9lw+1Nso18caLMJQvzinOZDx
R+mJMav2h6VjRWBgT30wMHQcHYN+mDIvnjv5+i8hnKSKsBgIIOTh7VadMtilZs7BGB1A0WeJqa1+
O1mgQtUtaMpDI0i4fgjZ/p9E/8B1S28wHUG1JMAS6guOPDO0vzQDZAZls7acSk3FQXz4sFbBgC/+
7dEqxGg1XUEFC6ruU8ASVc8MAUY1Gornc7VLQpHcwoEewikt/skoX2E2DHfJSUdBhBchSimkivO5
pjZW0jcWdghq8qjwjF5+mwnZSRdyegCC3PfmA3oJ6BRDr+Ruzcf5zq4j2s14r6nHZStG0rU2kcIk
4zqA+sOuFo6cbv/tC5WXy1gz0FmYrGdbFRe/rRUYoUC7P3m7skeJUAoWfSLUZTK888vTqkB1Zczc
P/Wy6epHXXh+612/iV7vaE9bHL4meVDuDxjQFy7jMpfgSz/0i29/cQ5H/tK1PJbyXRqcIqzgHgDi
7J5f6YvyBpSpYSX6pVebYl3OXH14+mBx/RKwp2gSj3yEs+UNkGS9MWK+1jNbHgxTqD972ZlOH02f
UswXEmkUqiwfMvABsJNhpmYnlY7U9Wzcw1f/BzWpXvf8yiRrshMBP9KOjHPzPmO6bpx3HiYTNrUp
3yk19RKLJgrw6nKhlu0OOhIR3OZqWF7U8ws9oZuDoeoIp9jZ0cXEE0UcxSj4BJ+e5fcrM2zCM545
vgr/r5BerrpItFRWlCQh3Wn3WuEVrDWt5FpcblldFNfWwIJDsuzFGsC7AQlxdrGLa4qbyufj+JKO
blD0fGzgQeFPmUHAWbFb6BsoBwF5vhbyORK4ahANTu4xBlwF1f/GPzAOY+RKDMXD/9BG/1nc3K1r
suJOdhoCbKzcatMqks9fEp63zdfZe+HMW8XbClCC43ZEf+Ty+fgFN07p2tY+CEAZV/uyVc8kwXMV
ZGrkfy2ethPRnge5SMoIP639puDi1aHEALMjyd7md8C9ciY4jlecHHr6Xe8qRgEcjt3r1QrjH3+x
BfP4qEYF9Jr36an201eL3dwgTu88+KEtqCUDV9rEDLaKkaympNKWGTmbLvu4+gVu1oWH/H2KIK6O
pDtGc8kbgfVcPVPHHd+gUIo5HB9Nh2DKEfFt2KZkTFox+F+MqCRbe4qQtabQSO5Ih8cDpewXQp1E
HuGs0isD7Iq6O5PdPoJR5rYbc1n4rP91/3fzxIdqoWGS40cQNm4Oh1zkvWtepTz0RgAnEql9+GpQ
f03wBEXLd/CI6HJ/tltYquCUeiSwSMBz1SiorTLyEJ1tL7//Nd0mp6WjOQ0c8TDuZFCrdJAzwytS
9HMzHMRNdmKA2JiGEKRYGLY/Bqsmd/T4WzgmbiVwaLDc5E0/2E1Q9RfXGJdnCRKezhSgXrxZ5lc3
YjSuF9dq4g4Ks8wTbZTvWMwHyoQif8hmxodCiWQZEbhxpbAduwDGX8hKxGWMnJNhrQXp1G+E5uer
ErEVMIszfLXO7DzmpsClWmyJzlZZNdF4xOM7Yke23jnlK7dYIsc8X/Mu37H8/3Dg7kt3ZQmsGEXG
fbUmACr+S1Q0yYK3JjYr9fcKZngXhzfaCM753r/zPh4y3L0Mptvt/gmEQO814Tan5wUeMUN/C+pc
lxs+n5Ob4NYE1Smcb2K6kbk+PM4gVhDG/IyHH1LRlXlitgkTt6YPGlR0eASAtptFsiLFOn2GtiuQ
7qv8HkSv2cFbZpa6vlXsbvXu9mUQsCtS7V5a+ejSN1kv8ceHvbyt8BJ1cG2Wu66TDCLgZbmAkTC7
jn9xArZBAsqm7ow4Mb+djZlx7MCZh9IpwC+BgTzxtP+IypbOjhxjGzSeA78C2xsEpqeKIyfUpLv+
zb4SVU1jZJChQkHfnONxnV7QHMzH0xEStYL4zWHlSGyhZ/PdNiKZClgrWzEJektNliBB4GUihaFc
k4NasX+pAbhERrwdwlfAsoqQTB82tCCGTLT3q5l3PSNwH1DZ7Q7FTMEODNeY2u5P/qrnDof98h3e
06Go06I6tVrQpLQ0/xtap2v29QNy1jA11Ajds7bIg5KwnqrDzeMdPuX1AwAXMXL719NDZhVDKnzN
YxeDJ2TXfvo3brXUb5mpx6e1Sq03phC45nb1FOERzrYMBkVxGQbRMVuhZlRfh1pYyFF6G26X7Mo6
sNPI9UmWr/47o/fOv8dF/yy/JTHcvyaFq5PR4p/dPVG/HYgWryjLMFjo7dW4fAdpFKmYhLDufi4R
0LK6XZQy7i2fdPD6fsU6ruECE3PzAZz9T8Fe0sfPBFt/rULIvEyh8B18Z3JTM3ZE5ni9TdvxGL3n
DWfSsUCTAmEqth7SVzD1aVe9F3pkTel3Kjs31vpUX+Z5224Kmzr1d/JEkWRzL80I7fqel2R18wNS
ipE+1K6PTJwuGIAlGZk/XG18H0tmmae5ElKrkzwdHtjqY78N0IHZND/Nyv+Il3Z8nxERIuecbUnJ
mvHD37cXajpV7XNjkTelgh/nQtp/iGCK9JlqArsRunqwjsdgrjvq/79O3M42tq7mH+T7/NDCQd9V
QPtNAsvKAYaPvlIuEYDCPptZzD5ZGypdk6nS4NL4JP/zJ8alnVVNSAhIJtwd6isA4+KzdxmRWzCV
daUq6Ney4nc5K0fPfUSV9yz0DCwRJp5bXejcgp6lsfVhjvoN9C97SNMRYEcy5LuKBJvceGX/jbrN
/5NqlsJ9bFpvIlRruhNMmMPksghr/XhHA/KCgGrOuR1HIrcdWl47lrHgwvvtIlt2QhUBDEyLDZiC
lmee0+iSlYKULFWXShbi/TSNXYV3E/H0uMf/Vhr95eb7mDiZJQKLk66L9250GcPWSOcrmnFEnhcI
lRGVgixbp94L4rVguFRxyWU4Pmt7Ea8s9xvhAH7mLszMjoddGUxW9QCF5/Ot5D02DIZ7CQ9oLnIa
VmMHqdyzohPCaHnU3oh/r7y+xWLXz4F+kgIsjvYnr+3Hmbcm6L94l0+3scbyk9Y4fgHBDyy0mQ7a
K6uSXCqdjOHrFErt23KgRQsmXF1nn7dIzNChZWLDFDsSGLlASFkkQ/RwfEx/rxcbb6s+ZwGnNSKk
MgYthv8Im+86DUuEZ2aoTXJV5f+4VwT/DkdCzBrpN0ZsNDc5JJxaENvctOHiwpJ0u3mITyIOTXrx
nlaTvOkhi7I6zAmja0y35t+MMb9TnIZOUt8CmYYweAlcz4VJArUFlYaCwkcMP6gUwiITvS2OPtKa
bPRKrOlYm7lDILAlbn7kTYEf+XTP1aaIpwS9sPPHg+XnR/WH00UQDALhMsY3A+GlIXTx+mQwJe+5
UQtfCsKi7CpnR+lpoaxN4+zkqdAFWV15QZzWvwYooPzBsKVZA6y3OE0Ana2A+0aGThQx0dkoh+Jb
cYRLK0X4FDTOP4/X/6VT3Fwu178KIMsfHvNGJRFrHO+XBh0X3ke7tDjCg5Za5lx9F2OpeDZzlmoL
ORp6BaEFvsB8PiE3ZNnxisGaRZ+iWtmb+FUaa7oFGFBG95pRRPQK6mME+cHzGRNrMJ3nP5rkfi3x
aK2TdyViyJRM+LJ37R/BC63Dp9Ndq0VOZq10hEwIVOiLEAN2bNhTzA+S2Ig1oWyrUww2j7JX0Yl9
BqHHIdbx3mfI43j8aW7B+qkm1y/SxQC9tBSagmK4XwGYHee4hRiWcli0lJkrEroocPNpc2y/NCVb
3+ul+PFr/je2VC7KnuJWJHBAntiat6Kg2sOGgLzF4Oj3dx8TtkGgoeRL/JQ28M2pn0z34MOwPe38
Ert+hfEfwMXJvrgvLoBJ8K5Mw8XP4OHfoACaZQqb+LI4Hxx2yqA/MwMV3J2EZGPYMIgWib6FmYy1
84T6znWBMM23O7xojYDj3AoRRBcsU2vuzhAK5BMAGIuOOiujjeSjHB9Ffji/k72uQV1DhhxfIIV7
kefWC+o3O5jmlvGu1DYJ/2jcGHM2TUm6kyD9L6IwsutQeD2DUX2+3SZphznBeNIrOGhpzv0CF/Ij
CPw0/q9nFgLlbipSiSXk+pq7JuvinMEZHoRW/6RsaU9ts9mS/zHMRSLs4MZ+7MwQFvpwa5817Vyf
r9pGif2U+RvDOFjArFV9a1/wR76LOuED2ws62ZsZubwzmO+CezK56GrKR/B1n8iQbmmnVojqlrnA
Vke7h8cSvBrISMqJZzhsyRqSX0cB+wdbAkHX01zg3ykpyanxjlY9h8eorV/wy+QogF5LhYBXcRhJ
WCp9Tre2j6m7tb3IUWrH2hho+Pk+jGpJiQnjO62XqunwKdacD6NajjCpd4BZJ/5lIRNSZekyhwTD
yk/VrdnZuaugELXa18UUhUqNjyygn3uY+7V32hV53v4so+rks331wHYni85vze4gXFAzFFPmmHrd
pkJjFQpw2xMsLsYWMnlQQYZZee86N7plIbEyXUGPmnRYtanPiBUFtzUgq7yPnm6sRg4jiwxuathf
lfqCTOi4+Ez0G2F4F8fLxFZWL4wYC8rTr8yDwhwtAzbjT2BVF4MJshTeYbyIoNzY6XyfauCiRJPQ
BsDHKOu+HVWyfk4hq1KZaSneUi5031jBNuEo+RBLgYCZBKsPxzuFkJbhPyzVFaRKdplvKGreRQYf
suxBZ2Vy45zQfHF90LgJLcmoUw+P3JqV5OrXX3moPWB3AWhWlaI7IQyEvLQraMlS/zXzMqyk5OqD
F20DMKNTedfkqSzZ4Q60lWlxR5P2PSgtxHObX8H6rdUAdqkSNPsLxsEDAlW5J3ZMwzt0AVnxaLLt
wQrBzTH86PGwNrJLBd5TV+ioWbDvKv/g0iXASgvBaW2frKveg1iKJRIYhV+5SHcJo0twM7QK0pHv
sM/OJMFYgMbTqHs1KPtMxEyU0zBEJMlnMnS7+ge0KH6tUImgNSX1E3dW8hXtUvSUq0H/garXwCTu
rcJA69mKx6+z0lTXAtkh+LauZ5hzRAkhht0slJNacqL3szySNorjSV9Z/nvwEA3/4uOACfS5o97l
857kxCJ0dWguPLDxMRG7N6EZzUl0OQsE56ldhIjzRWjFrzZqOLXJm+tVoS1s/ovueMGsOYqWcW7p
3TUb+ftG+oVcraMb047NgFZ+TRzHZE6fkToMltlhav+Dh06jYoOpvdBQhJ9PZii8aFgGhBZ+zqe3
+ptdra/Je5Ho+nuXfK29jjUhFldDEzBBW8CDIOiwpgqz6k67E31MxcNI8k+e0MuD+jSC1d5sUk1e
71NvEJ9fcKuNaW55OeW2gWCowe2LxmXJfR84VMgL9s43/etHjsSqmRGXBxTuvu5bxgKoM4MebrnO
UT0AW4vmzApcbpF6uIpSt3ZWXNz8HvYmgdPqo+nB/88vW575MKrE6uhfbNM1KZmW9Vkmr5lnXqku
C4uM9fb8KgPnJZp7934AzMVy0b5iFuQ/oQj8ZXuCVxLUHCwSRbFVEXv8Ez04HepUQsKjQ0qHq+Bx
KPT2ZxjArGGqOPf0fqUc45004uJQWvIL7pNu3XkH4Fs+JeOO+LOzorY/toAt6yhFe/gzRBG2IgZO
leAjQr06FEiLlEXzknF6k1jhoVTexFL2HY+HzHUIV25/rNOp0Z3sCOdjq7/xB+Yxrf5p/TftjoP4
UCebrwaTcGFnoaTrR5mYQXZdIWgyWNSFeAvM7bNQVSqVM2Q1ADdS04agHF0+otcQLfz2Bmy9M5eQ
HTnxfn0rW0QyhSk7QGP1Fc0g3ez2+Bw+EZsYxFiXxU9qQtrcPOmQQShRx9KqZcwc06GvgxQGnjdp
4QA5mJEqDTIz+fqUtbKy6avC+5gvFMtZ+1S6TBLonYuHH/AXZi8ixi+IuKyd//ACvSoGCm10QhjL
1pxAQKCo2OUCuFbuP5VjkFOrVME9mc5HxqG90BQpC94F4yJtYukyuMXUKppOGBvzF56/1WBSc2uY
X01Dh2VZ+lu2eA3YSC89JKeeAwf0O+Nku2f50piiGUPVApRSwIq4k3P4yEkO8o9sKsMhg43Tq8cM
O8D18dNseW78ljUTnnfGBpmNrgz57R+NcBXT3CDgqsUnpXYL+RsBTXokHyNlQyPMVuyObhnQhbar
ycoqmhvWfGeifuMkbTtKmL+9wC+ZtqtQPmtrmy20osKRrHC1Y5Q4qNwlo35eZ8tZH3SyrRMWtAHs
AFlxmxJuCjo0ClucKmovm0KySqNmNvV0LWqZMO/5DNs/U0o9E0E03Vpc3DaK7HtDIODSiMnV+S02
Rvi4MvNDyvn4RJAYzluH0Q98xGNmYJOKJQYI6yQ/JsI77pFPk5jNNWcd8BTQUOf2wBGk7HVK8epS
gKcnzcqBRs5325tGA99OpiTCbqzXEJCv/xAn0DNk98W9j+oeFW4HG8ey1+wFyHdDk9qGqjMDwPnv
yebl5uB6Y4AR0O8HrbmqPgL0eoFmC52hiBeMBXLGrVqNkLka2SmVWL4XaWiwHA8a26yHDNxhKMlv
YgXp21hTEUq2OLmzAwKXaEX4lr0GUbvPqTnj1dDCXEh8NLXfpmTI09NgEqCgN0I+KTkrpLpcA9ek
OzHuv2vjZJhDbEG2gHumTdUGwmi+OOxiXb1hAsZHj18zROFiNKRj/HyLOUCYwAfUyKdnkIj+mS+u
L+Dm+mhTAR/KFI0fG36IElS2+Z7uCJwh03F73ctCFXHaZkvUR4ubMS+1/A3w7HvdO22au1tqn0LV
3Uek4l/VSLKkMFKRvv6tWoFTb6Vslv1+aM9JZ1477eiRMHUBDLhhHHPLii/Pfe+ysWF9vMkg/mwe
FoeibTgYls7VCACgr8s/fsLrngmoQgRB4nxGR3AAKcvby2yO2bIi9seR172Uj44sEbBLFEO2+qGm
3GsG3Ng7ff/Vu2mas2WtcLvQCE0gEW+vljhQ21HOaUoDMxE+S8DUUL3WyL/U+wliV58fFVSncNTr
oRpyEQEWLqO4ARewZTEXwjkulkAvPnxZc6slxkCJJohrl9DK3xbjze4Iyqo3lqkY6ZCj9s2jqOvc
SbWo+Tij4yIVXzrVbtWb3qhsKiK6oDVbqlJqkJyRseDdMOmeix36RA7QY3kKm4J9VNyDhIyzM+zF
KbGAdCnuPmKprYmPDfYP8K9oV/Dl7s3bkJfdRDUFciKMbbE/EGHPvxrKEsA4r+5c1xvEEDg7bOWp
mwOj8Ry7K1E6hAL5+D+xchbUfpXti2VU/Tos1jufueEgJnBi3gVydbU3fQrmT+pwzbc+jTqHmASi
/hOt24tXV0gGvYxPC0QIzCZ196V4KZhoGBfLjtDdFh9Zq8voUIpJOEFSAdHherjTwOK6ntAGtOTd
iFrF25P5OtquVQFCozXhc1maLRM6DaTt0es7mo++jhS9LLqYP//x97NwB5JbnPEWIYflWnC0XILf
CbABoce2hDD2c/N84mzh+nNE2V1kASIkMvq23cLKtHbau+n2jyceOcWHqi9q1mL6bT60NhDhjfCT
qaDtROdTL7E5KIDgw9SnEzcuXssag3cmKVjZA3jFT8GwwUii3fNup5ovQya8YJ0D+f/LmaLW0/Qo
JW/tLthe2JFWkdxPZBuri6STWXb9yxpKJsrzvUBsYm2CFGk+qLoGH7oxRBWA2T5BC3yxMGjKNaiT
XhwMiH2yVxQ45p0zyxuTPxu/ft3ZX6Tvigs+M9kvutjB8t7/T2yZEjCWghx/Zd+g6VEqjYJROfN5
2nMeut4oD62VKoEbIwKrH0Em0TAsUQZQiIGcqDe06bLUJe02GFNIE//BaWioUZ/6dijnNR6wdArI
KXF1L/7C29Op9kWaqizfgRRQHQ/Y9vqoytHfzCRPcCnX8nuuuokteyqalw4aBFai9IsIcwGs/iko
O+4x/vAtRAA8I+odj/RF5i+9PgEFPLu+wIE3OEl9ic2BYjgb62p9TChzD3dLj3E1wuPaWwGPAaKA
xpzys54bdq/qp+MPmf99YAmGQIg04yTU0DEkQYXApYHgWsfPFfX5UXd77M2XG8SP0zapBNMrx0Ir
Nb5/P0Qc3haBqKxd9VJTdjw8mZ5Ltuyuoo4bcYvI+YDzCBkaNeyDwnKYeDPdat6i9mdclJ8C/Jz1
CClO+dlQyaaR/Du9KWdZjBs2OYBrgUQkukDGL/IRQ1u2qEPdmzppEwv6bFJx/XzRY3UEsc4l7rvW
A3VJuvyMJ4uHkyr/rMBIsZ2OLe4iPaltV9DOIsORoz8OUJLV0TFpqEonfOmO4Rjms5Sk2EGRzr2T
AOjmz9PuNSiCAz4QNjph69l6/Mr0XkbLQXPQJ1wAYHLMGPDWudKXBN4DS0QQRlemrNdzUx84Gloj
DcBw7YQybLY2ye4FA+CYphDxa6ZhGBLsmBtPTn1YFe9idpvkf1WJNfIdkfBEKAukqc0hELyXQLbD
E+EV4I+5gbheJmOYIUB+OpBV2iy7/44lwWLunBwBxFXTG//mkVKcmkVf18LU45v1ho9f6VJa+vVv
H1w072awjDEKlW9hN0qisQq8otA9D6COKE959UMzQg/1etsOejMNUvCQlAmZVZK3DdeGT0i29VEw
+BtPAY4rUi7zsqh1RiddAO+o1PrV0WG9oMsZmTTf9CQY2CMZcaO8RtIt6kF8wm+IWUWAYJ1e3bOq
7cO0yrJ0I4NyrdR1R5143cJBRc/07bikt3YQcsdZMl6wpm5Ztrrk8lwavLU0l1/v/55nqrw36v6F
5RU+VXQBgDfxcKznAM/YkSx7EqTqoAtYpbssCAYKQ1scLxYgBKvCkmb3bAnHJBjtgjL0PpqA83jq
Hiqjo62l/Vm9iBTe2ayUCdQCRLg6Gdwd+aq1wtsXr4gcmi12jwOh6pEM6JI0cJcUg6dAArqLp1XV
/IdtgsLuG0IXXMdEln0us3eKMffOVx1lAqi/xG85CQnrXtun3rq7ChbXqYunJBRDWEOySBFPZcEv
+7qA4dSjcSpv3tDlccBybTQ7HESQPYXbdzcIeOfRCtBKg31HrsabDk1mJz39i4rHz4IfeSfhqh2t
d5EhcNlWoG6EFtqXE8Haq1vofkKbVqefSNkVOd8VEWEEBhBiFrwKdsU9v0EMa4z5t/CRCzu1TZyI
om2WrP03YS1t0Um1aItok1YgTIYR94lb5/5zseyFC0i1ym2/57Cwu5dpChK3LY755R4hil1z14QD
89xd27j/UVVBJUzSQFRKx0P2DhmETEYoVo32qex3AJ7f6unUexqIm1KVwXq8yzt7IZOnk8fuWTeY
XAIwhHrGpn/993hEmATCtqWg0TneAKKR7sG6XrnvOwrzI9cKAMWXkwE1xgDMxtTvgr6YUtC6Qh+D
Wm48OrBKrfCfsU3mfiZKEYf1NcJ3yPtJdFn+ON1eheEdAxHxVEmN1ty/rHE5NUVilf7EQ8yMYP1F
QXs21yIA3fGVOj6HKIvuv6MqHV7Nn+PbdSnjPH7Yp4Vw+A6A05+bVtd6tDQyoPm1qbcSTpukNiu3
foyVKihglELxX9lLKgkqB4eRonGdtNDHr+UgTfR0WIqE9wUJZLsIF3sgZzi8KRCXZEr3nM2Q2mi3
9EZsEnm6GcDhErh1eXECGHO648fL25fpRABgqwhzFPZGSTqj+t9uWDifEexM9TM5ZDf++Vn8YoVF
p0aMDFdNvQ6I44yXGhUI2KEXOcSqSXko3XDl5yXaCcwWZo3pvBak1Dw9Baq4GVbHJccmzKGhzHbC
DrBy7XaYPW+z/CafSqUAPihuUpocQ369GRcx7O6cDXYJtcUbxg7iheIrMcUsYaBl/GWgC8WiyYyY
Jnm7ypbBZ9IUe5OfnSbWBnOLOV4Dq8qUSXGCcKgu5QQmZjX3gygqRKfyPy7V6HGZ3gEzQo+PLr/h
fMN15EEz1348WEOoLjiRLCo9m9jRNsgFpHqlPrM3gJ39xOz6T0itoEISEHWpkrXOVpkEtsCQkcZI
MVmlbpQQ59cWX0LYL/s0vQzBpiJwwBJPEwDcLIw8u5wGHU1b8R/Hx4K2JIn+/43ODLKHa94Q98Zk
19SAcUp8SXwaXpRN4iZOa/ayRuxaT7f+Inn0pciec08bsy8fnKDQo1fNHJRFzR4VMhykVymVquWA
lAJvLxl56KIhQgAxkQZp4A2qYFVZNatRa7v1oSYQrls51umgqkDV//et5/ynkuEzFRp3DIjXob4B
Pntrq4O9vVAk3CtcUjTcOA1ClCo9RGPT2YrF3IP9NS5r8IWWwyi03LDwE82DXOjMOXrPMfrS8gEF
5bOCpI1xA+5hwnIHFmFoYXLrtsGuIuHeBpBgP7JI9lXp1nMOCVGApKINvHohUTTi79vf7hrURkvV
cFT2tMotG7Y+TfLlchX78C0JX4gqLZ/3veiF3TWCY9JELtDZgadGpsYQvQAEHVD8n8tJ2+3C+kKp
AXBPmSmMUhQek5fKiNIEeWpEz2BcxGUmspUTW6hTvrI8Dh6lGeev1B21Q0NVKILFWCXCjm80XpT3
wBO+8h7/hD2o/4FiJBE9pXanRLmZteRiPjWtJjpE3YU1MYm4HMsN+QXnLeMbBpL9vjPEEaKHbutw
PBSRIQO5iC/wx51op9pCtBLfowA/1/KXfIHMEFnYqkOS+hz7zTbfzKpap9QisYlmDuNlVRRl5uhs
YXB8LisZAqQM+Z7Z+YZ2fWJEqvRH9BpxqbGCzhmg8fFtbGLY8AsfFYFNEhXk6MGs2upZxr+W/tfP
qO/2aNnj1KfuRmO5EDJ48c+iyXz8J7hNAzu/19R5zF/ldt3IrkTWzLQ70pBQ12QfTmU3wLPzcSPv
3/rFIT+jAcMj3+9vHtOvgi1GYY0dd0Qwam38uXTl5C3GzH3T+FRjKkuddb09Ta+Irk/eIXtK45e2
tfhn/DEQryhE5zPuZzRFHYVtksxn8lg4F8juJaDrva58PcMN9//lXE1nvm5xuEqLN+gGSbWfUPdi
dtUR8s1LcrcuvYJzSgmHlhw4qZlzcnBWaeUURm87U9Qd4mynwZQD5YPhmLgegK2xA8yNz5SmjIpm
CCh9il4bOutolVyvWfZdUj/8beRB9Yiouu0QY5tIcGzBOEVrUB7b3xnW1Em3akJoNXczSP/uUPRn
SDjY+pwV4ONDggxxDhKAw8szHYsE4VfZEqUUmbMfvDLkZraQFkZgW+nP/k3A+x+YuWMJTi9gH/sa
5CSGoTl9XaHfguVffwR36n9z4AUw48+O/Y21mEXL8zEZ24kBSnZWm9K9kFMQtQFszftJhu/ziR2Y
sfbO/j9vBkGWd1bTuZjqxm2d8VgAarqsGZyeu4Qy3uCC1HRQt/Z9HmnVlLDEdKmIpOSXwzSsUcaa
qZ6/H1PUE0n1/bJFbwBZoW4iSE5WZaUGp09SZ3qr5VarPwY9K+obwvWVM/gu3uvKMfVEV9BDjKtx
GmsU8Fx6DSBkB707Ia/4RFE3lrrZFJPxYxdTXN+u4gEFgnf25jQVd29ly3UAXEg2/U6dxzwlOPnG
unSUuc2F2+cmzrew3Gufsrk5voGiRR3v7GZf8qb6qUL07C50Jh8EnB0uuWhaF7yNpBHtcoVXhQdk
WjYvwwvoNT+JHRKCKIU11oq2ZFac0+LQkkpSvr81siWvftbXDHynJQOKMF02ajxXpDS6/NX64f6s
eldpB9K/aHw6oA8aIvaJAgFF2MESDB0SDIqD8FgMxzGXMVEA+JxlXX3bh6x1MHlKLfM1+md4bN4f
ELn84fhZhtbf/I4v3ui21qocz2F8pfobP9tdZBaan5Hcu2Z1Rk1AIBk47FDq9Bzr5KONnzV72+Ea
tpJjy4+/tpHb/+nMxKj11pSDDgpHE/VR2z9fQvgDttB1sVxJwdBui9jiABuiKh+psXUmwU6Q21J7
4XIoi3EykOnxtMI8kSZoY7pjLl0nbJlRJYM1jx1tRk3kLFAyjExMIzV8pi1NBPJ42Vc+6wMPVXth
j3zvFTq3p8Te5zKpD0zvM+pHDhHYFL6PXQ7iazFushHs55ze+lmFgW72RmaSgoe+fC/jWaoBAbxM
evpRYwpLsu1QmGiCMC9DaMVrMp1bmTXbBPFtBBFytbPvLn0bfPj/FQBFe5/h/MnhBxvAub8dOpFo
s4sqMLutOVbEp0jMIY62Lkbdc3W6kXGe6qI89g0gblFL5pHm4ycy07piZTr/xuBeUjWL5/sDTSwn
QqPMhyoK9170lA0vXwCwVw+A6OMK2An93Ab9xGbljh9ajQzjYpqFLtH8NMaVICzhuxC2gWMnQYaV
f5eHJMz3AkzPIOidcEUF29VG+/xlchCFmeMux1t1s50mJHbGQek8RKsvC4+p6GvpCIPiGSZxOk4o
6VD3K3uM0XHlQmUQg42Q2K7cgp9LuYgFE2mDMVvIGajiYowKys+N5piOUsiBiHbBzJlDlqIqXWjZ
VXKS/90mADRaKqrJ4dh+ov9TCuD7V1jQW35Jfd5wdHE5s1Epl/wSnRwc2EMiAEQro+xk5ub58ly+
htFK+PQa7g4Lc0s7YGHCgs+rmG1GRq1cmRYSQlWcMYw4jCqqVamd8f2LFHGWICKoxzWwxCQTpaqH
ETQuCM9T4a5mACScKsVq+0hczDkKKacQ59Pfd50KyRuVDv8Tppoao7QFxaMW+r6fAMtnPuRkn77+
qbtHMk94rH4y7tHyNN/oGUtigoqdtKz8OW70bftDbxcWMDGcAnfU+hva7t/ooXsu9R+TgJs4ANb/
UnrLx4Oydhgu7I2yTGs1dM9ZEKQ2pVvZWl59UxyB4lT+p5KQX7IUG75tMoxNIp/qukeKUaVlS6tX
pV7xKUGHX3jZjc3YOMh/hwzt6Yh/W5RQDcnvP+NSzeuUIu+NpLMtLDWS0bBKujt5uvJaoI032FC2
gO6oPomZRu6DES6gKEzYzuX7eIOp5H49KCw9GtnMNdCdDA6GFB4WBmJBeAW83+w77IsdRBXz90t3
TfCX81IUcc6sB8fak8HmuI2tE/PTfYD49mxC1XoWg8x5cT4eXtRR7k6xacFy5VNzJLcHqxDSdzvK
Rs2M+kR1MuiUhhpsejuhrGZGPtnDJXmwunEi3xrlB21VwzOFujxAWhvcriA+XTJYMvxrYDUFvufK
8GWSbYHl3LTtIesWDKqfkTokDkuOIjI7snxDqAgRYCQL1ldjRzZ6DH9LsOjUhMi2QR77+PXW+tnC
UUfNAKSLzF4Bdcbexb6pJKA65Pd1M8iOP2EqqLR6Av1glkVJmyhenu7qNGjxctZZcO0BKmprO6IA
QpKFtLaPFaz3Cwj6GIA0kOaxws+JMOPpEDh2N+9+CEAQL1rjlg1kj5EhYMTNMqB+aWsidnUmEQw8
bdQFc0hYKHj54lNAhIScvrWyfQYjcpm11L2D1k2F/x6MCL9ZWfXGPqFxgz/fjzKMjFaMe/D4RUdO
3cthqlPuel41otvRbWljFJF7I88JpTzP1o2r4Mus14ECZ4AjgnY1bGKi7NWzZovNMC+OKujxNptB
QjsA/xLrpkjHctGyTtKwfiGIqZ4W85yMRqWPsmB8orWkJvtb64JAYTJohVAfBQnHwSjr6DpQMwns
KSsVCTq/wFDThpNiQb9kLRr9LA9TtQthsPUrtDpaaorSUPyFm6YlzzGD4mAvJYErRxsJppHnmmhj
rQQa867RVFS8nXSaRkcN6uq/3rz6rBM3Tck4HGCK6zM6b4CETUslQqwrGi/f2pL2f3padcxDZzhD
BfNMe3S5ngB0yWfI74TA5P1VDUVVNBkVBse513XshIBOk2bK8zwU9+wE6qm5BkSb6PYosf8WvMv8
DlA887tHWjBiazhpN6LnaWsDCJagjlQ492qZeNXUpVL19FSPfmq5gkqe6xPpDVmE/KNhoLZjR6QY
Im5tPRhrwPEvhqwamXFrdDsOViPe4djpeFP72BRtaufylf5U+lyrXEHFW6nFHR25FghMArWm0e0L
bnpQ21yjFCMDw1CsGtAzeyAs7dijNvnfJTjuaMImHPBVZWBcPfx8B1plWd/8JIFwGwL+eKUzlEdx
pcEBxPKgCJBLzQp42vGtViJqeKX3jripUaV+FDpeBFedgwxEOK15sbRD4CtVAl8MSBG23MJe7wE7
KEq0wNTtFwRc+t0TCgv1Fn0QO0/Rc2+SbgwHa2WLzQANYo58nC8ea/269IJKDhiyN4Ya+RrVaPN1
jZkI9gSsfTvJuFyvAdyu3Sd3Oj8wZ9QeXwdJ9kXnTJ0tHubE29yvcxru76Qnm9yaMfWUARzy0AaZ
fDRmABDtl8rbJyyEgm/Ch/s6r1w9aGm8xuUAi0GbPQbXKJo3qJ9wcDfkctJHQr4MRvcAa248jiwo
ZAQHlNNWUD5k4qasw11GO7aKUuFtQEH7s4JEgdUPA76donXREQsUDs+/VW4TM6CrvtrQjeZo5yXd
yApiZfUjAKSDJXgelIhA3/1h+8zGVOTFQg35erfbTFWq88DjNDNICkB7NTtFSiNnTHGspn/Pp1K2
hKihsJnjmZ/JYG7OX9QcYCJm/hg8r5WkCbP6AkfrYq/sTirJMRKn2d67YSaITza2UMVQV8/0JrhS
B3XWSTi3jFtyLEV3X+B7OQdUC81HwhtLIupA4D29va4yOGFNKMQaUAXpcb7cigoeddhSn7zRq+Y+
dE3T7H52dY/3nC6OobWI5+TlbFN4EZ4W0SX+DxtHzjoDffPeesPL2qTvuwMoe5XkwHwjgWi5cmgt
gfufrnTVaV5bv3Mfz0xUkHhWKhRHbXHTjGm4zMXPGfWoneNld/bdX7A2wC1hRPHewNRQQj0O1Dm2
7AFhIhONlDgEaCJQeeMrWpwOkR4fmlK7xQ25zJ83q2roQRSCG2x1iHCkTb1bTGunnBlXum+Gz6+l
oCVwQb6DiRK4Teq2r0uMrtBMDGDH40qTZfPshNpLX9DYpIHZO1w6N4Wf4fNF0wBv1MNJMb8c1axV
pxKEEqSOb+iS5jYMeerWr5Pbr/zmLaBjifO2OGAWcpCen7dd/MzdQlhxwMd/XCvGHeQMxf/WCDci
+F2wGKo65eNb0JHRXEB7ZT0lNXL1e7brx2PmEeYLn9gw91YVYn6/JcL9KK8gGkdWucydAYrP7YiY
/bij/1Xbs6J5tMyXwXIYqbF83hHWGnt//8QbjVOQ5ZQhHNKhQBbzn2OKCuo2T2ic7dyIuFPJdtGp
5rCs1XpguPUz6Px5qSnXm6wGoiVJCH4HBULjYv35wjLaXXYasFiOeX2/VCM64682m2KOwpTYvH2v
i1RnzgGVYTwghLX6WF1stH3WVkmHOlXJ7dP+z7TjrWRSemNc8uErI6BQvxP4Ouk2Y8tS92IRfWjC
2yE/PiUYyHULU4Iq/PNss18YuPTrkZPS2xNi6nNpP0LDA/QgZxpiYvU7Q9X5yhkiRJ0IRv2ooCyn
GbehnvcCD4rh0Pv5ZtPSQib+k8mQRPSyfIONbe9+j8ShQx9iVbX+xXRr4ndpj+GCUlCntXazZBA+
kXYIynolNeOweV7EWN3XpYEM1ldY2LReHBIIyPwLWWUkDT3ROqAQybuWdNg+N+BoBMDVCQ/9UiwM
weESlHnV8xg0rXd0/rpCAsNxTP8rB5P0drxT9gPSd+pRL09OvBGFgm+hy/ycz1cgGX5WVhVOej0+
PjvyyVe43MOAHL6BBOVmdf0dkm3nFCx/SlWRErDtCCeJmxfTmfDXsU5ME4rapx5ZhwKmPGadCi4r
NB+ulTXENaXaYVh+6VKIyOiUP3ZWb/wGM5MkushEOEntIZeerbuxK+Ap91gmiHw1/foaHVOzqci6
p8VaBshKgSTftZ9EVc437QM0cZFy80bkswAhteglZyzT3bpaJgelgCOou90vE3V4TrqaaOJlSWst
Y7hZtFSJQ/SulksNdn8iUsih4iBAbw6Dic8WzzkfrWeDVqCpQFPeJuozT1huhpRER/Na0BynKNmW
xQPoJ+pVmCwSZJt9B/yrPfXo4Ka76dsILUrf5uidaHTEy0wulAl46aYrOvH8ZoaT0iLSoU7bORyL
O6F+YifULrnfUYXyzXLq26/o7byddZo1B70+9p74xObCcrpHgKiVR0hqY/qHEjerMp9UU7Xd9ysf
9awoQx/QDRob4mO63YO9NSk0VpV7pjMbe85Z+PCdBW/pWkWYCP07PMGgKkl5Yzm1A45jug+y6+lC
oFSrKriceErDFeGPG+b09AN+w+Roq9bqqIAybSdUEA7t1kOFLrVYD5u6oms3ZgrrUu2I96IVng5l
MxotEsDJhUDPR1/g7ShUBOPxDrANgZAgIX8/VKR7gbnHWbbJ47JSz0NN0XdMNcEu75tC57RlELcE
p74O27mdf7Bdj+5GfpbbQcu8xli3zSCeUb7N0qFMOcysV4JtXKuNSxOWx4uxOYZsYyVtuHkT6Ph0
SwnqwZdmsrpClK5Hex/kdvE40AqucLutIDBYvvTFv5mpUDH/Gr3gK2yWt3LmhAbBut5mXfh6x8ft
PEBd/PETXcyB3VTTwWD0bvMNBLbYC+sfEtHcGLyolznMd8a2xqFKzGlWU6X1vcuACOqSO9jUko18
DveejP3FivHaNBaLtQmbXQwt9c/Pmq9U/iBedMF+nvXSAceeNUKJwOGxyJMq2U77rEU7ncmQICO6
N5TyErfPC/fszscvJlz++SbJ/pQ16TsDpyTLxTr3i50adKGLPV8EADZmg53CZoZckj7rXRL02Ine
d9Oc82TjFkkvkDP+VI9/00Vhjll9ehk5iDZucDWJW44wlWlhK2af1a+38gnBB+DfQtPH7aunQwtN
TXfNKsH8qalmrmGAeh5E2EL7fglDIsNAUypG/uyjXoGqYgk8SznumPr3fHkPaIzjuEb3HN2zA1TB
OWl8X2lI1On7naWn/kUMzayUH1pVQZAx0cYLLfRHhBRSYOCZ0acm8zlmvXoNmyu8faLj2dvfrXFd
QpPwWJZ1PwhIrDZvJ0sysbJMVkne3sS0PkR3HlXv9ngxj9+m5k6/6CPR4r03zWhfspohsvA8p4Oe
QqN+ag8b41y0AKyVdr3RKJ2HB9EJ5boCjYCL/muo2d9tw3ho84p/1KiUM3dcXiHBRhR6hyEEB75N
ybIOhn1715r6WaKdXZLZ1whhQyGpPD7EBEADQJUWOLvA8bG0E1sgaEJTe7trqGcvlvEnXzN1xBcH
sNmrzID1Zdk7GGQ8A4fbYlHoUO3BLSgTgIntXJ9RfpoRspb3KX+3UNP3tu8PyTInJoHjOXy2CJKQ
nLmL/Pldwd6PEC6WSZy0t4ezrlXnT5ZzBL0smnBdI0hI2LzLLkpU5Eaynq1U4Z1EsLfS1TobvwXL
KgCXyh7Q2MZh1hfQkvzoRylYXhK6H/aoXkPAFIQTxpOmGcKbhbabAomZDRPMVeSnQ+w+VcBTK3+n
8z+w7bs2f4DlpsnESPeRZG6h41jbhOZg/XkLVriQwLXgDmc/m1qa38QeVwMpOs+zRJpQVlm4BJ9z
rXmGB7yPbkgbaIkmg1r979nQj2NJIDHedx7XhQpfPZU587hyEhQbeGfdUa6rmc5QNKB0YwoFHpOC
aA6e2FTja5wJjxFv8i/jbIOVmgzU5Z5hKiu4bmlNychmvnIK9f2vb9uYTEHkX/yfsZ2JXGKJjNjZ
MMBRcQ85wxDeHegboq5M2tCVWRWOjZcn3cmDZalzU6Bs+rsbdKBkzji4BpWOISlFtwHSyP77k3LY
H3GUxNdoVHXKkI46Gx6k1+omO5Dy0g4iHu8WO2VyLcVueUhF68aWUB0rDGmSexpwovtMWPg+NPfL
e5LnbggvFXsjPZ6AtZLVeM01loyT1LkdGP6e/urqAjAtzyaJJ30qMQXp6DqJnUAhtdE5RRTYfHyU
wLgPzTJJfo6SZQr1A7SYBbf3YoPJY0X1wuTgPiCecVt7c3SewW7uc6ge9QJ3tn9T+psIXXEjIyed
bq4vLULQudVS892scFCFIlXhVOhxfPOtckrwTlU92WHN95ZoXsGbq+Ew/4Amr57IHlP6inbid+9v
XVTjXXfBL/dNd1f03iKPzY/YGkEbhEE4Amq2mKEo/9USDSItuawGgv4kMpQWwEQDi5HHiyOPTlL6
a8iOsOm6S50kJjpxt3CoGsVNqDS6o8bu/ZpICIqpMw6XaN0iEB9duVKjxIIY4vPilmPgwY1KTv0e
Oimb/AtFR3De2J6LRWGYEX0mlwR3hnNAt4OtwBU1rkQWeJvMSo5IySVV/5ji8+G3kuO6q9l5vEaw
H5iWVP7MZAb7c9QeXJafXIZEkXBbJYKwg+49p+AV3JSlyD7MDTHaqVNeaf4kMccUFACczVPSekqx
xcqAE+V/fdEWNeJ2njXahwYGoHZn/cmIuBZmp2dp9zA25nf8xcqc8AHYVPjDLDZpyStUPlRUiC7J
wyuG9I+86kmO4doeE4Q5MnLNQ8imtzBxqv6ga2LZrXbn1VzyAr9NslUYPKC1D4KSfBVq0Q0oa3Mu
l+7k6OknNyjD49jvMMSNVzM1DUJDF6lGNldFSLl3si/wLXhenNyu/+BvKHj3hj9SyIMPNcYUc5L3
0kTt19luJejbY+PaMSZlcyo7/gfa6hJWIeiJ4HxWUmMnEJ7d9X4vKhYHTmKoIE8984g7c+Zfk/jv
awhdSeBPVGHQLBQbRw2Eq78Bf1EBVi5l3Mi/nGGC0HkbAisNZfwrNItBw6bnmoxQz4tEEMbH63eX
s54p9ZqGnJCGMy5L9WU5hol2FZkCjm17WwqOIP7z788sRzbN2Q7DGqTI6x7tevluONSEAW648tl3
YzhsbAFfDESfCRLpXcz4TbsfLVQkM1eu0xL+PEB7nO2lwp21b3C5OEhCuyqDObRRvLfRO2o31+Nq
gzar02pjZ8HqKMTqeMry/O1sMiXRKaEDEKQgUtvhfXfjCKegRNbam0PO/b0y3N6lOhCLUnHJ4MmO
iyTF9aZE3cM3WLHQ4LrXrHKASF0pxEeU6+6aHiUBfPrnahLaabJrLgUq6hhGHSXW8DZrrCZffPV6
o4JlHqYtdqN9MjceMxV/ZusPDMSf31VkG1lqUttfZwZDRf24Aqt9BCXTV61PnMVUSTqwqMxjUDRe
oPEcSA+edFRXMv0PZCB+HWqIZzELp3cfI0Pn5FZH3NxVuXmsy1XLCfH3poBszKFj0mp6GWEw+y0k
tJCFDU1dmAeoa1GtD66ZJjLnQWv0VKJOVkyATKQbwnFUdu5q9EeTIhLfqIZcnGF31kXoTE5CSQZC
WWCTbZv1ypMN2x17UG6H9HcpcazqmzooLa7TWz4bI00mvjFov05KPhnuV8HUH0eamgxiRm2AmA2z
Ww3q3xq8g2fU9LFWl+4yWyc81JlCXwmKJaPBjPsX438o+H/KkkzcKYyHXcchWKNctwavDMIWHQdt
hQBqDxZpufIxSgTwt8UHXcA2z1X0zZXVrqkyw412XUmU8jfqpJQ2Pn/Pmalri7mEqRJFMabdfDRf
h7spmYjuOQH1yBSHDbCZJ7gcDTUxktCDGR5pHl52sclSxxi2FaVErrq/vi+r/5rA6BTeJkvKC9aP
XgHXFzBwOkUSjuVB3kZsJyTNncH840kbB8DpnTctUDF4t0tApohcN3kkAGJNckk3hf5xdhuA0cR+
BK5MJ9GdCJGBiDMuQmzcW7xaH76ii1mEAlrXWpKym4u2VPqgtfN51jkr0+F5//VU86ZuIy25rRo4
xRO52ibjOnP9b3m7ng/Bq90D9J+7TSV0rehcB4OrqVOSpPJmi1J3V5SRPmaTOyA7XmZbXzkk15zG
oU43mbogXFXVZ7EQlHy0mHK7hQU3vniw1/vnfrbynTyNpGknvuWie4Pj+cVrgqQLRIcrQX5dPmh1
hCsQ8XCvNT9kRgWkehuHDmQqPgSjIOHH0NiIVZ2yLN9CgY5xt3Kemn7tMeW9wb802Vt+KFw2bhT2
OfAfGoo6+L0alxRdMCPe9d1EYLQGJ7LjI8jGzE/hRJxhhNtGh1Sp3Y+WR/IvekkuZofS27AQcXtF
Kngk/KDyGU0fcyMhqN8ZfZZ2m2B2oQJq5BEH2HlAxBQl63+9DK9+zsVJA73A3ORaGPYw28+nCysq
fLijqPlGOjeXv/mbztCKU+7TRBv+etq/IpQ19Xrx7AsXkHM8/Knl+SLvPIKZQHJ+nw1odms2t/jr
xU1jjtzmMil55yRXI56PJDem2Tn+F5+ZuJvkOhV+8pu9PHTSXoMipr0HISzxIGf2D7WmUGBTq7gX
DzGnu/efpe6zSjXE0sevStQMdwOTUh9d4KkPlT4M15vDc2eb/duwuwZEzqmAiB7gsKG+ovbx5YPq
BM1hkHc05HVzseWMBydD8CGpcAeEDKuyUx/WBLFun2Ai1emd8vlUbbeCMUq24KsMEYigOQ+31KQ4
3QybYi4UxxIJ8yiXS9GczoyX0HhH32V8h6p3vjOzEkob8nribz4gLKSCxYclaMT2wVBIPFNrzGAM
aGs1rky1L7gmtEFpmmH0guOw0y9wn6Y0WAJo6WxfbuXGeOUlaIaRuyzdN8R9AfNg9IOmcfleY1yI
BP0/iZHLMLBVY+kwYXk1Tz3nZYw10AyvkNTPvjPSs/WYzmDRevz9IlMzyBhUhAhrs0s23Sf+2hSE
HmRCARikcRlUXRByS27aTk/2jCQAxvM3ChcWHWbuhiNpWHKhmhpdMseVlBvJ1Reo9TmjXc97jA9y
wYhKBv3wBMrttXmw+v9UhUQLS0wnL+LyekOiYFv7NAdTsqOlRpBLaU9ifGawwbi5JXDY7HrZ5wTh
3Rdif3qAbmsdWxwjHNT7SLXENvZsnf+SzEqc5v27k6wj485ZvF892KNWg1vp7jntw86CyYDPrNAt
feCsHxOV3q9BzjROpOeGFdaxEp4IQuqMdv0Lklmmi94pLWFeK87OwYFapt+w9XRkx+VfacZQYAtM
NNsJ3eVlOvpAZgP3OC+4hYqQqMAcv+Gzy+cD64fgaMGDqXa5l4DVm3Ua9wUVgXthrKLrdVhu6AKM
8vt6IltqIxGGP1zdyVhduLw6qkev3mvXcgKinCaKoieot/kWQShTz6dYnO+ZLzQMZ3sxw5JzkwBd
SpZz8d6nepDvvAI5hfcLzkXNTc13VL/+qYiYw2QN3gpSXq5FJTqucNiSWZ0mNJVNairXgBekkx7E
yf4nLlrmpO7ls4gUoBPK5zy1m41dQSYkDOonXv5XqulSMqjRLs13t7lfSa6AxjPmSlu0esKXCLGN
VyHEvgkDzIyaarXfF/hLAUxeCoLxoCfFuMX/GWUcc/cqyJpAC2dR0/IntRHJmnrgHjtrj2LqMqi5
Q2KuQQ+APZlAoD8PBt7GBzdTdxHOPhltNdqNH+T2xBWJ2NvVN3QvooKmGCXTqvPe0SLptdm5ZHSS
OonhfFV6Y1RFW5+f5JXi78DFOGfZ2p1f9XSxviXm1zmPBlPAVYuryw+mcXTd7d6krdzfPEKwLO16
oyx/c5aaSHA3wlTVvpsZM3Z+EfJsWQSbdOYwlHUUt3DbmCV4fX4kYmOc7j67Ks3T1XpQEw/lN179
G6ex7+m81Eek/A57eZWvMx1ASrAvaWFq4vlk1FvMK8naQUj6zMyP1Ail5TsmWzbIETsDmRRWQXuW
nPBp1AiHQD8pKNugJqtlWl/pcZUYH/52DZP/4vBlVAwqu79ZinfL/ND7d5+LV6i0V1+bA5bCC4qf
QadXwulvTZNh+pORYJgvZilqJcaBxkJ27uecP+vNBPoPif201tjdb7TRPKgZJCX27IBfi7AfTlCi
nWhF/KZpINvm3bI9txSJgHdJMPSGkuVoAXrMYKcmRLac+PkVy1CEzGD8sEX0quLY9n/pI1Nykw/z
0I6wQIcuQvURSAA8RpS3+j+j1qASjFw/QwZKSLhA4zlFwaGOU1FPMLBiQKhq0nZ7hlNA9XBk+iAe
hblS/hfEf/VJA2MnatFbnEqRVxhjgWbW9Tznqk5YNQkDu4QC/35hHUNE8OS8p1qKB+uKFT0XifSy
diJ83y4aLUebu98BWmLTQ3guNmNQpwVAMgKxAXVV4Q1D2Z7XGqKFtrEaD/Pqvo6KQRO9JRCDJHuQ
Vh8Zmps/T/vbjdA1/pL/26uVUfGP8LimYeyaZ63n89jtQzpT4rqfO0mbthUebWiczHNZwQcul0B+
fUbwr03hhk/SsSXtJ181K9Z384JKPiYTsFgwQcfpdY8oTTEOxzvW4hI0+exWzeN5HqQ3UFvIeqfg
BORhnWOkAw3b+PxKAKxowqoOSFnwE/AR0Rl+S1fUUkUuRGjgxfukLTZ4q5ORkDHK+4TeFrYXoY0A
XsMK9cQldCZd4QWtSvZh061tEHrWcdCKPD0+wKa/wU7Y4Tme8JF8BNl9XbPx5wXLm0DP2HFA5k4F
mIUR18rTLoPMD0xk54ErqlZl95qsD1GSEeLS3fDEMBcDwEy6H6w47Svb6sf4NIvgxzzQlyR75ehu
m0CoOwiFCABxfFrPa4BZZYfWuLjgthV9R8L1VcSPqGxzeNbWhHnrIelpNcGL5pl/dftlUhe/1LHv
Rzcax9F7Fdwonzr0Ys/LNpSACmU4P2rqR24ouqYsfVGKq767Gq9qS02pP6WpdId3Q/EfZW73l/lq
d6h9xG8ypuEgSPEy1pRtJcRQQK0Swb9d01lvWEejARCHG/GS7G39dp5mvm7VsDzFy1lyabIvzbfa
4+J0r3m1g3zESXeK/WJ+Phc+yMliMkLTOyA+0xzz1BsBgYjzYpMaq6V2wfVwGK/yza316ZXmFo6b
PnCdJnucqICFW0V9w9pEDdH9XMoCF7ZpIp02Wljs7jU+Z6C1e3GVkGaISy6Ws0hJN3OiyomoE8DN
HlwA/uVDEHZlxpOQ3NmEuZDdBRkhenXF4+STzLCCalbUXF5dP4BPWMteEDAc7BZZBcheaRx5jLDh
V9x1qdfCEgAtcdp69NwIOvkpfkRGn0IXBDL9rxTYCoz+A9DLPVwvTPG+oBDHrBgs4zyEm1jsS/B6
DAqlA0XKOcHnItREZSL1FQ68PwFd/mJo1iIhHk87CMIdmgfecLELihXMRIeHs25WpRPQ5k3Y+MAT
oPGlnkSmMCvOFpTUicZYjL589k+rAKzI45RZwe6k0bV4DFqeyIWvGUocTEXSf0z4xZYWes6xpJQW
Edlh8Ks6LV3mfIiwEMYUTCXuVVS8yHhYD//huBMejb2Wrj5ohLApF3eYko2ATleZugfWPIXRwU11
dJJqBwTbKvsXnaA0Di3a92vZVlms2Kf1NcN8Ob8r0Tr9pHTWZiivMR5oFQAZ7JU1GqCVWJp0x5Uo
/ren9E6hjVJOa9Oh4nYDJkhQz6LyqutI4zov9sh2EECNSQhXhe46dFh/qiUNnoNs9GK/LmCVQWvR
MIa2nMpjM+DlvOQ0OCnRMMMTpE1X1T86yuVNwCEoQqqkm4n5EYQmACwnaGko12Qag+ANIj/Vyu4q
Wo/sf3tS35kxUCaT7bEkfTHtVGL2n+nfQTznxHl1PDaaylGGZvcppFon8NgG434iX7SPL7gyScqH
/eophp5s5gGcOjJEWwGdj2FJjECvhj0kSZ+jM+VaeO8Kl7Wb95E1u77XJcTcrWb/PqjrtHKQ68xA
PtdmGjhNap03r/Y1lTlf+aGm3vUPWJr1YucpyinGAmy9Hdt1zr2CfNPwk3P7eDquUptnn+AlAmKv
UtejEGElTonF4+6nHJXvgBmnecTQvjUO0sjCGabID4sWa7suoq0cv5u1veZEPs6HD18mgBAL55/s
gFO7tO4QdMDBApHYgzqlcKNK8K9Mvu7dA5sbNwm6TskwzpDixfI5rP066u5uVm6NuDoYo3YtSgT3
DFI4K460hjw0W+y++Xx96ElK+jUJv7DhuW3QIzbtJCpocSnDf9tVpHZYhlnYpZFV9+bc1j7YCBLm
9KQOEYg4U2pFG2GK0G/PEDWVLUc4tlF5fFOF97M6S+X8o+qkuO9ROC53NGKVx1jGkgH1oCqTcgtm
Tk26sJxH4RLD6F3H3z6Qk3ukU8ec8YL9kCoZBEnpV2Ef/pibrs++zdC+WgF6VXmVV/E95gL8NHfK
PMYEpZWBkIs/cBv70BCO09l6k0KPvVvs36cKqd3l82KdcCVhioELYOG6ayAcjKeUz/6nCrUbsIHv
fOF2KDUzhmqknwmRq6ZoF+WHcM3v8DShoQZjVWeJgELDqcmMqiRoDde/Hpk0dhRo8S2T4gXiF4sF
yIswoLYcQlvZlxmPioHhlUmalIA2ruzbFDTVG86Q7HQSmHjFNiRXKETuEkQWI0l+ZSpu5QNddN0q
W5tL+hrRY94f2uiXXZOgGMxVhSwwDJMHmWbrZhpSQWGwniMXF1NFs0DU0sYKGg635+wKIwWraOrt
pcGnGmKWigb16obYKLq7hexPnmsaDdR+EyUeUPN0TAWlDf1HeMgqkmRPb0+u6dGHzmeyw0bkLFRd
BmALmYrK8S/KHMWIevPWf/JU0MORS8fnOgDe/cLSWp56EIx2vIZg/SeZSrqmvE0jHZWt10KGx2/l
PqO/VETR4U861TzUGOMBXlJvaOxNtXDdaCv5z0ccAWiI7ABfsrlb0kY1VPCCn2637lZ2FD/B32Yl
wdIUy/w0htou+TwBPNNcTEoQlMGY+NzXl1yk7lX9DMSHzUSi66DyXAZl+G9n2MXtzjb0ZxPE5ECW
pS+CJZT71OEbxReqRsWrNM9bSLdP8BJzWEmWNwn6hcBxzJvuOcEO6t/PRIU+9tnOX9Z8kN0/s3c+
TzpwmzgyF6/AwntFOBL0EyZdAvMLCU8Fyg5KE1oQbtOFWtu1G9IY2tO8G99VZRi9ASrTU4J1EVYh
flZLpwdwMbZi5B3yP8U3wXqmmPrmJpU9XhpzIDviw3Dxp4wYdRBPEezswZxoanMxn2Qz/9ifdgph
bV4i80enJXuquOK6j7ESYDPIR6jKcAD2+XxhyEJoPJe6TDySlLWasQDX+GqfEF7zkKI8iSezJOnN
EDh8llNT47SyWUx9Cf/olgdDC7ILy4mGAWuEmPCrhHNGC4ddFEEZgBDrl22ZbaLp5rGhyGiJCD5p
eNpubVJY3qvWRAOZTH27rM/yiJAiXLFxv5Cq6UZQr/CJD099PYGg8T+Fpu1vS7gHsPk2empEQsD0
JT32bmRfbf2Va+BXRCU/dk2F26JvHdusMbc9JReKioGlUpISpQGa4O7ALOF1gXfiT1RLpYGsWLBY
v5XTm2+tYpQR8NtZVsj4fz4NF/bVbP5gXODBYhV3j2yCVRbyLWQdCMP/7036NE2WbJjMM9YUFyxi
MlcNCsdZVYrmQcm940b/EeeXs3Nk0v3W8kYoj0q1j4oxrPsReGYcfwPZUQG+DctUf1mGXYfyHIC4
2CFrSBqrhUs/A/8j7rUg7U11SVEVMkWLYAkpYa7vyD/nGViG5Dnl/lpGzwjwqTdDcv5z70TSQ79N
z48qdXXMPXWKoGhqgTisRBWsAAI7j2roBANcbohkX6/smVc/1oeqIPg4SWP+nsaBdznKnvKh42xR
YJn7IsREnpPHA13RHLOwoF1cZ3Qth3sl373po1Aj7hIOAlVEL1XtsKpc52CAyQWba7bt0/eMVmhn
S1EQedDq2C0R4nPyW8IAs4+SUHqkAQc8gCOOHqCeSKJscWGzxRjZ23GA8m+xDaQqruoeh6dXBeGn
ZLjHEx3/rwYFH+Yv5bClxIw8DvtlFmF9silVilMqrpvwc7ndSp6osdKoTDw38GW2QDMZWJwvoY/0
VjlS9Gqci/ThM5tFSU9RZPt1oBSIfi7kaS9+4XFDT0Lb7PZC0gAEcWokbvKnYh/2lN6q5Hh65jY+
irbraIGaiOlV6f5jBsr71v23jY/OgDKVdghZ4AM6/fMTZ93tG7//vqZHfSHIVOaCKYYsEHSXLMps
w6OeVw1zzEGrekjoxe6WfEIiwDyBid0gTOuzELJr9mAMolmaXsp2D9uC4cu9qEXrAiqDQ6p4cFzq
DcvbC1zUtLxx2gBGmtiI+Lcd8I1420tPw4D+0fM0FtWJguP6ouxyAYHlemhk1WXtk5Aq9hMW/TdL
VwECM4NlvVgzy3vGsZWEE/UsJwHjxOiYExr6Ktfa3Bi+qnz7SdnUubFdUWwhrgZyd32gP8dQuDJb
JDH7h9VWKkB/8hSZ8dcjThNEHtbPRF9OYt+led7/ysQ1CzS3AnBRmh6KUiYKY+ngrEoorWAuvemo
Erpuf2iXeS8yM/veruVCqQQiv6bfpcSOyN8n9jZ79VXJDW0PXK7q+jTQop6QfCuYP4U4OFZycwp+
iBb0cxRIGfsP8ZnA3gmNHqDPdNpruXe50TTAkIkGio91NnlFdZXFwdyyY8bh54v7EmGivJOT+ygw
p+e/En+NSnAD7171qM7oejYyL7pxDk3LJs9YYJ7wFe9E4ptz6TA8zJ+zQKgwUeS/fskEwx4i/qfc
5sFuGsPhn4u64DFWjItTYv8bEy7zKm0FseoYn32KAmNMEHPwGV+ITE6Gxd3UbT74nmXYLtxq3l9g
/1FEoUtTkOfJzcFxMS+t5pRsuyG6T0uCoRyzWTLBbEBwcXbK/5xpJ1fDQKSZpqyXHnd5bUPFOCxP
o1JH50ush1MpJKOlPAH1e3j6P1cCNzDp03CZ2LYfauk6af39fXi7F4kmGgmTYDaDiwWEVdfkoO6r
VAbYDxOLimN6qenKG79LaDFTbLvbMWxJzT1Gt47FhaBE9mv+gEIogBLXmIkuYAaD27m716mx9hxf
rtM+CqAtzw6ahAZIuXyRY3J9zEwGTbAarfTLCJk5x3Z1b8gDaBh1ORkLNTVJcRASIFys0lwv2vPf
DzHIav1i7U89srsCwaxTBycAZtv6goxhyXE7plkOW+ApKfUaKccuznmlr9sP+IVjaDjjKe4US6ty
pBYbcdCW31+CQm4YI6l2R5A4oKhDWZG27y7V3Lcqqn9N4BX6qp9mFPjZ0S3MpP0iqebWgw5ij6kC
jGSlpKlYJYPgDOndf7/2PMvk+e4FotyDLSEq3PR92rflo9xMGFnIR19oJ3va6JATvuBzOFxah5dd
UobzYTArjv9jx45T/1NzcSRDSEB/VDtJvNLLRW4hMgbpzJiheP7ltMunYQPi8sPZ6Xld3fQ6lOXZ
BHvSmyGGUpjINJBpE+C0jOlDs9zZzrPXsqHTsMiAfpvnYf/7+603JCpQHX7fLzU0QZoOl1X0qDMs
0e0U3BuO7MOqV5f2rrJHYsjLD+5KmiOEmAJ+dFRdJZN5EmUm9fy3QZsPBO8VrRn0IggzJwfzJ5PK
2698rWdat82YaSPZ1IYEriuQxlnaZGhfbvMiSHaqeSg2unB+zUMwx1R5IMVqbztpMzkE5CluinKt
pl0A9/BjHeeFoJxGQwoUCQbguevwIxyMZlWPuYKltbDu8k5hcyJluOi2dds6EzXqC55ZpfIYa2EI
Gsz0vLyTSv1kWeKW1duJ0Ctmy36FUeJ5PRM26xaH8BluRn/yx+2MVYJK8nWtGf2k3xrc6FwGqqgk
M56bmZ7vQ+wuS2FfRdVJjV3u2aZBxucZ0DCOfogXyFGVAlJge6HnI55R8P90CfQHTEXIWGCc1CB+
6to+rKqFof8uCuopeehUBjQ5mulzK0ZKlNfgaazXwgLhQRBwqRwyCfMWgUrHe55742bc3pVhg672
d++18ftUT4ElrH5VZDTr4qG1RHZZf27h38rDuh+EzLiQnR/507sR6E2rMorjiyGPVUYeX4mmrfoi
jhL9dGZo29xsXT12bhOp2Fx5pe68BYMpp5KovQ2uV4hnzzRxNZGzsm79f79RDwLji0QYDTe/L8WV
M3FupGa4tPjmtZBaRLGeiOjNDerr9GmGckb6pdrC7ZJc5cT/zizyptMaWyM4rCFNiWCaolvlaYGo
9Asp+jfzQRjf3t+uQf+BVC2A2CWO3j7bauk3+ms50UI7SILbH3fS+hXiMrMlA1IbrJMGqJ0Jf3Rc
5j6ol3mafC8MYkELhYvxfOM3O/UMX91fYgzEtfcHlWUqa7AmjuU4KvFOgZu2Rc95tI8NG/s1ihPS
TaOs3LuJUNrpUHNGeqkBtygLsN7CbuuEfsHdjcxNEmCgwyIITsSXM1HkQZnKfUHEWvI8bwe6RAGD
OgS/Uy09KgvOYnBcfUBSx7qhsqR242YFkqLenDZPQkOj04wJFKv2JqEeIMiQHUmcHDDQcLufbLoH
oVI497SS/HxzH0XOCRo5YHJxtSP0609YfnyFEfXlnL9DSZkcos7Hwr8mKqmbBMrgUiTL87dg02F8
/l6UkJMpY/x43aJBUR/IV7Tq3YK4Js8mFlspOe3ZkbCaB4A0NbbuC1+gMG+MIAPNWnG1syRJJAMZ
5+WlhBalWwtuZ189VRH5Uzkngl6ZVb3xte1X9fK5xY+Y+JyEBf90jTyppTZjEsOUnySNupPAQkXn
kdqQkUtSYPZGrVt/3A4BNKRB0qF4tcEZrRLagdegW00/BsfrTJPc9j4F1U3Ubq96AG6ipnh0z2V/
U8Wg/746cT6+s4yqorrS/XHvaEKoIbXefQsZ+JGYekvIpMyZtBajqAnIYt4w9phSBxr429W98z66
2axmElrYtYv0B2cJ4JdoI6VgJMVeXSo9BA/xQXHLhXoQSOPpneWt6XX1zIQb3zivnJb9Gy46BGIJ
t+t8HVQbxLTuUdOMrMyomLOQ+qaQKLwk8oHaSFKtxE+Oyt4aAkQF2oxDmnduTL2ByY6c/g0v3YDz
VGvjOaTepdOUdd1e2K5ocRK8zr0Uvui7dV3TVt5a1lrFIeeAw4s16BrRb5p0+bkjMQHpxU1VV8g3
FL7iTVpw5xINddafkmlmiLevyyt0tXABScmOopbEIeEZfYxt6h8bSdWkd2Lnl2EecAIwV/pOcuBZ
OgR2caNrU2yX30sVgDKUzCC2pK9gJ2SKa+vdmGWC73flD5TNniNa++NmB4E6kpLMkLs1iV+P/9Y6
VM3v71uoSZSimqJqbZAUd9+BHU3Y32/WlGC41Sl74NRuRpXr+NecCvOXrFcLfWs3Oyp0s28rgrAU
ABJrdLoU6pEcCxDkdT4fNLLPewNe/XNDONS60/5yROnicqoAJ6T11IKDJRfBospAqiJoVBzyqmTO
U5Nd+3bsdf3y2PqSPwHNcn1vy9ujD/DJDr+RvrPMioZ9xjW56m4p8ORlRXky8row9ozpg2g1U3kk
7AiXUPjcCaCofd1j0ie6gyUg3UbZCDP6E1g0qZ5Qrm8VdDPBYhBqIOL0smE9T0yklRRjC06Xn1ng
79U8xVXgs5Xlp+pHmy1IhI9mmR9ru/22Rxyj5U8wjv3HDqx2UpG3EgyhHWDYZ7lB4+q+3Y/CtdcI
Tl+RWElduaVI7iIsVKL9ox/2A6pQa6uwD2e9UHavLfBBrwAfamEhbvWw9FydezojS345jQnqkiC4
9PolwNZDCX6VlODq+p3e+H2rKYuwnHS7R+aiG7+m8JOsmCJ4hXJ5O5a5nHtEAUa43PouyLySNhTP
+IlpEthpVI+hC/RFF1jERsqcdq94O1pzE89u8veUiXZRELtly+2No7auZhQPmp4JPBdTDlmHJ6lv
v280V91DKHhSIi0rrKRiIN/VJTqYMtyT4xuRsFG3BzREUkHycH7Zoh2LjuUeg2mNv8ViJ4ny4Y3W
Wk4xkS+0SioqdJDRoDNEBiOpOF2i255ALz1xbmb9v8aUncj9AvMoURzJ0CD1X4QUnoKfuZ5hoST1
KqaE9tY1sJZEBaWJfsZZxHudEvdKQhCEUlclB47zk/C06y5H+qKu/9Z+EkuXX8JjmGd53kQzmGs7
C/hpvx3dov0XS5a3yToPeuceUMT7nmjwcIsOhzCVYMjFYAJ9FT7NY1wZfE1fpKBBd3wDLKT5vrAT
tqPJlexqhECbjNGdsZzLkfM2mGPSMXVipPGQLpFGL0E78P5hqyP6u4K4fq8fDhoVkkd6qQYP7v1b
3Zbf1zN5BGGWs0VHnSdLv36o/d6CSD6+L2zvCvqyg+/cTsNLVV/AK4/EFXpLXX5cEHxsqknqFSTy
A6c5OH6boEvYm73uapltyHuzr2zQFt93V75Aeyjx0qspnSVWF+fvr4GnMPt61colQ4rIZvUINups
zpLBqUBmH2tLHTlkdENupd4XMdkx7wZ3ODj5guxCTyq/0WD/w0Kp6hRbXd0eUuHtDQzAbIOIpXD8
mDjQAMs78AJW8UcZZDjVVtpe3iB+IdMlMGumuLe9mdyh89vXqsTmyGy55fJcQ1gJzLRhXuTd+GJ/
yuEtLPlghTlmpP4vdlglWo0FryPD9k0cqh6btfpgwpyMoz+fh/d1+Sr1/DRU6GasRv7bUYhfzcYv
6c6KTlmFiXFuoyZTihXAccqzjCGGpaKOqCFemhn0BbpW7Rk6TyBdEmSD/6eojGRf9ZdreKcnWvw5
mWOoIPI8YVmsA2aCu6V5jMb5cD38HylO8TViZEpRM2iBAStJMzJqHZ4JM4ZSR229h4CZyYzPUiSB
scvqY/3VUNCZZg3Ob9JWfuFzZoieMnwvEl9EMBSbxqK7hBQIGJWCNUodaFCZRE/Zi9PrdU9U+viR
t5OeFotxyMVUf/fx+jCGMKqJA98JCRSvSHfNAnyxq3RcLpv05Eid/8cWdGkkGVy5jjAuIM8ONVc9
hhMBynxKHXuMzLeKaG6Cm1afyErCHXOwghV6/Ub/bqTLCimNp8+znGpxjM3INK5rl+b4c6QgmH+x
a3t3JLjdOfVsfHSOLwwGhkdefoTz0Da6vqKrJEgCbm6JswgYqEbtBS9i/yBcc2sTexdejg5lXqfp
m446GN7EtpoVDbchiGsspEdPSJ1ZPP4RT3uqJu1JVl1/XOodY4xqGNk5fJ1qSFAejHTdXAHgqiHQ
kuzi7l1Tn1FqW+TJHkwZzAkG6+f1d6uEbsaDZ9GyOPdMPSZcwX8Q7sFyJXKlnoJ1/HHx0FSURK7W
jSr0Fl2GQixQp04gyCV9+gyf9a2b7ywaYYrDKLxPPUqQYJpsP14kqn2nV7vyJ506t6/zMYTn0snr
T1zJMOVe40TZsCSmSzZXMoyem8dacijzDLMEjhvW3J1Q/4nzqXIYLb7eYEJOvyYFvivjSHAFKZlh
iEZgK8uLTQ9z4Q6NN44dDuRycTiD22alqjs7BHjL35gPzvMKYQX+G4pfsxcaSE0u/S7FNYwVFpf6
Z45qrJ3Gkt58rxZQhe64y5884H4uO+FbVg76o1tncZxKLCWcBQEFw+WdqpKkzK8gIs5Z2NWDYCK3
JS97RjNFnB+r5JOrGU+elAg39NeJTghxtIPJUFE1niXe2DFCyQ9S/UpkcnrRT/yy0SGicRN9wk3D
ul9SEgxAzIM4eoNrnMswH4aCciyiIg8IYRqV8MGYsyVaexmPrjmaUpC1ZO+JWqK/xfvv74Z8S1Cb
IGNEXiuvos8KgzMf0RSq2slCXkVaqiam3DTRvd/mwoyGm02suUssLRfUFIXZl5O3hl8Witg9s+4F
POYZ9M2xIeviVmW+hnnPSi25pCGEp8pPrjat3PCloCCvFydBUiZ5kEq30Mx395OO1rmBXzQDhb0t
1D3RguRZCegpS1bVl5Zk5PzwfJsdWjaRePSKapJ6MOgl3JCEEXLWPLUPpU9HnO5ROWWVymjkjRf2
jNPJhjAuDBCpsEJoZ5ig/BeO0fW+AyBppWUCqHyi0SL8gNnI6adjYis3wWAZGmAhpzOHZ2iyEWco
+OY3sT9StQzboaYfacqIj3YFau7khvhcawnm9gi474W6+T9Le8/ZgDbXmFqxvmWD8NY3tbEZ5JFV
eunk65ProbLebrLwx+xpcDe4uawNIBrZWOZF6kCTrMKZu9MAF5B8QbQ+c6YpnhvatXyeVdBj85LW
ARrVskoUj8mxntMMOBRqUHvPIIhLaD3z9lkSArQsJsLv25DFXjwPtfropHgCrViEI09bh8xLcGOC
txt1WGXjn1kbVxcZxmJQqaQI0CQmyZ3HyfkA3nNg049AsXfQf9doYUSSpXXn7QAFpaXwc4Z7IiwN
ilM7+IOhW5rgyTSeGFSLqNkT/v1YSkeKVXr5mvbeleZpBTEMBjZruZxbaFSik9VFFb/qGJDqipk5
ZOI5HGds8kRuomnzh+D0rcBYI+BAoHpVbNbDVoIYLPQsmMqHnfgVtrORqW1o5s201SNEYIjFO9Yo
KkDbVneZERQb15WMYGTHZKJVnoIbtiVE6tON/7D2KWgWxJl9xBlT4iTEr03GvmkSSC0ac7QytGAN
NLh0Wd3CXJx4QfTtc6wGvDGAcgGkmbV8CoyLHbBgFQL83wxQJv8dVPVxaEDVkO/BeyKmmnG1MLYo
CeQbv9r8qC2fHpmT0OXosaRWoXnc8zqUs/j0SzkhoJ1Tg3SYU4hjhEphdrJ/OP9zgCDNFizaL6DG
dugRFS8lzod1HbGK25TvFFNBtxEnbOp8n3cKDyqapz0fNLOIYtM9NELqfM+dr5e/RR8UYKMElwih
YQf6ICAnMSJMCo02v2hq8gOXGos8dQDnPD8JGiGzGaTqkEWZuVrjPb9lPNhw8EcCkdolGTR2zGiu
Kq4YyxCXk30be7tYBmAwMcSuD1OMRjiPLvTxwkj4tAbDPn2rancIRQWymkXAnl2hJ25lVYdZMAk9
1Fixkjv1sRWzs9VwEY97np6NCylyc6cg7IXP1AuzReulm1KpDZtecenEzPYQGhdHY2v+tJxULH7m
ixg/UmsfVrlomt/WqnWtAvrH/lBpyVcvoTe35xEYHk8Ro9ppl3axBhWJUcWIezEhPQnjGaTmXiq1
QgCTfZ5rxvb5jSbXpNNODP9HbG3jsq5qcFw0Qv1FKLGnCCIR9POj268FFj4fgYTH64Gz+6qWHfmy
Auf5ZPYqxNihho/o+086cjgj1kens5PlYNRJPnmG5ofsBCr9Py1HM3geg39RbJ8o3C+5jlHSJc7B
5Sx9ixZxX2k4p29x0ZOVpsFqENR0+dDw5WFW+bdjjeuFdNDN0WTvkaLETyookafnOMJn+GFXjbcm
Nb4M3CMHj6+ORxRNn7YUeH5Sxcw0Es+m2VLGmnrWeQ4XK7rTk4W86u62uJfOUoLEkNo5+8Rv1WwA
Xa6XbzHj4rZGkTqLljec1Qk2982HS66xJthd++MEH5uZRC0qWOHznkDXdQC1aXLF5u2t2JG80auP
dG5g2FzEq/yVkqFmvzpmOX7T9LuVU1u4tYmfUqZoPbvIbK/S7W949ZmlN9mRlotxPMWosaznRTiH
gsK8PwgvL3Qi8b2/CgsJshNFRP1ehtnWUnWwJaR+d+WpXO6k2m0woDXV0xitCzSIC6pwloLMOEDy
ESyuaF79uNTEShpTrcAkxZza6kSkZ/0MLa2Fo7L4CKpB5qdzDaZ0hfWlp1e0nnCltNQL791fLAkf
tq3MDcjkalxFd0GIZktbI8oird4d3S54j47xPjhDw2kyZoamFKCRxj0quyORWK+YDIjnD59bqkI2
cqgLiM/vvafytMrwquLUaKropFjGfd9n4I0iQ4cvU18XAP80+R1fojXg/gJq6xGim7/RLmTJecF7
AIm6HDIGEN69TyVaOZDM0gJj+tFnYO5bLaGWc5ykbeeniX9IMxc/g6eqfK9Edorx+zl0FOSs/J2g
SsMv1D2WowO7AamYoqbG4tUHu4l2qhAnxbPEQvM40UJ34tPXBudTBbQKZ57RBAE/gTxbnzRkp5xo
hBj4Y4EbOKkAt2nfxci+FRjrg+A2IJDqOq1d5wrHyE4fZmh4Yr1g5fdKUYHaX7kjbI4yLxs6aYrI
48xUh2RQwd4Ad2h4Yo6EHryrCMdar9ZYj4X6KibmB/Gn9YIW+Pe6Q1c3h0XIRGx+/ewFnMV1CosR
rFI9xU//rgRZaAlK5W+modzmAIpySUidyAQvTqUtru9G7Lb7376O6uxcrreKouowncOFQ/ZcQEZR
Zdklg8dKRaxTTMkJGqpkiiLdV28fqiZ5smRgtvc3g2BG7kKBMIUXXiUORjJneQE0L+YCh5o8M7pL
ThyqQfDORDjnKWezrWd+Qm2cHjNeej9cJ5iDntRGqXrD0NqeIuuxSkqh+k9ijMJEI9Y2Ewz7129e
sAyJDkx20dc3vnlQUcskCPhHl4GhrEb5NJTYn78RYWX8UV0E3qwrhgOTYlb5YFZmORMAP0ZxhHQh
5qIzrwgkBozeTrNIuyh3hA1JQcjo1/vU9nPk9Ahqx8nv+wnorvupPjqxRJMIYG2Y4m7I2tjX6co1
TKuvuX7Pml7z74utqVmUFhH0kaNoYfFvAjMMkuuRU4WZXvDzK9vAVsDlaZD76PJVfCQEFHXLvWyl
D4fqiZE5jmqdrnnZ5rd/DfYaXzcJhbvA8d3cUxHTKx0IIhTOtgXUJYldoUE8b8fv8KGiLOddso7/
TtSZF4PujDDjpJasbEGLHYntXWI6eQuoqIjpVRPB+LxhGZhDzow8I8hScfN4JYovja9kRJ1gtET7
axjWWxpQVBDPdlQtP0TGzWtKnlPVOlGwflCiR/pvAXCON3+vPyDYOXRjb4Oew5twNFJoNhm8rmGa
P+1bFz5s9HmQVmiYz8/aPl14P8sT6dr2XmqRFSL36lal0HLENCgnH5+aWK1o5ZPQ3iXfOD7Dc/lG
W2yKKqcsmFxkt9IcrkhklAh8ZltkF6QiULxx9kV9kjVsrvZia4yYj/Rc4TpzdqHrkoV3F3RYeu5F
LnOBGap4N1ja0p2E6XQnnMmSV/mSJX/Uiw4yhDBRZ+EUVmvq9cc+7w+WOvZ9A6n1uineVO+abTHF
FcPJMJ8la1kSVAO73gLAbzZJVtmvarWxCWRYHQqmrTsifdOf162FKToEgwGsyVsjcnpVMkwu9dc0
j7FR4mU6lWc5REcJRm8zXKnsMbE4hhy2tNN78aFI2Q6LOhaj3H8jzjzDAhRVJMjCt0sl1phQpE0W
AuQHh6J09p8eOIggs9/CjsThRBpcUEgdqy2SfV6c3IoNB2Nyy76e5/ANIGO04uTDn17sQL9BD66r
QZlLeXM7deT7ZZ4k7XEnHNvzP+D7tyjnz4oG6TUpv4CzlGp1dscCFOfQCOtOPWbDOdMZqlj+jiv5
gDQEHsOPF9u63WDi6EzpmkbTUYPu40Nnlgm8V3t82xWODLjpThJdTscqBtj/NjVOGBmvfHlW+g7O
Q6ro3fe+uhFQWIzmcURFhx/4fl0j1eY1qnvV1lf916BO49LF7QVzcArFCc/gSxvJCKFT4D+hXAah
Ml70iD6OwLSp323SlQWY37YVziQyok9JqD+DAHOOEQp/qPNpXOE1f7JI3h15u1xlVK8hUIinSTnx
EwySeLXw3kzWejoGNLkDa9ExtA60saYrYWAmdPYCnvc4L02UBqCUax/L+SaNAhrRLVoZx/9X5k7V
SrJX/Q6xNgs+1wqPBY99GXmsKzK2plwZBBFrDw+YNvSguC/774Uooeyg/vlX0/2pTTM67iI+NfFQ
Y7tcn/X2b8+x06kN1+5Urh4v2i3Cukd0TpLcVhEIphQZAC9wrXMaqt+pfBgS5PRstMk1g0Gt68yD
MEgJp3uKlMtYQQsa+ObnRSIsGdYA/AvUhTy3BxLW3/pTiBdtCT/kp01orc7Nt+fri8JNbrxmo2jP
D3j6pRyOYLayMokCN9/aQaIB3KeucHlm/czmV7/v1x4OCD32ZI+fOn2AV5HUgR5RZIOpbKB3vYeB
sZ5BjsYgOHE6tRduo0y37j2BXZfbUndcfhwVE/4jHuoQiRemZ09DxrnIoenQPLxrSpYH8L8c3htL
GlL3tTHP1NzjO4Zi8KC19ERtAza75b4mTTiloBf3UaNSk9tfOcb9eeKByQYzkhsaOT/tVoRGZItp
+e3Ff2BaduR8OuLimkTubLNbMogbOLDDVH/H/uGjyCf6Z6YwNBYUeK9aObYYT7rZkKfJFjuy7yI+
kebA3a2QG1S9shPUo5krvsHwb3x3zlgTW7iBOphN3jrAeMQpi2QgVKDWFWBOXVh0D0tPjANuQFrc
646jqa+xho2IIupQEjVMjpVDRLOrnduewMP3gT0/iAL3OmKFF/5zxPUiGgOYDzKDQxWF8OrpAVE+
JebX6T++1lJ38L6XETGXxhnPInR+2ZRn8XLOc/s9v7emO6Z6UbRaniw2fMhLxEtPBLsARsmeIVDz
88egUDZKT/6K6pOPcP9IiUM1K4rJkTonYFcU4RimNlYFtCSVvm2PWJDkjlWDbOD3Yy5TxVnRfniH
5hBUrrMzp5SISyO16GJN6UsM0h6vI3cscsn8/6Tj7F94XlzqDno5jnjFZ1WQ4PS2YJ77EqlOu5Az
/30vXNVy0/oOQKvEE7uLCIySm2s3g0uh4IyRXo9OJvqE2AFQOdL+Qk8GmuiuYClHdJAETpMVe8Ev
RCsRPWyCgJATZUenIafwaofKDZ50DrUka83M4IUwcAjH1QYrNxx5/YvdSEeYMHNQaw4vkLFHujky
lw/6YWuwt8x59gMOeLW06QhCfUR5EhAueFMaQzwuEbZ05B58mwCue7pTi7qbIoiMOeJHTxtg1TUJ
6AKNrseirz1ZR05hs8ZWZ7vs/mNNK4k3QKUKWboYU5WOE2m/YOKjyfmeH4GR/jnmrvjqjTG4jSep
p92geYyPc98391X5/qNSXRVL5Ls60Gqh29p4hNXz+bHaaKoYA1QJQ+obvcVo+xLD08pjWQyhhJvi
d0LZDd6JdtrkA7O5nZm0THhpOZbN2F86v+4kKThqtO9DID+Ek8mN30XLn8OwpZwf0K61iVtOzUSM
okjnu1OdR0YskXv5AaIkRoqwVunAyi0NcnCtpLCBY4uviDYaaO1bxy/TWI/5ACUDlqxYSQCE0oQ7
1x083+yWsYYRHaoyXWCujS31y6ZWC4kCZk9/wRW0+Xgc6i1vrvyXTs4wuoAdh9NnAY6U0dWnaZ+w
a/z2W9YItScrw9qSRqkABhgHHZEOwdX9nq9t8inXchm0vnKmQPpHRVc7r+5VT0tRmPMFnhwUp/aP
g/Xwq7kMd9noFcTnts3jbKm/RMBL5bMzCDGRedE3vByaQz9WN6yVEzWFi6H9jQCKGsdIhMrmDW+B
aUwa+X2LLw8ENrLlFcZsUPyzCWCocBnm6btyGR/Ur6T0FP7SFG0n5Da+wfMsV4N389N8axxMfFGb
a4tq3MSQuXGEFNhnREuHPpcMw8y9I8KLG5kbzF1XA16nvycrTkLDygvoBaAV6qlPD/8yPJXdUfXa
NsYI4KXtOStoB3jfTfo5Vn165Vd5FHeaYL2lTx2Z6iR1hy5eDR3qDQjxqO71CJ+19P7pPIYCAyH3
1ZStwrJyDGu23UrFx1/0oP1REmgXwr6Hp1brTj2rbiOD8C3qWuIZKHWE96fcFPpcmBW/IPLlXhjo
+s4nuiEtJliC9BAneHZqoS5JhMwmq4ge8vsu966rmywg9oO8ShLaQB2BQ3y4XpZ6JWoq2wG14eHN
Ljobm7BS6QUiswdcpcKaOfGq/EKW8RhJo+02CSA/vn1uOcNW2KzmqTh68gHbvMsdKV+ofCPgOXrF
wyVsfDaXhXy/PTItiQRB/QwVlkCd8Q4Xyo09BuBhRLjeW2hDj9GkILBkzOuSZCqXrTy7qTQEuV0d
GLGlsu59C/bBLO9aceYIYCKFTmJRFsiw0MwUqkCdAEjcaSrlWv2BAvX48Epbwi6INShHwAoKUXKr
xbS3V7yCcnvGe6uXwoJ9IvcdvYwM7B86IFUSZcYEnvSDBf+mwjOf7CURLtG+qQLeXEv79+K3nea1
SReXUCnjCzsZuAPn/qtTIxqBFIF2chZ0nEuJKo2KQStFCAOwnVwDmyJgUb3Oat1yuNRi1SdiRaiq
FQnTaJnT8p8sLmDS+QzyOCJhu+s8NK8hesodu7dkNGOuq9j1nAVW7ZxHQEEBdkfwZRdLidkMvWte
esbjKYwqLu7q/r1J4yRPQRdHUPZjiVTh9t8aiyQz4OfT/gOWdhgUxd7hw6B/yFFpmkvwKrJ97ka2
lc+Z9F4oNFWcib10Sv3/avJ5gYmxlhZGpXKsQPe0LP18OK2pBFd1vPUdpyfOxTqTxsrTT43Hy23j
NSUOyTRMPJt5XiJ5/m9Blwvp1MLiPG+qtRBH5+4JiJb/gKraddxYGjX6e5ye/OWjf2tF92XI3o0B
2sTi0ctQt8keuWAB21rrnOSc98XB9g0kJI42UgdimxLdz6Aock7JfBRH/PEwtotp0fqf9rRZXiId
5PMcfWNIxqnvLLqiXGJSsQna00V5tBJ6LJSKCDqQpsEPo9fk8PAPqbb98DARLX84f9+BFgYg2CPA
NNkK7PuXKkuFCdkOriAbCXOUBDwQgNzfvelFnM987gEI8TCHBS9OrQHjTl0BpHfxzRmSBch9/ZU6
EHq+zAEogy8wBxjgwzKUsD8APrW4uM6pZZBr2ytF7u9J3wM2msOy5KdAP84YVNcoTTKUMP5O6jI5
i8RtKcqvhLrxvGsQ+4hGjdzqCbACTQzcUJbAJW5KvsKXPTEwR7BBLnJH9xGov9MuXw3jU/Q2V4A1
WgJI6Hzg9xD47Ovh+6G2roCtnIamZrw5xFNfisMrT+jwUpthaHAaoI8uXjX0nXVPPFOV/tSCl5T4
wkPfWRrwChYlB989g3EyC4wc0Tfk7GtYvP+/QjVizBgatFAEjwH/TuPDbZyD3YJ6cj2MrT4lPTbC
yzkz+PIp4xTgHnUqhoebd/G/sPDXE3btZajlaKF79aAaZuc4wEgoDFRfy19nkylVUYoSeNhn2ZTa
VoLfVDP8CUG0kJz3aeNF9tESoIWWrYgNpCWeRlVCYrLcPWJVjjwh5OGkZ2EDSWJYKw3y54cjezwQ
WvUcIsEMyMeRe1mGrOeka5zUwQgb2+IPzAjzHK2foFfH6rNBt/a5SmlJeQwqAWWO7jqaAl0bsZE3
QxRirgsc8D9yk2aZiIum8oWD6PjgD/l1mj/g6hvWGbl+b4GmoGYWeqmMqcufrnLCxbToJFV7aNqL
ZgnMaQcWD8c/2fHyhGRUxmFTvw82O8VQq7aV53EyG4/RZ7+N2yaY4CEq68IX9Da8X+OCfQqZZN93
fgIcSsNQonGGaOrichxXeIyO6vSjnalF04Uy/1sC/waGsngkB3Omz9++Qet9DFdPxAdbbE76XiFR
y0MsCF5FXgxHSBTcKeG6zelZAL/iNxF7Zxntam4xxLy01J8+JCuQTyIAuIpVv2KF2U4ldKK3eWzj
AwBopIVx1/oRGUV/+oizyvMOpOVxRxF+TAcSDeOTfPYj+UIV/CFqWnD+QHRgbaXuHWUzuMpbIxCj
MrVbqrCKNVjZsT1mAIonj2+YNqPalqp8AHcxVvcMjUyeUOddim9ABgdm2GHMjVy770b/5yKhq8d8
kWKdno9KMd21AS9YYQBpeGkK+E0WCr+CBZRMqAthXXM5DYZCEDZWddfIYVp3tAEG6pgDWEH5BXy0
haLBYQygV0rPwosMVxAZ8iZEysgX0Uh9C2835Y2qUOehjvDyJ8Tl8bKKO6oGk7mQ7jtR6+B1qqfj
UYcdZhnTTxOwCKDv4EahjQgMNkAKO3cbD+mK/ECIz9UwpoaAONZ8GFnlPBE6csCP9tnb027zAIuV
Ezao61lOzP8s05NZfmuxWS8UDvNUo5F5AyYH3udjxamy4K5Eh3C/MkX9BX5ly8IDUrT6sJUm4sSf
Q22G6ove7VhVnndAKWJhE2kLsna7Z7lkkIKVS4E42GpNIV5ZQqK0z5X7ZHvM3yZgEhUeFozO5A6o
Eln1I8kaQY2+1lErZY1UAhH7n02+ifxiaI32TO4ZEMNumfngs5L5OxapRrOT9Hye79+pMKoiMitI
J0M+jQ+nm2qGF1+M7WeW63HWUBvDqBtxlAEVLmqTde8SmIJBo7j7krowbWpz9VHhQp+gHMJoc7af
8Cvpg4893jpgwHnJhRCd3IEWn3NzrrBvCamXtq8lAaGDDiZXOSJWhiXBtP4zDwzSyzUiXeeyHKoL
z9r17o8oqeVJ46/KUgcZYrqw8X5psWqbeI1xOkPahU9TzL338W/rCyMgPOqOiX68dUnxQ37A7U1u
yBDxnzl0n5by+RQmi7/3YpX8Yrhd38KQFQ7Hz9WAdC1Pe4PZY06EiG72ymekF4+68erBIb8m6TCa
S7v+VETQzCt7qeFLNn27a0bbJpoTNURcHz5SL72JcgvZytlzStIYYoZjAteD9dn9P9ZS0f+81eLI
QJ+aqen4FEqWxIkQ9YjIw/87gXwa708YQ6SEHxyadDXyBMu1M/vHeHZmiWwnMMBkmNKa0q/rmFXc
UG/clLZg8+7VipLjf48aaen7gY0aAa4l6KmjsNhKScgX1kE6n8CAmsy8dzrCEMRiZPGCphlrb+d8
6tJekGUWaR2j+C+6OJwYgbDNvM6WWxgoyD3bF8PlpMXQfbFmSMPxGmHRv78YW5k4hkr1HM8/ZD0u
B+2d6BeTGOK/huQwUIHhOfinhL5J5UviEXqAZdaL5Z9QajA7MQvWsJPtvhXRBWKpj8zYF1qmqFtH
ITQOn96LnC86FFzbf1AlvLRXZL3l9CTQtZo1HUx6ruIdwXMFzAiRcVERCoSoLxjKAjt3RKgE8aGT
XMYCC5IM44giPD4DBXbFAmPDEeidvnrj4NeuWLtTQWUYpRx3eJUhMkZ8Yj/goH+kvGZ7cbGmhZGH
dWGtAN/GN/9f4yz1eC3NWatyF8328cphkhUyf8YSL1li4IFp1KpL/zP6s2r8vOmPJ/VRQN6SYiq4
Cx/1bbWa4T7anNU9ZuWyzgbQnNbJnjNdId/DxziMPiV02s0ejpSTl0WKbNV3unng2YaoqRplTdWe
a7qLllvhkJVjwlPgF/Nmzc1GWv8E09dJE8MMlBlhWtsmv9R9OdjxIrJlrdSOmuXbbEOaC0GsTTD+
yOGf59NCoUR2+DMdruteJMHUwEqIH3W5se9PSYUfRpAV3u+posspJGrimmiMKRhsOomK5dFc8+2M
OUux27kF7YK2FbcqeAGOPWqxwQLm3q2yM6kS0IGBD+mhrQoM2YpGdGKd7p68TvtmrOKyb+r2rgu5
+YZBkI80IUaxwvGjz+gRYMBGjd8nWgif69KVRktDMrTfg78GYdqm3SXDalPVIgfrdeNwux6Da5FV
xCFo6cQ83jsQx/sFZXffjdGNCy4GOyBGcfQ/3DyzA3jwf06/haHcbIBZNLLTsyaeSvbH/dmw8R2n
MsrRF/DKdc+c+xi79Xvpup+P+dIGfV1zKg8SCBi6VOtSKdU8S995OtT5VT2Dgy6SsyKetaP9YxNl
bJNntGz5Xh//lWfx+BH5RROxPwRy8ZGqDMyk5A8YJnsTyjQwPXPJTjN1gQTeJpNPUDk7HLSrKlgK
9GzZ3KUXUAbyx6F0aNH32UKTeBEXs/qlSvi3XxN1i+vHE/zwU9ZhSFLCLoV0fUEm4KNwHeTzaiYK
hqyFwzhRHhbHfR42/yEWOV/zmCpxW5BmtPg6FUiyPq6IKcRqzq9QOS8qcJcBnSLTOQFKiswv9hoj
/nPDb5u4c+zvJYwbpyEq5aH+WqSmdb3+bUOlHB3KXBOuHtT/dZAEkYy22hddNr5S1eJnWefzD+Uf
wRq9jto4KYUq+LJ7GoaimRgCABQFfpODgoo+60F6jgsZQiz2YxnCRpcAx8l0XHKXX7JadS5smgXN
zAJds9CNdQAgxip+ySjT+lQabVVDhE2V1J+A/ZHNOEpD2e3O+lIaiZnNUK2wORVjq4LN+CdBtbPG
HERfiP0DSgtS4kXFgMwQeEOgDz4H+TMJ9jtsmBFw6FH1GfflBgEFG0l+8EO8yXXyVsF+LtY2OFXn
Y9yyTmYtvnjeUmTgxXf75tyqc20GMAYJZ3TE+Bsf5HDxtqiMm2X/QkKfPJP8r7ovLfPffTnHmwH0
yfKIEII4qpkkpWggX1wmbLbLoCPRGa5z/5jQgRVAwC4KSsGBgvzpF3v5KK4uoMMCkHdKsv/M7fTq
vnUyrodvfhuwh++pTbw8FxmweXONj/i4YXOBw/JwqKM/Op/1ISKdX9DjvgofGUnMmYcjOH1CpM3J
6K768hoWMIuLycMOeuh4VeneB4ONS79yJXGIz5NAEQeyq/MQHtchTrnL0l6PUBjb9p492K8EAUeA
CWgUnYOKABxIK9kPhESLCEFPC3avzIuVGvR9WIcgpi7y3D9DDxumb/mYldDIApCKszwRbjiZQ/+X
YsSS+K2cZ0G6g55N1/ru2ZPyRsUW/N94oZVlYFNAw1fomsHjbLUAq5uAfmDeOQ5srgxc9P8ocNk9
xNp7j8N7hvx/5262zvis/ZGJb6Nw+oAsLRvfmoHwwLBIkPRuGzrBzRGEVctInG574Pn8WEuUAXsf
pwlo/JHgFEfzEbgxCu1Z7SvKTVkBuLtsUgEwCCUJNV3W11PYJPW5yqIDQH8VV4zWM/vgksyeerf3
8V+vj//dvJjo6Ltj0E7vWZweKvA9tuhEb97RftjTbxTdgBRqzYg0GjsW88zV3n/0gik4tCb8AsnP
FBmPpVH3EHtAQokegASSU+bPOgKl5yHECfHdJI5BDDoAF023ryCgGk/ebttpnCepHGREE8fqvvzY
mUJzoR6+AK4oSXdXBSfRQKneNVp+jN89ZJ/BAr263SluWJNJaP7tCByTjZ8DlP2Tv5LjhyP6ENTu
pvtfNxfe45bbgbjHWp0xTm3dABYCLSScGqOl7mO1UgT+l/J3yjzSwp5VOPUhvlPY06429FGf2H8y
hZMCEbftbs0qtcdOm9udHYUh643BzqtFsbM5xjNGWFLSXuhNr1H2Ggb/hMBp3Iv4xgIUwG/RJpkc
ROhF3MMv8lEFxtMRhNI4jct9uH2Nio0QgswJhE5IOFNvDV0rzhwRPf94MV7vpayAcnZ8IV+NljdJ
rZ3d/4HF4hH39oGp/KwYKtSXz2U7l38PQ2gVABiF8a71T+FfP4bcLp1fA3Tw/wIhtoq1TfswJMFt
Djiuvo30d5g5wBvmXT+O+sENft5fzEU8V4LaO9L9Xa15gypzoHCpBt+R5W+wddazStXo9Db1AC6W
NvlDZakiRfA3s7RBA7fPgk6bPhCSRCv1tz0BfkMsgybj7EvcoFrDZs2sHzt+do5zp/YJyBPrqAjm
eBYfs2PrGFYP91mRuxM2a6Jjz+2/AZSayMdnpGZvk+dN2zoSDOsYekiY9dRuqj1eQyP3acJPx85E
iTMKcSGlcaZPKW58Y5EprDpZT0e8fGtR4Gobui05UFznOVVcs3TldK9jhfPE1SWX7LQowL0mz22h
vp+jZgBFFdH4jVo4oierSQkDDrUNMOx6N76F+S/B4q/fOpoE9UAjQ2Jm+O2wczesINv/7hMzeV+Y
Q6LwI2yuMls8/YaJSXu7xiBB2cFfX3iHH+ndvzjgg5desQJK1kiGt8zjePGcmxuGJkoC1qHIbN/Y
kSFarY/CLHg0Fv87J7Qey0K9Nq07HdldLfhxmB5ijM+IcxhxS9kPU2dVQPNhAbAlFLw8bkICioq2
nCG/vN+7tPBFv4JNm/pyLMbZjpIiYaCCz2qxbIfOUQChzIeWOTiPCwPs0Ya2yOFgyRBLponreLtA
UKGqF7VKl52TVPzQrQolgFyi/ajPJgZKczzNAQx5WQ4V/H9dXSAO4W/YZJg7/OEb3vY8gThjZ0Ds
sUXv8+ukzkPzfBjF4pOIHEj2ZATYdOEGfpTXmtCzXPsjjd2LOe5pCKp1NefrbcMj5X3Fh9ZW0l4I
waRrMerccLjhvrdBYEK9i7yHqYVMTVpVAz3IpgliYzXxsydxW3mdYiB65hpVypz+2JN6gScjnS8p
75Xo5HPCoe8AmC8uA9nZVDnbLASB10JrZJrlqhaEbJc88PM/FPaaaLZ3GIZXjC5uVPNRGcz/jD+P
M0/dSt2MYfDg0CrvLTKRXyyBC9fTaZVYhJhfV3NuKOncE2iMuhZSh+F2/n1zj/s7Wr6yLvLkujYS
F/DqgSApxlNcoF7Fmh90o7vdeYxm4V3RfZtl4mjMY2aCdyGIGzs2P2vXdlOduEeTFRFxhKctdqr1
28tpl6GBWOq7CDJgCjcTVbyeX6fMKSfuIjjMxJi0zcOpa4nZ4myFlCWZyYhrUmpCd1hZD1StTzh5
+zE3XBsuO5p5J84isjcbqPybMUSZW0hZH8XY13JsA3iLPssBbKfDJzEWmnhpUqD+bAe55wugLsKr
10wxF7aYK+DZk5b/QOZFmHqzHWlT2dOWPIwqQkyoHUwF1Oi2CskvedDrI671Xtscg95HruQ3qEOc
OhQdo12Jy8YVWoPpDxj85opG1wmS2PvXHHHBNU81WwCv6Ivlk717zwijOzJ8LEeLwjkW2SiflqRK
d705DXn3nzBzD+es0UBlmbAcDKdunXwqFdyG9DaZAgwsqaaAsRDBMN9KMNRxLuyjaag6tCf1eYGI
jmkrS8JfFlK/GqnSYhS4ymnR0W2VZWdWQJMrVpvMkTT9PS+C57UYuTWNNlE6t1svIBG5vLwRYL/T
ZI7v9qaRIfFHC4Hy3YtC/F4lt38UhLu9lvBz+sqEDEuXJabWM5RnaWboDzF0lVXhZ2S/FuMpXakI
1NM1Juo+Trc5WEzxF/8rv3JLDaCHUv4rGOhKIIrvSAxicpo6iNOJIhXjhT05nRnS3niFqwmh1Fi0
cZUidg4yjTb9QEQPxHFIAgzpo68c2q6plmD4ZWolBqtjnnqZJOerMgf86ayb/4ruxwhGN2MiaXWG
CdFuoL/4hPYq9+rO9j/uuf3j7N39pWAklk+jSoMr/Ol/xREfWXQCy9gQ+RLWNitSmeK1i+6Xbg2w
LZG7Sd/Lb0HOwCCVuvSZsllGufWIkMIftWY27R/dpMzKkiaCL8UW9It5vIdFk9M1p5Q+01Q4rbrD
lJBScH8sQXZfG05+lpQt6267HFdgHpiMcQjF6osdc/Cwi2GvgzDLvfffjXjUYCRzw38nf0TXy1kP
tLg33lAQ+fNt9ifYlMX2qVbj/Wnc1yk/0hQfSF4pDXgpbRrQyKd845wLoJ5A8A0uRpDLgBr42fzd
DwqCUyhdt9e/pB6JbYiSIXlHdkP0kNGWhG5CrzgbjS6uu7u3OWIViyhhTbQYGXnQjfDnzADBg8gH
zF+i/Y0bbD8PpONjhdyDHQGi40o6hrbNl4o1gbLsAfqYCDlHqHdDN/HPKppaIqw+kIwyHZLx20vK
dsNQRgfTtO6fa7l0831UUnRZDHrW82HwCoiLquUKnI3WWewq1eeRU27ItU1AfGuHPjp2p+/dIcfF
YX14jKvIXJ0fo+dinaEnxFUvDc61kQ7/tfHDikPYUNJP4vRfo6D3O5BEElHRMBAZKzia1h6/qpEt
I0ZFKAs0fz8vTu8GfZell1K821Jqtpc4T0Owt7SqBblYLVST7NxqqfDeserHo8FxCBRKSbLO/EuV
+VtnrpreQ6Q0cQ+ya5coi34RwXsU9BujDQEEQfabq1LgYWvTkeANzzw7/DPCWMqCYcbgVI4B3EWJ
WXXpkF463eh4UiPEgk1phDv6UVruvIaMV4+psxjjGlcPtBRNfu7VQJXvQH1zsMsV8cK19Q2JET68
Qju0Muyu3MwcH3O25SH99aLkfeiZOnV2t13WFUhXWB4Nb65Jg+6xvdX4W0aBGlj9BKsWzGTL1edy
m70Wrry8MVoNsD5VzrYGopTpecVJRxn2k/XSFcFiDqUfJOQ6v5FRBcm8dequh97FzbWI0U8/rZ0b
V40PKBfahX2Ap+33ma2hV5RV2mFgnfzcGH8dVZ1qqYBYLaTX9ovhJpltrS4Hyk1w5zJ9fSH2xjF8
HoAbI2HzY2FohPJ3W8+pVZi6UbjEV6VvYYE6BYzfH6hd4N+AtEdi63LH/A8qMjd0xlduisKYAvLY
zg/hscGyczAEHhq/o8a2Wb6MpzH8fbkd4Go+B1PcsLv6LqlWxFXRT/3IbnMSFi+k9zZ71coOeSYR
U6iFKSD2Ve1ojOOjlz4AxOurueh78kB05BNu7gOkL7nS1HY8sDEn1FJknB/V+2i81mHeY65sps9o
GuOPduXW3MxqTK71+FkxHET3Dfen9gXe94PDQQ4BLxr92vfKos/+jdvQL38ezl9VTpffDHgAgs8+
Gr/FA6S1FZw7tcSIn7i7Y8MfgyiWUh26TXKkp+MyfBvmdlT/z/+3meHTnw1HNxafTHo8JerEdw/B
WeSDAx7sLOCzOkzXp+/mjdQe41303r0MHPWJlFsAdEhxyVWb1o4T5y/q49pXQVh7Ji1CFjPXoLqW
ZYP+qonbLfQrwB1YSwk9dRqpNZpnpjX+NQUt16Hr1hB6vVioDIevYL/kZ9R62Cf7TtHc585ay9Im
XeJnlOQPqvLPBjwv4Lfny5JVlvpsyUkQsEdfSQxeJh5+Qdq5CPPvm59RfstuQI3K75DdwtTh5yJ1
tg/uPtZJ7fQ/0gtHPDNBBPDpYmgWFlaU0r6E3ktNDxy10mves8G8dIEPg4JHYbsyl2xJneRj34g0
UHmPMU/SSqp/qmRZGF6/M7PYrWaQeXScmGG5I8dhxVHMH4/K+jrgYPaN42NIU+56IEbhB8MRGe2Q
R2fi0Gk78yzkDVjQHFtmr7Ira3AR3PBleBTJ2z5kxA8QVS2H+AARUmRaIYwTKEwmUgDx8DNrXB+7
K3qInYC4SYYxAYa3qpIT0JDZdjLi7K9ZL68IpL75gNJAZMW7edQONPrAx+Rnar05AF8fj3M7ny6N
d2fK2LjbHFU0FGCRHQSaZ+P+OGWHEvQHwQPbDeJPA/GSk9yoglKmvlUCghaVbHFUAQlo9R5bCC4O
LvCFjra2NjJPd9O2LAwXj+ED2NDWSdWO91iXYLqg4TKC+Z7bXJjMAvJwbrZfQa4GQ6obtYCqibyT
oRH5bIx9VUdBGAN7EVKMotRBHtNQpIgalIbFe8roPKuwrmBHEMmV0q+/mak8lmCMjXXJODsbrASt
I6839IHgqiJou9qf3S+SW5t7llCZ9UHvioZFyiu+wdRyHh4kHGyj5D8N0luDC51vm+gv1AgkHVK8
N/K2FyyXxwtNbmx70RcyvPKqKYDS1vPymil8QTUZUynZUk17fZ75oNeOWmZq71ORL0iAGWR3Zc0S
lvyat7yYzsqHGP/mzBgLTtwg5gw4fxDEgwUz/Wr9xqelhUEJ6fz1vMHeNNq0X/BfD5rbkNhfWVyP
ZlNTuuaia5EQEEsKnki9+y2g6koPvyfZQisdLHJQzJiaM0xGxgBpHc+sICGBnUahggDv9UM6zj4t
JejfJiI5CrSbCUn6Oj3YRlz7H3mEGTlUZm2Xl6oS7YjGRNdL9IkFtRM9w+GcObhLKJadfG5Bk2hv
mM9d8My6/tCEPd8jZUjQH5xWjvptmlwabs+9drh8ImArZgTJya95643NT6UTBnQ4vIaQlWQoeZ+7
nF0oOGiqciboOAuVDp//oKLZyKh6ZytKyz/sS3e7D+Rju3oUMzQeuGci8UwRcU1W9qvVsprtS2Bj
dvdRy5SzXdkvr6peO1fIoBH2pDsA4qcbwa8cyDbsWmGuMjNkpZxzNrE9On7I1DRj7rccc9FDkXUt
G9+IrVKLgkZySnSs0RJflU6arac+ne1sfgutO0SbCaddvldfYruTsDlEERXJYgVyoTrHv1aZjG1r
vnCNNxz5nyGsi4TATIxwKy5IsWCdRbzZtdgQa4NqaBPjfTPGJq0KAJp4owYCPNs+iTrY/9AD/xfj
8LqlVf890DzELnjS5vCCrUFqc5lZ5hwH3Gm50f2QJMq15fcJkuwmGjNyKUibI4up49StfKvpBuw3
3gZ9wF7LQUty3Hn8/ubVf/uwD60NczMKLVUm5vlra6d7XNBTiFoCIuWh3/pqjQBud3L6Rew4P4yf
R3G5V5i6MCXAFtFWibW8ri7PspwAZdqU6GQ7c8yivDlaq7uKUj5nVrMLiyVbOxzPuTVgDCjxnJF1
mXjHSdFG1swWuxOS/bmNw79Bip3ENXGRFoJDg8op+nazH1EjstoxjyFAAAXf5QzLNFqdilKH+RxQ
tJbgfwG6MkNWpXn0SNPRQW+5SOiJwo3823FcZnzppNLOzMBotGMzrODd0whTtoFLdhPH2VHKYi9U
a/j9BFbQPpliJE2mfKesQ9+cTheaDAjl8kCtAIyqUToLw6jFrCLa97b6eip2+lzOFwQr/QQebp7l
nhDqVqd/XBMUwpXjSHg5joNyXEO6fHazA2qzCTWkqUvv9bc0vA0nc0DlbjSDCf5QqAoqmmm5CgCc
BWsTax+40o1yWUNpnSejPGYuUAlzdiVtkUgBMWZBSBa8MqvH80CZots1Y66Br0DTat2mNcF3QUyM
nWijoLXAxRNlUTNp7B4YzAkr6wGKO61CY/CPkU12NBcU8gsdNUX+mo+bCap/M+KIMG645/3oXAdB
oQrbrCo0A+lYNEzolMmDZoN247A+nsvjl/VWRbjXciVrW/WruVMl/Et6N2x2z3XmETs4O1nxAbKs
aawsfxVt6U73aq2xYrmRelUXwU9JN7Sr4Ip9hOJMnNY+7DmVZU9fXRHQ3qLC3wOB5mW2M7JNnl6u
oujvAfo/19CmxQPERltvtYhpCGigW+nvXD3ILtHi+k4WUU10ST7Pv8IeloOfU7lNSoKHiGSMry3M
hd+DLBC8gzhNRQz1j6rdPrpap+brvD4e6N2HLBsTuNv6G8PnRQXOGoQOD/Ax33tPsV9Hhp3Di+jm
vKWnwHiaRoap7JG1qvz2b2PuNG9BLaCBxKhppQjcdf1NW1/qXyWrGxArM25VCbUyoOWT0gLitSGX
ewDzt0Q4lQ419XfTfWHE+l3QlAmU8yPh//WeaCgYLpA4O1DiETCxKdCVTMDku0r+1MB8RhI1CRa6
fmhUYqwm30B/Yj6qKwSl+uQtIv8RmaOjvg+QgTxEvNrMAHjEbv5GPXIhflMCHaU/zPrTBlU5evcZ
hOVogNH6Xu81C0FdrMSP0xqzhFxlhFGTh/v7K1cpq8f86LRKGTHIDAWlZXkDyxXXnMxi76G64dH2
I9lM5eNHZ0u627YauTc6A0AXK93a8kO8J9jbt0fjk5OweLjZbv5bohH4QUqRjjWphovJ3zQbh8Mr
U3PSU86kk41lOhmMs4feuN0Bt3CbvbxNJclNbDKcYmA9gTBr+4r7jvLYyBG8yVcwKr2vosUdfgFI
2rfieLa5rFX4c9EqAZQyPYmAf4zGB55j0xZcpbKluI8kmKw5bEmQ/egJndPHF2YAxe/ZW/hLnLhn
+wDycnYJRRJ1soDwt81VqCJZg4vRmupRZndtqedSYLbvli/2mQiudW1/UlCP8ox31BgUocsrJ/+4
226T/h3x2SwSpxJSmxMeDDd4xIPxDqK8nVyDe41S034HN5VxA6rwQ7e40cULbdGFE8TdHawSuRBf
PFlKzBGA2j/0iPbQoiySpqmMSDfclc5Kvew37DANK9jTKr7yL9vSEXRMmg5AbuhhQNgNDotj5hC4
QN9s2zSgL/DTLBrLD3dLZofAPyIa/LAvghF1vTtpsEsaNJtjpO6/HEsZ2Zp6t0bBScP80PAYS2Ch
qmqXy61USzUSi+OQ9iouQAo6HVMEKqvzVN5GByifJsWUKiitQzOZafGLg1F2vcEKfcCyxCSZMXL6
cKp8IMTINrKVD7SvGesOKXZaRTWd1Xtcha+e5iEgyj9AfKUBnvUDjWmN4eZv6AW8fkyzfGStkjOQ
LRjcEOheA4xrEZRMmjgMjWntxyXEr0psp+KY6sYg9+nBYzcSHX7K7x9/nj1JKrZvYQmp1HNeqMvg
mzHoenBdb6tD2HbPhkLVa/m7knHqknYrUuhD6c0MVBrTnATWSQtDa1Jj+Y4DhMy6OzFydXNIFJs1
XjQPQnY9PnsFv7nTgHy4+IaATgjFkmrdqDsdF2nyBsXGPS9pqH7XAyi6uq8VlRTQtr4QYtZxdU+H
zoDRH8AzYLmn+Fe9DLKr6FyZB1gDi6JcAamegrT4ADE+5LpXcExydJVW0p5fwY13K+O2CZRMn2CU
ktcj3tEvS19zdmWgSCwJdfgy++K/QeiyQRS5YEyXLGNClM7U/DspdCPWWJQE/wP6tri+BYPTGgmO
kqrUfSC0hFGZCyU4cK4oCE7EvfGzl+1MWLwhPsQ5ytvrKboznTtE3e1Q79jr6jfnP62uzor488SS
WAUWqZQNWnFhK+Vvm4BHez1FdotSLft1hQkM3MxF9kB3Ry1ut0Um3slqfVHYsQtL0tFUXDjCcLKG
xCwLZu2jrJeD9VFbOgTB/rlvTgABEACdKBc/kIYmiu+AFuK2XdpdoZrUxgTNKQ9HUX0sV+QmTLWD
DeQ89ZUAUjScxlscI9JWqmEupBcqh+vqYK88F1RJeXRAOFdbMXbPg+MphR9XvqJ8XvueFhiD8cz/
qEQNxhc5ZB26OGPl8fCRuIFs+4xjCXcW5Kbbh+ie8q+omNFBWnpp7Ng8QdaiCs1wYDJQYGyWIsVd
FbtzjNkdreN6HrzhxGNUSNSCGUZuDHvFlQXmjsL2kPxTD5pJMRdMyjMEtXGGw6DsNkRIbQDHYMv3
FbDH0Zm8XyZ8FsO7OP9i1hmyGhz35jzTF3vU7EyVXhI0hze5QBkDMnsDujYWbT0LtiNm88CkObFc
ha1qfA9Uvydiii5Gk68aYyy2R4/yZgnSQ35IOpw2M6vVK+tW9b38EwHkGDZadHocT8Ui3FDbup1e
Z1maboVgHqKj8j8Sa16hYI74PL9+poNKnUqopW84WFYHC+EM4GYhGgUbikTj5arfOgeiuBjWnWPm
0FvtiyIy1gSJf+WJLDYHEMI8HaHzxLZHxQAyS+o8WRjPYsGbaTLRE8H0E8EF/Zsi1YnMpvDVD0l8
td2U3SAoEdKmoGaJSuR4NWOWNd5CGdflTt/GLMERcyUBTy7Arw3EIAMk75XpB3iHzRnD4f4UT+JM
/FzaeSQdET+qQl3P1vnA6nLI/mAtHX2CWa2rnoswqidqubUpKqgpDNDRxHa7Qq4VqXWA4uN6zwh7
dvDu6vgrZHYspmKFiliaU/OPlc8jN2tiaYrO1kKL/HBPLsz20AcLmgjpx6EEimDhbGOkPgEIOLkt
0CWvMatSUs2AnSTws7lCLGHvmbSmKNCZ8waElP4e8yIQZsEe41HgEpSlb+b9GRCvSFEdVWSW3v+p
htujkAZ0ph3hpqRkgS9f6BNBpYUbjNUUTCrytP1MCHeU31bPszh7LAwhGQuqVPs+DQ3IexIORamR
u2DRn7cv0NrBpdPbIugrJjlPJOhjfp8IuaVbYrAKqKtJa/1ajDrZwkqgmFLuUaCUo2W9pfNrCD0L
mIS/xdOF3ieFCyXDGRGcDfjn7AS2BIxaeqxn1TOkAu+yyuBM2pJ7o99roANzuCqec7aKMsOE19lM
KE3XjQSbTO5KuLmWn/OdFDYD745qnxMmxA9mFQAxPKidwu30Dji06OONELFOrQMq/gIk2b3nZulC
t/UgwLXeVlKR3QGdrwtfXSTt/h9dETyFzMzYkFpoa7ojPF3O9Ndy2d6BEot+TNDD+fD6PzkeWsvQ
tRj+X+VwKCAM1XsWZp1weiB19dUNMgZn6NTJ3WV8pPc4mDg+F+MESHlK0GtNGqqPoLKKl6YhIttF
CKNTiI79ypfZghDM4+Ply1WJw6DQc1YeLSXpYljBp4KXacExLlARSc+pb4/cMwTY8EcXwZoKsept
L1dGFYNw0MQP7LkhpCHC7MpbQ1qkiHJoCCpHvgZHMnf/KaPnJ0jiSAuo5yQBhtfltZxmUwu4UNGO
JBMrVyLlInrgUfiRN9GBQuum/mlq/QXkwHipvefWVkRYF5MZLM3J0qH3q8zZwA2+xN12/gYsu9Aa
0Iy5DN1kPgfBMXiFzIhXYH/dLusgz3/Ksu00Vx2cV73QhMPCwKt/pVDtbE+7UQt3h4YHD/A+35Qv
OZVvnBHgdkcnbquoV0EVII/HdhNOnhyhwsYjcod+ucm1J7qV1mZihQPp6YQLO/WbCuaI5bXytxXF
VgNdHG9z2eNqVVGD+a1QnNPbduX9ZTS0pXx0RX25+yWkQ/CTvP4QYCnTu4AY1CzqFwTd1DES8/1J
d6g1KyXA5wSnYyyCu8YakXt6oQguKt19hnKP39LxnKnnaZOnicidLzNd5Xy4jvXOagITu/RAgSG0
zODtM3t4n0QQfxvCZ/Ug6IflE085GNKcnzpotcbarBth5+c660aUMnmvUVtS5OH4/DWyYdaB+GD5
RDNR5o0l9sH+03Su5wPBTfutM/VA3qEE4nlwcUkRL/OQpCYgWt47QSFH+gVyuuL9F7w4icye19pj
w4aSbqaJhRmhHv0uXgpZj4Lfi5Q5Ebh5bAPamM5sGvyoEe095J+5gdAGmWfhgycO50+SP95yEEYM
96WTS9OleYUnrOEk4ZSgpTdzGKMtZOYtClsseTUkh8hoDE3L/iwthR6YPbWcLZhU7TLBDhaRlnEn
6OQG1aXjT9H0QR/AArJBLA6319Rtf+CWXq49lRcxgQj6Wg66DGPsuAmiMkpxDYFqOkHqLbucnQn4
4Ejysc0ZyGJtC6+b8BcABYXxXOZ4cZW99db2UP+xL12O6K3zEwFdAvl7nCAGT9ZHbtCXX5h1Mwjo
oU5e5quWIUxSyP6coXkGGJ38tdeUeSRk8ON2Ma/+S7NZBOEi4hV58C5HP9YeWWKLoxKsfQiwpwFX
dN8XP2/NKuN00nR4R1dTW297QCET5JY5Q3vcYeN82bUn9lvf5jJXCG3wwJAdR40fDMQCfXxWVzV4
9bXRjTD7IMqKgvP4rOwCB1WBGaqDLAoUO3cO/QkYDGrHgD+kkR8VcHbEGQjdeimqM4IM+8b0N14y
VurANS4kD4XyYpQRp+eud6OdErC+GT1gEjPaLz3jeKGt0bIn80OfWp3zrlCjgAqkFBMCTC8ymXBg
InX0GM4Kwm7Jh1WLMubEegGWa461tX4qvurWCs0rXLyz/zxCyVvfQoFwpgIHxsdFbHrMcRyW/t6M
ZLq53TyCkLYfRI8FXGOQYfZgbPNqU8btgheKyEq4XVQmG6vS/Z2g5rBtJhqXaCTUl/l6Kti1INZD
jRLgOaIHd+SX45+1COgFmP4TKudIX+VoN90SmEnmln48Yco/RDAdSoO0XPdUKL0LHFblpm5Sl68j
hOpYX2hd6jjfyJ28wnq65IPf/dWuOS0lruSpxwCKOY2OQFoOBDbtPFDZbbkjfM5dZkOndYwyxhBW
njh3NoyVr9qWWC1tJyZDSvaVQcX1/rpDoycBfCjn+Rs/rH6sA+gUk2mqxaLFXYJXT3dQwKbSYiav
L/7qGKpDlUkhXcZs9Y1jljj2tkxIY2pg7GZUNKzdjlHDUhfgCr+UQyJqVH/nNfmC+O5kNYPwI5Rh
lydQudUI79S1VX/NRbPpapkuwnDP2mmoHXI3kmKt+YK01FAXNWnHRL+KWuvB+tG+C6B1bJ/cuboZ
+Eo+L21Zz6UFV07ZWsyL0fc+Jm3dgTbOiH6q+P6lWNB04YwUZ7bn0OF2GlX+PW/YaYaHHne/BkSy
53tYDfsPzFOgUTC/Ee2muERzk8/gAI/VyeofGjDa+B1qmXat9oWZ4wghRiFXAJcmqoTwEIVmimbk
k+gwBeCjagWEVz2uNsV7SK2yNACaBXfsFBURMHWpoUolyOyPHn0ACprzKRSky8eLOX1qcaHE05bN
4DsR2TN1V+RUbej7XZCWbRQioXrZTGb+hWbMYxRFCOiXHHOpy3E3eL1aYLnU6uKit63Ec9MEjtAK
PU0uBXQzS7WJvkWbbFCe9aqxL9inSYYZDVQB4ga0InEz1j5rdplgqYc3GWNi6HP48EqNknWPr+Uz
MS2hm/6Z/Mz0C8QmRM8kaEUA1edUf+M0Cn7u5xmGsolj/SVxDe654S6mqqRAguqUz4OSRga3Oiub
XAzMLFuSlXGhChQfB6bPxzpqObQR2BxIvan9wWpgpbDoz8hFCfm+N5mFQifysD+h3ZOYo/vBEZZl
BHT9/VJVdXwqAQWTK8fZytT/A/+pIwdIp3l22gaVfZVUjyZ+Cd7ZD5fzx+lAefme3QDR7SvmMuxZ
b6VXe70v4sONxQk8vEgv0ns7Z71im4NGaZTQg71ZgP1fzoVede20qAjFCIxXg0jwXdh5AlyC6q6W
xEvbTlac+sGW4n3xWBLncuUFiY+vB7cT5J8aD99BNjeV8Icj8uu5jn7d6WNPIPh8QFRr+JR9CgFB
roCJ3hr3loKqclt6hv67VFwtZvegq2giyI7DhDOzIqExuzZPKy/AsYpoMgKv9mD97rr3u99MiP+n
+0YoBpdpU0cbdyYvQ3W+AdKDTm+WWyDLQg8vX925eAOKz6Uuqh78ouWvYnIHLEXcDyYIIxA4eOos
SlFyjzvYu+VZeQ4+sPHdv/7nycUDlVKV+xxM62CRjM1qhJZPmyiPokt4x18zIyzbyJ1JCvlY9DcK
6bi1xPpvgj6gUEAmE2TzLWIPfDdyjDEjAlr+8F3haxsMvZswc/gqJwsDq3kd2TPvxxKEViyDfueK
QLJUau8aRMuZ/W3ZgpDNhpB3Uui/DC4mKknv4mqbOIBQCmC23bVTEVxZTZOj8cal8HmQ1aqxBXf0
wjlCpsHQvEP+a6w0hZD/sZJ918Ks4+37PknIlHN7Zgun9s91VP2w7KHnY3rnFZ8wuzF3IL2AKS8X
U7bRQIeWrKO8ZZxL0hRLGuS2C625Orv3M/UHSlS1yXPJWW1PVbqM3GPFrzV+3JXTM9RMz9DhXPv+
8Xq+kGlHztJnJBoK9HpDdFjDDLXHkaxRRc/rpDg7U66w33VTJPrqDO5nuvrxIOj3bIg6P8Mytbv1
lN4PjiDSuRE4Xe5W7RLOT7aSXtcnKuQ+6N06oDFufoYQ0H9es2KzR6HMiTtTgVzh6W405FPPzHp3
TqqAw5eMCaa7a8njDbsbL+JySsV6Xkxie2GWpi8hf5Wm8fWtMOvam0L6Uy+++u2ZAP234MAoJ9J/
rLrWGr3Hqw6ZKM71l2GctidAgL5phPix+i5DXZDPpbpgLn0GYFcjJImIwg7560HiqZPUR9Fj0i4q
dNs/9ZPBFlQKlh05vuq2S7KvwYTCeEN9DIO7FCBBdO3hkhqyW1sLCkY3mdKwyNJpAW38rx0Pe9bd
tqZzphMyBOD1xw4c993ia3r3wvAYAra8thKsd03h0cSRkCqD9XNRZp2oM6Wngt+DSF/nwKVc/ZJL
NsehKaMD4g3jkjX7DJ2lAKATkzKleIRWnZ/gIHevLXonMnmPkggYOAnNXwnHQr1A87hf6Zc95Foz
7VR4WvSsKYfH3OhgnEYdV2jJXMbSk3gl3lFfOgy/BG5uV3GlusNqymxgK4cNoLJhGbEBbGbtO55y
YQ8xhAny1cjoMi/7V3cJgEPGP4CcUx0eMrdBALZGMyn1RzY9z9ViqCn2JisY2RO8CLccPP8hMMtb
Kj6OxyBUihW3QvFUsb2uYD8ukFDYri6zhHOLdlRUQ5h53OsybQQ0vTRbXJZVqo4054yC+7XLIKRZ
704FeP3IsnWSGD+Z9cb5ZWtKDlSSgJiBXiH2zjfL0tak+HMWxQruBjyqmwK9Ok0u1Lv2G1yRuAg+
emyxFkPPxhTZPq67khcOXUW8KIoOlcBZzeA8Dmar7GdYsd+uX/8G3FG0bcGZ7jqh4FVJa9uuJ7zb
zagK/csqRSfoCnZ3KkWGNlsHRnUyhlfcQDamdpz5V+nRHZ5C4ii3YTOYOMki+VEiQfbWKTseGbRu
4i83iI1tvQe3mPW5d32GK8ac6UMDAkakbNJ8ptaMzHSXeU5+PRQcHEWkWfyalu94xcAG8Gi+P1Fp
Inz/xgR7aRkp2Lk/5ESK8kkOM4R3ugqFexHTofQOJPThVmi8fxWyyozpM5ndmjNdf1lsGJv/B9gy
LwYPdoA5kbEdgoroh9iJ4y7fIHOL+hMEJX78ntfo0gVaxAxWYG2W3lJhCbgVwTYl+6vpJEL77l4g
e6OjuhoNPl5Uu3ZU2P4k0rIKKHdLJjwjyQc5BBtgZ4kqaQg9sD9hrZ/t10OoKv0GkuYEy5PGyaZm
P9QCMXjAN9Fh9vqbN90JMtDAuFc+OaUs/XQr8MxtOQHa9Rxd8rVYxTf7YEA+Jxt3hjUCb7uEvsiD
ElpRWJ3XGqnnPbMeOIwrw/YcLyZvsAjBlaTisO7VVUuWHienDwkyQoEW+V234Y4y+CNIgnCO3514
BCMzyMhfIbgbKvhrkf+x+akf4CmKd93Agn6THrOyyVEwj9zXWhyHn2kxOfzOgUcpPat6T+D64up7
k6AROGqZCSCuR/xr1llr7SFGeHrgtCv4Vx5y5rdy5ySBCM2Ro0kgFe/VpBC2dESzrJguC7B8ZaVt
Uy4oeGW7OeZFRsoGLrMfFSTeXLaYqtbFsEtwz1p412udmvFe78X/YVZaeBM2oHF/agCa7CYiC4X9
0iHlJ24QUiD2sSdlMfZamYyUrJ6ItJe0M2dqNcEhcz2M6ufFj3y7kkn1R4JzpE9nBG5/zQJmn+9B
HHDssvuWSoL2nPOrgy/99nX/0cIonaakoWbm95V8Yp9nYHrel5DMM/cP14vD+UkIFO0xAfvZpcaj
MhivigzDyZ6NbYGyIgbnoSdDyro16U6+SaAeMLVNlV/gg51DI7MJi8/gbj45RqOrfSCbdOkY5D+I
vXAvES/xq56jDTOcJEggsBHl9Mqt5meTrbjIZJBMz21Wsv19Fk8kvexxDnH4NnT2IRi+9bIjbXRl
kCY0Lpa2pf324QPMz6fcIpEUo2e8W7KeiXWIQZfZtDfuHVgjhdaw9abWt4F+Li7/IBwszz+J45HP
RTPP8wv2wPAbsNSaFVTT41j4koWHxsncUHYO89dpdagzxvIpXrzf6boKJZzzNM7sfEQksyNVfcBb
revQ8REqZXbakUbIuhKAL6wSgBM3luYT8S31XD3puRs07ah5AawT3e1jL+Ydus23Ul//cF7g1ax6
5StjStlGbMAPRZsixon1vswK0zzfFJJP6gt3tKvPLRotTaMSAAWGS6VJ5Nrcj0/d4WYRleeOWRdd
n6/DadvxSkCZD0BS/sTKXtCNZo+SP/F5nJYWTXtISSsBMDQYrZoQLzexImBIY4piMiCWVFVJtaic
qBeMEHsX2wWvITqTIo9KPWFOk5LqSg9ZiwcMAP4aeA5ICOyNUJ42xmRC43eu4w2RXMBtoWnYBh8L
MSpHj85iR7FUVrNqkd71egisVNFLvHjRUV/Dh0UoxhXbN+tb9IHv3N0dg/bRRig1weL4AWVPG39x
ytsVDLn3ucxvlsn92+UeEIgxAIDDIgteYty8fe4BQBByUXPE2OgeocS3O1L5ckzjDWPtgdv+KBdp
xblhzPZEq8Asth/DfFPOtRl3+dkm7GnrSEKcEpzM0J2khc2qOLFl/LpzPW53ARpbXzHQrQTKiS1n
gyRoT2cpM+nEgXDuCXu73JEmmioZ6kUtoC8EwPgrzt+9mdIQwa6bjaN0uyPklZs6ZpvroxZmEEmK
kzgX1CQuEgOjEikEsCtm/0iSuq5f51BrNED3+CCf/9IJawCmNk9kuWMYHHmtEDjjxKLxMae65gwa
hjhqmV2nXTEJlHWF7S3i0aVH62xwYtUCqjYzgdBDNtCasFF6T9LmPjhNxD1ttJoHtKQZIkwaNcrl
pfc66b6XH/+H4QCK//z4nU7w2d4Fq7ypTsBAw+nudfg7HX/2IssI0Ywgbc6G+c8HB2ItDOcs0BbQ
2spwGnCePgBrP6BQzJjnXAYh5QfN/+1cY2C6PNtkKPTrc2kpzs6Alx80unqeEWnV7vmhnrAXuUyH
Tb71rl5OIFnTi/kUxlN/MzCaYKi3Kw8d+LpfknWrWuPuvpUXK7kHO85kWuo+6dyI3E1J0u3UdV0B
22m8l7TbxekGdUkXSsfBnL+zii6XZ/qLz1EWfDI8rq/PmEe1WifQYZPkaRVTzfnbY0n+ukLwb+a9
eKZQme5renJY0/VVBPjWKym8I4n9WC2r057eTaveDi6i43+SKRlHTTG583yLXUFxjgjHPjqk62Ye
fVv+O7JM3b6h0ybkbpCYvZiXcWNjBBsWdK3oFG7NTkvENtQck1aPoYlO+BPa2wfRz3BiBoYpl+kn
BcDXHbnItMLgGsnHdnnuxw6faZW+bpgQX1xeU0cmc/wbVfKk602ap/I+5xQhxIGnLu1Ih0USH5hp
Bljh3QZXpHRkKf/ro44b5ad14QnxG3AU9AxoBaUdQGLvs9/pa6XuG7vU5752DJl+LBhvaVkvugFp
Nj7WDjSJwlB+3o4kilcd4X8/xf9+yW0Mq4yJwQ6hL6Ih8kRpeWlrN9HfwA4bzqyL/Fy+zm2Dxide
BNJgtERAwVqLfePVHH/7ae6n2DY3B4OEEFmBibQPPFNlAYN6t+T7UH7/q2c/9srQ/Pj1SJElPYDi
AoI5Zs0dxPnJ4NLkO2P63O3J0LtFtxbm9Z1xgtDzF4QtbGHNW3PONqH9rwF/GQynojI1HeehzHSX
5/FZMr7PLD1oavi6EBAZpDGQdeRF6UulW6it7A0Gpiw1ufTZP8YTftzicrDn8iIioW0WGlHZZzlM
P7Lf/LLCHjmunkW0AblQR7q2LAiSuqtjV2OXhZxfyIHcyoCW0Kir7+peQdiNuVCvdvQ7Zcs/ChB3
T82/4b22gC8BNx7nJtW+oqgCRD6y8x8z7N1DTrBx8LmyzpXMJ6VXPmW4H5yHdGxApI/dYRz9Pjj0
AZDzWnaq/2rkPA/juXZeLvVdw/8WlN05hosqQq4pdYrR5SYUII5lbzsEONZYgWQ1303Yv43CpKDW
gjWZWC1N/IGUPdk+CPf9p/5RjzGZ9CnQF116A6yw58Xst2gvk6uIDnECsJw/vbmtIH1iKA2JKoya
IEOOpZJvuHjlEtMR5Tj3/RVIUVI359PSSHKWw+60uXWFsZiMGAiUVYUcfFOBmHd5UcInR3h0yycv
Xai971Br2YJ6l9aaqabShs0C9n/l1P6mbtmD0KAbFi/jGL3hFW99LyFMsC1xSNZIerc595dzIcfn
w8YKOhgbDN1BAeb2PVmFbjJW/dvHYIP7VvcC0U12LRtixJUdhd3XdxMxE4pKxKzEE8W1PwzVfqfw
DL2js6mIbmD/Zy8nHNrfIzykwF61kWaWHik1qaGG/RJysT+Daoy/S1ENDdBRhPrumz/nLsJoELGH
bU3gjF5FeGMsJj+4HZ8jpVBPffO2jVeYgh7yd79tNmum1qvre4LWjmSfqTRPIqomJ+CBsd/OXQ/+
9JmXeCV/8TzJA1EYireSXlVIlh8DagFlXMbNtX79efkY15olXfRuB664DFcC0xmFr5duWW5aIBb5
AmprWdQA2xUj+7yZb9lw9vi6L2CSHLxeGGJbWnCs836r0nmgCNwVyP0S9VtzjJxCPRpqx50YS8eQ
/xx9CjPTUdSQwNPDbrRe+l9wMCpKWstFO4dAPlbi6iK0eCOWhyynqdJrC+JpnYfMJXawRlX6cgp3
oJcAZZDcnnNLvM4qUU9X2x9csBz60x9KXVnLDxVqEFb2kk3BvhDegfX68gc0buF0LyfE6g0u+fuU
R70A6VdadClhKGR6Tt/LCNGvWbOab3A2gazWE4vC6+Ldy9qE1yqrxb9bb6sh0eMRmc6Bm17DZKv6
vz9eOjY65zQc9tze3my24Msie77ezwxfr14A8X5jIIC09uWHs3Sztko8Syus1W+Cw0cALhYL9IA/
a0Kzcz0IeZPVZZYzXDigLeBMvG23GDiDWYqCpnnoOHd7tw0/VNZuIi4/F1k3dM/fJx9JKv2z7txu
B0uiPNY8JpGzkx/S/qjIrsQUQz9O+Nql76N21Tecn7lUrJNMHZhV4nCrfZSd67x7uGz1TIx9q/79
CRILi+dF66oIKmIDP8Cg+2mIGBO3/HPvaUL/x7E4Uydneviu41EgFTJOWGPPtmbS3YV9+VVgBrLq
etwuyri71ymLGkY6LdThXkPqhcgyKDNr376Ld3a+BkpKMB2uQIu97POjpUxTWioZ+UXs7YHPH9dA
KykmPliw0AHxEB6JpbnhW7+Uck04GbVAxRIDAXuh/r0MuYctVVzL7kMha3xZvhOzMcjUzdn8EDqU
Mv/WeUP9A9L/V33V1HoRY8huyk+PPNe98cjeejN01C1Bg/bOM0KWst2Q8v8mCHYrRDjJf/9XxkAs
whwgxjESnDAcdeCM/LW9Sshf6TH2/nph6tTNI4FDVHYdRFH9kSPusaJgpx+P0V7hzcOAE2LNm7ea
1kLzNv9DVis2QAAYPOKgAo3Bpo/eG3TW76Epjx5m62KjevUHt5c7o2sjgKVq5MFKKMlGs6vWAOXH
WaJCfXQDRGoM/jSF7ucUhA81sDRzPUls5Yi41f12ZfIPbmgTuZoRvrq7SOmMonlp7OwdGjxTKd5V
r2eFaeZVGzICXYGqkIblOPZBVdCjWc+6nRKkokYJRhk+L13rJPczkTaQ3qnMcXbAjSE+mjf4r+Jv
abSzUPhqHEGUBzI4EJpjTrJfT8f75Ah4MEUHouGltv7kCTiY+Efpa1z6I60w7ySGGj5e9ytbX9AH
j2ciMwL+KXq/ysBAYslScsxxt9g0ZwyvzfaJ4WkjYLmVRq1P2cFLB5QIWleftBsA2SExqqDrNCnI
QP4jtnDeKqSVBqxAJXE/KLxns3TsgtCj6jVHLSns61o21wwPpL2QiYFOuq9i9UP1aMy5ntsH0pqK
OF2AeFHpwdZmPP15iOLQljlHVDdfAbDdfNTwl1gmIM6HoRdXPsDoGPZO3N8QN6PalqZGB1QVrwjX
3Cwvpr1Wvtsc5MZlfTEe/GDR9ued9M6IMn+TySPJN94gpbRLcrZ4heWOikgOQ87y+EKm2clfoNcr
Z9EEDHu4THN30uB0V1iHSloAuNKpcpWLQ+duED9BYmhuflRjV3YzjJPDcJU93koauAYi487Ka3A1
fLilc5VYHI5yvYG58OMalpXAtq42oRcyIb/Emi8kDGAEqDp70sDUjm8lZlVR2uv/wBavo31Qaihc
lkXeEyvezLyMFqeWe6bsHL2USzFsH6UxT+U34ILVydB2N7eUQeivX7hCg8JjsXL/T2wpmg+Od+j5
5+YuP1bybjSSLNMecb6ltk8yMhBr54xt4X2mIC4iM6NoXVAgVfY3g0KpDHhu3rr9RMHG9WSmV0es
ha2dOj5VW08w0jEX88EPZk+quaVkJpOO7o7OB6yOWeN53smlua76wP5BbgYVZVa6JSDZlgr7wZNA
Bc3QtfMKTZGsMWsZtB0Mdr+Vx48bZDK+rzBxXQkgVigzUxjZfVK792ubtUcv+TrPCzf14aWKM1LH
1actHLdskWMfD7TgAcmmZG+iCoBQ5743ACXR9KMbXEUflpitfhnR5+8JiLp4L31haNUmNPWCPRoc
Jc/fL4/RJmVaAjzto0uEC31X5Yjyqxsa6yY6MmspywE5zpxAX4w2DgSNv23sQH33p3BGOmH5MxE5
n4MN5Kb/EF9Jf4G5TGg0Yb6tEtm62/3qbOITN7TVouvChRu3V9jmUDCMLrPH7cNuyW5iTFmElvrh
6/8pjcJlkR0aB85+h9i6E/vpE7XgNl6a7SZD14BkucVgvkBQhj8juWzlw1LU8XAodml1I9F/1B+d
Zf3974rjYLG42L/x16y9TdzI2c7owW+E3emrVFt4qgc/zYoAZZqm/+76vir84q7TwYmsG9rF6AuW
r49v1/ix7svrJT3AOrp+rF6barTSeXHHIZB5GFMHs4RtXzyeiQQiMsoccBZDwWIP4x/fAVluOEZf
z2yLqK+Od5jseHsOIeOyIMaowzvOYFqMhBacroChPCen3oBwFM4t57+gJImDdrMfJFBMisiP6vji
rVN26dEmzJsfI94nQhK+pq9x/vv3oxB1OqJeWjU5K9v6IPqNw4AexAyl3++XnJ8FWtbAqJlN6lwW
x79XeMm/jkLOKTG0QAFIWzUSqJm0rLIjhRhXdVihvVLecZ83r37I/+lT7wPIbh/X4QE5zaMNT7qk
Aq0mnGF1fSXnMTzE85TzhhxqEp62k3IEE9Soer7x3R4ZJcM2vszaUEz4f7PGJleVv618WToeY3oZ
I5YRVAZUxkfg5hcA49dba9Fn2aCfzBOHr+MLnvrcGiii5hqiZxnv9YS56LR7AjGoWO7qH5cQPN/q
Qo1TCjXGAgAKWvLXZUhBf1ELNJiKIn5u/LB2QCshKMjC0oBNvGIvNSqbZsyOZxxlqWif37So5EmE
pws2sOsnvFFvYqtgZIVve6JUQURzdVf/Bk3hZDhef16OxJh+er5qdlxpk+12HLg4m3aeLokAlA0C
5cscqOgxWXLeD1HIiUCOD08njJ1AOB1SVi8M1BTRNn9LCQ8ibD2fDdGpDs7AlxF0Zr0fygHV/hzY
nPgrOA+vVzmS0oRi9eLrgK5LFtbwyFupjHE6Kxpi7BJJlHuL63fCIwaBM9HsA6sYhzij5ZumINmo
HYSqfovxbpA8FmJh6TCvCifW0EBaUp4Hi6y4LWIMBIZCgWIVyBF/0GZOMqgIoYprI70x+Mr9yT8S
mQHpbSK+fJfvnQ+eimizqv5ztJLJD0wsWii6nQpvXAz/NqlsKACJagpgxmT1756jO06/GRai+otL
1qNn3ubMjoi1kko5Aa5zUCCIHEr42FR6r0D3gWp6/1AaRnggft5K13Cd2C6LmCNHEWbcrP9yiHjS
GnG6cK/dh1PyvYoLszv83ZItq9bnFYMzutF9T5x+TUUknGec5Yjl9OLHCP5QrOy1vAQu7ojr7C7J
ojz2wMA7Nl7JQN5tgZIEtr1aZM2760QiPhOGfe7hPYHw9rplfpNXfidui8bm7CnRqSsvymyPfCXf
7qoRPzQW6WbiPbPXvbSOmlaY7mXYT1nvEBozE1KU8cIRyMbLyfHkGlf0lKTwrF6A822oKofjn5g1
RAS2ItVmvfOMJfBkt3VDAnko9HywHr0vWAYaJ0iyxK8MpGjGSIAwpWuosf81cHmj0BdAMjo7ZpzP
Ofqh1/4k/m/UOqI0kEDrnRlqKVDVy0xfRI5e4d0xIAxxtQ+61zSWUjsbAt7TzKRL3/mLL/jvTUfl
tNg9TXJ4hTxzopPqRpMJeDY9DGdnofTTw23cWlIBQYy8N2LvifTIGZq8N+4aYd0sHJ87ADoaTnFb
a4r+MeN6qj500pmEfSj22aPBQDLlwQEP8cRLp9fk/IIdo1ZmuQCasvmiXR2AqFI+fPQd/Bf/qAQl
aNeSO6xzmwSIyNNfFaJ1mo+Tq5czNqcPC9KtstwVyolVRkAZvL0cv11Bk+QUNeqiHwkxMGbdruhM
ugFZAjtXh976HD6XYVnojUFDAgzkF4HP3hQfprCxgzA4ay9jrWFm8gw0LgCiVAc2CrtXRD/dmzb8
3rojxaS+iZiZrTMayeMn4ar0HOXldYaCqUJU2xExnY/a4vr8PkLy0jOGbM6RmK+8JmDEbxXKvr1b
0mMg9ztLcm+oUIj9/tbtnQOpMGT26PSzajRQhjBDywbEDNiehm/yoaIvG2kjxwWHinE7cjjvAjtB
jVxM/bsogp0nAYmMJda1zOPaHne6yeyjYv0WFOzi1wex0orj5CjXWkNveXAC7YlAQnu47YBZpanp
D7/z0F1VxUGo65/tmcWfTFdI9QCELKvgodGpliQqQJeEejBWSj8MNfhAtMVRARbjMeg/xYnpl8p+
wxnfogVa5cdfWVh/0rS8tdvgAEd+7nyAQQydNh7RVetZT/In83Sjq2NvJrLG1r4zWbWgMhs1IPeI
mDq7NXVI4lGdbd1d1uFLmR/RUZumPjuAwenwOvqT68gXjLy/YesaVH6DziIW6fWzUqqh/6UE7rZg
gVQ9ApOWDdM6fKoYWvY3fmFfcQexz3FUU5L+R1+lRnM7O83Cmh59rqJW7Imvmrl7a3zPmZ08Q616
1NtvQH2Vo2IZnvrofAtoH62UoVTVCRSQaiWCxuEy7uZjpmkmYfxoZ2STtWR/vnNtMnZMhRtBzXol
ZQOAL+dlQ1rMsrwnuSNWndVA18a1sqFyAKsvm93+zXDPOP3ZC9MOnBg9qwfFap+0+LzxmsBocsQf
Q8Bqb9HoueYVQRcEmDB8V3HsuHRk33DU7kQD35bW/GqlDvKmjBpbUdkmAIn74NESzSsE0v9nue+m
3X5Rg84CIrtWFlHQ1HhJkXFLo8iIlH1eVui+ysNyCPsIBpumSSnT7kut7T42SsaWap6wFmZYDOyj
u70lNeYBUUDcdytPjjfbUpyOzL4WJq2+T2rWNQdJDRnyOMceumfQCUCfsDA4NbcB9Gw9Rc1yF97r
+INQHrHeklDW53TOn6qu9WSpi1OPbp36+0Hgf69QYNnHydCvH3E/k1famWaWcMd6pk+Aq8D1wI/z
W2FT7WA3OkzJJxiFvRIinu/r+82A5UrcV3xQaDTso/vt/zvdy4Yt2KLij0Jf7w6AnD4BZ9deToZL
Fo6eLJbG0ijn0oWjE3CxYMyhT7yNatbdStwhre/maoCbf/VF3fjYjkKfu+ZsD2B3p+HUC43OkKFe
iRrH5ug6qU+Pns9HDL/zKW83n/RXTzshZWbYhvMSOxCM/ZU/LlorfRvPakXm6+COkO6Be1PFD4FN
LYO1ZGZNMtcKQb9tNkDnrdMokDzi8IgXurKNYLKGs1/QWVYTchuHYudDb1xP32YMJo+OXQ5DEcoa
Ua3YMAk0CKtcb+ELhEg0HM/Ez+5AaLLc0MiAeFfan+1c/3N7WRHhfHbLp1Yoeguxmuoeo7Wxafo1
xWX17QhF1py5JU/v4Nk3WCYrM5frUWDgRQmrZfvd5eaW6djyyCGA0v6zWmEnk8Di5ei+pURqwVap
RFLSyXMrLdRdRbndRcew99TWSsAV357oBHREDduH2B+5YaoikBtMO3tXrDSU4Z0EHFS8yg3i5zIe
kbC6NNQfr7EAQ1hHyjMnfuPhh4ujoAKelzW+2KFg40vz3kkVOZICBE9DGBLtoiRrWY/7ak/y824g
lH+Qihxnh+YT/khDpifL3B9SOv4nYvjNI9C3YjdACQuiH47COhYbT7mRH11LnJ0ZiOQRTSBkuS37
ypkCaUAZcd50tUWXg7kNzwP3k88YgNe9m5fN6MXf0Ss/YKq9ZEOXJ6oZfrShcUtxn2f3Kz9rLTQe
uwEJxgZOTskKQfYf0WmAqeZxR0Lk3dZCiP1pdic6lDN6LPqEpYZm1MnaR+ci6XDYZ4siZd56kwZv
MQM90j3/224adktck3/jW3Xka7Agm9jGJ72cXDq7j8GoPrXxAtasHg0BsO4iJ4NOp14wacE/Ettd
MYvA90RGxw6lBOm7Fz66cS/dXYMLuKyN5WOKKRDPUqa2UG/jveRdH6hzXJ01G9ZGwAZzIql2ahNq
Gl+z71UUClwqqE6mag7b0OPcsEngof4YSEcsIdhe6HIGtooNZUN5NuzL0DOu1L7uo2IDxAQ8HNXl
SDzEYigwdxnaXqQ8l3kFnN2xdD24JZwP8yrI2qt4TteEnLDqy191jlSTumir/a17qh0xuSDIiXKK
/Uqe2NbyLTHmB7iVDQ9yy5BqEBoxY0r4gFPbVR6H1Eq1b9EWUSi+S2YHLZBt4OeVgU21VajBbjpu
8Bp9lzFpdtxpariNUWY0TVVqYKxYYsyqsHLGKYEM8fD39Ne20utlwFgeraI5rFqTzcBUedU8ebfQ
qGEUM8EenaTJG3IZ0pstP81mHUYgm9TrtVUH5H7kpEBtDTaB29FRRsyukC1joMUYEHGyTo+AK5xC
gfH+d6I5e4ZqF1EZZYEX86kGOgur4EhvXLBK+bmZf+P2LGRQJjxqZQC15cpMRP0UeiTMKo2NrRTV
JXKkt9HHwHS5JL+TsWdlNPm8fj/EpocKDtI8v2BctSPqCensV+gqR89lxHTEPIUuiZTzPuezdfyr
6NQnBIoZ1h99Qj6TPiP9dt9+q0VkU0HQ80G6G3KPG54NRvHWOMi0PrgFJNRaia7TMamsWHMi7PGH
mqV5Bd8lPrNwwxQs2O/xDBPRrgWJPh14UPeKLzNBhv7wk8egmyVq9yL4LwCbiO/GNU9DpoidPnxU
EMHP8aU64xuRRymguaB2TUnSoVMsx9qFaQWUVedSa1SRmPeGr/Lv2GiHse4TASTEr+9lw2vzdQB0
1A02ZijU+d7pw15l31r/EG5+1CdMBVQwve6Ca76LNTGHOvjX6ZAMa8jcrP6qKQTI0hLSAR1Fys3N
tQgYzR2dPmGRicz9Uz2Agb6DCTriIRfdgecJsI+eKLNroKxnM7lC1Qm1qOxNZfqP4/uhs/tuHX3a
eaFmR+Uk7AhywFIft2Lcf64f6KA5eZnQPY4cF9o0KydlNzWdNK7M7MReGHWOMRCg6j2YdWzB14z8
Z1mYqZIIlpojsxbVLTmkkZSeYyVj+X9YQwL7fLT/V6cZ/VJTm/2FEPzW/AZcb+8rFUTa2W39/PuM
IhX+9hVjsxvBkWbd8mgZjotWd7Kn7u8AA+mPyWOpmUkgGwXDcfZvEOgS/LvM9/4hJUdskB2TXETm
rTM/TKGiWMh3SRf3RcmjGVUmaWh9aefuc89B9NBWaXDElDXi3W309RlBnVQ8jJHlkIGbBahqI/36
yFC284XxfY43imU9rlcHzTh2fguXqoiXoVNKlbxG6VjOaM1jz3jG+q0PA2OshXG4T5QbKl8VteB3
3XEuqD3BHDAqDy8k4cDODnau8RlgFIY4NgRLivrUrldWR11ipL66McpncBi9wx8JOLSSDb0HJbZK
MVU2ErTMQUjYF1TLYH2SXGTY9AFjCsSHmPbuVOOXOn6mWsXgd+ePbCcDmj+zzHMIaIJb+BFrEyDq
tvTZci1KHBiPqJzGaCKePiQCWfb66ODnfNTI4NGgs5Hy/ZWqR6f+IpT6BvkiHC+7iYnSdF1aTygY
YCCszpkPoMMB9s86fUY3xawarjkiFM2qCZ/0PqJEcJojUnKB75TPv3252/v+NlaPaoy0JUl37a70
M3mpg0JkwvcR4nEpfkBez4+x9yBtPmjHg4fK2/f5RANGauMyMxQFtPIQouCVl0yW9a7YMXgo7tQr
9KljqAou+y6sf1ezfd713ymEZeC134HUrr6kW45vZE1eeHkAfLlwBcFkZng42lAltJ1aqpA3FWJw
AHUzm9fuqZcCP/JaeK6m94ETCkmeGkYht6lh0YsBaOcbAVwYA87lgDyIAOmjna/elGgAcZdHLAwr
jkfsUklAQefaFdGxS9fO4kE4JieHraRwdvs+MYmpaMXtxiK3iridgJ6AiG/6cJIWiOOha7/PGLDP
4UvV62SV3NqxQyXH0+IDhnuVJ84T8TFKOTeld/miy6Vgbu+O5SHMqJofoc9klvo5C+7tPppyyueX
7PPMYoJxpa6B3gkik9spfJMfU8aqqFj/ZWyWQuAJMGhiQh0SmAxwGK4Pb6ehuPJhNy0MdcEyzfyK
007YlX69/tqwArzWWtZ+RbUCBGrq0sPe2PS4Mrgi+PpCsRTw1NGzY70AuOpKBsGzxanlS/udyoZW
t/DWy8ojd/hqsHnbR+TThKVSuascf9sC+Y4pK2ypneV9LGrBlcTs6udn7LTc1snnVV2UOjInBGLa
oSnTjsBGqLRckNBE/0y5ku0FfUNd5S5dVTT51OtK+7lacN9kSipGfrEgna9TAXyvVSV1WVWGHAm1
0QUevjUNA6xfqLmlBDTYQHz1UVBzsp0/7CGZsbdEq1Fbjg4GS6cqXm4Gl3+kEAmEHQ0JFGqKdu9o
XZIr4h9AgG0TVSQ/AQMblcZjZMsVykuknFggfQnGKrn0Ia7plq+95MWe+Ta5ojpLYX9VPaUvc4jU
vhdxQrqCfXn5Q/wiX0IzUtCAb5oXTCNH17cwH7+dTwH60loL04CjVZe6ll2TDu9HmpCRTfs0eB2y
pDubYftx+TcuhsSXX9FAKpiTKo0vQXoJBsKh/P+ojCFYWypO3o2PDwa71mKsuzSp1vUS8zfN5Jpa
lwNl0LhDIegPrX9BU8hhroVL7umO9XkByzrmwNn0GI9LMH7bBxP6m5CpBPPxNUKV8JjsI+TGof1P
afcDdWk0DxTWVe9yQCd6wQGcu00diVtfrdkYfH0c6KlUWxqFl31mELAuNY/kccbDMbbGU/1LCjaX
1Wt/yXLC+R/UNGT6wL8mqzsxa8MIDWLb2Sj6HOCHT8VAlyIBiSTrWXsaynqvRmWGS/uY8kka1Gfg
ps4QIlD/Vpc8BTFW5Vx/NqfGbh22c+C793gHay5ZCgq5nJwiwW4EEeyhf8HqOGrXvdc7O/kLfkuE
s868/HHWtPjTJxXM5DEx7TbGUfjre1AmHJv0CTLfOsnPEsti2lkiQn5ykQvzn3syUK7i9lSWcXsY
3gqvmanaE9bm2n3Id0ru6qhjVm13RAOzOc8PsENC744ZQ9MXiK31mvMmO42IHYxFWoRwUXaxA7fh
YXtkcyE35kntrwUh3lYDODCSoItK7T+qpShu+IOjsFdFmmpBQTFPffiOKl7ucF2idStm5rFgQZHu
rIoI41TC6kbYzH2PyX1gVbbuW82Lz8yX23FIQLjlJ5n96jT6KuBvbeFOnvBuzqlnqYkgxC/ZDXE+
KQKkKdSgIM3K5goT7ONkyhlxMniF1ef2/Sw4wcSf7BFkj4goI/P/W3Z2xKpXSSDWhJkl1fIXBuVW
jyUW8V4LaHJxk3IzGLYiKwZTVgYO49a9+BnHPoBgdpvE8Ghq95fKqcOT8UeRkfM5pfBR5cPRbDgB
qQckWmY+GODlyR66oJwABfeNTtP69vyhRo/6lKYaVzmf01T6DcXm0Mq+3MVa7VWbLFTlhfBnkp4Q
RNBRpVeH3RuSzOHIS+OZQsj6djV5iaUmHsY2v00dNyfqpHiTHwlwwovdjLoi6CvA7sQGVNyVzEUS
gPjlTmgw6uK+RQQzdx8JdOz9MRuWdbh4FXj/HVL2sabHbRHAFSchdq3HvIgkNkexUsCwCya6go0o
r70fvPlE0ympuDGQ6hTH5eL6xbzXnHNOPrIxzOM56BuUwwOaZyXRR5isDHmJJfgCKdnbLZNqz2Nd
vVug1u5oPGmmk7htuPzSB/UG+LEHB/Q2ymUy8S8yeoFfprppN54a+2xls/9LX+v9RU8Y1ieXG+9e
NOO/iVQAkTJaxWwEBL/J1j+eJ6QYGoJFQ8UmglrzpnupARArdW2311smpduTPX8M/o9/1uol3wGv
oeSr/bVGqCYscJeFtPKPOKG5wIvVA+YxKw5D5ZaC63YmAL2hFkycrwtcpBleuwu//QgDWCFaxeKb
1PvEpY3J3IwAHLE/dwlVd+daUw1Ejz2nJ/e+LtoD2MGkengYszRrdHFENzFKX8WjijVaptqQkhE9
L+x6Ay5gyhNkBZiV+5LwQc8mVKmb2zwmxqB/VgPY4y0NkARIBaDotzPQal/NAuT8vRqvpXKDyaPt
vO/z/yaHyttkMoWlYRc1mMPrgCS6rKb+i5dE8OgMS6Aq1y2XBmebsWOMCr4lLKSTf87uGs/K1s3D
zk4neoMTiGfj6LNAVv1x1d1uUPVDZzkCGEbjC9AYnvsr+jloxrpClUTzZMt4YtAEWceTAOEAIjGE
8fNYHvuG4bLNu8dPzQmPpJF2eR+QVwXgCCzWrZ73Q2zteVJl9hozuw9aDakitHffOH7+6NEGv02k
YZNt3Vocb13AYEZ3Hn63VqUweONgK0wIQdlo07uKeks/iTufBUFrgh7Pdpj+qY1szuFWLWIlBR68
cgEnZlYkAE6+EyRyak4w6JZRxLm2sgBfctH4viki/80dQvGWAqrazuUgntpuyArVWMZfxuD/CoWi
BGnaiceeMh+byGVVZpmGsdlFrGCewxU0O7zeyRsA4+/VfNm/UQY/Qz6kEPFERR+5qZon6vXBKa6y
v+4Dbrp0sLUo2rPVsSRL+d1hKrwsp8SV5HzqoD3aD8HgDYuqQVMuPyrAqaElc1WMbI0br65ee/ZG
+5QvihGN7xkuid7EQr3XfXxlns0NwZ1xqoFupeG6W3KbniRe8cumDEpEvKmiXH2took+dTC2U/+g
bWR97mpOxoc8olEpKUfGQwoUQUG19RZPx/+FXR+yCz8ZBTr3yrIASZG+S3PJBpYG4sbLsW98ZAw0
Lxwx2HNTmGiyzrQUj8xawXPZ2Qp235jCeqrPNsiy+STpYNygFK+QJof0d5YenO0VTTFufkPXeanH
rJkuV2ig7MunkzGliwx4haMCwvTJBZ0gLEZy1wwUMEdLQzmFeEwKnHHRNSxgcTav5EW+6PZzwkC8
rx5+gM9gPH6CCRrIQyFKac4UIZVe9dppdGKqQjv9aBJQdjtC2hn8BlCj6vyPktEhCUim4IAxEvoJ
EootbzZncY7YcRH+hBieXMfdgM61Yp9dzjAn9Ua6R6IJPxDRzvqiBNDZmF1AGYg+Eay96AtGsypv
FUDLjJITDMzeSeZtB2ksFLmtIRq0Ez0orGZkhIunwwjjO4pVc8+8BN+BdtEor500vV7U78lN7Qoc
0QdQMbHKTAPsvmswrgjV2ZKpP8EUjx/HPFVn+wEz2R4GEOVHWLCpAtKb/Shr8OAHEI2C7SnEC/uj
nhC+N2HEUu1oDJD4JHrxSPR6XBeTFYrvtX0SZlwCLJ+l6G3vfCvISgBJ5eUbcs91ydtuofbX2G5u
0zcdK18kRW0o17+A0Nb7R0ZqFpF57p7OhSrocuGLJWNUF3biomxauFZIzLjauvaoT4+fGErZuOGc
Vsku/UCYVp6pz3/htPATL2LPn56Sq8WZWWeCQTLNvnUouTzPOxt/++GQ9Stcj24q/bRUIlthDc1H
E2T5FI6ASK9klDCjJp9VFobDF5nzQWtQ4lenLwDk876coCpPDKGAJ/kb08KEWkUeTy82Pld4RLlK
p2eeMNtiw1+X+w2XaSSaBIJoWDVgoSHqu56ML/CYAdwscFk8iS5hfYnC0GqxEyIp3fdYHYrSSE+Q
Q1UgrLBvWdOAQ6LY0KwAC0E3aQwGHQl6BVU7VK27QbbFr8Xrr7RAch3ZnUADgRdi6gCYnHuzFHwF
KbO4v5uLgpp/WZjhZ85BzDBuSZIo579QFQZjcYmQGek0WOxoZvgP0Ixc6qC8zWYFJmrgBmekr0QG
YaZ1btDRkdHXxwtxMUpqRbf2+I3JNFp7ojDucpD/wCism8x9KvMryTbXfC1F2j1kTeozpX8DtTYs
bB1NiUAmcv2Giy45Br97wNmUQhpK/DNsPRfjb2LXn2z7cvcghCugNiylP/y/YtUGX0zOj9oGDelb
HhgixvWIn5ph3dqu4cRXjWcLRwRMEOz+ITKzumcyVkMe7DDmZy+6hno6D45iNKVDAJUVhXdB1Wlo
ZchyurhJ03Mq4RQs2yToCE1VcFzbyWlsFLQa0gftk4iViwKz+H1OlZ1fsUR+PDwQijSV+TfoMTm6
retwjWZ4o7JrGB7otYyNCGd6pL/9kar5JHyXuW9W922HRaPLlh4niJPLbh6TQQQ4owcPVNJ3FBlf
9NxCT5kbtwM+Xo4oU8dCUiy5EEE5RHf8HFx2YyNYQ65NfRwhSe2fwx9f3EVDv4zN6IJk9g40j7/L
U3mSS3psnUUy4LljTyj408wtSBLb0nkAauZLM60OxHlpc01P2wX3G/ujIZ6B8r8hWQDaSmGReZPX
7QzcVFyJvzDJXlVBcgXfYO1ecIgCQuDjucvXMGQ1ff4KP/AsS2UWbMcpeHDCj1KiLH/ogXo9cULQ
GXbJc2aoGTPVSwzgoSao81AnokWQi3B6dhOs+8wo6uN5eAlfWKPONiJeqrkKb7Qe9Vks3xBqb86F
X43LLxDWmRYDMHMCu7GIfRnzzWiqWAihNXBdmv/MTeXaYtxZwdUb/WZ1BhFurYvvaowB6z9EKcSn
+/qGMtCVZhOyuDsXu5nECq37OT8Yj3W/XABV4cymi4X3IrrH2dUkVlFVOZcvxl0GelRwnfSgomsU
WWs6GQrSwUpxNi1PGlaQOObhKu3/WpXWiRppxiOFokRUc0immLN6ym2KnponoEw92vZWgiw441Cr
Q78QKtPtvYKM4NwlCB+BCzXueXsVm971TNg8t1YbqZmYX/wW8dSGuDbQ0+DvhbYsxG9JChGtg7t+
G6A/m6Rgc4hz3ZvcpW1pUS0lDPHoQiU4sVRiiV7B+d6DHU3M2WAhQpJrUhxLMtJF8Lasf7amhMM+
iS1hQ9Aj6JjmaG7UP1+1wkqCziu+u2BVIGN3cds2ZDDYW8M9keaN49Myi+7zsn72Lin0xUeLZfwd
NUvW41N3a1qpznjcfBm3dZVc+po5m200E0tSCS4gk2O0fDScyoY7LsMIMqR/B9rmsat7pyz9bvKk
7vPPrQnyJ3xngUEf8dDpd3FUzbF2Tpn/vfXPX5drg0X5dWYqxLRLyYeBsWZEZXWx3wU8pwXBWxUS
582J24GzNwAPSFh7Seb3hkCjDQhOiMvdqtWsOmwRyJMnxkIa0cmTpDCaQ2DRkMhgTgDC8Lul7C2F
+YwSBkiW0DokE8X0O4Ku7eKGWwsdrZ918SKG3+DHSU0awAsEaqSDLU0eVvoTotelVlVwi3V68Ava
ewb+/DT3DLFw+DaCgXWV7c7P8B0PVjnZrVv6IBWQnhZBKfmi0K3V+AdQwyaPzYSF07Js/VmYKIoX
TgaB+Y3rmaQW5ktfJ7fqeOQ+FHcHoiBDdhzdPlfn1atcdW3NzDALiswg+9JazD5/z0S+JLoKBNWu
UTzJbi3vAe7k8uAQhRQhhFKII2THSOT1f9GzTO66t1bOu+i1tPUlDyCm9fxWg1pMA0hO0i//W8DW
LFUIeKpFAFJXrS0WuGT6lVRW4t7o7y8eMvwDN/Gt5Az1JuoIBjcgTSWFSaIyva1qZf5pTxCHB/Pp
pcuQVDiDsMKtDoR+uOn6vT1KVOL40VmM+QP8d3YXPaN+/ApESbSmXVG2QbComGZ2pJ1DICOJ3yDz
juBQiqQGZzBO+BDdPDV3wmeDPtFhS7fcZuDCsw96+ymYIDAEiIBXe9vSUMap0KZ8kMSH7dBAnTV9
Ok6mXrftgcojA7dkq1Y3cU0gz2+Vx4oail7n6QD4zMYtwiguwr1FahtECVC79/N+jWCcztJo9eo5
wGI/FfFr+m0PWCX04j/Vw90Oc/p2+JCj0KpuEj7tr7jai4AXvJfun/Up15xgsznsdD+oxVF9ERBB
quSCR3NrfyXKujxa0XRUv5hXk8u7xh/FmgsXayhFNHc7UELl27S4nrpN/u16kHUT1xoROhpVQqrt
IuISB/DwoEg/fOFc+tRC6KlvsZxyOsePRLYI6jOXp6V+84SJeZuJEzN7yfzRhu/WKUrz40sWlOHi
OCOlXRJhb5SJ7LcecQMcF0mdyABLnhDvv9XSyLApamSEn1tbV0+ua5Z1lTJatP2/4DaUK3cfnlV5
cjj1kLZuQAagyRyBNPU//2aF8YVPZGnOmK2XuweXkPWLCgp9hDQpdj7lRnaQ1HUS3kZi0uKHQGhM
CbdJmka48PiDcbrV1q7mQJusxZ9MKNc3g01F74O5Xn0jKPHeK5MaJqPCXb12CzJh67FeMTU4FMhR
QY1MBC6mQjvZmJaE/HlrSE5mjjEYmD10CzRVpOQuTjg7zIJK7R7p8Bf+W28k35zD3UqAY7kPv3BB
UgphvQ0TTWldlpx4AKGcbbWnmXaWxZhSR6qi47LC1+MD86NKTUu7YF3PFZ/M4R7YXq3yHW46aaju
Fa88J/HdTfQla9mjWepMPmbizp43R2+IvEfFjc/PqvruBAULSVVxKMaMXoBMeo5BYxRqrN4TTMOg
XvcdH7O3IJ2iwfCi3NfFQDLoQE5mPDO6SEeUpzXQNM0ZLg6x28AFi/O6b4hWwG4SuoIN0kWYOs/K
S357HsBhRkmaVwUlgLtZ4tTlNtYAXUAyqWDfMSuP7BZsOqpEixi01SjdwWTjjh47o0+8Kk6LgNit
MsfXf0X/22y/WG7y4b1WsM3zIE/yzhJVg5zVuTRAoG96g8+IF8YFFdmRs4Aqoh8ifEC2d0Qvr1lj
RICZ0DatkYOcQgAIRCOcBn35uCS5DfMqNzHcxaPR81j05k7LWdQpGar2L8SpG9nuHyNj2eCyAXB8
vdQRxr2ttQ2EY2Ceem704fTSmVD6JXMUxrCg63XCgpw+WrkPN/f6DrLteUsu6GGjUaSZERFfcKNf
D4Kt65MRv6oPiFCkrkIzsj2UjE+1qspAKwLlj28xgWUsV8W80UKprJyNyTVJ3ynKgXPLx2JMSSkZ
qXTJQbn9TIsl5tNnEWw3QhqNqZaO10zSg8dfAV94KiqVe1NZ7kG/htK9Jt2OiO7q2ox50K4ijY9E
X/ThemVgPbSW3ryZOR6XEvoYkqU8oY2DP8XCxejQVlQqc15/CFPOIR11CmGEF8MDc6Fc03x9crD5
QzjpLzZ0lj+1nC2idY3gj/+jKUi1SFaOS3CB8I6HEjn4NTiYjObnyXuana0/17p5HhjlSeI8QML/
Y4DVgCDbcKYnDsMkyQNSLrq5Qb5hxAv7xQ3jTWOnE+IJ2HpVrSi5kszeEf4bMu410rdUwGKEZpHF
CSjaG4G8iFoKZy/Wf2R28WtbtboaMsG6e/JM++/qnhy6UQop7t6Dw5OQntaSxVRUQ82ww1mEN63X
wJAG5agbWgZ1/QSpockZQxz16eQB79Y9nHZCMkLaxWFb+SNcNrb8BdEMt6gbeR7edCWzWou6ATMw
6HKG7H3X+ja4Y9POm3WOpkL3VRAkNw68g66SZVdth5hMXL72JCDOXoe2SFliVHqpHQkg2OqtmRIK
cJ6QGYxsW1l57B48CmDdHDgUfNL6YY9ZYZH4IUFE4gZFBE8niCiIIaBMTpGjTQ5PRKc95NzVQIFb
cWqJhXIX0BrxLKjqMpeSDlN0ZYu3k3NeU91YTNr/CEVsgEw8zpqSAcx2oZ0QSguHra3qvqy3lJ6Z
ZSp/Ij2AKFsvw9p1roBfYEwHbSoEfBE7cchTztmg6c1kUHWHmgl+iT4vJWsaWatgIVzx/bz+vw7N
MR0NpnpZTX98pts70CVjBzPmjxHv1lTfztqJWqlhN/ejncfvOED8UKcDiwWib7i0Jtl3Mh8dHmxT
SW8gsmlJpXDWpIi/htLcRnxyD+ZbsMHZ9AfKWZYWED17Y3T3yCdii+4rZX1NuefWiX4m1OfPjd3t
Z0ddS61EGL7XnvhPW6ZxtnivsshufNdgRnoNtGSKJYTDZMvfoCiRK/uGKqJR3W8Ww0RyAGaRmSEY
gtbRhlQ8JbULn/ZPwbMt1qcE2OXYrvuaCIgjsWuSdQO4Rl8lC+4hz3kbd6OWi45BkQUA3/TkZW1u
caXy+C7XmgdRMycZqbdNQ4wvfChRwzDEzjAa/RAKvm7UCSjfpOlGBBAZBIePtWcDd7iIkR3+zm4h
XHu6e1Fcn4xGPpUqQX2EZte5X1WyVKx/QRB2rBWuRsww6/prUpnuruo7uRO1JyKkg0KIOpdsjoiX
BpV1EyN51nJpxcdeYezmoviZsoKqMrnbPjmyYnoFWYUHeMbk25ecmVBqQF50yuzdUdo5Sn69R8Rq
b1I/8bjFFnG5ZmBZs/kdkAbjcYUh3ytlTOuJdpfU/i7eaotVK0bt9D2gmaVymjmfry3TKMrqn+Y3
kHrSrvh0R/IQrz4jJgA/oVuE5hOouglXY9HLlOL1LPqPjpgK91b4AkVLLxG9YqGHipinpLccnK21
yzSypA3SuNmcaduoPZlMOSJBDDPqQ6F1K+/SoR9ebpHbGRRpvIVj07a/A9+DJHeUTK5PPIPMppRD
L5rISyETlvQPCnthGRJ+Je5J5tm8l+rn5MM9//1ZRcgI4gxsQMqsdM4MgepQLUfxGGuktuZq3dax
zZmh0IkJS9jtN7gtVO8XgIacnVhnlhFSzislGIrwrKiwKvYFzonDjJZa38r/SCh2ZYSmmlUZP5to
lmHHY84i+qEp2lGv7y604VzsjAk3xb99vSNW94tytF7gNCMUPl7EubJWoPz8XAGGi4FpprIVJL8M
7LG96WLZJRXRAkdm7b1Y1yUsjn8l1HjA8nw24uODlK6/nnKIJLMALcGlRSzL/P3UAtgqYDl8Tl/q
hpqGw9XHFNX2lBpfwsDNqVVu/brC5UHeIAEop24pgJ9jxumRuRjoT2BRDkMxPEiWn+dxvPYGLThv
GizRXsODZsBq1kSolS0vm0/qmU1h2QqkBrYtl+anFgpVE6sDSisXBtDzaVNFQajxWRhHoeThxwnA
4offd3PJSL0x7ZP4sazkfz/FG2bEtF+1fyHpBex5uBw0NTo0Ul0W/ffTz6PKC5yo+15Ssut6ACIc
cex1iHq36net+/jCRdF0xyP2TWxe2C7Mu6Kf4GoyQ4oUHz1uw/7+t9caLHQ/TM7Y/iNOCmaoOrd/
FIAHxWgVP4m6j9QNibPB0cDnl1Xs2CiB4jLEohUfpZjbCb1shOIiJHqOzZoF36WwXhrdi0zkzNXk
Vmf8UzPEJ2eKEh+J3g4cewWcPO8ceWi0ifDvluAcGVXT9wvREXx+dIGLd5h+PFhyD26EeCP0qRNq
Y7QKvdGDFuK8OeauQAtaMnSQvbbn6dd0SGsIj4GteNoTbg6NfB4Jd/NGMhsT3pEO0jtOH+5bqZ7y
ngZalfW6eoJot9z9j5osP4B66ruqDyDqFzkrhcrTKk9MORbW+zH/p4pTkqzOemNclfXUrX2fH/HQ
LOiWvrhIiShkIrj/1bWQ+ZoiBPHNpo3gXVfLgW1CdLaekhLa/r8lrsN1YZlV5Qet87oWlYhaeg6T
79s9andQ3Q8ea0uGHm5wG74X6Y03kXIs6pvZZWxF2YvzE20t19hNylA1pQppaddOPMZQ3dhcqvYp
3/YCQQwiL7n8GwDbEnRvAnitcDUKNT89coeL7PHYtbG7aY8xb6SmfYi08wiZGHslZUVfDoJdPNW/
1vD4qOVIu0ue5L2/NL9i5semurw/0D+2221lrV1b+4jHUY7SaXJpydlLqEAMQaMvuro56Ic8LSG9
PvynSyyDmGIRdhI6tblOPqUAOzy1vXodJ9BKKDCt++DsJcuoUzsPd1G4yb+EQCmQDLpllRSgJwX4
o7zbHjInBAjMzGxpFnrM10p9ogeQYjq/pzCmH4mOhg74dfm9RNOR4+PqFTNyjnK01mINl/JRrVQy
IVin1f8ukmrFZm2i8GBN/xatJHVeAtM6uWSH+d/dZKsprIYRPFmq86xcYBIfKUybZFtY0Njyveib
E+UqdZeuO0XS1uqf3gzeyl3vVooLehnYAHlXmXkgd3DHHK7r9d8Q4B27pW5xjho24IPWBIg+H1cT
2oBd1jjLFZmF6zwSYE30PDTIXZyiH/d4/0u2cBHwvXaK3n1DvNfsQ01zN2TVLWHyc4xwon4yitmf
14ErQVSG6whC8EBFz6BDa3HOVFyo5NiH3frLS5HMDuO1zYH/Pb8fgkRCgak/h4JqcRHVV8DJnLsr
napiutidWvA2InzWqdJpS9GCdESfbD8rG3qQeb15fxhCWe7Za5lx7Hj2T2s0b5MpuD8+Ix0V8B6A
VRauPS5xEq2iDqiNklW6bV8KnQXDtFMOG5yZXKDcsKDWrEIYaoli1hCQFeCawQ3b3X3arQsFbOMH
cS9OrLEqog4Zg36bjtTaoCvTieuss7yP028XUlp1/jYO3SxunfoVvpS/15qI6yZJ3kqE1Yac4g1x
f7971clSVaKrsdLFkd8Qb+/SvpBQFiyeub7++xgjwy4CqhNJeLP36UFRjxD+GxiDG9j5iBLYrKdl
wQXsPidgOf2MjgD76MJrE2mmWXR31ea2F9Rr6dALb056AHp52j47RiOqKXHWZr171nnLVaurSTDq
GlgutlLcEpP23uKksqW9JArpPot5GSpxt9pipSL6ytx5JfdhJD0UwRmnlk814WRY7pbGlu41VgCC
TQhbWRFX6ktgo5AN+Iv4+pvuIAnAliTreMk076P5gGIlxv97m7Vud6RkEF+SyD2jFWS7QpGdn7UA
hxq2dX2mXsqPTEOVhWQXDwbOYELQcybu8s0WPsgkeWZ98YEscCbg5O2dyKjAT/rWrwBOfn26/jUj
egCJe7yJpVmrjj4JX6+2l9wC9B+Moj/7HkkEnSRGGrAjbBxE/sMThffZcbT3DNDYKXWUFQ/PUx0+
pfJEpe8QZRShaodDVibJ4FB3DAQoEWVR/5lvu6xSQzKZ6jnWmjKpK8ghwu6MFZoFZgA3V91BwJ/O
Kd3YGXr7DRfpDUllEYlGWL+9EJw3XZXpmoRUv2ZWlypp+uOhCqaMw5/QKQfu+jbDxY53VdSwXzbQ
PGb/pJaI0pV0w7aY/Fwa4BO/7Vq8+Ash3YxZvNK7ktSR96xWV5ufOnKNAOBwmJrnwAyBobVlzvSy
B+d8M9jhk3fFMiSs/Zdimo8fPFiEaes+4+CmsNJd8M1KUAv7mL9odPePLA+SmLRETVuMq7q8miNf
AUr3dseDrdE4kr6xfwqSodKY3fMO5gOK407uKJLPrzrL8ITWtGAxFsBA++FNIuI9trhmrtsNWYoK
YcdfudVmTElTqRRFpU5iaK43UZJPm5KLmTBiSeB+8tbaPmRK2pxElvlhVlCNKNdmbzBpdZ2xjF8F
qyovXjX7Abwr4TmwuOTgi8CHgdZhT3Vx5HisQwpExEC3Bi0wiEk1hPuPlTLMrj3mC5ZkTV5/0m+A
AVHz10M15P7qULKVKwQt0zV4OIkIpssUhrNoDACnI2OXh1l/R4QVgCN4PHjtQIcUpHCbZE/g1YiB
VJghoYtR7z4hw777h2fKIQnUCyyS2u+z7RUDT+a+xKG3ewiLr8dlmC3B/+1d2x7NplyIe0icwD1b
sUWJ3SA8cwUZ2arFu+6ASfKCHQVPt5wBgWtof0PUynrPeLR4rkFnats2uAndPZMnlE8cbd7HlFM2
0Z5eqnJUnUsoLTVfZsJ3AxhLjbErh0f+ob8ZxUDje5Gr+N8hR9Fr5GM3awgbD54pL6yCpEqPz1tI
lC511CoBaUrKgbb9h+vvdRmJVkI0VSqrzSdWYA4pOS2K3a6Z7YBpN+cJptIydMMpRk291+Lz/EAC
KNrEv5H7QIxdqntfwSdI7QdTG7hLddt9DZUVmyuGvtbQ7ywMzY2uCeKMis3JFluL7+5rN7z6OyeP
PxMUj3xyJ35gJucZ6DfSTk7f8RHdz9qCLpraVt4hxt+Tm94lNwmxa04hi2kdiaFpCMh+116IHdSx
OjxckJdovqhXZVe/elQFY94OA9NYPOMKzCpMqpyVd11NlENGhToZGq8XkTGQCqYHOUJ/mYRGHwQd
F2lZHMe9ydoUSIMYGmggfqXz+ZaqesxbLzq3oTvCzzUYtywrsCmKcpKmFOb2zK4cnSquLDgR+9q8
oNpZQoqQx15p6smlyus4ZnridgPxdNwnu3wqRJZ6ss7IGMrHGrPRCOjr/ZmTfBrMSAP1UI6UaqBy
I72CxilcISKBeAHuvexRIsWCN5Q5XzuYovSLiv1rh/6hCUVy4OupTdowcRGowlb+A0DQLxRjqZej
7LtamoXmLjufUR+n+tFJUqoPkqdHAI4FUQ8NIxpwVx36YWj/sI9KjQ+xruPZTUD9c7lo9AWZmi7d
//s3bqu9YOyhjeJzL+K74jlJLGF7twbQebhpaBXkxo2o/9xhTRUhwG8I/KCsulKErc/e3LbEJeTO
aFgyZB8v/xK5yieQVPWkDJbPDNEdpBVHNAvZTNia3ex/S0VMnvgGz7dq+AgtLMoYEbLwW6CARZ03
WVmrhX3ryu4GD9pZm8Sugf10a6Ry6czpJJF8beNHz3iOCB/TnvlBxw7Jv68JhwFgknddSuxO8Dc1
Fn6bo8fUQBOSNKg+AIP2VDUr5dLOcn3aDrKGyvv+pMnoz2GjqyJee7U3HKe9wYpzn3dvpbbhvoRA
OXolRxZIVYb5hyOgT/vkRRXLTlpNxChQ1253JTTp17DvY/CFQgI8w33jXElp6Lm8K8OaG7xU9615
JydiLzA20DqOAsiVYw06MQNGy/sgIJVFytLYjRO0z+56N4ji/FegBzTQm0f7Ktcx5NRNQ+2DVrsF
J3dPkQNF9QDse4/jEniQkEnY7c2TBJkoZnfbYCFj5uNCn+ORL5QNh0s1i8MneBfReQDK6sFV7iIl
pSbj8jlmQ1FR4494R+/rf8ln0cxwdI+pnYLGvHZGf3WuRlpq2ntAGLiKSOhGdf0idqejEjNVVljz
RqEtsbtm+s9hauVgrK2R2KSWkF8Va+zQ6gsgLbC95npIShA/XrkMQQcCv960igpoV170rFqXwyNe
eKyXFsTifpN4ep9AUOFTjlt/tyKufz0EtvgoRVQfjiPZvj5B6NBXMUOg/4Eung1/qoxLJs4YrrWZ
cgN8fgZVdfvEN6OawH4UTLo0gLGqGJUCablEX2xlsF/hc1OcKMREY1mrxQb4de/ASXmDxraGUHW2
VISVuCXDsGb3pMY1Tsfjf7lkyv2hPU3CsZRpsv3DHXJ4LMsG9j9+yF8biUiVF24il1icNxDmWXm+
43tGGUox7KIad87muhXRGHcxkpF35ZZPIyiA2nv9jAs23IsMT9KQFTdhueY5+b75A3DF35DKfjh5
TTQQJax3+lULZv+JCmHpfPbbaDsUV32FG4yLtv1vqkRyQhsN+W40ESQWV0XvpzkTXda7V8BXwzDx
AJnkkHp/gsfmgyFODlLMIfPkLF9M4E7hgTaS5TLzoTgN+lN/ordZ91FT2fIPqh+tP4UXW1hfBfnZ
H+m0y3Hbk+uWNMAyq4PIl4GY41BygLQEj/VpGwzKQEW09uQIYFhgjWobSjHyeS9hJHWhyKnQKtZk
Ca1ZRTB7Cnx3tW7cjgBZckAxQGlW9V/1Dd7/GaLqBMQXDT8spmPyJek8gJJ8LGQ9ksHc24KqZhEZ
9xldLst+oY/19qr1gvwhaORNnMdjYlm1kMclWLJph/XGYSLIDjSf2UrSz/UhNNWCbesQZfYBzGT2
QBQSiLOd35AEBP6PXLbDsozp2EgbVBb4prGiNIrAcf8IOTx8f05XCrIuHteApznEkdBUJ9buocLS
cgEIdbbl0Xcyfqm8z0Kxg8Yn1XyNB2ykHUV0GKq3yyYrgJahCOjzNexBiHcmuNYXDuvpDb5Sg9vO
1NT5SvjsGJpyIYgvdSuL0pilcn/l2BL9JK8Th9RKi9wRcRP1MW2WfiidFgHrj5DTApEqXvu1yS6p
qCcK5F66hCKLqiW4PiE2eK5Hl0DyGjDnigtXnmO0ojW4PF4beXJi2kCEfSxASflTVsvmwRE3s9QV
Gs730AZ2M1ZmCrKVZsLCvBycKr80eilpqj/8Z762e+Bl6oG5q4RcYxbP84iLYNgLjFJa5mPcbE4d
HQYdxtbkiq49zoetFpyLUYD0UIp1I1GmQLzOgWCSdGLBbCEB5voo4AB2YqhqcA3or19yOUhb57aE
C0087woxf6vmHuYkigM7j9zgVzlhIqo4eqhs/7tLt/lKnCgtuRgzTqqYeHdA+CsTxZfQCKtLqDbR
6XEh4h3FzmYV12aUU3/iiSrhJuSCM5v/xMX9Y3JnLin3sz+j4vIZqr3ao9jPoUl5ZUgFejm45iBX
AXiAnN5jeduV/T6VMcJOkJCHJZxCpLqMJAQYYahbX/AFuyqLG+W1nCtclnS4YZh/xE2KHHy/6c32
BGRuCemUhGcJODNpQnO/oECBLNp0rgQwPScqj8NUsCsobk5owrAZS5LfNhyB7PbkU2ALcfyIqC75
EtOpLd9QSE4vfdVMNckyBMvhy/BpcP2/67lfBpCNu5buW8jDoP7ENfo8h6Azx0oKe8mpcb3cSzYt
FY4wvp+7je5SYbgciz3ILn0LcOEQZPdygF4C0HV+qyE21kK924X/ced9lbqCONw0Vi5Yb+O+XNY9
8dM2nLOUjECt3stwjeiWfo3iFwVUoeG6GbX0SXxul/WcYKxCL1iUlqgKxsl9K3AaZ+Vk7iGoIkhL
4wGCkKtj2aUgwZWcZTiH5in08eOOhbukPb7IrNtdO1LKxCgN5Y5luyURpzcSbA6eTU/xO7uNJ2gY
KLLcta9/wFrKVyQVsWpMVkUCcwFmgH3luriXh9RevskqxTQcnDdibeh7jnb2zbgBW2wOOLEFEslq
FuZfbh+EUE6r5hRUrTaat6bdKP9TGdN1jefy/5tVUqmQ1XhIVvLDo4lkv9EQjE7I3fGFbjI7ZU1H
mYA47fBoJ4xWim0VOE8WEzm2+izQkIwwVQAvU5JhNEdfiJxkmnxDygpmRVRQK7kDPgDZXd/EbnDP
UKY+H0O27FopeWrjx5MZI5Keb3yC+isN3RLAqaBAznGIrsVu9vo60gYwWo/ucBd66tfbgVGgzd8E
7tJ9P0PcUMBHSbZIlu+XTdnyGLGvUuAwNlic/BoONlwWWrWfxqy4Y5U0g903i8GC9Qc2OqxNxlzL
Tra6lzaTT37ch1HPR+WHu5ZJl1VzTdTT1FECx86m0rxRj09mbu3qM0fC+B2S7k/40eSdap1UnHIJ
dCQG+7MVLqHs+DznqtqRo7kBIay51CX69bq89zpNKDMmOmAA6iqdB+gZE0wuZ7paYnAVEfEXe5Pk
GEUtH+9XFMoJv+r3jLrzUNax0vMYtniGTkAuy4o5FD37KJfgaOq7Olb9I824LHANCAtCWvMjsfbi
OwkV6l77nW+MUt3DZ7pYsS4iW0B/UB9uy+0gb/VtETGaHzWE8THm4J9aNbRY43S/z9WQUGNl4DnP
TTSHvfbhIo13/LSsXATqltJFteCykK53wE+1AIqaIQUH7ygQMkGPN1I9X9hv1eBzc9kWwH+hI8AF
CUfGe3LTsL8ZrOG7AiOXRP3q5z1LRCK8OBt0CvImChtgtvdPyMcAK3hZ5JgY4hQiFa3pGNESOxjg
J32iOg48lhhp6bfNTB/C2/rUnVVI9TbnBKCa3xAnUlTJ5upHo76NEBh3t3NIsbxivoognx65ixDA
/UgbZIjht9hesUiE3/IaJvC5klwt2FxFQ7sJwkCUIWXq2G61vU+woaGeAKKs9FyVdwnrtHDrq5nX
tA4zj0u0ul1djmVp8ikm+Kx6SJDxkBrxd1Fs9TKiOKIpb9FJaQ7ans+PrcEVoG5lVnimy1o1ydal
nbkRmgfpgKgiIJbMzP2azxDSulij1CCvovZbZqL1c0iyBC8ninBFcMCk9S3Mv7Oh8nMt6qxpTKKU
CtOhkrYui87gFkvPugg+sUFyx/mfRv+kQZzE5iW+z8znQOAlghmRKIqv7p/gdBb3J6Yi1idJRQ6E
SMdC8MGoB1DI1iKmn5gfrjc0WD1Ad90tjoSXyA2U1SXm1AHeYucjm+Z9NMJ1QfeavIqwDOOgKBix
GGmkHjmfvYMoDGzpg1ncZCNPVJzNvmVX+U1E5v2iM/TrPj9dzmqYEtLzh6l9FL7Fv61OB/iIM1tA
gc9FAL67SaPHjqwtXWZZtY6m2NiQqESshVCLdGgbZkgGPy5YOr3hOrBhNbpaH6uwFiJ/kUDvIoUC
QAZ8Rc2eMQv6B5j9f82pU/00qWCYkuVxOMjvGAIP5d4JGOSGg2F97rA0AnEGVorQWiti5m28kOKh
eo2yJVJHnsAeXKK/dLZmQh5mLn7rn3FTNLv9Y55Et7XpXVyxEzEiUXI1asnG3DjBwLP76cVj/qyx
hw+XGXF5JzDJEOjZFNE+inSk9ei78GtiHvy4Ed0MBtVsYw96eSIK7a6HpYLHAaA4AmSAHDM7CfG6
DDo7aymKOjArwTD8LEhhSZ+HXgqj9QxtMNLBzYOySnPGPPpSPGL+k2RI+tlcPKzIUEZ27lLBiyIQ
OoHcoFMM4INcah7ozrEbcEJvJUOO4CWbDSDvjou6UUB5P9RFSNXp5tz7Utc3z0zRXtj60/7PB1Y+
7JOqpWvw96a/R0HKtagtV2vo59FJ7vOTJmuAjiBhgTD54RdpIJqObVS8E0EDmCLx1zY0J/oksi/e
Q8P9RktGR67Jm0qQ/GSsAoxwFXsM9V12WEACGIajo+KSGmw8B1gFjvjUyaLH+K/WTfPsfdrP1yVP
EMubNrNDx6TgGNbeLWhekt1JEizeyOpEKnqBCSOj32LJitTFc2m8B2qIv0Aof8ozlMRNYqsDnAnh
CxYlsJb+WMtl1iq4vt+k7/bW2fNC7YKYBUBjHLpxycOhZIQWIk/GuEertD660Gi3Qs41AO3Ij7Fx
AzmlzuXfd7ZySCFVjv7Mgy1y1ofa1m5fhy/oCqgq+uOAGacVTkKFJkYTJdgESdoM6cfWNV0Xz2Cz
HGeXQBk19LDhAkoKeLCq/BhmsXpMwby5A9RHwh2WmqZCJQPWI/v88JSyy14phmaVkKNaNY6ATH1V
eO4Fd23XviweT+oYekrTCy3jh+bbj+Vt9Uj3GPtus9MfCI/q5vObWKlWAHFsBL+NooubEHBIf9RY
H8vPxthuW5Caq3+tZ7NBYf3B4HLDhoESgSVQKsiQ5PivqXnr2DJnfxW+GtqfiLSJjhdZLAI1n6CP
GZqqSX3vrIJ4GWi2tWMj/PAO5gwbvwVFq39XyXCQ7SLVSjgZQHajGRHrNq5OGPkghxfkTnmqT76S
m10SInieUNEgxyGVDgeExSkEORnw/rp/B5gbshlhjqVOxtmq2b6rrtxUontm6cnK1lzVwp9lFB+b
P84gBAfZl/qY+G5+geedE5sRjq5kpvd/2D80PoBjA8X9/+Ojlt7cXh72GV5DKVM5OlYCdQfmd1TA
62fJ1ZFQld9FcXckgZnQWDq7fd/b5D5avCrEQp969Cs9tK+1hda3uSGuUi1PI/L5KncaoLmBOfxz
IsqXqH9GF5SqDFrWKe2Bid19JReQQi0j9z1pQe3WrHuN9RinNLVK6sqwdsM8QlC1mzVsVEzeSZwK
coP8V2NnP/nDZnqkbI7kEN6UMqy7wEfOXKU0KZMKfvJ0SS6CkAkhK6YMJwps9IzD3NPl/XzCneeS
C9nUnyr/8XQ1njFyDsERg5tx68j/fqAhke3ONDel3jb40uL4IvklR4S+RHDXYCsVIdB5NM/zgZIb
Kz+3AVmJtQpgdl5uk8gZft/mNniSgT2DZxiE2U8CEtGQYiLd2nqcIYTv1S1N5Uc3vt0sP3l28KKm
z5a13VKCtR4VzlaJN4Rxt8iVJP5eDfJX4oCLh9piMXCMFXEHl6NvanaW8VEmYzowQ/VXafrTE+r9
yMnBYEQVCDeSi9CHzvQcoJ06JbIU2D1ZupPaK5abuqzXQfPd2EziM5tlggf6YFwTyN88SxhknvLw
BCHipEoveLChl5dXPFKk6p2HrOBcDJ6W3/z5P4vt6tLEFzT5WYuD7wdVgkw7eQGOqjHzRuUh7S5z
LKjUL6lvpdcw4X20ixCRkUtdpyM4TYNTdPzfpleA9sqcxaDHIP/kLb9EAml6hYWbM14EK3cfY4Tq
KvSXgUaM5mq5dHN+2Hgh+QcY3QpGoMsZHe4AaHPma5tVIwS0AdECHKLfX/xH7tuewcjFzCqVi7kj
uMxH6bq5WPMDq4jrfJtKRHmNgHldkrJeSZT9SzOwlz3nQ1PlsPJCYbVHmtyO/4oT6c/kLrWzrBbw
ypM8AloiT0dIPekozXbOSQ+EBxGhbQz+zJmMjReoecY+vrSSn1f8Ojxdif3iWd07II/iiAhNMNLC
e4rgCfUkFaQpu9TdH6HLmOYKIPE/6ZPKpFfeFJHySqn9lxPw6PLTbqRREQwNQCMbwrl4elOdvEd9
Wu8HoRZuwCpJmCuxdGdQoq2fKZOyzRtvDfyx+d5yHF3J04RPtY3M/vCbByiuZqpjPIwT8DddRmKs
5lkWZmppYTnqabU57hiNgl8d2YekahvJURgIJ+mt9KDTUowMCfayvl/+lkSLj3wLTvMqzpwATI0V
Ik5Oq0dXodqH9NoGzE85W2Q+FYtCr068EK8TkYHuB2Uze+pyP4nMq9fo08ZuqekghirYQBTAftFC
hGs1I44t6I8KEaXsxbV63qLECHKUBsPqYP6LH6M+yiTghydi/a/xzlBXfrCrGRapk6TYSKEtV/sJ
Ktr7SiapzQRGX/mGp32U+ccDTl8pIEmZM2YTOvHMziuWqx9iaoSbEM8fgIFKrKbAIPm2yD3sYbp5
R8BKG/s9zEX9wbwDlJSLjOZ466xNOEx+86uXbnAgLT37R0nCgNi/OxmGnYrIP2xcx3/BRgKB8j0B
GiKFo7qBdbJbZBEkJWB9nGrYUBNO0+H8h3LlLx1nlm8j13qZrM/QbIbWDKLauRxlQ4pMb+jiVP1u
MaDMLZQhrDhuDG2IOduUFDjEzJc7AvQoQYFMlZ8r45POUHgDsthPiN/3QOMn0W+UN7f0BxKEXTGt
l/mb7fl9N2yduNBJPqLuwHN9D6R2cr0ZDtV10ep9hmCoMILBROtVaFuOhLvZaIcyDBPW33iDfioj
BO2uSmlwp/wIF14vAyiOFh83HsqgqIbgBu3YWqbfIipKAoLNmup4EH+MwrKoBtZq+TpgQ8K3Nlwz
bvnwkULqNgBjbP/ohRDBtfb4E6y11Tuvs0ZAbyRfgdI2aFkpnHfEw5VkBuu4R+CPft5Pci1r6VfX
Q2biZbztdLqPjV1k2CUOSV165cafMbOqDuYqYPtaaZPdyiIkRUx2gJdGH+rtEBT/sdywj43vZvRX
qLaIMrrfyTeqq6zX9N2okjdWJtP1YETBqo7+M5lEMbvOGsQ1UTJXGmc8svdECV7NB14bd6XEPwiH
Dz5Il8XmL6cZkJQV3PwBqIHJBEwDAHowIJN70t8EKzY1nGZ5mV4B0bEgvANXH15v1Z0Shr4N9dEl
TWKOKxwEqLHArti40boStIz0iQjd/RdMgAdIX2PluHereSs/Ep2Imt8LPkvfcFmxirPdJXQrvCVO
mlrZkYS71lDS646u3mq7ugjJPm8CTFk8if3EDyGw65eyIDhHYqJuWEcrPON5AaxEDyaf4sRkNzdu
en9aAQ+3/QCgEBi8ZXgwwdbRL68+NIIvLEMTh8e2DpliWnbh48Y9a+120fELohe7XKKHVuBzVjkS
blWZtq6sdxLoIPN6WW7BuJ/tb7ZYjSa8uOB62/RFQVwLBCIWlDxl9xH6bO5ZTuWRh7RIzVFx5d9d
OD9HZhKfgnqEG2nM3kuGYhNnyQyi6bv3Y4mk3Ai9GEMeJ2vPSdR0zjZlJYS57g2WHl3ph8gvtpPX
11dz6TyvwDUTAkkVhVCu8LWXfmm52/TSp7+Y3qcrZ4SKJsyI66ZTYVx8nlIOKs/099Hajye278aR
LkXQwoQ5CnNsZhNlOV4wfmKgdx4HX6rchqzmnHO6gHsxIHvIbaqJWfTNUfW9f0ZlPbGPXlij+dXQ
ttu36qgggtv0N3smsRK3ZCSTJKOoEgT/0n7958KxSS5yoPIs6r+CpsnYNrZqMEfQFYieBBGBO4jQ
qtZbgVQuwYy/KhcP8x2PvrXE7GFoPCFw/e+26qL4pykIRhzf01tcr9ZOaaeaWa3i/zNQeKp3NPc0
8P6XhBKq/TLDnXfZfgdNLxlUCVFAZhKfgmPap2G5E15Pg/hZPpMj+dF8l5Xycs73+sl4Ph26EvqX
aPBWv36yPuxEpiRpd7gc6SGZ+8tx3vD/WUouxAa52MisjrmcKS2+qWWZMY+zOIOAgfOjHYo3O536
99XJxJI9t+ijFS6npfHp5KGq7OJZ3YJa2ByZIdtWBHFXqr3VUvJDKlCFJC/H3t+bHYsIuLwtiT31
VIbibCjoPdG5XPY50JMDk4qWsdf3uT10+pA0BL2T6yQTsQsCLkhJDkTBq5ITgSMYVZCAtzJu7bC7
CLSL862ubHMkSkJvGI+hCQ27cXvfnriu8To8ZhWXHEOmGQXTzb0CtISMCQpN1isPSBdhqJ39Kjw2
O2yxu+8gHR5BvNMNtmRvESzYuDTgEDFvvFuGcxX6unBhWm7CpyUYHXua6TsrrsiHJfswUlDDGO/8
om5BQ7ezq632st5MqQdrOYr8hm5jcWhpXynkNqro/yitOVaIm1gJddrcuFHbHxZdNXbICOqa4P8N
OktA4azJALgeRX83d/Encd1CLbkLQoDuyWEGMdp/4DnMl9R7PH8yL5MMmCvQ1UcTtrfv7hD6QeAD
H4sGfnP9V9uFbD9PAWSotm2lnNYHH8pKnyVE4nQ1xwVkli6dPGK5Wh4hI9jqIUwqAaB2PSZlG2yF
ngz2l6paGIbkrEpOMhI7B0/IfXHA4UJe4fOGnIaNzWeJPXGPvi0nn/yhP6mITO/CTwkExqVSSckn
cAvTePnGwaWjHlLmkxeqGGKlCiMHa4aoXMwNUIfh4H4VYJKqc18pdZHb+O4QlBKFt9E7xc8OnWXK
bZf6NTRC4g2vVT/3/hZ22k95SQqTVzB+VpBMo+qSlAn7QLvh2OTeaOA9vSKAw1JoQepIRH9AfTdu
rAu1wvyuYnbhCxoNOK1eqoKuyxVrqnQBTNQ1+5nzc/f4B1xUOswTbVE1ZeGnjeRLHnAdils8EQ2X
2AfTv7MuUYac+IYsEKYLxMsyA9TDFw5aQcijSww27MDEOEP4pYmEL4Ki6ewTwad4vdTIGcIXgWtx
xBAkKOEVOhpv/fFwFwBeeUy5NoyQfhj1VvqmVZ1yFwg7YqRbOmE/7J/Tlp0z22au0rdEHYKz99+0
lw2xRUghBzBhH5C3VHsp8XvsRTcSWOCYrDO8nJ/vYHPP5EKWPrNJzo0DESTggRyz6TZt0Y14Uw5u
PAS7R+/QE4bt38E9uoURntf/3B5wJOz81oJT9Fk7doeMCzoGJC64dWwRL8wrmFicQKHBuqs4SCC9
67fyyFzo0aJB1LBVYFoGVTGSqcwte2MptajbnKFKhXosa4cvQZPKeLPxnUqyGtKZ7GzTHG0zNLBr
Ph51WyfM27g54z/stQpELXqdJ4tUDWI74zLKM17RUFdJkCjtfC5hMhW+wWu4bGCH695sKcIpuaNQ
dWZAKYe5mGlCfguDjVElyPeAr3gieobttrgkYvhles1I8ZpUSQSeHDgCJdn/OwV9OwoSxqlz9u2c
SoexmeetufEogpkaDU7Dv2A0PpX93W6/WzZAXrQi+7eEvegjeG2g3S0WBes2bGaMxmt87RZaX1Je
LNIMv6LhpRl0fTU8VXroLUeuOw0yAXvc/OhyK2W8/iMVFPM8WSOLPBl6zluA4/Iqhh3ykJKPTPwJ
oY3BEvU/GnQpj5N66wn4bRMIbcBsgJZ4EPV89y0wF6bs9gHmcq8K1Urdh4/Nmk1iqxzdwJnSnzjF
8fCBM7VXDJuWraMxPpGQP2wcgztEmQB5YT6lVW6uA0PFPV3sSpA1gYaDfm+EPCjmtgYqCQH4YwWO
cR2TWOUW3POPIyAW/u8zXjJMDW+KPvW9kmD0NscXpHo5hAZCGpJCWRZ3f4EzjNFqAek4W/SELN2P
9xlvvIaZLglRYQqqEPuNT4E7yELNIQvg2Y+C/Kbhb4uRFjJjFU5ne1YBh6D9+yi6XpQmH8zfDpwF
sTeGTUeO7DvoSYp1ClhG3yksbDu8pbm+GW7s+70aEImMuJZu/liX0Hfs+3jl+mpscObNuLUAzX49
yTTeVKOoAPM1A8hMi5QsoB0DDd/CEUEytjvxGV8wMDLC65l+nzRDs/QOvu1jAhNm8EDgn4cIp3mN
DLfVNxB+nNDZbONuvFUgCTC84T0Bi8MfLqWXaA22pcuJu/mvglkp+qLKl8wzfe59W0kUpyQPou+8
nuqI5lk+VDb0KcvIseg3hBwmN8tWKwLLWIwklBmM03bJz4VP/bgCYfHCadKqIFlCKTOoll2YRQOm
PJmwsRQdzCp14z1BHN/1UvffKD2tzBWnA9z8//3gIocObClPrDJtEV3peMe92x7NBluMKOs8k9Qr
LP2pKPaqsdp9OFcVwWWXuUbfu/q0i2SlS3ecFlmlfk2O5Feg11ht/+ZrP1nDJJV4AofgbIl+alWn
ORcmFQMrCI9+ixtmh/ldM9iZX3vmauX/PNEbbEOOoZCdSauNc6jdtynJLa9N2ns6gjAeY7f0dkm6
RQwL2ID7TIl09qkk27+29zR/gLlC+z163VUBSwCfwl6GLcRnvc861aZjy8F9KnHbZxjrcNMQIIyU
kcLapeNsuZW7z0HNmzwDiwOVqZJGiXIr7XQUMwArxtGKHOs9qVGhaLz4cnUEEimUIZ5VyPXcDhKI
q8BMrbzfItCp2obYeLz9vnms+9NnyQ5hmvBwiKEHJsn4mJODCN3JL0VQPKiBukmCb0TYmFXZvluS
fOVkM/R4ttgzcxoPShMXtOaRQcY4B05NzxobNg/gtW2gN44YHm0/mK8JwgwzsNKj55JdrTOHQkoi
gFbqYzy7y2wAiXvYFg+0DHA2cRGeDiUjuZsI6W6sKuhW0wxTL1QrA+h7A/UEy00rTJHWXZLJVDjn
CzLAg1ZIZQirKmhbPcPhLoS9BMhSLpRkBc/5BiuWpoeXfT0z0nQMsmn5WzsVxgYy6U0qhvnx+hzH
wRqS9VtTlfaMVMAtw231+0MzsXiNDmrMNPBv0F/miSpsY+16CK18dzoE8if2Q3Op/eqzrHrSCqxt
TKjchp4Np0gm4yih21mRc8uB86aFgY7SblKygaK9RIq5kgCBAT6bUOoP5bwxx4xD3L8HtjYI5OWd
jUmlOxzD0xixMR6PF2oIJ7wMl1ZrwoXIYqgOQuBXNBfpuxCqMsfvSsT2iglda8cFQa9Sq9JFSBYx
/Jx0XTdUyKItFbZNqlInW1Ap6LZO+SdrVb3Fa/mapJoLwvl8o3L+xQqQT/UEZUvj8u5QWnDTxknm
hMae0Ns52uUzOkyeEqzraWaxO7Q3dLdwYMbReyMHLCijWPgzF3LjKJ6mcDRfPGNBj/ZL1Q+jJCxS
ytwp9QNxaJmCDpBgjNPpK/tamygt8Db1axNk4b1uVWH4LCEn4kyGrWzcUI90yIpHvmMtCQvepdID
84jErnZt3s9N7eH+QBWSR87RfAgaJdbJjty8bSZij4uD+sXeZ8hXu6BJLZ2gAUttrz1dAkwdVgQI
nXd+dUqMyt8h7n9CQHnNHWh3IHPdRnRo1ZPwbwILVanwMqaN/+mzxePTAF2mtX6BDZ4m/xs/qQV+
3t82vMZ/sTLyBKPbBu+CKbc+pLL542NCUxpQrO7Q9LqScyPYBST6KguZ9zFIWX61fIq4PtG4U0WK
b6xY1/Ki8haAN9BK2XwdA2cdRV/z+Ki2euTNAyA7KnS6ZqQ2kLEBgkQn48jhlnNAhRg9CsoLM8VL
j6abgNEoW0v04OQbOhusMQocuaM/hxJ18pzit0n2oizBK9HYEwZQScx+o1pt+tMfxEqz20AdFzDT
pYiaLZiaybov7JcqCiifimc5KlHkKSWB/2oj/d84X2583R6h0SW0m69YpJjK/ky6VHvb2yK6mSPx
dN9Sr2ylXxyhgI5mHT6EVuB2jHba+GvlsHtRZhhpIbvvjDzQL/ZfFe3Ekl9cYL5wwC87c65Z+BJw
ShzumENS7/3RD2yXt2mCnUO/wGxln4jm4+f3VQRiR5WxoAx90FpfCpv43SfCg5Gw8mEuQVw3tWMF
5tKqYeSG+ca/5wjUL5/OWqBJmgxGau7de/Hn/sb99R2j72tqdyGNW12SU/CWwl1xhyKLB6rb613P
GjmY77Bqvk79ZvsxKPEcuEDvoKbi4mEgeH4DEdbXiPfW/r4tNLWog6O8lCrXQ8RD0BtfHEwayBZ3
EKjGbWqIcsNFjAKzax2I3fJlQQ9M22jpaQQRnFqn4yEdbDZhhgKXjZzrzffr6qfKeivnE3AIn/pv
aAaAKQHKIm5SDiAusg2T4fJlnfkcKy5pJQd+xUd79L+cq7DcMMtZhtl3BPITl4y3iNWdvEKa9FHJ
p15L+HBtfUU1+Y4uIYsKDzzpeNYvAV+1CZ0P4ZZMQs/f7bLlimVNHo7bf1maxGuSIhH03BF9Tfx9
1Vto9CrhmtBbgmIbjND8hglGqnpkzD8Bpa1BTSPR/IUL246UP6gyjzUP6AVAD/xh/mGk82xDUUHB
u/9jMwgWckYg80pYZzucXKr0YCn/wPz7JoCdzh3xB4WFGoeE0dNg6NpUZOhdv6F1iVOiUC+hlk6J
cTmRXkjiwO3lJ9ag/f5R3bUC5n29yen0fJF3mcuUptRat4TkXgv5mbs+BOGSIJbQ+VO+EMbzpefr
QFWswahxSWfT8kNRTklZlCZmsgJ3AO8+wuRXeG3ojn9JslKT74HL4dYLsuQotuLZ8u7+P19ZFkEU
tWVg3ZMJ3QoQhgPPo0m+tbgtEFgAb/K/Pkuqfd5vBr3XpTrnP4cEizwdNVEXkHONAjbA4r9N7X6M
TAluOk16AKC3rEvU3e6tX8VPry+ed7xZk9PhDBk9oOzyc5mgwwejdgyKU44GevTM6ytB7bxOBfGE
dqFYitORILkHuGG+YtLsBX0la7Sq3js+CehHU8hZywPa3AngTj7XwC3x5fGubd8q/KyBCoqmkG82
vTKMGH7wtwb2o4I+MYzUq9LUmeQ6KVu8Jdz0blA1h9qrxOzS7zD79ZFi7iQxuaOXPVGx8a7S0Ex5
/tf+Z0S2d9W3fyYxp11LfdqhZYyUDPtf5XS7rPCJc+wUC1uBaFYa6xq9WOUQwpu3ifacTv7zeMS7
VCQwM5paB2CC4KoBgQ9NnYH3aeLXeRu5us/N1tAg7Fj7S4mB2bTe02XFLSzAhg0V46m96p8w/57A
DRdABrcgPmILDPILGpQLdFnleODbjmnW8sCxWWRQHYEyAAObNnntZZ+hKiVVZlPiFruDhlIMjKr1
hw7RxvQnD4oh9m1+xv7XbM90Wt+JvGE8GYB48cbVL/zqSbpoe/f1yKrSj4n0T+1Nvlxg6bxCQsTw
ETT2SL9WyoSUxWPVh1xfuzTzAyCHm4OrB6a8uSWeW6kxcbzKT57qDQ1K0PljFtIjCqCzeFkExMVn
pa43daU4bPgUjNz5ycH2v3ZR45QXlHgWH8KYvf3wiqQalE4StQ+vdd9teU9o7fywiKsegjFCl2Gp
1hptrQeOGHrQhJO2QFZE+JGn2Bb7dVKhLclQW5jBMqcvRk+0MLiy/4gcLW9jyX5DGTpqssk3zUD8
UTernkm2NWMXXBfF9wLt2mHu+WfbeIhfANj4vtOGEsqqwjmzh9pDEa7BYTDc2s7oLd5uHKoJltOF
f4/48gZCm2oVyVmZ4nUG0sz0f0FI4YEqpNYIJBAYG8gLZwgn9hKnYBOtAPvkQ9O4hvDay2QTixAT
4Q5SKxiwQUo9ZWM0+oQ9/3X2vQAfhOfMZRUR6smmFtdOECTn3tHImjegMzGLsYA0iLC/bsuYHPjf
f2YDMKbA5GRYXmtVGTXyKruA4djkNRqKiDBHOsOPa9pMFcUwLKTljazOFAaISt6fn/YWJMs4UDTS
hCGLIqbq+aAHDIGCPIWtTCAFdghi3wWhOOI7O+w9dbqVQOfD9NiYDbtCKUrifyyRY0JFkjgKKo7g
/c1+fF8oBPBcYnyrU+ls025hJYU5Qeco3YRbOc0w/FRPh6UrZ+w+PmyYEdeg7SFxG+kF49XHG89h
GLlrIxQeoLvy64e6SPVPw5hRw6RgzzhtYN4DQ1PjHvZTFnESnkOuC3t8WM1Q3YXmc9arGlzrmbjD
igv/MMBVF1MpePuA+1D7b7B2v2n03zJtfnSVmdOufPEZp06+kSf//gzEWMT0C+8KTTPROQVwDh7v
/WEtML/+4F+LA/Y/3zQoRBF0P+tj03DyECvJD2XWAIUNkBcUQDFjEt/xrdjzTQKH6JOpP3M027ke
sxbi7k2CARQ4GmtVEMp+nEC6GttVH2/bIXHRPAzht48fAeozTWj84coYGkDt+/WUsjjh0wMVJDoE
cBLPpiZsnrWlQAqhs9J1EMy7uWE9Q99y/w6WzURQP8N61ZmVD5fm+pgfNv3ck4RZ6QJVY+7iaib0
KZh1dHAUdWoakMRhAwfwaE6HZoBjrwzVciNLNc4AOJBGz+6tkGwI0FohHKA0gFiAEJ+msQPAMoSM
XZPkfHmdkPZz0QKeVHOE0RzRBjyY26KGjf5e1iWR9yWAOqcgpQpbWq+9b+uVUI/WWlPFW3oB35Wi
0oCtHjsVWwk8/JLS+0IPfrM8cue6YuOm6ryedr8JBx47OUZ4jUNOWaq3JobbTN4tROdyw/9AecmM
20nRAq5IoOEAokkQpl/34clS9xUiYFLW1/c/FVP5Rkh3D5XU8JBGO7wUeOxagEY50w62hIIkND2w
3N+O1BEUqV/TFoIVNIyz01IBpwD7AP+TcEnzRWtQPvlO/2YTMKBV3Ns6F1EBP89pMqeg2oRuJ49x
NHGwwdjzPtw8TQOK+ldx0czPdh25hR4DpLP4radhuCfHnXCNxmAaZEzdJFmFtMSSQVjOj54BKHGS
+YDxdFYOEPoRC8xadmQGyhT42Qp+jcemyrP1wATgPR1tCYdlfodn2s22TfQVUNQx9D4WKQQBXZur
DLD82xC4xw3atKbjx81BR29Asp0ncG5SHnXiqK7hlFbBTA9+5bU9FtaTq7FFiuFqHjrmaPw8lmF4
XrZzeeUkZEHj2n+s0RgjPGrvD/zet/cvx2peTrmbGTBrL/RbuZ/EYEMjC1I8A9LxNz3AzP9cjaPY
rgE2pE6KlurdfHL7uGGTED7AQJKi2fhw9qObRzWBll3l334U4T6YcPj1dUmAHPUTeSgnYLy0BY5a
LKoS3/jasjsstCJDzIB9OlMSMG9N90gJWbRx7mwLj3QvRet2x+i34Q8QpYsRU5TdkXAH12bSyY5h
2T9RdHESyhVfTEpRg1ZFLnn1eAomA4Tyckh1glCkfoG43nlJAQohYuVXcEkN9GSqmsvMZUIQwvAc
edoKMfw+o9OqXDolhMr5J40szwj6poXkS2tlf3DVnY78g51GTZLcRj+456WlIftTqNBj8zkXDml2
YxkLH0XN0wySSr23vUHFQ4Z9GCdsgVODOZvd0Rd6PHY1jmCNpBcElpUmq7r6fTzdmpoOoeIG89+x
yAv89hu71SAN8FApAPiwF2FbsmY8XFDGs63ifcqMlhr+HPyzvupQXGQXpM83+bchcxLe1EsOc+9p
UzctEPeMgHGHUfUALhN2rlmVvKR/zZkt0RK/1rHrOWBXf2M91MVhDtk7c2Aj4Ns7BX6ePAGLFFD6
TQFeQabuNdmvP+9SJd3WyJKAWmsq8f5HKEY4HoGR6pmQIo1Z9K9/hWNZyVjKnuZGwNdoDPtwWoPy
cqX6l8vFPjzNSq1vaTus8gy031XTLjrV4NWjw1M/kYvO/c3o6/2MzbIah/l6INRNlrd6S1KtsEkX
xClAyTBkJDo+CNDeI6exi5KsauWUX3pknrS6CXo5b749GNAaxDp8ay1ZDjy4knJCRoaca1KcoUTK
YkTqmMhVfFWhF03ve8yDlyTZX9Rmqst1X1k70lgUYlQos0UU+MD3WxrfH+a8xZxaHLTQfFtmm35a
jqEoytT4cmDwb+lJ7HRusyH20fZ6sxQphoo4ebvdDQ2EoByMTqro2DhR9svuojR3IOSuplfHmnlu
vcdtPcgIforUtehP5pZAs6QeJ6+CX2WB3T7iu0zX/HJmHaYXVfvF0EPdvaWfdEZ71HfdnU7QUjLb
I0Ybc1yO/sZfh7Ml9/RCSXmaRzWD/ztGuEBaurWcMPpvaSQpfd5ZCmG0odf1R9Z5hBjshbrzML8F
Sl0P/OGByJVpSnvFTRHelW3JaCTIdj/eXwqe/NDc8nK8Qi2vW/WvFlw3qHq742c49miTQjAWuEWH
+oa6oTx9v8zkJPZPjvf4j+PzGw2VYeu08Uc0AxqkYuZJVIfwaYEmYXrGs5rqkJY2CSrDajYaFcMt
ZXdkEAGjZfeBrdjC4crnkJWuCZaOfa6FsDDzDn4v6cXx9XFAOF7fSqeoRRpOGHNhEdk/j5BFvoKs
X+AFud8xSxQywfGcshLVyqqgJ4a4r0fWAflYtuRFP3c4gZMOUTwhR75l6fmx6XvMy0XNHVwfUJft
56DLXAESDJ+xH3DMP0Qfne2zQQvY6nzvqJlmY0QJdmxWvBIe+eMh4phm22RJibn9dpRCummpfg+i
vJYzWEnCDNqoVqH7uaQ+/BDiAQ9h8oo7rig4D5QL6ym0PvjJmRaV83d9WuniemfyDcsR541tp1DP
LHZ3HDfRRWO2CHHnDNiwM+3Q2ncMe23Hlz3dafiCTDeJnwLV7MAB5hw6tyVVHbYgmEv41oNg7Lfz
96A8AeALhe76yE8mVGJiG3L4k6IIU+wjb7yJV3NGrUu28BHJuhdLIPq+5ei8VW0OXRxeG4PBu6ay
K7aCROWQrVhrmMLqBIWDpaQ1AYo1NAmkec8/JKNDWvYFn94aKX1761IXtnu80wnf9D4gwYjM3c3N
/oRW1ofbhv9nr/fpDxJ5e+esr7FDK5fRrQ68Gh7xr6W68W7mXIy1dwLTL2+YTvkfbO97wrJ/Bfyc
ZRpxYs3zrXKdIy+xSVas3WnyPKZqVYwwoIUtEyiUd0MeHBPZmSdRP1R7Z7FLsk+VnWj38j6Cqitn
GkfzI8Z7JVNL6yANaylygnhySS1qv+xKWO6K71mAeoABrOPmqhGwQt62j6H3rmQee3/740ZDtJdF
mymIpWSpJ/6uGV0634M9OCO9Osar0Er7+z/WclRexCWQhy6NQ764fbUCP2wXodOA88WEyB4xDjGt
60TYcU4Wgeo+KRbu1BY+Fk0TXm8FdHYPM3p+E3UWLMonAlQoGghq7OHpOiwJrp3YZljsYCvJdPpm
EYUtaXn9W2ukC5h9WFNpjX07qo+HnEWzqJAXC91Ika+CRmWdpdtr0N15iDllU7hWmLRJxWMASN+r
6N94izLGxj+y49Ow9MM/U0VpFkLmDleeWlpvMDmsMpE5AqImZd6ZAED8xcJf7TM0Wp8RgYXFBSsW
8MU97MUSH7j6JBGRI7bN9eVACWcC5kStXEqZByXIZHqZbrrrni7MgXSEXtorBJccBVUorLrP6CNi
bc0kZN7NS9clE9VQb6imrAZ6cCcVCnrXrM9DGw5twfWF7U2jKHij4FEiDIkYST+H5Ign6tXkg1S+
0F93JzRav0ZieQcbSnJTj7oHhfL+Q/1rn88zMLQuF4N7sVzUgJq+YbEl2q28J+GOoItl45aAJQlC
krlmtuCYA92JuavK1/5ROV3LvTOeTNai6GR+VAnABt3Ab2zWWONIbL6KeHAEdODM0ghHi1HfsE2n
Wq93k7H39i6EzlB2XjgTtccwY1qn7BKmtLw5cdTyOxMzbgjvD1EnzFt60FVdR+HFRCSe5krAUHmP
aUyGn6cHoYrU2vr6+Q9kjW/LOXaiqW+GiJW6lU85wtsdWKTWWpog6pLslwfoV+SklPOCteJphl/b
yKktWsx+ysnVsiNXNiHPJwN+3NebPYMaFPtsYUOwtjTga+gL0enF/eLlDZmIR2mqe0Xd3HxKbDCZ
66conb5t9oNDyXHDA8kkwNyirJZRUrxToYfzLnlWQnIlV2vRrW28mpdmFcW1fxEQ+4ZZXi4mkP9r
IkKDPuUlC29YJyn3OuEjgSJc08I9PNCq2ybfu1tYtjWvTJFG8Lv2okgmYRLBIheGHdiWuZzjDYWy
Hf6+rmTM8nbJ7LOpJRdimuyt4Gqb4O6+0z/cAYMvRHfLaJvxgkC+Th3CEGfTMGoP0e/sP5obCTay
vlUNMnAujzSjMclu3QoXZa7ujCZiXxTIEa9EVJY2l0NCcv1gxDtksKuF1RPJdIlqY4Qlg3GoULlz
Kqn5+Uc1ecQqavCSBPznAbSmD7Hvs8cvTPg3es08JaqqnquI89ZYCtrSPBiNJu8+Ik/bY0Svt7RK
Y1eSsPlbfHpl7BuGdNvOEXsbkNM9+Sm8aPw2Him+/b34wQfsmNhjddbE2SGew1RBzVsFjQsZGG7A
oa/7D8JDp9UWCKKNRG+sP7mL5TUR3uozBcpT0yxcps3x9TxFEROvg+c+MekTeMhD/iy8+pz1Jjbs
2+a3BjO+6WbC/ENWm3wY90/xyYEzwZpWAVUlB7k59w4r30uIyGNZkxUjfU80LUeHGNQ+5jiRIJEu
gNmFUzrUl2eUhjfbDmN3yxXR0VyoqWPKsmVDpJaeUu2jO5YjGry7iWCRX7Ynr1GPCGtcDN68UXLP
YHjS10kdiKWHzags/DGbX9V+gVS8ijcCe0Jj0iTw6T8p1ucxQVDJfk2DNiJZx+BZEzuAyCmseGs0
34R7IlJTnAcAImCnOIZ9DNm5sz2d/RTvjdHaMO+zLSOnl1TGm6/p+FIuzSnt8x63YMmJbkZx4+/R
BB41ojXbCvBs+7hORXaN24sO7SB/GnHTMz5mGZOqi48dE8nnLUp8tCLaUK74NlgrV6R10LVtZSII
yilrkOHDLb0UiREo/9uUcUa+EGfws4VvcS7T6bLqOm3bOg5aWhFBN30lAdf7FB29u0St1KJmcOt1
5z2KYICtankI20dBcpYV3RVGI+OVKr42UV5FjN69cqB2f+iJOWIYoFjrOsekxrxbbhjy1vXHjfm3
6UjCPEm5CPB+qEXcjNXqeaXwu4XaRenSXPZFlB4sNhDq7wL40j4OVrNzpFSI3Vy3pWR0KndO4vGK
mTm7YueRLagTw1oyf6NgQMUGgMTd3efhEcquEWasWxSpM8X5ZaFMnklGznFJT6B+NF+JTb7NVEYS
/9B6nTwlyD6voZpbOcwh7YJAneJsY7hNy28zBM0bJzVQyKEYXtoSU/eCiFg6w/0T6MMcFgrLiJfi
GG8PRKgrlYNuIYwaGdftHueKu1qFH9FLpJr7G2SeNZplVBb7NkyR75QAztkd7aApXbmWBGluOso9
hRrvPR6rwp7hmed7H7nh095glpiQP2Wl1wu8PD0cMkxIxqLtaJWHkMLXz7IenJzjAiu+a78zFEia
2utJX/OWKOPjMn0GRAQ5xmpg7cRbSHXLMkMOPcJzY7zX7qPldFSmfcjYm08RMfQdJ/d/sp9dTDjq
m0amlIhjxlVM0qVqIBR9A+uVTHbRY0SI2e69ylofrI1G4G3QhEwyrDKhDNvbldKZ4X7xfkOyF4I5
r6fOquPOl5WjHTP0LEzq4yCEB/hcyoiAcsYaaWoy9WWYEfdh7jI57lM9mvVXx49iS+AGUtSYd2uz
GryUxGNakDq55tlwabAcHcjauzsIpm2KKR8QbnbnBS71FcFSWso0cT5xbEA4c9Ver69QZDsHLrio
Dtbqafv31GceIMedofWIgrgP+qMYflc7qu0ePltAP+JXe+qvOiIfQtMUzPlk1o7ydwedLMoX38ig
091xA2JgC794GsBMlPX830qfCsUEyy96CjXSjzonc94fNrqbT5iuYXy09DYxnCO1D9FmIRzo2nJC
Ozb9S43KwM+rGL1GnTXoVxylKDXVvDTtYyfow9KlgBkBWurkBnCwxWiZQjzQvfWsL2U+1OyNduvr
5WdcqFRlsFLdHg0c9ShwQhyvlP9BMeoAkXDO/QPLONUDJI+lI4m4eZ5df/TULm8UO0Mh/gdHa+vJ
WGx+MQk/MxWXZIHjFt7TbnzIYNWYX4OJmRRqFU5UrNLR/+mkpFJyMeWLtoCDQSBgk5Nr74hOee+w
3qFzxFtkxhN+on03dmkJjhQJSX3xU0YTARdVpVDJpLiyVpF7ZAfOTwSDXH+7K0kY/NXV601byOdq
+jEsvN+JGun7idltRSxn/MVagTlrjG8/xudof2YqrvMig+dmG2f5M1tvXs+3kO1P2SNTRj0fRIum
6CUVKbu23RK6KaZo2VqGCD5LgG+bSA+wgYMLPkJXlzSI28t96MeQEitg3ihrLGcbLnLkk4nxjrs5
Y88itdjku810AGyVXKayfehTE0scncwSmyg7lywzKHvbDG2j70rA4AwbVOHS3jpBwsgfRTD72pY1
pBpLJeJbT1F4XAjTC6PDuuvCQtsO44l2JLvmd9H0qoGt41vbsTCMOkmokcwIlGGYyEZpGG+X5TcX
UREW9uxr7vzN+nMsRLPfUQYZf+fbWfKcOl9F+dYM1wUCc9ijz4UUaGydExZBANzNDbTTZD8TCaTX
g9J1etvxXwwUqlc9bF6/+rRF8WHQWYET/ZmHJfVarlC2T6dXD4qGiPCeNP2mQEZbQ7fjaxc/mDeF
9Sp+lcb5ylywUO3qKIqWpiJxIq97CgU/8htvjpSNPGvT0mq4mvEQ+p8tXH1ATiv54UT8xbVXAMLD
G+Uaw1fiwXCswIbo958QUbVw1d7yzfgikLAZm62SNh9Y06V20BilmtzaKibyktyq4L09m+9k2dY3
KxXhKh6fe5pPFPn/G2wyLGQR1hfu45WCnvDC1zMCk9xuuJ1t2QnpMd1bXx9Ot191gNON3FZ7HTXz
qQZXqTKn1lWmFSvURJvswzZZK6yz0QcN6a85BNOffMA/Gf9XzSEWSZWyyCJ3Pjtwbc0FYOjP/lBo
amZ4dseWOEjSbkfLcsRdWG0Q4jmPH/kE5BlurhUEjwsMMuCF2okoQNylj8olojCJRsQ60cRqdVtB
V/mfGYvhVHhgvUShVEuORn8/uGiI/oqfyOQi2CGeGF/LW1OhGQfgJ10/xl/C07G71TDNuEFAdz/s
58nBovD9ULk3j3REPrE6gkxqrzvzV4NgbZ+6nc3jfFm0JwjtIKb2lq+tmDBSzkxp/GFpsCpgGG8n
1Pb1H9mTDepRaYlZeHozCaJlWJgrFdDJPWsDUdnE9n7Tyi97nigkNR/0Wai8J6L51+c8uCIWP9FG
bpnvcEkRakJAFkvMGblRTivMSccV7N67gGEjNvnSSvGS0OuoyE6W1Dvy3nrSeNtM68iykx9SNa10
yjKji5gxpZjf5MuhJkQAJxyMmqqUTKyKudgd5mMGjPzlcV9u2v4bPX1vGHJ32Y5WKPJQwvMGcJbX
9X6ikegTWlFto+k5fcVvCHb3hn2Ti3c+dZbpl01SJZMtoPnrjYpx9J/UZ/M/OpjQ0UiZ90mGyIBw
i2O7LvI4o+UqNaikeKA2AIMiOJLHr85YdPs18EMi+/6IL27PwKp1J8THa/mZFftFH8rLKnqZiOma
1h2Ve0d8ZkmxunZs8GFBRhr0joZGePmB+jQs/g2JFe7T6hV1VA07nHCysFicaXQphhUO1EfqKu8m
rNHux6PGiOR/S1Xh9x+KGL1bWkEoCxpgSGsqWApiov0t9ma+x+oPKCWlgoWXqiIDc85W7vXiIoDE
UesHfqKQv2ZKmvANJ6q8UuzCtvk8eEt1jtfOKe3ZaOZjp353onfewAmCcTBfQ4CpLeLJJy3ullLR
BeRvVJF8mrTLT4plsAk2XgAna5QIKutbKh2Q5UBOy9uoYWJKR7BJ/SqKa0Pv9sp7U9cC6AD3XymU
u1S6d7sp4IgbZ8mdtaPXbGjMt4rqJFqa89OC0gZ4odLMiciP1IAK4mS+rr6/obqGSD+cl7iMbL9e
9mjZoT+tY+CLe6Bcv6h8EA0VUqGCByDY8/oL8/EczEluiWYUr1bOEYz8xD70D5/fMq3bzzUhHF+e
qVVEcbSYm9Co6PckNgoG+MtreNF4cF9j3IO1J007TwW9/5cratTSOYDLdLBUyfGNZXae5WRkqa7t
XJqnjknwRRZllN102Mt3btnIfDYydCaJteLfVuXihdyM9dknxkPzm0JaxQrMmujCfD4Kh+0mx9ig
zrgW0I8O5auGExcYOoP/YTlWOH8BRrQX+lDd4rHIoEEimHVa/HnwGPTXJ8gXvcLcR0HMvhmOkWDu
5FaTXFP3YBK7boy0EW/vcCJNANpSQFwTIgfV+WAsQy8UdA2Qzp65FvcvmfYgGHwL+kACgmijCda1
s0g32na7J0fzCvzt14/RQ2Xs2CCt8T6PgDxfBBrR8MOIVf2WPXpVf28PZSN3+H279FcXVQ44NIm3
sUSxGiRNfDDPXzdJel3W5539JXzQKLCrtgZEuL/OpEVTR3jG/W/l1gVR1F16KYZF55mJC5FcM55Y
3odOdIjeAiWDDbiaNQwRYcxOk9siLr79SDH4izFJOxtg6nMWF7Xj/sDFgTJKDeXGDYpM17VqS5A/
XyPnOAf1RzjKR436rqt5MW8m1K4sTmcluQPEAaGN3nIGBz4gGTjNJjL4XMDlk5ofB42w8+ZUs/9M
OQkhq7cEJSMExN4/lq5o3+m2kVOsMf/Qz8+7kepi8mYKJkoJ/l6Nko36jgRbiUFEbtvANJtmyOwS
dksWUYELXyE8lDtrJubTFOEFdgUBmVmoOOLVIHbHoqlrEokaWM2YejT9GvZD6DyFJrkEMCu9bu7Y
UAobwYdbx17IkxGXOKNoxLi5c5fPpoU0nWxaQk+U5i08l6O0p2Q1eVEqPfbXEZ8hUnM93u0oyKot
LuiNBbaxur4simze8U2JYuhw45vTWvkyAhNvPG5mKgsguRuNFqIVK8w+FLucWJJ10kOGAqMux5ft
UFF3mVhRAW4LV/hZGmKSi0YVT1I21VcLFwE4r44e5hEwj9jsjlldg1RAqXwZz9MochoZ2pj8iSI6
xfiNvx+yRZjV5YVsvynRxRoLCYMS22IP7J+9ecm/4HYgkIOBnzqzCE+QQRIXdjFz1Gq9MqhhH3Iw
ZNeW7Rc+kX6CNsUCeB/fyeg3SizCbpWOqo5kpFmtGiU7yhr3XbjThRD+OnZ4taAPvnnVHNXsSwXc
DweeruI0EknSgVHzl6H4fTeqG6rbdcosyfZxnh6Y7wwl7vwFHS78N167SAC8YQzF82RBSRXBPGwm
nIc5FNtjYveSInfk3NDGH/Rn7sAU9eb/K6Hm2wDkWQqjuB2pNYFaTkJKySnbzrD1nrMg1DRyjzVP
kVVd9xd5bdncCLIvhlvQT9A9iptWNZ6YIz6MneNFjT5xAbQCxquVckO8N+S1SjY4aSMnxuSc/RnN
MiKEWywobKaTqoGoK3R8Iidlw/GCHrZZ9pEn9L/yscNo+F3h95+lFucerMR8m9QFb5TiGhWf8oN0
2cMf5Xdn2p422ND97EP9G2P65aLOzzZstJqF7sIbVgsmUtY4sTm1QRjKSpizfdzXbHtFUwLp8n85
X6ijlpclhP0hsGsvg/sCQg1vrEjV5Q9TclDu2yVYhTAK8En+zs4KJdZWhCaZfuyCUZYfcWAABSOa
3L2/ZemCju3ledDYLdL65buCU4bWw3T+L5q4B+IQxMEJK9f3QG962pCFi7wT3w8+Sl0jREtHG1uS
+b38cLm7OKUqxms1uaibc9o2VmR3urmJkblJJ4xCyw7C54UwZIgyAka0rqXLh4fyOZopPvM8cRV+
y+al7EI8FpyBf9l5YrPKvsiKz6PlZHLw1+vt8ybvYwyQlMdAnmMzgNmBK5muw+ncRcIvvx8ATF0u
ZjG4q1CSsGrMpz6EQ9IiFdugaGxjpii8rLQNacSyJLApYH0jnAJj6uBvPpVGCuamgaIIzvNuIYhe
O6WlNY7sxjE0DQcZfmYXMOuOPrw7lJQ5Z0lpkrEUZVtfKqoggiDIKWNE/0nt8AyftjqiPAIZFqLd
+5vSmehIRdXa3+zEdwS1/yp9r5A17lIRhBDB+tbCi5oB6KTRqrtlxLGAO557IUMBMtXRIWE5rjAp
ej6QXWp6oKu/VAKoAV/Zoz2taftdKcTaIev33xqzj/mIcxHZwpdwzva8ymFPGJ0rGk4oX6NiT0iB
P/RmZcvwDOzSF/3WkjvGHGYptP2EdfmKq3yeZyKWYks7uk3Dza5RFbQ11wSl3CRsQ99haq6ZIHF+
NbIHpnMPnx1wpCFWy4O4fRGCFUI+d30hD8xbbesv8oANgaWbZ5QBOEl0p+neks3ec0pJIU07MA8Q
baieFKwq4fCudpN0PsuwooP1o+5Q8Pb6E+yGQAUmAau1ySgPdwsbxCKBlaxTmWV5oi4z2IV8X2DH
1Pa9F2K2C1j5eG/JN0cDJO+GAwJyzrvQ4G+CvDpVPAFPZuJgBWFGwGBq9gRqKQyOqtzohF1NhZuf
0auYNPbCv4Uw6WV79noJJ0caAmWkm3tscInTzQzAJteKaj8eXGTsKkLmXfXJ9nXGtI9gFF97Y2VB
KbXfl4kNgRKAQAYGxWLInjhbtUGHjQykjQgp8vObFdSMHDdQ9Jp8JlNauCf1ZlFK2BSIMowhbmKQ
6m0qtA5EfN12ePzjtX4Ed1JmGTNLmxgTOJD4N8UfT+o6OVrwUuRiV5IsD3JRE4X1rbirRzlfukzh
wLdg1Zqi/SgQOPtfrqr9ck9GRdlG4xyvAjLvG9UvV3dG0Ol8SNwjHXfTp/A+ri14XpvbHR1AkINv
SkXSDcpbE8lVOgJ7jbaa4PtYDptqwGYHQ9+zUvvvrxLliZTGhT2V+guqQbj4xb0nSXlHTzw3RtG2
TAkIWYuBciUbmX4ZVje/LfpqC8wUHS+J+IsCyNwsQGVnF1EroID1THDw1GJNyXHVO/BLnG94Y14I
NA7O+le/G/gfTJgHCDJZ1emAYODi4JjW+iBb3T1h/R5zn36x1CzmDFNCG0dmcPOczxTysd/EA5ow
SQcQMVmNToQlbKoXEmJVdzonBaXrg4CKxxLGdDB0fB+CAFYEnvkt0azEECPam4kBmltX4qqltqyB
J26k+3yxmW3DCYn85x5xyXgmHiXD3VKVZwD93gVGbIm5GE3L4KwORaVyPWPDLpFGBqw6TtIJSaeD
ojklH0/Fg4gXY23IxNnFsYKqwl7dBiviRe7dDNPusmSZnhQPwXcYhHp9+ZQKgNLqPmco6mQ76M5+
JY8pO9r32W4rIb9zCphVlJcAwvJOrMqehCgxH5gDo741Zdd1fY4QBahilIcJMjDKMNk5NMFnG7aw
lIoRpdhPgR3XS9+0AnOo/0jecypS9JLiPLwUogOSn6r5MEmKS0cGD4jkEaDoJuYmXsiP8JbaO0em
VP1uHqon7yDQyNAxVSAkJ3irhVJ7YwZJHCbu1viS1pn6m4S/Rj0yQMljNC1d/18PO282hec/15h+
YHbykVpTiC9xdFqxYODfbX8j2GHdnrJURKX4QekRaHdt+MxOpaOXFUrOXlfyjY+nbH1XPPEXDzv+
/Ts2aur62QrJmG1eKJ0LCUx5DcblMvEOEFXONwGFtI0cVb1swqwZ5oRCSiVeAF9myslmLNm5iFF7
sXNEzIf6SY7d04MWERSXBvmguBCIFkdalFLmzgkVwwJT7wqkqaZXKZYnI6P/vbTCsVlOHuDYxMb4
J6jC5zvw/Q6eU3Z72kc6lkTIOT5hnvXZ75ez7zbQlgl30hyd3Jh63k2I/NLIz5d91FIP3XBqOCuN
oBpmcHTEujF0vI3Mhdv/lhoAM9equQCG7VIkcoO7e/aLRKbYOheI4TyW3kaDzIql+xX02lA8f9Yx
fxHSHEUm0RGAogaPqyy6VF1NTanGZX/THrfs32cbcFtXTlZX7mRvCoTVPco/O+p6Zj6E2kVVOn3t
ZiuV8yiNjwVvH5RyOLR+ER50VN9kwPo2k4VzbiyD/RLwMEKMr/gIjYO9C7s7puSz9yGaTznN+KZC
uBJG54VrYotiPRFqtaUnuP/oTiplUD85fpuMqdWf9p7h9X8lQJsPes/NttDJQ80CVJZHO4zUHKBO
Qa2PFBE5Wrjtx+veqa66wlnxeb/MBSGz6RGUoLKFZ8IyM6eqDPwWV3ku3QeA6MdhDzQL7UePRbk4
S3dmpnbr1F62fNARD2Z7AajxWPA9pifgg6Mow0FfNmKdsgka7fJ1Ba271xNKVh0hScmqRPbN0bSs
7IyjbICIcqkzuSlpREaJksjUnC4gBsMLU57BXaSEgjWDiqsl7NMeeU8L1FGAfb95f8oX9CFGkSat
Mie1888XX9UiNFO/bzpSdkVhu5mBL3P85siAKd7LxEB7k8ZFPSAIAuI5Hz4V0C8aIKL1Nq5+cWH4
KPcq2WyMlYaUtRP7I1ailqjquX6fhrA227BsbWgh/UpIHQYtcxn37+rnbjkonjhB752crBDlkLYK
NL0HIw/H0iAY2Z/7139iS34PxBBLGcdcm0k/Ltn5M78Bk6uGMwKAfy/69UXHTTGoZesTMtfnGJdh
UUhxXxHNkYXw7Mmg9TinVxSZ4Mo23LecMMFXQ9xlx5WdckcKSJgh+V+LTq01MJZTSYF8n3iP2z4Q
/pxGXn3uThv1ib6Bjk0wuGsql8MaqHKTdRbKI4qzeHofTmxUnQjLxYGz8+ZekwhBI5gQiZX0h2Tm
ydsxQn8gkDokcbPYKwFIKd0iJOBpEIW92y81eYpxTcV79CKcpH+B1XCBRhGCZLFKw15IfhXl+MQh
GMndSlL3JK5xqJEE2YhrH5RtBKPXjD2X/WEk4v9U0GWPwqk3ArYBgDPmaJKqocsUu+9/DkIC/a23
XNAaBKQMb2VrVt2k96s+tcP3clkB/H5H5MdxS6Ki8sAmQ8v8IyACjYpKfkVoQCwrmm5aoutWGm8V
L1DXyXnQTYJs53w+ztBm/aG/ry94fJw2l5iEIcT2M7OO//usN1CB3UKFa5gNQwY4SGDwYIjDAl5e
FRQfPf7Ypengg51SrOr/DNJMhn0JUhFnHyrPiOHwlA4CPH517mV81b8+a/2Xtw88+olrYjfoqnUd
ktBRnZBhpJ8b+LpiYyyDRs23BOrw9shMZ2Uy8HyIPqa/yrkhYT6fI8gi7bUNiwB+hfgcq09iQzzm
fKuUeOsSzY1awVdqKVYDO3Z44l/6dV7pF6mIr/3VlgGSC1G5iZBkvBzFwtm0ETmuH9nqiTubyBai
hgDwwGIvyZaAE91hI15KM6gJYx9N91j0j5PD3NNcLegm0+K9fB3Wh+FZnUtAHKGs8HqxBC7amWCv
ylPrUGqWH4WOKTXJLz/ORtLVtpNPQZLh0lNUn7MIxAoLe5LY1JCVUTzUceotJmO/6cQa/LFFgoG4
B60Nc7CoV4FWObMnoPw2xBIdx4mM7Tqm6kdq/U57ooBPJQtGu7zym2YWwXlFczTWFRKGlW/Rh97a
696qlEmH/Y9sWclzz6HIL9Yo3BioJ4rXgo4ACwz8csKYrAKlmv05tSBXYsVQ1wJlnwMXo/H6uG4v
3TLMa2aRrlHwZ8ec5Ii5Xabi4UP8WqHdWCuppH1rcRuu3+VZedxLA1G4sjodp7CTdxoIK+jtt5K8
WXbp0UbwhdmnAY4XNB5z6KQlWtHgft+Uk+qi9N3u/xX5VxwUk/WBKUdxl3enKWHB9l1PkrFlKjzx
3YrLHoHb7yJNaaOmJn8Q3b3np2ppcAVlNluWGNN8Ug8XrzDIWn1tyEW/zH7+v3hlsHsXEywx5NME
Ib+6IkzbJdfXKB70dNBhMZFuT2snmt4hXzrTnRbHpHBkp/wUKnzURrKeicTKRRTXHvJvS8kundoI
zbUldj9JWz5VNkZCzY6VDhe3qgEQYz7WOe1t/vFlHKYE6Z0lZP1t9A6xzll9sR0NUljplIrYOgfN
j486XNutYrU1eN9oiqlJwreFR8JEgKEi+YoY8pn6TDxId8iqSL9ixBpUz0QwjJ2FtwkRPU06fx/c
r3F3ujI5reFiI4u222lg6U3ZLTC+KmjqBYpHsL1+YORXFGRmu77Qc/MClKhvy+m8G7ex132/FlNq
eSxC+H/zBJUXGC6Ob6Px3EgwHTdGe+jinhujp4clho9sU8IN2Lu4mYgOwbdcdDS5AUgaz/IZZ0ZN
ki/bfAYYOkTQujZh0WX0Pgj9RstVmj+/CIc4Naek3r/yuYfBnmRr3qZZDBzlCbaugdJSPKZKCt4/
dRbDWO2d8va901GesFRy9rWpZ25W0w3s1Lq4Jg4r0YGjNG8E22jvRUx+O3WOPrZTVdlPMI6NSTg+
jCsEjUlXFIPyXv+45xSYS/IHZFjdVwC56WJC43TR62yoXXa/NPvYe5E1vmw7q9/RwW7odwtaCefH
8p+DWT4AZDYBQbzkJzUJhYWczeFpVY8JSWmVMd6EVioAzsA77xp9G7XbbR5hAp+MZWH3EW7Xff0K
lGXosbiOsnhBQ0bTLHSRtlL0wAv2kFrc+geYLyk9dkoAfh1ZxHM1ZPUyq4Dhk2o2bw8xSsWhXKrN
Dpsr+cuvIqgf2t+yPwCNJIqDp5m0UVt2hvMRYLmgDdmmCT9Fj84ruHQeyxry4YDGbGAuFskkfO58
l33cmr42VvAJB+uUc7JHXegpYOULmCfWzpzIVO7gJ8IizwOqr0zLq1YkWjxALk+r4X4Lsk60gYtJ
WPJ3TyuvRnXXfHi2H+XACzIn6N4E31mgfYYxBkkubDJ3W77xs0m3tOC90gPMChD7ZIChB9VmJ/aH
BWakLGjGWa9cox1/EYgYisOtIgQU067Dwdkv5+RBpFaWtN7TzKKL5smkEw4RjYhR7FtCXd6F96P3
Uc3c7f5nbCdjWy+kODOuqSQWlL2Z0ku4TfzDQDIrykNi+B37LpqDdnuRzqTjFgoLq/8mCPduQ8eJ
ZgeV08LUj1ucXN27sFrs0u9WGbXVRcWtn89JVz5NH5DttUdntqTtwYK+gRoB8DCTCm7cAYSdqFAk
8j5dHprshapitmhgCwzGXsWlmeZdLkMNvURim6lP7pU9pHFNlh568ChHLxZh2dVvX8IRuT7WgolE
+5aTFeJ7PSdIOIC+E2SUsSR5oZEDBP+RXCRtMGqVsfKa9nTuwMFETjE2Od4ExIGjh/2ZO5doJNgP
GT/GkjDnBMXmzHTEAAB0PqyH/M15DSmb2X89r+zBotlMVQaOEgRfAeSfWZ7oe/3xxBMDxMHk7tW8
1h+4itksNVfIiwoQtHsLUrAs3vHNLyEL+4wE6aM6cHzbl47zY3UTjH3a1BSpiP7vHUchDe+glFmJ
4WivSq+7rj+P/1XTQ1ujnE0VEP16fGyh/+q1E5TrUhtfpzlAFD85Fhqo5wCov/iyz9BjIjK39Mw1
EZO3t6/He2ohuFnwGJNvqzbzurgLhNVr1hScm4Uq6h/kCu6rIj9WBBhIpyr0C6POexMc69hRI2h/
z3I0vYXsNKa+JQDaZXJqbanfwvM0wPlcHePi56q6rjTXxz0lNZlSwF6jxnD8oAUsVaedLDPMTGt9
jFqvYmsdKpaBMQc45dL3IyKgLmkSJYpU0zuLrEvTGm2U5RVkNDm27ddxl6l9qJrRA8L9M3/iMnK3
NtDkh8KZwEkS3lgFQRfTqjCaMCldAdPaCz2UVE9Nc/8tr9CEE2Y2NkXAFASgNsLWW0FjM3SKJBzQ
EyQPPIt9/9MoWeLlBEk5/UW6083NuSyI5mmHKTZ6Ix2kENyGlDZPi/fRavxJlG44Kr10xwFQHTgQ
c2ZoKto4Zwu4VzlNsratbtaQj+P1H/mWtLpilejLrp1RmKnokbGNL68FI+zvdRhj53BpLvwDMId1
+dGGfVcjsnCEEb0sDmv5tAeVoDWg4Q6Ovbmdelk0lh6wWA5mcE3308N0eJZMW4OAhq9rZiseCJJf
sxVttiPpiRxpihSoUNYVzGgWijzlzfPc141SoJ1ktGEStVGqBhpmQISUlpQQSEvS/jqqu+5WGz52
c2WTJ/Ojm5dRZUKFYBOqP3eMdJ3iivYbRLKaIyEFmHAqONskmBEcqZe4xYMRo+WfORVULF9HTHAk
exiiB+JqIpfWJwixgkf+O+uD7iR8eEz3HTUmuz2aCRq0HE7LtyHPd55rh4lOya9IkZPj68HKl9/U
72aQAxCaDgkS2LnL00bSfdCY6VCtGe3gkyqJkOtoavjJKn0qlqkC29RCjPW5bpJ3qKemkbXvgVG3
zg1/jOksQjmb4wC6bdL0O1YyGBIhMTXKm6SE1oHkADdA7hgpREWvnHOyacB4aNqV6CIHUxTqCOZS
TfU/0oxeDHaItlE1Kl3eBuZVHoJ+FE6w13X//gTfDJ3Db6PKGTyNVHgM7YbRYo8zG5Dv7FNPyh+z
zIvSI3RRWGHwdbT2i8ZxW+Jop/0fsFw/aJT1o3tap28L9U807lrc/Mm5uWqIot/2hupsun9wHsJY
RennsmcZGOOObO/XgrjGytDJMREEaNq1q77+QwKjRcCbSc/3mZu5DtY0Ct5gr565dA9oSRYxlZ9D
f9skOVetZP4DLV1KUj8oYgPYgvmdAiGiCFuZz39fO4wnsoraNmYOIMZ/HcL+cS/FdWaekHslKPP/
ycHSVZS0eXbwT1Ql00fnLqcedqRUp0Tg8cCqs7CEphPL38g1vCBkiY3C3DClCyeGy1qnySKqQ/AB
rrp+ZGtjO2orsgpQcX+E8N4wQrIX4g8JBq9aT7YTzgGXq1NrnPiTZ7fqnWjlzEksc4mSJN8gHkNy
SBNUrTakU8dybZrM7BA35iwVp3j5/vFyhbu3I3PDftpr12RihHhXlwjdNWVcx5nU0dBPQmwnhunh
ilaYbnRqgMp/OT9KUtZMEOI72S43sFIXrvoIbZOyOskm7TX7AwB8W9NZ29ypVNmhfXInq/oicOWy
daqlld3dts1WupDHn2juajYKMWg3yBV3ppy75ykM3V2FYCo1xcbX9D0tBMIXAgbeMBmPmZ7efhAW
TGUmTFjsi+PHXJU3p3Cci4qe1yiEyhDIrEMo2l5BxvrdDawrng/M9zhNK+Xq7iiGBJjHGDbW2een
QOIk1weL9pIy9PnX2QCihzX6SJQxUEt7mSSPULNfJ5vs4+sqEbgn5yUPBW51qHWhGBNsoVe6Qano
mDm9c58baUW3G7Pb0y2g7p+CKjgvT6sJznvDilk9ikEP56luKU+vHxWotm83V6soZPWCUI+xPqqN
qaHN76Maute3pP6x4nhTsygJDGaEC3C/GinigQcnH1Ud5fta0fx5AvVub+l42a2lcjHmGVyK3zYH
kuIhMUvXrn/gcXFt7OJsEFjta8/FJ5moULY6qnWg2xce9QE744O1IZXXZVOjp8U5eO0NCDceyYYl
SvoQl3yLHTPWCjXnLwKtjwp+83izmWLAHmr6KmFJxoctfglbgRhVQOoLqf5aHt42Ruhf8oJoKBL7
2q2tqIM1dchFlEOpu1IbnCdhAZtvJT7o6YvAeSDlUEY8stQlZn41TppRgZA1MGAGVLl6tIwHSrgy
3Hpbk0g027eE4vLUrNyOqordWuAnxADkeBUKkuI0k+8a1GUXgSgilHPxs7g8t1PSvDh5TXiS7sLY
hFwsKMq8IOYl+sQ2bW3Tskc06EZ5D3OiUbBIqdaDQF/yqzbK810gI8vnbbAegrXjfmYVy1qy8DZN
ThZPuHuyRjG1uQikWRIbOfTpb8dEJhlRCfbh957K/Eto07sUEZPqjsVmQ07JDlnGsqwaj+sXNW0i
sDDrV43n40JMLDZykqvEJl8Exl0ucv3qah3JLhj0xV2XuXLqfbcTxb92eIMQqyNOrcVSAoc0N98k
g7tHDXUXNBK9UWlSV+u7V1yt2wBr1IK6FsxWa43pv6WO1pMy7RdUluj1RvJK4O2RPZYuzDY3KVeU
2b0ijr1tY9R48aZh+9lCk1AmT3iBS8D4J5dDFv48WNhC1r+MuxGouRn+xQitIHlvyRisZnWdNlZh
XWG9rRThfcZs4hVXpH8fUkwj5M0ReUidhESHdluxN+qINXdG3EvLLgi/oi1kqlEAFWJ0/qHsjx60
sj248Yum5+y/o0ujBq5KLUkowdmmQW/4cPm8gmtJKqIZvmdWX9lDvkgkGPQBPAWR9fq0SWrG/1r8
uzVBELZU8HAvIyn6y+AQesnJoV9l1Rcqaue9WQmlK5ffqTBT+ibqw5eMRwFh7lFPqp9diL57IeJ2
dE4f8epVmuPWynYaFB0c9h2adoLtfVbiIZzk98c83ZJVE7+PoJOL0CEB0dOzfd05G21Mfr5Bi4sJ
NPjHTZE9D7DYaY11FRdhOFdB6RSRrzlKu04KFrePuV9FyWr7NkLen9n3QDEF4X0vFHURpnWTcTRG
5so7CrzoX5ly7Av3r/pReSBGyIpX5+vpf2pwYkOG4Lduj6qeOo8oh031a/wytzHP7CjzWA1uQiqa
KuVdx5sbEAKiPq77zorRsV3eTwW4axmq9j53Mz+b/fOYvb9gvE28GR4MRIByrcpa1nBmG1BijEYH
AXEN/zft3+Ov7YyxqZBLsNI4s1OI38UfePehyXcZGfxDiaAUFYDRgyJD9k5eH2nbJLuV9flc1ITk
CbwpRHjokjYDboIi7z0eQ1TJjua3B2LKt0fA5QhrnuqMAVJyLUHPiitqW0Mf0Ix1Wrv7XLfJL5PC
a3yTU+AvisBmcZb3n/mEjedUUvYHQo+MnR6Hq1QZ2YMKSGVz7W75X8+PSfqEO/TS0lAxgVxNWsXw
5oL3bUp/QszalSxHkBLi/Ysl5T1bWzhME4iD3gssptzuL57HdL4p7/omhjlt5+oMk/5iak2iSRXe
2vpM6VolAmQp0hTfZ4E0e1UaBieGuiuajDXw4D6a1AXtu/+gH5IotE4pMgq0gh6Cs4f6Pw3s+vo6
cXitdnatE4QA5qVHLGUaO0pmPjoNQb6mlEeVNWvRYY9d/nNCv+KGgSv0CAscKiJg6F0v1YwWuGop
q7oHvNfye678B1bNRTts3RvJE/Jlh1XMhwwrCDSQijnpSREqsVqx0qJcrlCfNPamrNtSdm9XSCUl
Krs8TQrjyaG4TXIa822OY7ztFOBgATH2zaQ9yPagEvNBoaA5O7dk0qT9FDpSNw74SlI82h/qLLjS
JniYK38f2R4fSueHNppB7rDFMojOoUdThz3XTbXGVqRTJUMcp+Fxbwgav3Yh5KKNEdpQbpZps1ZZ
fpFSZ03z406H1wWZkvs3d7KdA5+VcLyjaYsrXgWrmlbvCq6R5YHAeguWNirIjm20seH/uWHWLTsa
4Z3lob0Dh1pMQQw43kzmxz3FrrJEh0QYCw1kEplzHrj/mC3PJJYowvhwPf59pdubHr1TCbQtZHgO
llNzuKXSOlOz+SxrwulPoeTx3dbk+xOtLMDghl7gSEeny3WTid8w/txoLOqOlcY8GRnoFKC8LREZ
gMS6vp7svaZxTCRh/L+YQeubTuiGpKMJIs1l6FAt2yrq5z2fNLgJTVuD7k0i7po+vg/oqetcC6yo
5cOtZBKZohVWndBmpNxZTlH2gixefGs88/KkVqO51LwpHWFbsSRJ+UzEcz2Xd4nTEfrtlQjmAu5o
JRx+tJdBGjiiZ4yzszEtlz1IHYvy/KnUYoaqA1HcPgD9U9wnc+uM9A+fBdeQlkpu3CWZND5J8OA0
V5VLhsruqZouIjVy3JNBfa4oJ4nLFjjuuyYwofvO6fMl/eiCKOaQCYurLcNBaCV2qbLHBvM5u/vr
9EfupIrrU/dpAezBrFPDAHrMdpzmyUAmsVx3nqsiJLjgN+Vy3Ws95b5ca5yYZwThUMoaxTqFgzDU
gC+eDCgbFpCXz3JKgUiaa0cML4Uq7KxorZ9MW9WFOSeLmqeloVxRJyT5dXKvCu5MYlQJDYNctsFK
MJVLEI33z3XDmTWvLL9pjJpvmR+DHBsXQT6KDHs2RhVjZ5E+by8VCeTP6Y4tbPYIzc7ominvNva5
jXuMt5WnEBJ57nKJ1aLEENF+1Byf+Dcgg5CCNlHS9QxoNqVztagJHU/xyPUKgZ9b2r5D8Iwg6Va9
bGSijNhJc1bDL+4g9BYSAp7QiTwe9vHE6tDBFjznEBSYDU7U1hT9DO3IsBdq9p97C+Gt9wHLINFj
KDa9RP2L/jJeo4EXOQ5cXUhVM+pgFsQZ/YI6TMXPJ5ZghYcrW6+9FLb2ZWlla5FmMdUGXVpSKhcY
taDFUdPZJSpkPSbbWWuMJd6sRuboGcEdLzBAmwrTF+UbDT0TYVD9fV2/YeeYcZm3sxGexMa5gCEi
rYCPKKzM302/tA15Qb9h/iWHSegvK7q5zZnoIo1jGfsf5XKIl6pcI6kr15W9GdJS46KPEc+jTANl
IDjH2lvWaPGh/eDgOTgPokOwetPmfaVZoHD0eN1GLl1GCeTCopZMRRB0n/7vkXndu53w/xYztJi3
xgZyxif6KD4y8lem964ut9NeodpG3gXKY6VHWF+NzRy0Lha1Rb6sS7Au/iZb79Nqlwu/k6oeAVWA
stENpQ0jg1cLYLAaH4EhrhQJNWgFpLsk7TPrXDVkR23m97w7QQFAMfVMe8YFj2nyuEEk4sDfJqXF
2Q2OGyzigf4l6Js0Mput3KeVgslhi99Zj0SQVUzqmDIrJT9IhHS2Qx5tModlyFzmueor6w8+garv
j4J9u915tcBVAFAw/v1ZqqXH4e8mBLSowvEUqm7fj444zXOz/QybZa3mmShDUK4OL0UhoG+tAFKA
k475lEx4OKDbBTjyT914Oe87U3u2NIx0iRkpLaGTqrtNKGQmBUpcAykAUhkuL6zXxGew3woEtUXe
J2jG6+2VDNJweEMjr1rgcP/hcXfG9h5p6n8MSRQITWl/b1fxindUOhbljAo7V9YOTRjbA0PCFa2L
sjVZu2LU8nbpQoOUkWekGDAU/7fZKf0QzhdNrwQcjvX+qZSqvfCVirWZftUSgRSXp2ZinN+IX9RK
DCUOPvQsqyIPihZIif61M1UfXwHC39dONDzHxL6qTKa/3SsTwy3F/FsLTDltyZaSWzOvJ/xV9NIr
7hK4nSE/FalihtTRuBfs2C6R+rZEiJGtpX5g1wFsM+FXxUV3Au3sb7F3O/hGCh1q6smGxnoDYLd/
SvWNpjZ4Pw5TZwdEXOaIMcyO6TUYtcmo9N2fPqytBd3bVQhXlv19bl/GjEmKaNwM5DDgfggZ/CtP
L/+WKSWDsCkpOt1LE5Kfefd6XGRnryH5rogm7FA84ReSEr87aflvq3Q/4moPEGRujN45sWR7G1Lm
rKCh6aSi/bBRkevkbVDbEptq5oVZX+k/LfGtCmP5GXSdDf8CcsKjd755zdj35kZZnNlPA+BO/T0z
1G03q8/kg+YuxPhXVtffSHx2EN1FRQoKY+SgDigMBCjdLpf6Np1FYqswOskwIQB96k88SCTVcIdf
ApPHqCjf3Tv5CZWtAkmdl5AIqAVsb3GS4zbkvQnuIB+GPqZagg0PU9yurcEttBfWSICXgEFJ8Oym
cruh2/GYzWPxZzEX7XXB1d80za7kRZzVXeAp32YE5PsGrE6g+DK2r3L3Y2syiMOxbNsFLunWyYm+
1ie1jB5wTh26OjNCKfpmEwQgZs9WQt932/o0cBLxBTn/a886rSafkm7h+PQabvLnfPRf1axICOth
ORRzbPwe5pONUaR5EBu3+jmDF2ELhfDfSGLcb7bewIr2jvyJdX7a0i165t5zkcX8ErJ7IJnEZYYf
SCEC2wjoimA6j7iJbXWhpNkrZ0PMTK8MQ7Ike5D8n6G5+aOhpDWWoso3/fq+iS3yltYN/CJh9Ais
dgoPrEB7IdtdANDckuZ8Mvw6Eby5YUiNuZlfsZ94tDxGcdgLG0WAUitXcCBJq1LDo6B2QdSHau7R
YGrFGs4akdcIQxuO7Q04hmNtcy/Ok3T4HcGVHkZbh64N/gdTVCzppmtfYUuQci0YoRqqaC0qGW5O
1KhxwP9C90EXO9BdlMkvPTgT3MSS+z2zxtpAGbDdDURGvBxl2t4H+7onnmj5ckh33tnPTyiz47dy
a/2oJMTs7o1mq1c12g534zBzPjySEHQjflIi5iYbeggvOStEqMZRMZlawBNcsQbvfnC+guq17b2X
Xsx9cCIc9mOCiBUvURkmHkROtL2xAmAW9ZqwrZie5QOvsRIITwUeeIAlLJEqBIYd6LYqIFFyjApg
2woRCbZBMqlX2aSNR6OGeGJXDUGB01+C0fNQiqqG9IJ3EqX326ulwGRTCYWopQMZP7epgSmw85Lg
B9EaFS0m2Y5JcYkafNOv/PZfc9ZrUNxKwDifaSIVfdBM9tGk7luNgTYbedR3GxTsHGo3sx3nrOQo
MV3W4j2P1u16pEyqiCORpGiVQD/IApBVNb7ee0cGm49wDl10FWA9JTJ5w+/t8SZlecoy69xrPs9Y
iaN2RXK7x8HuAZ+xI5dlcw5k8p1W5BvWGinO8hUSbLuBO9vAWHoLF9B9WYLRPdHlv/5dsV36zfIf
Pi+xmaFC/PyZ1HPjMv8Z8hbF1fIXxXsA643qzJAm3onY+Qwx4B+MFcxFQTNd1FGayaixPEbWBZR3
0sdDRBv4s6FlVWQIDNy058uVpktIzjFJqE0Cq/o7Dkh+zBiDrQbYZytxIgGMc2KTV+BEeRnel4KB
kQbVFgJlanx9PWacCa1qIynM0NNg6CE6yjOOQonMkkpB/s6fznYl0bcfEl5hSfuamCuAD0iYlGQm
I9+sDpuJiMmj2T6Y/QgASvoan/NrtohquGv3dKVD5Ioo+lR7U3Ru/B2TAVraKPcSTq9TqDmUu9tB
BpHX9vJ9B2pASgGhlm8FlS+gTu4z4WSWODe9r2EsBul35tjqk9B6m9JPWLaXCbakuSr9y1mdPhS0
2GRqaVnyCC3GrSXcQfswvvB5qsy/v1gwLLSJAVPFVbJm2Wb3lA5bjW58C7e+56VTzpp5FSibLPGM
RKG3CLzM85Riu+G//8ZmpihkbolaaZRJjPBCC7I9A+WiLDyWxCzBC/V4QrUVmlY3qSXPHDxdYk/U
7kDVUcIESs+LqQggZIYsubptXvqdnDOUW95V3No56WAtRB+O8HK2sJz3FXNV3hVzJKIYk82Q89d/
fqOA2AuKgGKUmL1Gquc9pJhO4FshzbYs/N8G1KUnBSx8PCU/NKsZCVa+4TNqPqQYMM7SIfh/m+pz
1Fqr11i+R3V69j3Cyc7NmEdXrbTMnJCKihNeNMZblj9lnvS6sSonKIMlPdOYfTF2DqW3Y+VBDobJ
Q22xnr+L5v4hi5+ebeXQSopO6VLDCnAmxDIB/I2rrU48iOdG0ODo1HGvxoQtgv2PphlwOANXd+Bi
y63gtvNeOR5t8EY+QgFaLOANGyznWYn4YYuuoFum+zjLoLHK6c37Rt9nJ7KdBwGQniYVUmd/+9Mt
SDi2Vu6n0Vd/+xvnKvtPfW65I+qYSP2kDsVhkeo7+G/wmNLIgxR1t5EetrjYviaMwktRDUPe7U/B
1uNSWMj7rcJqNgXWltYzz89+AXcIIyW04D27WHk4y3Y3IkY67MX/KNipOcvXM0awI08eIZo08Ppy
duEIzFCpoypwo/nl9KMTeliTh0CSE24t6oihNEAOwpBlNYiMt4r4gGxa6EtQvPGtFlUI0gi8OIIP
3OFUOiOkq6H9r8bve/p2sgm0kUcB5RIcirlPggMkaucsKKXLx/9Njz+5zdHfVd08+O/Jwd/sgCzC
lyAa0BqsIQd+1WKMCJExFiMW1Xrsu9gb+msHoM10a/axA2f2+euCaOjAJ7Ub02NIB/HF68aHn+11
0slZoLYzGjWfb6X5uuwpdqniGpJsbnj3pzd3X6wlAIQM87xDxaU+FNGZpxWczGlw72v44dCG2Qo3
HLIe9CWWLfHE8maSdvOQWAiqHbgNzhv2ZPiMvF1/0NOLB3Tywj8rJ708brmRJuNapRNpvUxtJxjT
Utjww/mOEqB3nrgCj5t804Uw/f+W26JuFmX+hXQS9S5A2g18agPLH3gohWAkWjr05HeUNbddpqjj
oGXXyDrsIUXrLGGb8O0x1EXR+7ddVUWUDsIMy5gPqlPlD6qVY2v6c2nEkZ+jmP87fAXQj2cZGkgZ
mbhvESLcRirqWGf+QyKtFNgwav5chdy7TZRxFmkjUUubUwJbrFzluCpoN77zN4fLzamIa0MfqCrP
wbd1bXDETYAzTivlGiHTFiki+KKzQ+dmXz1JVucajF3I9QvlFiA0kgpg2spWxHOTCdXQg6h010mv
8Jfs8LoPp+4XGoSMKDHsT3MRogFtS7rLaj5v6maGlqOlBSo1qJzOS8on4LDPGVDX62Cu32YDN90y
N8xsb/SkW/clHGbY/dRtWujVrAnx7FQ6ZsN6TyuE+5M396kuoHjTC7inZFH4fKatYLLXk0rxTHx2
aoEyZaFvvMbTXfkAQxV9NYdKYvCpUn4MO5SKn8hjLuy4/+QnLNMItrIec56xUCQlzB3Su45eSbPK
OctV+KF43DqLI29bRXMb/dSt6pt6J4KHBIoa7lDn6pQ9AaK9iuZuoRo+NOL2JwKXKrMsv8/YQDHJ
q2Cpcw5JTVX5VIff0JunXHvkKSKggbwb91DDEQWXrZ6unNvHMzEmDtytJaMgowS7HjCsJd0MWQis
cUZ82IchIrgZg1n+66V830PNgoA+I9YiGJve6h7lVf0KTmVPCJxBOzd58y1hsdKzAiT48gD2pFwE
SnFfbpd4S7SdIerI5Bu+Wx5LmrR5l/aYT9dwa0xa6NH7RxNEeQWFYpyFo/6mtY8tVl2O8gicaTUi
ECt0zWgxnZDr54nDsLmrSp6gILpyc5xorovyeYIgrhTMsHmhfBQ9RZJZVhAFqlwu21tBAibuNVXc
CRGOJb6lgnFYPu5L1sOAfTJgp33HYP1Q8O8eVsNKLXjsLRbo+KK2vIGil+CNjwdc/XlB2IFF6WYs
ZDoOV++sGjnbWV+MTpoVw0zgDJb0LB2mPZ5ZDfHF36zYD74RTRngku+6j3uU9rS6HrJuJc0sE8Zy
cbZcH7b4xKgnKWDd1Z8ehVENBUJY+Vl5zu6fkLSVrroXQC0AXVUsjgHAakH9ZSnvj4QAuIgobpPb
QMI75ZF4VIlHhVULXBzp+BemSwv8pEE3QQjEml4vFS+F4DXev+zoqztqCC0gf3+hSLMRap64czS/
2WVwmORl9C4uKtY/76wQq1jfNzci3Z7FJuENuBZJtQ6ENwtDwW4aAFkxQii1Ut9LHyMTHvdcYlGW
bxwB7Mj8YQbAnYBdj4xOBASNRyxVJxrkFakw6kpAUXKqtrEwpvQtS6YDBOQOP5kkhv8wNz4UTMVS
WEA5zAYPe2z6TleatGKg1ViO5ciW9Y2Qn10EFHXximrPI/oWbrQ+7j/jJmr5UH7X4O7/+/A3RXBb
dHIKiv25ai8/zoTJj1TlaPm7MP5bbQVqCHV+PynlrkvqsuJy9+IsuVjXQ77ySz8tiRH8FH4zvUM1
A9NH05PIX+ZPPgGxgcVy96eYr8MBpd/4gRne/c5vQ2E0qf+cPXhTqLWZrrs8qpfFjaJKfTQ8fL39
TCC77Slu7bPQb/hSDzVxjSZHduCcUnqMSH81mAqjY1MGSi3FVPhNMuwN3aQ9uc8BkY2pb7F3uhxs
+c23XOSfuGfc28j9PK0j3MuTRF9PEwTO5Yu7vuCKvpDqy+pbOSJvqPPALg3r7Q1Oy8CjezO/+sYv
hqGD09Pea/DUZxgnkSpYg9/dKhy5hJ5RNNZycVGvm5V4Z3nkIkatOWV+qx3gTrOqCFqBu1u4Nmuc
c6UhUvIKdJed3k114o2srbie3gPywzKLdk1+5Nexaouy3WbvYgggYJpvvd9cLEW/T6OZ95tbX/jC
cqVyTF8XElmB0Ym7m1J1jRGPfy6UXZ1Xpn0BO8dZ+LptYNAQn9k7Y7Ro07YYtCTXrksbHa3Ugyhu
uU+l4PVWhHpDUeO08h09FIn2T3xA/lxi1Y0dNQdVsmhR/eMxdsWHpht6leOhowXecoKIY9rGvJKI
WNaFouQpQt9WyFnhldNcZ7BtfOQrTK4G/a4e8Jh4JhRkjwHI4XmLD8YLs+qiUK3ZR0KgBbum4icu
nVgYOKJ4fxloOAnqMHQYWr5lgGIV5LhXW45atUehhla+HjdZ7OOJJ6ctwn3HzYwjHIvR7iqHMeO0
XVY8hzD5vt6IjWmQm12ycZ48un3ydKnmbu0RXtEwTnQpHw36hCxuaGuF0IQF2hfkBo8sl+/y8UJq
TeC6YM/xHO0DcVDwQxkf24ScDC/jPGd0He5lXVEb8fIfOVxTe7uGIJXxJuBp6jhVNwU2p952uiJ/
uLTnfRByqOxC5BXaTkkaFMWR7zxgsd4Ydy3SzoIFMrqhBfUDN5klJPJXNZSIFDzx9RhZVEzruEWr
m9F6YGAAHWy2nObyFCqERLxmxAw1SnzVNekloByBL5Aq4oZFw7ttcM403XtHERqwBrm4PEiJZh59
7HnVymFYmYPtC4u3sGaQ4lJiPTifGdtxeFUSlbm3/GJTr4yYCqvCEi1T8omym1pn5wc6y3vrWDky
h3VMVwqLRzAti4c1PC+xKWg1Z48cOMZZX8lJ/uxOj4pw/L7+cX0a3z1AOIO9nPsxacAA0PnY1nzZ
US28uknLymbiACufqwmbS4wuRkFIF221TGEEM2Woh87iLHlzRe7bgEuIOWZZLKSu0vpuo4P2DyAU
/4DWHRbh6hgNI/5r+onwbGzOIww4IknQ5JbXUtZ0Qu6caAkqsD9drMUPcNMyV0Te8rxWX8WuNvQb
y06W8/S/nQnBYQZU4Lv+9plzO1BPRo3R2gnr2SwDVa98EODtbLbFc3P88upIwigGmC26YkE+XGtD
PvK+wRSw+EWX9kukmOYwNSvStXeA6pD/6zhdsoFaBBDhjQXAdsr6APZ9xmfx/U6IKDsbnvUqXo1V
3Zi1cHcqX0nie0VPDIsJeRCBRxv15FovIZ9WRHvvmxj7dr2hmHMXT4BNS+8SmVQDb3XpcHn7WMjX
qYJuSO4pGELWRZtP8hnlqXq6fATGLAlme12vrgbrYcy90IoCciORWYrbBhEITIjvBsNBddBGvqyT
xfJBNHHP4H0k6a5FiRhNnsIMyU2ejXpFBzSESw5VTBOu2NWlw52LkaEy+L07Yp39qspwr4Eyfoe1
365Byj/flNYJll8Xm0VNmny0iPMMXjlEK7ITMNNFIxPU8e2P7UXTfRuNQG2BbfWIKhDwZxG7s90K
MuaRyjgMAsOZCoI4Xm8IMRans+nGLnI25Fy86AZqGcXJOfeHbEwrtojtUvVuixUHGprKkjRtDtwC
Ss3V+ggUGLgJZZ/8voh3wr/3k0FbodUPtJyFnfnq5sErLUUtLevZaZ4gpzWKvpTRi0TErm0zPVP4
Gl3oUfee6nLCA2yK5iiCm5ytrnwA0t3Qp7EbofWU40p1eU+JgwGQVD5vIqFXSWgkY0Yx1T05Nu3F
PosFgRoMMsvHc3EGCO4NDOxz3odG6T5NoN0DDuoPz7PzcM4EytFWULVfsRuKJfx9bVXXjkP429bl
sVrYBKU2a3ZscJExrhwFAhtfQVQVRE0udBaDpq07+7UbLvljZj1Hil7uC6yij6+MC8vhG/AqQCSw
85v6VPGfoFNG6qa6e3QexhSRhCaCGLwZpBF53/vnbs4hyPV/4PQ1RafE0K8QGXLLheuaAujlL+MB
1z6gCPopABQzzaXCPxDM7Or06ELl0hKHoWhHh4nYDwCLIq/afKTJfhaPXYBvv6zynCzNEAjvkXei
eiUEc0Bfrl4LpbBGK4v0kBSP/2ENWV6rhVZJXg9doS++OOHWvTa15fIWrqwwzF3sgi2dXiu4w1s3
H5sJVjBMa9mL8Co6Jpru2G5jMk4OeKNhxv32H7z6bc0yJ9uNhBnK3N+aU94F+KHM9qvsHjbLHwG9
msxcTT+SqUhrr0vSw/6GJPILIdB6JwUKtYW710CNP3ZmGdFFES/Ec6KMLVvuJZAUR/zINURDhiJU
tUigHLbFEruW8pgbzDGyDuq3nWievhuy7NgaBM6Eog5y1KvzX38LGBcYLgKkaaZmL080RHO5Jwjg
Z7Bz2ccxwRYC3l6dZ5QpgVvwCa55BFs/Xl98zZnmwWU3Jv5Nx4IRfodaAlhKromesxIFxXc0JreE
sYaKyJbFlqkg3qUpKfxjZSZlFMk0U0pukY5vRALj5nCsY3nktDaw4LIO8q7H7PGHu8CKjaZ/44pX
pwmD8F0Yooz3CazlctrRDG80w7rJ4QbDk/MK2lBHZrImL8Vtpvh8c8fb12+8zFOC+5dP2HwhJVVQ
JxgOx5denfZfTA97sSVshXWwjMOXodAKA4Z3zToOCAuL2onxe94f/y8Yt5QWoSRGmPAkzNqzh/fT
zB+6Cfpknma6JIAgL3IvWLHhuJv4Lz8KdABra5/TaPB2JreYnv1LSW8CSB0oVbs63kTO1vXAAUj6
rn7hpCOBb9eld3VK1odV6BZVxlhCDrJv2f1X78V7rI4Csgpk+615Tea5s2gQUzI8HJynROSznU2W
UQGcRfQe7ZqA3rcpYHXkeY/kCm0UDNk/lneroMfzl5x7CPzzJG3XQzhMjVlh9pzOl07HtsUiX6io
+44mwCQ1t6G+5GvExMsA8oY6t69ezCe8/9SVbpPmKyL7mzhGhUUIcWsAK5fj1362SlJvS5Xn63V0
5fuJcwEIqPO4XDhjmHNs8x17Ta8xYdKIfUV9hdmfoK+QDY0awzMogedFrbjXiQRWw+cProzl0GJJ
+G6APwZfphXbOkmcE0hipNKil/n8HNBRhSd/wQ0IZl3BPhekOukgWwAg0woN6/vet5/d2ylqc/pi
m35q4g2VGma15sZevlnUa68+pAZEsVtfuV1M334rQMPz4Daah5NLFt5JjlFg5V+Pn/1P+lCCVxdx
yK2GfJ3HPjbrM1j+mrNQdjIeq2byora5PNDZ1QvU2faW0A2Ax0Be1qcBEA4MwLdxlvoHcBtQqaAL
Kn4Co1Is0j6K+11Zj7BrgRSx9H++Sckk11ULlOfcT9FsUa3w0IP2zljNxsEbzKp8yJT2vqcMqRmC
ZsCmpQLH8zLEKbKqjA/91QuxU/hzBj08ceKCFIuexAU2hsXo8a8hr0E1mRTZuwjS1/rI6RpzwUVA
4s+XFCopE+hPkF8CNFiJH3uFx3AqLrjr4pxWMqxlgLDFFVw7QtvFNKGwtgqyQd30Ghbrr1FI1zsg
z6kk6rZzWxckZ+dN0ojxY1DFvBC9rFmwh4ivSowdcpqfaVZptN3U8eLfk6gL1s1eroX5jnq7FpaD
EulMEMvhnycFodTr6JngPOJdYATTPBwixTudmOFCTIRAmqi2uuO3tyyt6Y4l7X/3kInTt0D6p4wG
5gMjanQL7g85ExeRs1C2HbNJqCoZUvADDVCVALNpM05SWswMT4EO3OfhVzU9QsUF7IAjbW8z/Y/f
rtfwpVgHlg4og3xZGMVaMOLkGawpE5gh0TpuKXlHJHb39NQtQsQk8XOemZjy46CX7cMrMWPsjHoY
mpS80YU7baI50T4XIk7KeZQ2bhfTEySjyisU4F8x1GpeKSUay9NeZiYO1S7TNJltnqoS/Rj3HTGL
FPIMdmSdJV0aa8oqWrtnUN40wuRxDBJ29Nt0YpMeso42E1K5C2u5InLbeWpvC9velwZ4O1L9FVkw
mvnxiI7GuhjSupvCI4ZRv3oS95kquaoNk3spqMpQxpBVoW3h/nkhrk1Z79GMR8c16zMnnDvmrK9E
WMqhe7L5w7Osy07lVr9L42KoAqW2tDpao69bd9uRTDTxTHy+WyMIxS7fMDgVr8ssutXa6hZoT3Kd
GcWTsrq6CfvDFhWIj8Gi9NG//hOScWaYRpSl42WCkCdovhDz3nESLPjW0rj1MNxpU3ZHgYs7Q3VR
Hn8gVRUYPXjjpEL/ffp+byZYL0RVN9TAiiiJj+3mG7RSGaNTcKllWsuJqiiZzrGX6ARBmCatmq0E
8qpuuVfZCJYyCtCIZN2HCp71pOldwFXXWzYyIjYBl8RbpSm0Xl7ThoYXZ664KIKOBc9YurdT8J+c
R7Me+S5CW/QeGuWtrCePmCbtgm4qdGjL0WB8YqMACqU2+l0sFSKK8UrZVRhldon44ng7aSdsHpsf
3dSMKFyREr2eKLruxMYZKlX5Ac5GO6ms/QQQyEbsGdizB8rzsWAAjHTLRuNemL4o6agncrTtLtUW
Qhtf8mdalaqTWUm9ZyDBZDaQ7j2GkoB196pqfpHdHcGHRfjPlQWnI8fA+Dk6gIPvv/dnAxHvZUDL
pQqhDrPkt8YF+jaq+H4iCW40PNr2tkfl0g/oUJLakWkm/Ze0/jGjyMraQtLx7a/TvFF5QyqOQu6I
fC5jwGNlBoXr/Xl0SqrD4s1M2ci8oo112FGibTwY1MT976Uh+EE2FTM3kcTbQmSpiFddVZPPuyiG
EunDofbD/rmXFjn2Q39HLjXC76khlIEMs79y0D9+9ph1jPAyc9j9wSzafeRr/DruePL0We/v5MCG
XiQQOZbE7c6CJMozKHXmkH1ldqQmPmR5XNkRudJkip881KtikzMI3BZYnD3XXA6F92vzw0Gh1OmW
X9kdHC6S0FN32X6RAYnBBnkVHBbtrL4/ysAzygcBm/jKJggb9DMvpbygmfUrW513z3LueaJZxWX1
bVDfPWkjMMxopQRwxK48sUcWYQMwSLVXF2YjWRW8sO2RSFGuwkfvF0KVX8YX7DPuoSvm7aZqlOk4
M3MbnchBM+ggQz3taNC3ZVjHjLxaxqc9HkL+8W+UmaoHhxhWs1oT49hnJ7c2aFFQGi9ewd4tEgPK
XC/MPFS3QZoAgkNhpN6YGEQNIuwPhlZpgdtajPMIB6QFe592T2ZtXiO9AvHAbCtCNZFujDirlMXY
yzNEb2C87cSzA6rtKB90+7eEtcEpSbCCLW5G9Re0x3WbcLWAG6hyOCmuMD3YsfGHVmKoYu4VIxZK
0AhQSFu9F76H34x2K6mtsEHYgmXXkNYMlIurGqbkpEKcpV1pK+PoYfXhkJ49YVnqNwDBeXztt0xe
ZXCNN8uDGfyLqojfQcSkqGSxNZPmCid0ON9Es1dzevsnh1GUhfYvh9YkMknCyH2XjdIFTq4TJr2s
OSycB/iBnmPlLb+R8fbfJXksOr7ExPyVo7hwSTgxo79pLiPBIH8P2yJM2JwBfCxrhEIc/4gS/13b
9D/JgKrCwF9Nq8dzDbh2ildiXqr5LGZzAGcj7td3YMT85enc2+77AgaSUkKF/MafyLAFoaNvO661
9RUfF737xqd3Kpvk352W7ivQ31DMybsZqeReP8MOsTYrL1L9UFN0D16nY8Y+ZhAVsLpycs1eRxzD
QY80UidQtQr+YK0oiJDBgWOS/n92O/nBAPuzkIZWmuamAsihXo27IWCIQteI5M4BZp+Xvduff4Z4
iT9BByEKADNNsurMeGC7fkpdu44M6teUWnr7PZkySj5F9b1+WcKgtjjVkwpoTer2E2GmfbQ3dULJ
exY/FyKNbFPKA5jJ8yExocatWJsbPqnsK74PU4zBF7KU592cJUJGxlP6UA028KiAusNwAeBjNvT6
cNZOuOkX8OApen4MaBJmDktfTXbfTzjyG+K5Ha225Pvnq77rAxeUIdGwEAcU7PPCYrB5N3xAuiS+
kh91YEhCF8/zdpAqxmPOZQ8fLX7PW1TvG+70Uku/kQOARfSDmkqJySPgapFCAMAy0gBa/nCrCGOS
tUca1iWpB85ib4mFBHK/yvOOhiCf6HinfXK9SU0uxb9I4KpO3HetZKamGaP2Mmi4qIW7/5TPWHH+
u+uLFzpi2weJ/x7Eid+N1Rs0eIH7rc5e/YWM7xW/8OHlTHNFtsGi9/2GEOCjfseTKPvtdVuI1bnP
1LCtN8BO3naBvcQgZpLVWly1I5mVHu7tRsXdzzkL6sjvaUKBBFRtNonl2ciR+UnuP9giSdQu4EJN
SqkcyAFB59nW7YRmoyunUfsbROQlH7c+PS0w367csDvLp6zOiW7YpE9IrSSWsZdznAtlizCme4qm
bmcA/PvawuzEYk0V6X6p2yr7/SUl4uTp+A4xdiE0I2YpD+nc/ZVpYDuI0D/t8m+nS+10hFsnEKYz
IvezXCgHRKk4CacS4GFA9nJPazWpPr+hShzR2x8ATh4GMUrFJFTstfGAXLt+21b1HvXbK3XlqUHc
BVOQvHXhEiTJOP3rZMzHoKJ+QzJqUek1jytsZTklklnrAwdVImj4rE1CUASKgBWSbFwlQQ3h5R8+
BMzi4utZP7g5q0345p4i9vbf6K/fVxFgAIRw50kPamEhLd3KF8TkqiyXauCIP8hTz3HBYw7xnZaI
2tw6jgaQRL8czHmLY3oewht9BdN4/1fltSKGpT1zmKKXINO7VhusdrGtfFncZK/0cw/ZRBG5ayVV
0yFV5m4tMqqr66U4OCoAh2ejBKq6GqY7RUk3LI74uuqMEd3sFPFkxoCh+2lfcjQYbFH0Q1CneSQw
B18wzkaZlIJGj8f7ImbUeONBqyu58XnPh6QbwvIipP9vBCPTpXo3+2cic+SEQVkKmhQ0WMwj188q
ByAqOqw0szn2ldbTqyASSuCVryyue6a65w5D+KARscCsHFGVyNc6bniHorda83ORynlMNWrKX9A0
bPog5iIA7JL8lsIvqNTZHZD8+ZV3Ok4i3MWuK3dwI61QmUZCmY1qHViu023jn6bQZ5JcCtnAHr+Y
zpMh+x9+YiH0L5xTlQZkPX+NeLjlk9bxjGeTcW47TlNaO7/ftc5TyZBGK3qbzzI0xAbWBf749Hq8
qD8FQc+MsY18exqpKfqZED0DIUAN1yfy0yEYJIah/KEB9s1CaM47HoHO4v/AhWM8aAxjn0Q/MhUy
HOxOOsqdX7s6DDWBxLdDOLcuWYSEn03qTaVJhM8359xE5nb0ciKdBxLS2O2oYOkOOyz+9izqCddW
ISkda2o45qEosSGCxfVdKtCtD+3YXt7SP0VASRdeC76VRM5kc5FsFpBL7HWgBpvspRWAf/G6Pwff
ED9zOqx4960+1lpbr0fuX5JU8DwxNWMUjNM2nll1HwAEY+uuBc16tbUHwUQWqHhWdcpsThw3chzT
cIlRHF0I+JWxs4ZQ6ztRYs+0shAydhZW83LMUvoSFmbcYMrw2S1GkVSmTbGh3/tXTw3W+vJ5Le+Y
GrXpEffr3UUlW+p+82RtgDC6GmdcNwOc1St7yS3l+hk7G5Lu6BJ54bXAlLif9w4tLfJoSjndlKgM
r/8k0M8zdysq5JvFNjHg8QXpN+b9lArcK43SvsEJwgEdtU1M/2xHzlyQrGE8v5otfvfsuTCxwHRB
rDobKQf9EDn736Nc8fEyUqfAA+zmZE4hoPziDeaPaI5YvxoQCRa5Ap2dHzHXkvg339z1RQnYeAS4
m3LNyw4A/yr/q7PRGr0IPCVNHWdVLXnWucba9X+ycFn41F3qiC2msAyQgkA6DIevpYKL4S+qAf6j
j6fAFIErw9NKDaZRLZF8IxvEm1LA1x3tgXpSi53lFrRYoNE7axjYyrpM89qbw1QpPpb5GQ02p6wo
8pIhNWnw2FiJyPHBZx7CcR1cK3CIhCNH9MPQNEOALt2Y2o/JgaA6TFdLd00xBA/Wxf93TEefLNZY
u6up0pgDx3qVmvWCgaQClKNfO0+a1HI8HY+WWBG81O5ly4mEDQ0b6raQnJ+PYYit7fgN6pk3cII5
sydzlllX/MDlq0A+Kb7S94SnCy8ODgEtVuAymN4Ct0wBTWvWQrdhqTDESn4QEh3yuVcgMT5DRP4o
0gsZsQAjpfLvF9TQPAyHn2U9PXpSlhESjsjiEty0gr/yYZTB4lT4mYqmy1JKk30raAgg09Csln/s
l8ohxsntxY6/Nni8HWUAhJVrPvf9IJ3QrEzTLI+t2SdLvgg5Twrph6OG9SI1t8Os5b9u5x/gqCkn
0v9iSj4NsW9ApcpKB2HLj+NRds6X898FQhgBnYa7PkeqYyANC+NfkF6vIj4fxrbYNySFfBEbn05u
wSoSmWqdlfGGySLltUp5Ym7vicuPAKGNnnNtJZtZ0I8aY6XZKbjPsXUqzT9/ZO/zRv3qxH11CnKi
APv75kM/eQBzg9uNZKLVLR1zJI6tMMzWpmyCvXURFYIhcqUAmxuwF/jBzZ6F+HKVVKiVs3grQgCP
UoSXNUV7mGqvQfUPjhxUkjP0fhLbiG7kBxO8Ah0gfZAxnXzDOZLlf7qTCxIjcyEUNWPM5nmejcFp
UrvyuTFVxZPsd1uWAjPqAOdSLq9QZa3olyw+h5GUzq8IIgARaApq5VsQFWCIjz8AXlipTqle8iQe
YLudCAZT+EKcb10J+MRkn7/CQ5Dr3gJNxvBEOQbmn5BA24j3MaIrQbtxQmkV1QYXVcG1NB1I/lnO
7Iz/+jJdxoBrzGiibaBSJpdlrNvmIB9a3tuF7eVWiHVqI4z9tZyRNMgvuZuYcTj58ZQ3kBW+xRhi
yDb6NS8sJZUIhVMQqZOhhht3njsgS0DT2wYPsUwPLuEE3j2bi4Y8msppIsl7MGp3QFpc2m8GKiap
tdyFBhUVWiC4EmHjxrizl6ly922mBtKeTvIFWXLbAmXn2Pdr0GLDYXOYqK0ywbcGoqxkGytD2mJ/
W8kqhrQLu91jQdH4jvybgooR35nXeTKswapvKmPt2OFyfuvtzdVrNYwDS1A72N7HHqI3DHR3FYH3
xjSv1NiAAriPJ26ZFZStWt+3snvkxF8kuJv0JEcL84tllqW1c24eTDt0lzrKrrLhlZWInfJQgGtT
ilXEGSKj+XNjccV+lLIEr6ORfbkPpmD/mOOHwf3d9SrkuZsoQG93ABcOp5dwXPJAVp1fgOPlEAmY
aS/CyFsculBUylrixUX8BExcXsHF7A+M26TTBLjuBwbFO/3rozp5G2VUJTRJLNZuXHN6USCy1AW5
WBuZU31q3mr/7mEzCAmwhgFDVI/3pL8ywd01IZu9Rwl0dVssy0ZFHh0+tBnlSq7ajulesWhYNOVd
gbsnhAIoGWYiZpcEweDOmsVz2TJdGc1Liuay6cuLYp2bbLBz38m4RaNKWY5mSJNi/vzacaSimGsR
kZ4VJbqM+rs5mwWFnZraFvCUoVe5OHrr7FIJxKqSVO88JgQvnfkffIy1jH0RSDesLfyNe+VrPm4h
YanFNwgib39LtWP4QiFAMgcf/WkxB/5DTsCZRt1knDgSPrK5eGgu4ZsT9c+ZlA3Id4GQAiAyESgY
G5FqqQ8jKWgijukIaSzV/e712dI2UvV6tNHq7MPpCMXCQpCLu9iCySm1Gz8aats1xKVQAmilYWBi
UkgqKmX/0qL8iTt97Av5vnTAwS9IEOzcavtRWLXFyWCOf7huH6UThewaaLC9PwBQqWBPLzinGLFw
8DQl7U2UoaHkmO6OrIN6FJXfdFF/xjoilGiwqzDMYJX490CWjKpHp6bFOQGSCxdGzrYDCTNSWkk7
COeDhlikV1JwNwrgPTtdWwYu2Y46oPMvF0+67kE5oi846b947Z8BbnIxDngyiE0sRDfA4UVkeyAz
nYAdkTNq0HF1U82Sou/cw/mgsqvamKB2iOnoI6cDELp1jgT4O/iFgPx5WL+SHSEXi9JGIIGxIvxp
OCpC77HASDBvDYdeAV39Um8rh2i2fKY1zBZ2s1AWAMooqhSs0Hf8z94YMmZ+mxsJ8PPsJ4U3bQrR
hFjx7BUkN99RT5TPXN1TT2oHx72XZ2Yk0qREyzn1ynIshuDr2Sb++Bgi0DabIBXMWWgW/tBmwP0/
kvwQ9AkZr0Rgf4JlLOYh8zse9xfcvJ6zHdNE+/O7IbEjvHdubl8NIS9z9D55K5bX00Ek0VAxrjkR
cDOW3BNxTkJoVM/Iwb+4JMY68kecYXbzmay50gGzzZI/TRkFnp5D0HFJqbGR1FNxbXR312LFztkI
NW1xlOyxetn3bGY8r/9kkKBUAWntbwH7br6ONe2MVlRPoDCEst1zJkv1A/gEhjZFTIdNV4Ym7nDy
ge5MnjEDk99/gy/tvfG6REN3X4cehbIiu7YNb88TDAQlye4k8AgILa5j2kOiA2oZdSKKfIvzbL3B
0HWvW1tmudEhWvuYdS8CFnax+9rejxP6QM1TlnEFCoQ0CRybQeIBS1wqkEaBNJvCk7LzS2YMZq9q
fuC8GpqHl2xOFpn1vd+fbu6L2gWarMELJD63xzITKCirxONgaR4LiI58ENbcgjGm+0998ujHQQFa
jLUZl6u6WzIIMGc2aBGtjf6pqO0uSNI5gm7r11v7LM40h3GUe1gp+W7cNIMKjmwdUMcjTZLJPeTv
iLREq3RwgPZ9rf8eccmUPUSWKtuubK/yY0jh/hXnI1xpE6uKbzE69N9xaHmy3N6F4SQ3X5uKWT/a
VqSJbqnQSaQ/lH5IDLRFuuQ3VCvzzVulBoiw5zXhabOoSAr5rIj5CfIuUBmucGUEZ8pBlSbCYKUl
NQl/N37U+DqklNBbkA249CMcVOJjDJ26f7MhalLisIu/5uzVIHhtTmpBSAu4SW+qpMy6Mb/DfrZQ
/6czvlBG9IgM1gv6X1knWQySXWMoX5pg4mUEFt6SeUWGBzbJO7WKPUVE1hdZGC6BtIuR1ybthHHl
yiiTW+wSzlaya39u91TfHfUtCPoz2CK670WZTmhDkimRq1bOYITYF1yqtWOa0hOF/BvnveawzD/S
hc7/MAcSjue9/cs+V6ECjoce48fI3+cHR3lZ6Uv1BgN+TfUjGtbGOfxwewa8gBMb+u8HlHAMbpz5
0/RkdeT7titmcBafOjGgGx7umard9YeyoGQtcO3l3fuRuAhO0kOkQzrM3TAeclJCYbo3sCFpevx0
xTj90wCPeUckely5/V8p4RAdlpJr/PKHfyP/6zZxTYuIpdfnRYtDI0orpZz9y+wHlv+ebRNRN8fg
mN9kjwJZI5TWtJaX3kMJRaTTiWRbX+t4PhtwHDkqtkUCBMTTHYhlfx8n4m4+fEpQ8W1Hgb66uqsf
XIDiBojtoYlTKM8GPMrUWlJC77P1Z3aWAyJS0aeehNEk/m79L6grwKHQjRbYYts77McTj6r9GfJM
pQP75KomIOVZk22JZabtq4NLnWgRG9WeDEvY6NPaqisw7026gFZPlv8Yo3UutN4GL0VNhXzD2ArG
2ANP8DnGzAVkjIrM1qHmbDCrtUuFOHs6km1zUVBSu7mN+KPWjVrERUHgWotH06odIoW5ryLCJ0pu
sK8WP5eBlYli+Yuw/yCdYVi/1EFysRCSXmgXQH9dMYzb1cebSJwLJxL29zQl14nTyUpGaOu8bmuo
4TlCuLxU6cZG9Rl80waFazfrRhGudE2HHfCCnBdLALaTSrTF/WHOb5a4W7aZXCNTrwree6atXXte
vKW7TV1tnxl7M0B+gr8aKrmv5RJ4PNsU1AxhuIWllsJfeP+0NkyCE1LLlOjd4q7QPwj6Ru+e6RWR
XvVZwQtfFWG0fdzdJajz7iSwLAlg3xg+KXKFZhRfDr10MHaEwGDQbnhQCOnlz/hnMwgcMUD011Sg
xQrxwZ5W4X05bhEOErv+gCxaM5E7JIAox1+bALHdlr/7vvxdKBhD0kswkba9+07WwN82H6P+z4z6
v0bOoPz83+/d7PLKnV51mW2gUIsT5F+BpYrELSXHkMkTN8VmB9YxLS02i6WV7BLCHc9XpLgJHG1D
V6inO/DZ4i3J8ebYkQ+u0tbyP9fWzlAMCB2MoihrINUqPoa/qdAYPBvmRLoyspDrEMEy//El+DGq
L3I+FkWv8ghtThy+2y2Dc4TA5XtNlNtXcZ6/FuGuYREqly87jyudj6p9RLXxk5vmg6j5nvu9sKfb
wF1k1RxpVWOsBkrKE013MJRAcIJfCha81UosH9LvZvQPNrPFKvCLuu9aIc8rp8iggfK2HxqKl6n2
2XKm69u6bB9KbDxlkxJAEn7AKURQELK+SbBauf1FXTjJZ6fCPvT+5+HS8SxLGf/1TJFeEXrPfMk0
SC9L4CgGvl1MZzUVgrmo+Pg6OLA73CUrVExYtykyp09UA3vdwRGvTZtOcLRob7asKZXLa9QpE3E+
sUqAB4iCN7bhz6A5tW7pj8GB4JSki2KVuEy0p8XbrlqBXM1QWFngA3Ql2r3amG8GFXTxzAhU6vtu
Z/x93x6wfq3jXK2UmMZcxa+xptn5ZeYJvLq4bV/MjefA4GCn78+ZeN1z63/sXn44RWE11kXmGZdB
vsXbyAsmqgA5mrJk98xaclCO1d97nbnWZfpxKwO3Z2qBhGasMycFpQyki/M/5GN/DX4s4J0MwoOD
o64fLIgriPWlvsbPYdGqrg3qHHnyj7yaU/73Auk7YaYCMjSzXghT5p/8UHEi0g/BXLVshIeynU4m
H++y2C7XyDuRhsdy2uW2I1+OdhIYHRc0gkZ3boWFyqiREKQZO/A8k1IatesqhHG2OLgmy7qx+pW9
HYvwfMCyc7n2sbY9V069ST8Nd5JDgq6NgxuwhE7OpQNipM/JGMT99uXGRaYOzGYG7TG2mmuWiKD6
ACrexA+ktyYdwjcZuxc4R3d7n8g5lf2iRrS+l9i9EZnYgTnl74rlRWqvJOAehewrNm/R0f9ZZ7JX
4Soqcpo8KeKi4oT792tT0F6TZi61ahVPoyafrp0tOkImaxp028DDYFP4CpC2ybvn1tkf9HULpMUp
bOLVc49uJ2r/ltFFwe5UhcMpEC4oqAZMyu0fWDmBue9eZcKHJ7vmbCbtwHEt2s5fnLNRkDa0EmOi
xoWWlBNxw8AcMXbRuRq5VntUSYJyiDu7LYvBRNAed9vjZ5YMExjWvHOR6vuPLWstPTaw6U+149sc
9zQxaLX1Th6lSYqINK93KHCOLNqu6NSO9hiFX5oG19GuOH5/2h6AjqgRup8wg5oUyACxZjE5GDm9
BMOSl7rHVj9dBsDEEkBGZcv4r1vPPGxwsnwnu9mhyNxhpugQ/ze/Pz0k36/XhXDV5jTyMw7zge/n
rYIDXo/Goi9h0vPV5E1uNg3Gh+OZsqTjOQGc4V6wjOcgQLNkZp3+5P29K9RWcAzQklSTKm7WNH0y
mS89RA4gcdLpu93P7/8laVGWHXYNdPJnwS4EHAh0AWi7ooJCCM4VPwm1bi06WD32npOGkymHHfEO
k1YcnbYtf6TB0iAvJLAVOGKpoMJBJvtU/US/Q+1Y2N3w956Drtz3MJO150UeyaMkzcXnMHQWT4YM
uy3HqgfJWEO+tRKXrXArAo8deg6dlDd9iuPnuqbam7y14ltSpdM49c6XgVqsmULeEhJGCoZhfix2
wIR/a3xSBjyHLYPxrU9NDg/IDlNmK4HKnqKz6N7kFm9GOfrGjV/UOhRVauvRnL0JYQwNOfF7lEKy
j64cHCVe6GIa6+xhCR018055h16FukEVKuOZKkrPCziYeYD1FxhLY6MABVCBA6iMp3RRLnxKzwgl
lSBsTfb0pwI88DZw99kErgZGtD66Kcg9+n4GPC2roMsCDcvEGQFNc7miX9/U1nNdLVSqTBML3wXm
MGdAdlkad+Kt6SBQ2T4uSERZIJxLlEymekY/7rTSBkdC9PKr4Ozegtokh49rKiHjGLfkwyEgJKCI
2dTd76488LDLVLIalEwovmtWXonhPTQQfpLq3wHrxW5ba1K4tKa7flISPzIYlAzjSYS+Aehkv63K
jCUeB2ikul0hRGs4KPN/xMpwPSXtNCihxGNihIFK1FdsVaHfYiNupPd5+ZZfcGn5+B/SetDw15Tq
lPZ+fExWoJE6mCAj52rNTuB6O7R3+zmRn6oqjzAJc3Y6xOAPL/3rnLaGZOWJ1kTtDspsRUxuKWwb
tT16rUPn67rJq7H+Dn/+1wbpBsmGVXmZXp0yE1F7ag6KVOONJ21TLKsVITq3vBRGLM36itrktNci
iCL3KunDKBsm7sAZTeALl69rvK2/yoEy3y4J9p8xQeqp0li3mJEfWLWTRVRClpXQP4UCKByl0Cgd
eofI4+zml9DaGXRzml0Ty5xpDJIAB/P8+z3SKZl4ROqLsz5ztChvs2dSRYbDcWfvbbP9SkWkxfym
NKNE+HF3wS/WEEPeEEkiw3izSVy52YaE35m1dF9McmR6MxnAtptCVeXT/BkbcHba4ljwLC01mVwQ
hYlbclHdd5WxW5jNB8m+gESugSovKB07EUVlo1ObRm4dvGh9HGSARlAEEPPxkNE+rZ2qhya0CRFj
DILTvZkr+gP/H6LOSG/XtMMzfmgVRYkxkU8uHCb0xM3AXLTWpoUtT0Le4j6FUJXCKEK9ySTmXlQZ
jJEFpL3+tVVgeuNOvmS1/cewlUYuUDiXvl3SzNIuVZqexgOyA06W7S+AIFPa4TQBZmsOBVfwT9PM
tpCxVrcAz1TKpnA4qzGZeBjzaLA96/AEAhTKem6mnjQDhV2QgFzKIGfuV87a3TyBCK3koOKFAbP5
l7bAYZ9qtrpJlNbrocQhqKM/Osxj1i2yIRiETVHAveGMPPw3pJvE4q/4v7bJh715Pr8rj0an5IO7
ptLq6bM/IWXe4QkVQ1fyk5euqZD08HRvjz7LhT4LhLg0VEe9/f51Rn9jn931mY/8vPn5LuPAMqoN
rr9dnELXCiJfByXHIj9AwjHOHZDKULkHhUEmhQKoKmLznfODyRCkukjfpgvdbQ2O8PuIDYmobQfG
yTnZhBccJELofiE8GiCKhEY1QfBfo0woVfri7qrDO9GAUL+ZwcWdKBjokvK6K8U/rjK8yxVjQWDp
kEtxf0N77rqjmqHdJp+EdYS2SEqPCqli9TjHJAWS1WnFPFN2T01XvQhQC6LmvWeY2lh7ULwi4wAp
INGSLjEMFUfNGq1nCeJ6bBIyG1pZ71cRjxqSADf2a660HOWZWF4dAdc9AfW/ekdw5eM1Es0wq8dU
IXpBfY7zVEUaEJf97qeY6C0Qi5Xn0vUFRBptEcSdQ/LwnwMvrlLok7OLGT+cWQHJmkZDTQipNEPF
tIMUzHPIYohIB1ZCIB2KwtsuBlcgasXPkTAaxyscRZBxzeiGf5WlxKq/q6RFSaCTHrpWeaDkyJrp
nUsTiAoFvzJZ0tVAAA1DiMBva+5leobAgbSlJxOtkfkhJ8Oc0JNcjIjv1fF5lQ87GpgQpE0S2HXH
nfBAinsRG0BzF4mGq1eDexL7NfbvJtyMvShJm+seVgXWm4nFU0X9aTo/cX6cyBwt/JwGmOWC01MQ
u1xJDiFwv1DmJYSz0cAv1VPKA3w+GS0/sPreVhH9R8GVbPVhvU/JmwwnBLMYbDmHZDdvWGy4Ig15
tEdzZlf/FO6JQ7R6OkUxmsxfI0qjhxWLJ7bw+rqbGrSY3ygiaLq2j7bKXHK/ievuUpJumRL5v9GV
eszs8xQOTgtlCQZl2GGkeo7AWd3Hoibj456VgmAvqnjvgGW+y9Q9+A1y2W4mQGjBRF70CkdQ48pc
1jdTCRgDkKc24F1XNnF+X6CHkZoK66m+rBIYb43isUA9WtejJONGQjwevFX5vduNItZQ2qcVVbjx
60zwJdqNc2y9eDSRUAellK8RQRoPr6Ow+eYKKs9eq8uX6YgZi5Z3fkj2GtUsaYRzOxmcuZQh9yBi
p8/mLowApVM+QiHjccFANCCoh/EBACAk8mQZEkAq/gF7MQz0Tp1mGTZ0X77AHg58TnpbIi3SgBjs
do5JcgNznhJxzTvk8Dipez4j+YLhNX45JfdBh512kUuSo3Ng1/1hSwuPpoV5cTG97t8rxeZ54ye/
KzfAKhtx5eCTmXDkHrlZYrsHe49hqx4mzltAMkWzyR6mUsx4pameT79EIZnbGFy4lXS2imLRuEia
gegbtK+lljIP4fE3/qiqzjurOD1ChlopTsgvPXIW8GgnXpW5NIzIAO6aGvuDc22VMBmzsBgozlWo
RnRRRPvkXic+hYrAlLIStaBtliM4Zaiky6FdqcpJUfcX9oNOb/r9jerP+RpmRB5LslycEB6Eitk5
EmwHBzquQCz4560jDcM7h30g8hdB50goPXaiHsPt4ldk+HTssTgIHorPSuQ4Wjjj8tkZufaejFF4
rHayLoTzAR3JVZoGWkLJVw/ct2ih0ph6ybGAnY7bg4EG0KSyPTk0yDi5OVdJibE+vw1Sm9JwoqEi
p3oSag6UB3+koYLdFZOzFYtUEao+XSuKpQ3muVxDiEn3cS6HAIP6Zsg+SoLnC3g07vTNpyqSdaOI
P/az7SmIFjIhRxXSmwYHbcdRGYUyoEZ0HTPWnD55W9nyBOY2ic14lKaqyWNIFRNBniOABVUeme0K
Yg8QcmKfhoR263FqcvMGVBphNIFqtJHD7SMBBZKpu8AsjW9t9qjRpRVQjE7F7kI0Fplfehdi+2lU
NF8TTDUOjjpiugsZ/jcAr7HDjLLA7C0ewkOWKbuyj15a70FVR37ZUNqzZdqB9kZ+bm9xWm67K4B4
LXwK8DtjPro6gBgbVJwZRWZ14M4xGZA3fVBwC3a6vz8VWirIg0XbK+VAkhLEW8LajGoUO+gx54Jt
GGLOzuoRQhAy6gFU4wcI+/Y7DZxB6UfMkoxDWRpSk25+RqGODbwLAfWg0ThGvNvv8sCfC9nMJUVO
n5ewRfFmpr4cmlJHSq5wC5lVjTGiMNmTe/Sdy1rjhYAfhWoH12mi3Sep/4mDIYZGFOTEMJDba5cq
lyJVsykS4AIJzfqZ/mHzvy+izTY0yD6tMkxDizsIDLvVdt+qUXqgIRZX8pFgJGY/lR25vEh2rnHQ
G3G9Iy18XtxWDEiryCWD/zNHYuI9ybQl+gMjx9fe4awIY5ogHkzsm3NuY2RS6uZYOlElmy0/z4U1
4s4ASjOl77DpXgUdlVX3HLMVGU96xBzJtF42Y8KtRZTfxomckuVOeRIWk7rwMXzv5j9t6mrrBzaj
xjkN5qyk7+qTGNtP/agyuP5YFjSpI26p3w0RxvMhImUCq1bybZLYyTsSi3EvFJpZtLKbwQkCVUZc
55IZ6JNCMFklEd4im4NoEiICKqDhLx2/edynqktYP9YkqyOKTWTIxXnWwj+DAviHD0CIGujwb+MI
rs+KclJRrEH2UR/Z3KFUuNyRohKwiQC0z7W1grmGQs6UWSNlRUy8kW0tQoW8u6TwyUuEVI73pYpA
VHd+cFCTROXzIqbsaT1f0cBzl+qsHE+Q0/uMYtcJmpKnetikkMNMwpXDJqjNZLRn1eJidpBo48IT
GY1UrYjG2cExKv1qEIf+w/mvFCnHd8G00Q30OW7U7AvRoVKWWJJJeqdTcjDzf/Lrya/fGcY2K+iQ
Dx0b/QePk9YEzyEnU8084n8IqAySQgKAhYT+OLezGZVbD8rDD3q+CmuJd8D58GNlKEA/5BrNIkNq
3cbPKo2lHn04gbdyRtj/BzuRfYKp9tzmnAIi3mBbuU+0nxjgtnpIicxHXTziDl8UVF/x13Ss4TyJ
zmLrnw46034yV0JTYGWNcClJoXjmbzS9cZmVZnKWthyX59hejZbV+D++6aYtDdzb5e+elZUNXO+4
WRHNw36lZBI+SWjVdntJExgKU64YfiTasLfmEGy3XJFn2ADp9WmtPurlpn9tZ60/AWM+hS51VmnP
Z6yirgvDuSsXevQ6kF7ZxwIIySX3iothcunh6QMw5S1UJlVAf8E3T97/CeROXbz+nq/9hj7qdlh4
TyZcK64mWhuSsZpIZTe5ovyn4ymo/tmIx/FIjG6GqvrvX2effjL0q4bGY+KhjYzF7ULFKaa0Bqi2
bfXCDZst/PNxkdCPXcDihgJ45HbSJtjc5duKlLHa5uYY5cARlLwwLHVIaPrssnIMGWAeZaxEyFW6
w2atwKenzD6nDushvGdE5URHEJGRHzRQMgwHB6qs7j4A1YQFrRYQBSupqt5JWV/0I5zxFYO/KQ3H
qak72meQaxbnk6L4J+NFtiUsLbYrkTfNke3VZaNsZ155lAfyvqWDtzUxn3+zMS/lYNiHFOFX9NNL
4fzTA57TgR1RpVza4Yaki4huIFLxx9q+P7imWJPuJ7le1rT1xWyLOISbg043/N0Hm1e/bKLM0MvP
xKUrfoWPVa6NE/tJI0K9jdDOe76jA2mmXHQ866oS/3unQ/8wLshJF4yRwaUYfdvsI/o5HQRMx7DO
l4bxLGx/9MXuaYVLkpuNxQ0gZSfQTmaRwke7bpDNbThekNJs26tLz2n6u57kDUF/8TrQi2p8c4xN
P9dxKkF0hJ8Yd/Xv1omhs1y3RLjvsWRVQ84r3UjVHkKCDnKZ8wsBXr9XdSS8RvEG85q5IdGQ6TQ/
9+74d9vu2rFWt2C0zdkH/SrnRcxAXveml+bimMX0OF+BU8OPiACS/RFmPxiCSgPkmnBomgIFvkqR
gK83RicielESZBItDwkTSzwDf4ZQAfDU7GbQFuJfvGtNUuZ+1KFjDvTSNM3L4rKhhKXVj1p7+o7I
+bB50s6dbXTKOn38aQfQTVZMDuleIFmAubfLjdg7ugkS3AZSFw5fnQkAS7b3rPdsii8JgfQcHeFl
wjRLWwaVulQD2iZ0pxfEfbObyup6e/A5KhUZRRF2R4tpFazgosWk7I7hUdDQ4+Y2gBOFYnZupxpc
+Amate3L1roVeC++yWi02E0LxQhBNtz6KlCNo9IteNyK0pJoVUmbSBv+7ZIFst2ta6rhkV1+n/tS
hTlPg3TniWD4i9o7SF0VlVPh4okKgVMeJfyOn8IPIruQQvubvCqcRXNmNoB+WNQ89vNKass4JSxF
d5J1q8cOZ/loRR/Tx4HYKRexSLq85Lg0bDs5X5UfVUNC2ytu9h4ietYAWbj5fq57tmrx77VStHN0
C1Opay5xMpsmqTXdCMzdjMbkaEa1cs7w5zzuG/UFa6j1KtwUvhPlNy7Acrhm/4/pUTaYX/+mY37t
KbOINk/9kGwTIPpkg4cm7bAcb4FWrADWO+vwLMkVdqBKvf7H8lyPV5U78lFQXourJbx5Ma+902cn
K3zqNOdyEQU96qv0k6NTnZneDOcLTjydZOcbkirXdQawiOYM6StXBDBCtFsTdqVtn8qPqxFRckfq
11tV/Xnscyr6vKFxpapPHJp4mawtplFyXXmBQZ/qX3OpKC7knE1vFZhH1cbaIOofgpJpIy1Rva8s
s1wMR2vjK5QDyfGUuQqZFLi0JBH5/xJc7lOtXWY6V3Bvn3AuVnfi+fb3GUjb5/blbi9hw0WkDVeR
w1cQu3aQzuDw25YS73440JknofCHqlBRgO9t/eJdqwlya2DhtPOquAvWvisFe9Ba33f6z4A/hECT
9a8aCC0SficqnGui1/nAL8LNj33Afeh1Y+zmE19fSXRYykRhmfLAF4/3ujSPCR99QroPZzjXewF/
gbjDIe+mXadRHIuYsTaIauq3FNgqWHvaUoG1IZ6z3HlilD9gzgsVF+iu8dsVVYeg5TzBcq48fJg8
njDuxYVOg5thzI8XqPNT0gdON08cicZLNrJAz7NDP7swqrr7+uPLSvagBuZllIIqBSYw1bMLbfoO
XxCVPs9oKwzZE+jlBuBegMzKb6cuznAzzA5LJeTolaMi4nYZDy5tKlD6EnIkXkfk6XNIVATQ4mmQ
5Q2hXq9jEAjzyHgx+aqFkSN2Ahmp0lY+0SA2lJamOpBZvi6qKbCMC4BoOQFOMf0hkM4P0Yv3Mx8n
cyZvFOY5gJKQ2Dfec0ftbIuHreWIGEfEDcGmCDwrQiMUHP3KEqu53jeS75GtPXQm/CsZPkdYj0LF
zm6z5tUzzkGTsLqpV/JCwH/NlIJC5LkvpCio3sDepXEDw8YutKqNr8MQxtDYzFUes2ujChUTZMNN
5sVAkVuf+legkpFyMP4elYFpfBcYyVOCzzP6eB+LM0fntKr4+JaQQ9W8q6GNtqlKZ8keFydnDex9
QqNhuiKKruzebkQiI+ves/s0avuhveK+949hkm+qeBv4H3eHxKKkFKkEj6mVWx4bRTcC9FhQd1Ek
vOvErvjfqbTTj/UJxlyiuYHTcNfeInLRzaIblwAQbUDMRzSbn6gO0x1Ify0gSqgs+si6xqgAwzZ9
iTI1BWEWCrJhOtbJmXDupvu1BzST3tqyd3ceNFVLvTgsmlxr/yf/A2J8Tygcod2UkF9ZhAVZZtFn
Stk4h5W5mRPG3+eSwSLoRAugWIUSwrhpXPQ71pROC4IXWnx1Bxt7q+4LUg/rcbIGgBO48qYe1PJd
PL6A79H75rGQsefmXewlmY1QqOweTtZxrE4ki/PaA3ij0+zz1RQRb/yAJxJJXXhDWhd2s6Ja046U
i5r3ABkjx7tQS9du77JaVsd4lku4TD2KUJM3Tf/nurpW7BUyBERGynwVxCi/G2gFD7GpuNtnsliI
/dbvp4fnYNn+4Blt4uwKjjfRvgqH27DS+D3bHgKR+IwVbJ/Qs/eSwyZSiOorWB8SOhRH+QDcxjiO
+U+ybz7z72pnWn34PQI6X95tINLMqsGIgdB+ZCTWmZ70hB+lYTPfUi96xEBRcVHzX3Qiw/z0oQGx
QYJjt4edhTcL0LH7OeAkY4woxKk+iikBY5XmhAqj5x1HIHHrD+2u1amJhqH5MDH3x/yDWbRLUxrq
j4QTxod+ilXLtrpJYAb/IE/Oc+28/5nH7ToVT6PHD0pyHTT8kkEbladtpHB8Lj2UEiOho37APhBc
oGH9/2iCW1/J/o8c8a8ZNxsO/mmn9m1ELENJGLv8flKrv7H5ZvNyvjW0K+IyJZvLLfrPnGgxr74M
TNsOSE03Wmc5wSIrM4JlVvqgV9CcEgekCeLhay5FcOQXKhBzkIvHVZN3AXjZ8sRkahr1oy77Gmsk
6cou/VCY6LgmGA6dhFdOlvo3iMJD55X2p9F3Kx/9TH/sRM40qy3J5+fONhvM43bHtvdRTSR7g6ni
b3Oy0wHD4Ouq8n9VrObXQZ9O+hUOn0W5jTQDPu3LmjfM1d79KxKfUe9XQpXZddr+wMLM2xNNQX2/
g09x7sr2kgjrq8w+Xhm1ukLpplsRG3fNsQ/GwDhPE3jK6S8h3VAc63jZC/POGvLkZYFYgMPtKEI9
PJwCYRTZI+uNO/xjf/g2qValNcM4ZMKJpDMbJha9DfaUWPWTJ90Nm1rn+jXAv40mNtBZs79JVx91
g8HuP6nWTnHrzB/axNQsRh3DLIcOBZn+bpkmuRwLONjs1pUfnm47geXHe2Wm2k8CTMibaHN03/m8
PlRvWH3pt5Hj27L1161V5xaLcgYOG6tp57utSKh7dOS+Y4yW0B+UKdS9k8xjSeETnKanulCFkB1M
MgjuYInzWdGxkeWAQmEpsDDiiqlVE3jxMPtfXRNPUd2L9V4QGh3XfJuL6IAPBqSF+w/Bt4uhKczY
c5MrdszhErKeK9pALWiTaEbBA2h0Jy/9Pv6rJIVPq15oMjMVJ/cxgTftE4UZFRohzbYvVRWRCshA
eEXry1OOSPtU/Em3PAIfCJOTXTdfa+rIjno/pgNlKHWGsOeWn1vYig8tPoFzJnLBBWdPQJwMOCzO
QOH4ZRS9YKxee/+zzaZewYtbKuWQizPfKBvG8P8ZeDYVbQPxtAnBQb3U20DBYQxd0UiC8qO/DmoL
DpR6PcUhMKNF7tFff0WFmrobzWJ4+o2gOgGHSxbZkR3pnC15UUn78iWGKR/N04Vw7u9DbsrKjPIl
xnsr3oFdkQ6DQUVx8devBebfDvFluzqHqrYsgZrnZ/QKvC9v+btvUhVVr2JJ3ZEcfREse774SFV3
2K+uOMNlVLZDUfcmoq77olhOJU/seaClDSe3rcOg6LvzVKTDhHidyMXh+Go51z4ZI5XHqQvntyTQ
HBssUjgV57QxEOiqBkOT1kotGZKgDODmgGP0d75o3p+rw289S/uNtN2FN4udx0FbsJEf10Zl9qHe
RT5yvUEOI9DD6BmXq8BZbuOhHyDYpe/D9dzrZo2/paZvhMia9KNyrcrLriN/aeTDHP2JRpE/meou
n5cnazjTOIkxanWJNnueMY8fDQf4LAwp2V0EFLnp7vtXNSeXJsn73CGpvhaVBMEges+e4xNcLUAk
O62TT3Im23LUMMswlepB7Hn2YQk6s+238OiXD633lYAw8wLlOqEKpFeaJyp893iEpbQiqeHRERNd
69DYmNtDGLPkCSAWd0T+Gy7abPEyL5/RPCaGzbFuZtB3ifNkXzhC3XxliP3eXs2WjQtgY2viq9RR
qWqexZlFYjVdm+wpld7BAgjQMoeylVqEcDhY2SHn/95Qf5XpP1QJmb+LnBNYvOX8EeHgxZxgwgSu
Qt+L+vPd9KB4Mvcim5gdLObCzvr4nRZIpQFK3chF+6bgtR3LOQzTcjK1/PfefFjR1JJctDx6GaHz
pt8wv4CKjgK69RHd0Ca+JyDMl/N1Uhf34+UHnk2UnGLENlNKhdu4cDlUdDK7moLWusQ9qqjFcEyp
GoCZnTzmgboo+O9j7aI0f+9sVXq1gCyfVo7yl4bT/q4Jqqt/HKZjHzLu3XaWCPT64reZ9zOCgFkc
b/EzRN2UAH0YclFiyMwpw17IxTCMu/QAyEEU/gbdHqSAMkz4Buo89kJ83TP1xpWM82RjUbe/24kQ
k96ehyq5LFmtJNMwWoQqYsZfp0rBTd5Mc0H61VdD+NR3ncglIR4opu4g5QV7cdcc+bDf1T7qtX2T
O1zQMLq8GF3Hcx++ZRtumfSrOMKqi/pmtqIbDRh6YNi/E/pvirHFkI/h0yh6CSmy2/tg9Qn3wYv0
NoOORv4OOkLGGZTxoGG0cy2ko40q4bHhZdnxh8AbYk76WSXkdv8u91qHJv2YI3AqGt0RpCHgrFgp
vAuMEOStvdhcck9HewIs4VAtlIHrWH6Zwyhu10EooQNVgKvRl7/xuKXOEv9pUMrNPEzDgJPBj5Uj
Dg4XoZXCol0lKNV1ltN4yl5+0CMlLog80DcKJWJNAVCPpdxTHnXieeySeyrBiMvLnjWJYKBmkQKF
7/qYd5wiflzmAh+qVdquXLIa9+xDuBaelgYjUmZvjkaInezfPS94D8m0aHhvZo1DHmKgd7vruuU5
3Uvn30T3uAfvu4foF4I2H6dsitnpA9LSM82lI6YdGW+GKh3CqRHUeADfUd8c8WA7ZniFBAvpZR79
YLnd4dy9KPJXjwagAivf1+SBDMmZWenYU/PrNV4ulHzPoC8pIUO/pO6iMgARWUwLZjSDzMmihdgb
e2StqAFZ6OnLwgKgFxoOsJD8jtKV00hezJOGj1W5VmrpXOdT96RZrj94nXevCTDu2rWq+iWRveSd
Qn5yq8+J8qcY7d60hf09jqi3L1dX4K7qCU0JidBc7OytsX9McNgq04nHd6U4JEnqYoilYsuJIVsW
2wHm5ZPvqSYFOl290dbzi3v8YAoLEW2fMWe9f4r8puavfeCzECllPwarDzXrRn4Y+M8EY0wbfMRT
z0J5fStAEkmjTJh5QYuVool+kXw/WllFCYVu0r65fp8rmAyRd6MjQDbfeXNQVhFPtx7/SAF2YBXc
ciFjCugkF94mAS6I+vBmlkmaPUsIfR8xRg/iSGoOfRsM7PBQtD5v8f0hr32urRzXFoBr+0A1qrYZ
7BL6WZtFKODnJGyNi5kxh8S8mAgKryeHzev5pyZHeT/STIVxRAUB7qLhXpJJqQ56RtX3REr+9YYA
wan1QloAX+tUxlUw25ZLWQxRDtiNdwVJ/CGhIp/gRo401EKk4jwB8rrJfpACFNFG3wSdILb5iHYj
jz1rR/Bqsir+hYR3kT9tcv4U3CupGDGoR1N8eTAiFBk8VpjLPgv/UaiWxiT+AwmciDEB8hq55rbx
mGFAj6weSotMhnhYkatWnCsyT2DWAEdsyBXNfVgAZwkgkCkF9tKGmeyqLMr+T5I3oy6EPrPE4r4w
h4klwD2pEKwb1KGd7lGRQZogfrSVoa5je5T4AXZ3vnnLA5z6u2EJ2DXkPOiKzeDaeP+39+MFMmex
oGMUUyvHt9HjFE6SvlzmRO+fpQnW3emi9CKNvUJhNVyahsDcUGo7Z5nBo9PGGXPYt3f6SUeAd4SW
iSIK/xJXCHW9yBBdHqQjOTWW5FiAL4nuIjd+ua2qnl4qvLMBi15uRI3vnNi48uDcL3HoQrdW4sZ+
tJ9+LjgY7WGOFJcMAXFdLeTbMGQj+AcgRUU/GdTCWr8+VnGYtMixeVCfn0nSGjxhIzLVWFIKj3tt
Vn7r2ZR2ndiD8nVsP1g4OCW5XnWcO8LGA83tosN06njY0xccSK4jZuuNapNC3j8tXCiLZ/nNVTWS
C7rYK7adjhPrORfKRyziuYrQZNPkTuMhA9/2MBlJMQCpDlcVuFOvX1TpGBwqUPlsgj3LIT1MI6vo
GQSm1qX3OuNbb2ny5P2cpcjjCjifYw1+sgxk+ubBhpSpEC0QmF5cIPrHf7LYGDi04gSOg4JnKIvy
jW6759XR6zXg/H+SyNO/s6wmaKlvj8EAhpqT4MeQqCcAZyDAPoQnNhQkYTK52o2jXl0EY0GOvU92
928dBl/u4LQxrOSL2pAvR9bj9zal9GY8zVoVPr2Cb0Madj0f2LmIrlhPkBVT2sATBaQkizjVn5y9
zYmjKVsykDzrXGBPGQw6EKBQ1Qt0VxaTnM8zXNGERYhBm9BWgIdTgnTL/76g2amWnWGm6Bf0PHGg
f68jED7ALFkeTKqrczCWRV0Ahct3irKGy3VaLz+NKN4GBmn+feATFsiPbBWToDDPIQDwX/aalojq
IOQnKSHHeFE3XXhq8H9L8bK7mpou2YX1YPyRbLkJuocYSMP2uqB/e2P9UqMSJrUdW310H3qyztg8
8UA2gXzI/JqU/sE5NuzyMNhZmCr7w9D+7gz9+Z6+xoAOhJx0HuU+eDYaowyPliGkJKGIaZw7MR8J
6JgOeyPpYfY8LrHhYQqKWe/GcNFb7qi7ytVqnQngvi6Ts0Nm7+cqg+DMp2NHnyu+ERlqsKYcIF3Y
IyWJyfpNUbxFQB/TdWqh9CzbuD3OzKvuFBlk6fBFJdU7FQb1qTa+o9O4pUQ5spPShR51YymFQRS7
oaHVgoT6vJ9QuoqZRD84la3UGFSpebV3z4flFbknn2H0HnMrLWNJT6V9Ei1RNNNcg0RP7x3aJFXZ
lLRyYGeYlsRkmFky55DU4yv1flRfHcucNsZ2puDUrs7jY5Mdwr8oVDz5ER2n4FnR0Q21g/6bFkYB
HA3+yUdN7V8udCnjr2inqXDt7DhEAqnQpyHBY2pv9Gd1peSVQRFVM6hTF+EB0JJTKN/g2w94AoE/
fCAS2WBUbrwmNeuOefKt9noQgrj+1vtEQcvekJevhj1zygHbKd6PVOO+vMn/fIiDGByvUhzN76cc
YqehEfTnCo4Pmkv0ZXHgjZ/uYGoR+yETgadse2QLbwskNh6cZ8+TsllMJLmndJso1MlnhC3H1qjm
khFf+8r5uVM85aAucn5rxPSCqe52e9KGfANglHv3M4Ybl6yhQHc8V11UB4Xdhi3jBR5YNKcilXEY
PvFSaBpAI77nv/k/3Ug3QNsNw8JP9+6MLCpWopu/Ct6PGh3MqL/XIAdA6+PciipqQEiiC46FcFUo
QBYTaxWOcQ9l0mf4gC1qIisU4ZxfNI5P9S6wvXTXcG5IZNtdT4pz1m4KZdoGvcqoGHFggFFjutOl
oK9a++Do4zl2EvYzdbWhB6cZ05LQOfTdQQVfCUW774WFEP6JbN6rro0FQG6FBSCj+BZqe8Wo4J0k
fVUHT6yaPvyjF9sctbmhACY6lsK9OyEPLylKV/bJBdGHtKBBejScNPr/ysoiO7TwzSlGSTy1w6l9
qvRQ3JRgdezMzT4oaitxL6T9L2UB+CMxrRfSxEB3yxDmWxNL1T6ikGZqSoV8l59K6C00eS+ykpG3
7E3bIOlUKsdBDqPtpXN9xiqcMdeBtLBt2b/3Kn+IoGa+WwSEXWlk5e8/Tgs3/ynEWaQdXJ+EEoE2
dhOyS8/8/ERGKeH/lFlkmBMOOMG9XvcSOQhiqgra4yADTAoTD34FFCEUTOkD//yEPkplk9alQzBo
d7UE3JX9z3Eq29LDEEXjabrGQLUsStM+8Rp4x4BQ9NkbuJeRZUEYcU+lAvCt+QqofrgJeDwNA7Ms
f5qHw7BiyrVY7sSolFcpjhvpkKn/SQwg2qjgdz7Cve/NP/OsvDeO5V3DKikCZuj4CKjNToxwyDJ2
Q6BIXgoJp9PXermdMu92W6J+NRffaMeLGCaNKFP7N3O94S3mJsNu7knnPHaM3M72Lj8OJZ3bMPFU
ZxMThVMiF6L7bqqVB0Sks6z2xJZ8sRy6eevRZcsoj+0eU1iZ2o9nS1cRcyzQK2oP0QUU2Np+Nvqh
o4ipfDFjHR9oPF6+0FrsVp/sJSai3y3iy3QOxjJYBsQzHZWGttwMjtRlIsaLbzRPBF1Sjk8gYJmd
Qub/0Mj6rNukKOKAqYdy1yP4SaKKhEb7Iqiptr7vXN64BDU4LCVmzml/VaqD89LF4cMaSSz+O5YQ
YYfAibes2veMLjTnyim+cYr9ldHHpsLf/cG+U/I0xaR1m2q8dLjZInn9UrJxWgxv8sgW9DN+9mmM
JFnsqEm23XTrU5m/DTezK3EJ7BwiVXv0V53vExVD4fiqI8kr0RKCEEift8PuS0p0eMKfltEV4hxM
8Jlj6XU8aE2CgZaOJmhVZvl2QVHKUWrd9Nzn6/Worg4omJNS6ABIdofu+eFTOreOBDog34yqpHZr
a/4Ml5wpp9JjVygPE6PTsj6njysrtkNfXRnorhzN278O9GuQ1L9SWvhNzTSgXrbSYNNZtvYkBB81
St2Oer5EGpOv3rUIiJE5qWJRg6awmN5Fk9wdeh5CAO8eQRxHwlvoVzKHMrOnGPyZyzYtg+Q78SlC
U253Kx1ZL+yzHo+3E1xAOHx/YFW0D9rdRAAB5xdmVmhYF5vRDvGlYMzRZO4r5qrVBkDUTi/nWK1K
qn1Pxt1HRxeztVbagYt8GG4bRkOntktaLU1gmvctdoFxQNweCdRMt0S+sgWKCsfxFMcPfEFJywWW
4pXzHsJMcE0wbBxMiMg/4pLTo/tMQ/Be+Js/VIeR0y0Ek3bSqQyKSdWbhmkKpqTc6ZylHQYDhRHK
Amhtb8FnGdU+cFJETMA+J0f1k0vyxAIspPxnqui/hhe/Qr/hAofCS4Jj4FKPLPrItwszqy9RhBjW
FbNCISaoJH7qiFMEsHEoD1LEOEfoLoWe09DvdQB+bYkXMgeeKGcOq2wEJ5Xo3G0LUtdrEyywDDzz
wBOSWVrTMkgOsfs9xAj7yyXkRZXPmkErCAyvDQg99Lna9mXrYP/7CcT8Q+q7MOK3WE1K4EV0/EvC
8MEuADqgwYwPXktLGyDCNj/qa/NLaU5clwod2Uhd2+p6Scim1f5E2Ml/wGZIZpcsStOy0T7DB40r
3BqbdRLP7zfMpY4An2++ea8T6qByR4P3KwjMpw2hm27P2hD8PBHT2h/Lf3dbFZkhJHEgl5k1kOWM
89xjv6LzcZ0rARnVVSu7n3dUpl0n7Cmtr9TYcwuTFiiQ2HrwVhwpG7N82uEcRmHbA48sNokI8CeP
Ed0PExt6ayboW17cPTNZz7TiOb+FHxKfzdfnyuuq9LBzU1UZEeVzgxLZohpTBKRZErjhWFKTpTb7
h2fZ0YUGqwYQdS9amCKEz6u3k/+SN7NFHxMcy7WBY3vyX0OezHRu9pyJijFPXY7FOmUxZ4ISnZTw
Cdg0lPNSBqfe05ZbxP3mlNYYWxrxOHXTW7z1XbzGkDfn1SOEXfEWPuHvg2/XMSk2F5twXARxcazN
glyFrZZPSnOhVDZ7H63SfNnMTGdx647/xXTxPPO/9Giq+C97ib+1Vlnohz5vAnZh2To5KN7KzkJI
6/0c8CtFNKL7NcFJwhFJMvuW9aFnMwNJDsMtNeCUCl29ThWohlyP40DFt+NQLTM/0GYdSxcLLCMv
T+IbbUy5GHzJuXdJnVRWf8LifTsLG5clXRrGPFF03fheVVHlgaWG969u+ajADYQ4qwwVkdK+W9iP
i5mkxXNEfih6jtxtLPa/YxE6sNwvqdFPoK23dhH/SXoohNcIWERIYnn1I/62lSYe35QytiZ9+YmH
gUwaCDwP5yzWakVRCDxHKOKEfSnfiwLeswuMeQGaPdMjHaCbH1k3REidCfcp+1EXheBEHelUgV5/
WpM8FI6bysWbhifuVdR62xjZDcKRB655q/YytnB9NbCzgyt6HgEJZyUNw0EtomDkS493WhexgpVR
UYBpwMyDCwUuTtU4Nqcy434T7DE2GTx4iypmjCKXRVRfHkKlvgRpzRvL6Z0CAtu/sKhvwIvTj49R
ZqVTdO6HdW8sUp8naHNx47Pr1qVu+CNv45KBvYOPLj78zhCBW6pn20+4PqwcRJuuB0OqOP1B984D
q8z5qE/ELHdjKOBWkXs3SUma7f1i92XVgZopHcAcv+0jhpdxbGQ5xw1b3WJrtHabus/50vEYpNJe
a+2ue8VHOaqzo1iDkN0f7XSr7HDMfmpfqYCPjgGbQz921zBNB1vwJ1Y9XLc6dkz1UkhMEvWLUdnY
2nZM7TGlm446kF+v18vg1gkpZ+zoVBDR91gUg7+yted7rw0lV45SZUuFkL825/gGF4KvwDLLA2+g
8w1OjyA/AAHaXuYeco21MhlLI467szJc5T+cl+h+eVn0yCdnOL4Yqyqe/q3KJuPRSkuT5ED1NR9l
xb/VVDDz6rOPC0GQGsx+CEUr4CwFVlXRFMNMgB7lHpXj/YWn+Fd9VZy/rLnt1tLFGv9wMj7N6v31
Fi9e8fzCx3YDLlhK0xInVMB1uKC3jnHPrE7lYx9DaWv0wsuSNNfqTrYEM/L8ps2n3sInWV7tvR7H
BrtWTWOZNZPHMwFYe7aVD8LyTtLOHk1tIpIoewBMyJBnTwYFAqhIQAc+qiOaymjmSAl/uH5LiACR
20+A7xOlmYZQ67jwGz2yRuq6KdokdXu+08K+V1/GcnGEWcIbjmIt5Bkizmofh8QWYpKq5aNe18wG
ngtymf9DQEY5fM1ZN9/vY+9eF5i19XM970ohMEFYuXCgQMbrkDQQABvA4OSVBbEKVQdn4kxVP074
lccrqPmZD641eyQLLywsL9UgJGUjIvVnhbZKE0QXVK7dBXdNsT2F9dfW/JOCCkJNenHTqQA0tKKv
SIyf9ZqmqOxLvyX2wXcI+ort9ENBXHS0lm9TtN9QZMJmp9SHFdKL9lIA122RNQwsAmlthAtluiO9
Ghl00sjqUz1xIpjwKsGU3BiCJIjPkirfFZBjseGIyabpgD27BQ/z/wO1bM7ufBU3uG/uEc75YJ0f
EaW8fO/n/Bv8Zm8rckEC2nYy7u4OX5hvXCuWYPjhBMlrkABDY3XBcktuq/HSfEwFWsd3AtUaeje1
w5+rwxzzHxxq4b8saUsEdLN0Dc0t/I5JgKVBqUUGmeCiw62bZJXcP8B2FNUFB0iuVWpQ0gYE2Y/2
aDIEIZ5ijFF2QoB+qZV0v1R75k0GJYq4JpDORVrsaunIEWiY680hsNtvfzb2lstcso3ETSgz0u5q
Gi4A6mwaldpnRbrVRuFIrpYg3z+8oU50HMHp6lsYJSP2YgQuyxhuMJ6oA76OtYzQlu8fIa3gGM7g
dZD74CHj8TIGyosWNm9wm49hY5hCMckRf3RBH9o69YcTOzqwHTv+BTRUAX3m10C5blhPIcM+32Pb
xLCvKr8/Bum/XZ51B9bR8Ep0O7NcfTlsbFHbb3MqxN2dIi7NAxIPloiVNw47+n5kzPk6iV8qSbOc
7yCdJhSRBjp6w0TAnT74/InEI5g37DxPek07KlzcRBqge+Jp37cEcO2k2ZoEC179Xy7wE7REUWBo
IlIO+v6nAdHIHXgj8GJTKoYoD+JW5x3QbMZwwEGYUcS1BbWnQ7pHGx3LGt5A/y4mQJNt1CgGkWGG
yumgxjmzsASwWGYfThmRJXGGu1JkBa0I7BP9vQ8PK3dMb91X5KYBpm3X1RlI365SeYKhGcGP2RX4
0QDS+8JblQ8b3NKclvufSfo01Nn4HUyFTF+INXU+XObGkWP4X5QhnPwg9NW00feZTTBzoYoNMBrH
V8CJrJfW6VLbeyV9/K221UIY7X/0ctW8RWkvCMSBYMjNemw+BZW+fh/vez2ldv5+HVXhjw9GqX4Q
kLDM7berOsifKg3NbqyMUV0td55LPf1S740kJMbdSYCE9fyc4bsg1Vcg/hw6Cm5X0AgxK3ktfiX4
Oo2s5hNo+2790ZSiqd7NrWTtRgzeyqgvh6d/nUdan+OwnPQRDhXb5kWODtGnNcowGKd/II24n81i
bxxZFUD9aX5P3Iq4spWApvHuBaM41E5cU6F8BQZ9zNyZrWx2GpDm2gqqJQjh0/WMtn9czinioeFr
zkiT7u2/sTSRN4FggAE/jnFWswUvS9+MD8BCmd6LwszB7BdkptWSFAlKJhMDnJ11BkzlpuOINdBr
6HBZ/3Q7fLqxmi3TIvtY4knE1mwDphKlkosfmPsDOuLWschcw4wa+kvndrWONL5K44uJR54gohte
VMbpta489wJipyhFOvZgsJoZ1pqIqDc8obycJF0lzo0be8r3m//ZBNvG8URsLhO9UGInInJ9GGHJ
gxQCm6EabPiycZSwoCI1+PBl705xubjhm6fAhu0hJ5IqPYhAofp+jYfEVVqYwNKImVxlbU1euCLE
uaB+CHVbllmBAz3xbf7QxqqEkD8lkz+1TgFFSahgsaWVwICUwCbir7KTjIrz4lpjJir0oiCoPPOi
/QadRaA981QC2hy1QyTWgNYwJQV3i6q4f3TkxM4GFKssL8iR8V55rtoesVaxmwuFq2hEKoa2GbV/
Gk2Gx+F2t0s0bvrlQyJg5Tf2xrzEIHlgtW3o+QOwcMzahDYn9YM5U5LVSleVwWPwwr5mK0cU3hpY
wT9ptGv/KfvnkFB40QYnJx8bk65nOxnp/D7j2Z3VXvkVndrgQEMoi0oRxsJJU1XsTxI37c7iXWm6
KGXGH4eXS2L4wx7J5j34hTen32E2xPcjsH+AsW2Jg+Tw2kIHoRtvA5YFFB2fuFuH5fEY6YAmZD/e
psBMMzcxKIJXgFZA69am53s5G+3Kw8ZUGeeSQctYD5oWcxqWOBOmB3K5xJPyILqecwK1gU3wpEVf
RLiUOTPW5L+HUI0QjBw2PQ8eH1oouAk1aK2SL6EyyeWxg93Bej1Mey/NWB/vV5grhP/R2mwNLaI0
xSqWY7zfofKqQFgFra3+9MGL/4ok0okb+ZHeik5LoT1hJzbedRQRovcyniFrmfPNGMDviek1EM0s
Rb3eM8xT1GH4eTkl6Q9sY+vgv0YaFHuR6KJGOlUpCDL8qgLvKhERmDWNH9rVZyUnX+tG7QQMDcMt
hhhctgIvxI+z5EbwTU5hxJeAGbvhWnwf/qr8Y7BQGAHll6VvNSKZMDccvJmcrzG3Ln5nzUHrvjCm
SsOvJZzQonmW/4eCAzJ48WIJUPcW1IJbxSk8ijh6Q78zmSl+5qgA1V9p44yRBCfXMtlNgJz1e+Ad
4TI6M4B3IyTv9WsEAPmTDBq8M6v75Uy3niHfWRMSni7VRAzCmdNl/x8JPorHwRpUebgX7luK/fjt
IqF8Psexw8zJ1K79jKY2stfbKF38MeX5QRxUhfMrk//pB83I2cGLRz23tgEDtzmRQqI3oIX6Idk6
FdC77BtKtHp30qVIoOg6Rk6QwcLcQEnx0BHRbJgk11aJJ6IFt2rT92FamfAihTQoA4KiT8bw86jD
A/n0IhZhsZZmHMaGgNlhG5IFlQ2exxXp5hsQYmGOeMqa2OF4U5u5ZsDn63Cl3cjNrBiKxrzO5Ecl
qlzTmbhrsyPQC5tp7gmKKxmMTfj5w5EuPhmVlMJkXJIn8AQTdirh2amlM8YITFH1HZdug1ZPBHip
oMXi8Xs5uit9h4Y5LFaXpxgspgZqKzU9DWvv44k9/6NQ9P/+WoAhGyKVhvGlWyo+c9QlOYhvUElb
pmQBJzU5Tkkk6rfZ6S9ckFg1gSRfB0IwaUgwKzZHEELotdo9Dh4ima/4ncBxu84yDPEYuNQvlqTY
Kf6fYEEIxiAlWb5QRjcXq/CTUzh/DYiMZM7OD4O0XmGUWM3Pgl/9Jr6IUUZTLnRDJlxcxc8Y2XOg
yysXXFy43tPk8jr9y0KvqBpxB8GGYtPN4WuLYDQD0qxt46fvrhXem1JS39PwViH2Rc1wAK64DDFs
jvt2G97UYRuUFoDHAuFQ/poeP/swVueufQn9TapQ5olktnUHRY9lBa3RqylEvzC2GEEgwzHfVjpu
8iGf+04eM+jtb1e5WJllTnnG4pFH28Z+5/2Fsxl/H9DfFFJZ+z1VFt9RhC0SCy4wGFfdG8+AYRJI
EUgn0QxS+WVRiQkui8jcLHP88fickHmeRWq0uOyFI+Xv2eQaIi4cWR3Xq/kkj8y7nVYyx6FhvDYc
oHP4MFOgkclvjuklnGIuMkO8uU83PedsQeLhUfcOWVk2bUtbEvd8kD+FSL101DQXKBqdUCLYpmIC
78j31ozgAGTg4yAcfFJahU16FyNhm3kcai4CxDWg1oRWCZ2bCNGLiZsKs1yvtsx5PaKAjXvFEVPD
22Kyjee2mREI0hFLV8tARF/1NEBjtu6D+qtfwZ+QeKOywGph0qDCXaKkX6otzD3vXPEsUpl2czyE
mMR/71JJ9nVkL/xuU6I4CvyRTlLpE+bbLecWW5UR1ArtC82f3W7w80ZAFZfqfYQeacNdZ0fgsyyF
jBhbAZv7srRLEdGrNzSuHF7dpKPywWsqF4skG4P4wCerKjHqk4YQ1+DDw9ZASi2k9EK76vM5RDMs
WJ1ztMw3kjfTuuJpn7siK+RnpjzHjk3Yimf/cSjka4VJ/k+bNWrkzucaTzVW1yvgTPNaHxd+wmo1
Huon0tmrCCIP88h8mFWtJbtwBInh9z3aRpI0T6UHMHHPe2oGiJoI+p12p5eUSco5wlWSAdBbwLRM
v571H7+SRDVlCdBSNuoZRZAQqhm0QlTc1OqP/KPB0BsWS8J4LoZH3TUkJe8hjMz0rLcy3ccbFeB7
kVxZCiNpf72ReMLMtZ8XtkVY7fB+juV/bEcqF7ixh5ot/FNmsBOGnXjK5wTOEQV/A/RoRttD0JbI
2N2L4tCxjk0G+OmiIbWt+K7inC4qEiX1g1H3AJr92+aQpCcsCEbpmmZTgp/SK40gbtrpjk8lmHnc
bpG8v4Fokj04vrLa269ngnUuVc0rtSQH+r9XsUUua0FQBnHWHFEOdJYbZ0uG0yW3il+iqnY4oZgX
gq5CPzBupbdyoYeun7GHg9oyEgZgy3WQB+zQdh8iHNeJpkha/HY9NbA84j64omOBGGzFU0OvrI9d
LyA7iHivAwGMTwtfp9bK5kp3bK0mFn/O3OScQrajOwm1wTTYAHqVjx42d6+Q/b67X6o4tCIcwpqK
X30KFFneTwbP1Tiu44R/O7S5NJT6cIFNBvf9IjmwP+MQ8EfFRESN8zHX6qdj8ubFhcF2zB3liIfC
VDUOecI9SUYVUWNPTzo5r33407deEN6J8l+yZ5WGY1z6ETX/y4sGr44Sx4ik9LnKfbhc9ECDqGzW
Nle5XHsdd/TEWnnZ/8E//iy0p5owcjP+ezJ5LO7GU6N1MZx6+hhnBJR9seeKvyvMNxpnPXmBx5+v
uLj7G7OSK2CVP+CyEbEB4Lwn7qKJPgqLWTX0MMrY3d/V9mz1BuAdtCVifgvKuLR7SnpNd4ZIXwmp
ElR0NW9xzxARd6otA9BqQAvU9wIC47rRhv0C20hNppuLDqb+ZY2G5xX82n7EPDvqSntfVDuBISHS
3dC1M3Pnt87BYduNouUSK2JbfM345VbTo/z3eFIPxUN2qL4FCli7TYslJJCJWfY9hV1hDWOaOQAV
cRUMSjHr7RTNlHeVdNJDV4avZ7H559fLQky7mO5YtXt0IVCLUAYfEHmZXTNUsHphuK5M22Lg+0aJ
53mLy9noJqxKict+RBowhUwk6Z7ZiKHYN6HFejFJk/3ZJpESdjNZ1ArS18t+UBSWXO/C+uppYCSQ
tuQQqOwZ1WSkLnxic8fXQtzW7c8vTZ9dUf1f1M7v18m9WXT8f+DQ0IA8Z45pF3LGOmtPN9Oz+K++
rl4ttYz6NVccrRsmaKyYnnYFLPPRntQGQoKl1804hvMgAU6W1yEJhOMXQYHBNEuEwp88ouzcw9ed
FCx9Eav+P2hvtLTDxltm60JSL7uRfWaBKCUCoemiJzjLbkb6xoYksoVw3G023HCFgY26d/3tBpeg
ICaiurWuRm5xHSNUf8yAUl7tsK6l5R3i2gPPGyG+1NcOOXDFlcjLzd+iWvZ/0ouWEz7y3lGZbj3J
K+66mKy+dfC3oyaYiUxPFRH2PxUXlrqldrFgCpOCECeAYYzcGcrZegMeiGgKqnjLc3i+Uieq+5ef
cgLhI3F3fWdbsqOmKpXOE9/q/AC0y+lxZj3abwCZzM+UUKXMk/MrbzVNF2UF4IwKe8siwXLnrfdc
u86JbhK9iiAucpJ8ZVfoen9DITEasH3WeMqCvqrEIu2SciNlCR73CdeeQGugrTPUFpYwynJuMWU7
Sivop3IedsFsqmRcAqPs2rYoosep4BN+JekCsNZ7Aizlg80jUqEJHhKHEW2wsD5HmSX3BvSJ2bPR
Qrza/DQxE9jKEu2ODPh2U6euKdeh2zU4RVkBXOB9NSfoa5P4owdHBMAfSJGy4MBAGIrzNU5tZtqP
EqUhjxl/gsrMRpysZq6C2hz/8mDqZ0E7VYk7hVXaSZ2zmRFC0s8tocBMPdlptLOF2LkqRiKPsWRB
gyxuDlHSiblvqhflWjDch5X3GMhUNIamIATOAotKAR1OGB9pVdTp63QmJ3+EupJbUW28Oj3YOe5B
IrOpr/Q0xwNcPHgoV1k/MYwQZxqnBNnTakgsm5dQiOFVoZHvKnCvpeXXMPAjaTzjJ3+/D20DA6C5
OyBDtkL9Kmc64lnBRDH8OrLk5xYfQoZmtrbudWsDs3TIzeN52AJ9wcCa7aORzCHFK0g+2KRxQBCy
YM9zKnsWWCV0n2n0GcTV3dvrR6m7+HMTLrlhKb7x4qnrn8q4VTC8LFMgry3asScoQHP++2Ix3jlX
o1jQpQILdM+0K7yiPRBdqY2hEXyHhoKvHgxeTYJU9iIOphYJ7G8iNLMalLWZclNT6xwkrhck2nGB
iwOUUvt6AqMb1FHd01PllzrI2WrzhIAmytE88tI0/nP7ux+InKaKzWspoxYeIFtnJEJAFec3lLv3
qVYYLB4S7e7LL3+wDe9rWVYzTFNeJ8Y6eFV4D/G/MbWaZSr6HEpL1DzZ1GjaDXUXzDLyKjvEPvE0
xoMzr1U5BSTocQZimvUYAxcs04lyl61eCpLRtM9SN44e13JHYPSSwNsgjkMOlvw6TwIBSThYh0EK
e/PJS+75EWws0EnCGk2MH1UPHlwsNv1w/ZvVRoHuTY9go0TYVMcwzS5Y91z/Bqn4PimYzzZ4HBQH
l6gNo9J9cY+W6k9Oo4A0sXVcBvhGfZsWGdvrJpLM6gzTPod2avQ5KNOEw4nDI6we03ipFeP9BdA0
51QzOZJlJsNpXJsxJlGcvtRFdEU7IYKLLld8qhkSjEpyLRmHDKmd8MylzIFXEzWMZR9RVfHxgp/2
zUsOgonTDKhKCvtQu2wdEErmRdPQ0RQh1gBENSM3O/HH57tWBCJPY32yZe2xkf1Fb6jKC5WNyk7Z
1ceevKGuouql3DQqRuCUs5D/Xkd3KCzBujIJE1VVh4VmqPoraG+5jEy9+LPqrAOc3lNlJYYI52N1
zXbW8v7e3j+eP4pAwND/+bCytoi30HXLxiaHt4Xm77ZaYVzSXLvoxnnBYcA7y7N9gYTloB/51jS1
0ApLq3BJX8KXcBDN3I4iSjEXjpiSISyB4YEmZfCiIB0gS1JIPqzmrDVnHvsI9DYY2RJ+mJe1Tw+O
6qf/noSq+EUL1w+ZNMjuXECw0ingatsVmtn4BoaRl4PvF5yqDSJMZV+NTWaZRs6cgdp+WL/4kx4J
jH12THlTECN3btrhwhxU9CQ1p0VWoFjDl8CwgOLHBcIRdmGGkbRJGLBBT52g8wpAo9asnxFm1pOy
HMQ8y0x3TCvog910NjkZEymbZnxIomtsSmAi0sj5eoeueBBxK5A9cKBrhbtv3TdvFlMqhOgyvKEb
ci4bVed5fGfif96r4RnS495Tp/Scu+3TvnKn4beLkOj2ykCCVZ9IiFkGLZ8S0YYBrF6A6on7igaG
W9A5XvRwk0DvcD5vY+SZBFJG0ULBWlUDrKdlQAOgyzqPLvvGAvz6uQ82dEnfWa+XI6hvIGzhSMkU
k4fjk2srRcJfh9cxfvRiLcas4STlSbNN9+LA0Sczf10XqGQ2AkZ87LDC7/1dAmquExj/79Kfy6Ub
D+9aqbYpOnzSIba2d+9/qFNBCUs1aeuHhMQv0F2+Y2qpBz9gXNmxXzMG0CrMYhL1AsOUCRWAhied
g4ckVQp+94DOqNt3RkELUsQjYw0Nsbm8fbbvrtOxPwPknh+rZ6/eJto12b75CyX1tdgvTho2nlGO
5PNMDhyIOlrJVUuuyXUIgu47e5aNOoS2HvkAhtv+LqJLBGA3G9rLkyV1Jr+x3YeVaKDtifeVtLqG
HibFyDodsSrpXQhQqKHY4/fnKD1qIefKTnaYRFRt2n2HwE8WCghO/1SyZJxgX4XVGGIaxqqJC0+5
6uGr4N6ZgXaoIJnsdy+l0dWx9K1Ll8cKD62JwCw9f5Sgy3aCAcOggBxi5JXuQvF4w87Abg1OsgAm
lbFhMaWLJ5KCtlC8fJb228mXlG7puO3/+hdQOAZfGFK9OsM299ume+3e/UqCJcubP6pGBvO+NYbj
kq80E1Gjx/L39rdo0wy92PfqG13zCJuGZLy4JtLrXRgMC72x6mlEWMbFZARjKwQ6wHcW6L9pnKTk
FjR0YEyzT04OTwNkFs5UkGSBQd14vf/9t6caLsxMV3On+5S95ErLMetFH0rxZ8Vn/9VUvKtF16oV
Dog+tCyWspYY37gaVz1nzNr2gNE+ftA2bxzthW0N8qXJ7sPW1LCWcBT+D+ZymHY9qEUj3jGRbASE
DzL1Ek19hPtZoFdTTBM5l5yu+XcVc6G9ms5PBGhyigI6nN98kk+HKb2UoyW2RGzOLhjYli6XPtUc
ITp4dAPfAvvt5coEHHLkws8jgezadmaCTSWgUq4fcccrXIRLs+QMhNJK54rgKTC+lcCGMAh0uE4K
aQ8xtwvtP+u+HnDl3aRmfQ4UcK6xt7WXGskh4XpFPtcicOIoBg41iQQ1inbullER/D0Ri1U3RABi
o9s6hdaynN0Eoh1RUfzYp825+PQA/+WSpu3+m6Ve5e0+Y4o+pMN3tLGVtRbT4U69JuI+3HCjKbfo
cl4YaesbDRuQqumVF6ugHVnBfID2+0UOla9dvP6HUZBCbpnr9ZYbCVRv9IU5X6uG9o+hi1O5VH3X
ZoJUFNadaTgxHiH959UhHaFkpbNEyGEnzAaucXl1xQaKZHlSD7GRI6ReIrMYUlMIdeeB8EcmmxQb
fSExn5nRe4r0nvkLMNWEoAmPTeT98rC3eRvFtIGNExCDmqtJ2CB/Hr8pxTmzBj65ZOPbZq+qBeyQ
rAjXR5JDmXiABd/wBA8KRDg6ZDfjuqzopnjhv2xQOa4VayyEq9F4oYFmj8KsOmZ7Rxh5aOhI2ON2
XTYFEpGWul61NK5BNmTWjJsWi5SCtdMd9gLD3FeugflX2jYZ9R2FvZAHhZ65exIW1SMzjNmLIhTn
ZR+A8RYAbzJ/LKCUqPMjVr1Bkp68/ba8fpp6s9IPG0yj++txWBtWR39gLWkzYp/V98z9R/SbCv4y
0HELqUljcT+XSBCWMA/u5CIgPH911l8QgomXCGvN36Zj6fLetBA9+aO/VHOS25rsBSLROQtc8i6C
eDOUPlbDeD6aFLWtZ1uOymSGyosg+JAcn2cPt3qDH2oSrPrSmaLTiep1U6+Lgg2u7W+Z77CsjEwm
zkEvJ3lpiYvzqbQKQ/5RBABeTOyprScQ9WOACQQUfKlDU+R1BiEdqWwUhdBOeEpzeYOptYX0uiRJ
uXY6p1vMoMYmf8K35vLKL3cf+82k2/SeQtDQ11WE0ua0mmE4/fw0bkIwKLh4bjw+BoFU2vyPJHYl
9UVqUaA6t4sgnm0W5yrRYY0UCfC5IEzL9rzpLKAuLaJyQo/h1KNs++g+6RSXXjDIxbVHrD1sbwIp
B5R06iuVjQ3uBv4EIui0TibenICV31CscbhE7B+hfGtjRa+6OZkfdI4ukZF7gxmFLffEZ68Rlbk0
dBJwidFldhRX7RG14GfzFUqXrGBRZ3mhkOA9nNUfrNeMIOfkkBXEK3J58tgedUUeECQHDJbvyWCG
58/vEKEFTcvFJqhnNF6FgX6CHyR6bq8IuImtkMzp15ya7CYHYGny63FKCUcTbZBCNxcnRXj+VSel
5tThzHQWAdsoD2IGVBb7E0ODAFP3xuWlwV+myRGy7QOEMHQi1kYFtA4z7E+7/XP6pSDDZQFlH4BU
EbRKbPuhs+P41MtY7+K1Veb0rrSuK/6tACK9/sRQVC/YH2eFZEL7+rLk6q2bf7QCf017oyXsoC2k
GxlGDQ1si9UpVXTAX5Bhx8ayfRyNN0U2VXPx9dg2vsvnaTzya09AgyCKvd1OAgFXNZ2OaDjddbvO
vmWPpPlYcfsB2lx4sOUGOj8njG/0GrwGqwRo2IIYg1xHrJQcdED9bNG5JuJtzvA6LqFIBrIAhJJl
eFfrKlgfY8iaPZcE4DamM+vOgSjcI86+onJSuGJYYgm/HpzY98JqGuUQO1LhRQsaXAHufBvglz8M
QKpyX6BDCZyxNrYs9uLu2C/Q3YTecyDS7q5SAus9V+1WfKp1izYouVxIpkBOyfuYNtub46XIoj5d
K49xxZ/629O+GBzNyMj+608L7vFMng+3M1qn4Z43JcZ2oIGz6OpYEsx7v/P2r4/K++t4oAs1MRlZ
qjEYUdv9IwMZyvt68JkVL1qI9qIYkIe7/RI+q7WNCsetbTtzpMVWMy67rTPJBnKofeMcBXT1mFwc
71hA9nalXNRsaB4OvYeyG011VeGEuEvW4HxDR51JygOnJxxRDTewm2BC1kxwCoPs+KvxWPN4ASI0
8A/DEWMMtGLuZWlTXsyQad+VqpTZ/NhUAm62Zt7/uiJnh/hPoHzRozQ9LNJmiWwbJX4voybitv1O
HG+eZzCWS7irvyrmXyPyo5KrybnzhRrRyAZdLGVcgGdvg1W0ZAQcSYp/zjPTFOloHVDgzvQGPmgv
9xInQTptvOYPxFXY+xI58YIphpR7ge9hp52rZLqWHHiyy6oHojf7O1485whA7hZfgFsMQqUU9l1Z
HNxpSmwqzFAri5FwknTvY/GbLNfvF48SoVN1o0cp9N7l7VAjDD/Kp8vyON6l9mJv4LF0wZ3MC5K7
3QZGHJaN7ffspCYsryD7LsV3UfICY5brcPt+DmrR61nEsyO77b/lqlmc9B7K0LUng7sjR1vfqEpB
01SpOTlCwKvZZGIOpQ/I3ibIO5HHFD+th+aoRpQGEdV9whXQs807rVgu6SqNALENHIZQAfftyJIt
E6VrmlVOxYdFicPs2JH5Ot4bmaYt/KMYinYNUSeeR0oWMMc7Gyi6kfvX09/SGNFSu1uofKT0s6PU
AxaUQfWtVmZPJkMgNb9DKcGktS+mbSYtbHKxTiw06sZqdvoF55+IT5cFrOWJbfr3k4gJ41SxufFe
uj2VZuwmHuR5GIGDGqLqzHvTU+R0AfosZxCWVmfkDPK5Vg34Q8cL4RpUWRZFiZyIoBM6JOhwbjDm
OStBnVkBpkEY0pBtUF7TYK0W9tr1UEjSmiCfL9+mq/YZNcMtKMLMU4LAtynGSkyF9S6dxHM8Hwoa
QSTzP69lZJX6xV6K1y0s1Oz7Eq4EW5h5Q3BGsGpIS07vUm/HxxjdO0+jpNrXFzbNM1aHojDiafD0
/npuhUtLSlIeFJxZehFQAadhUim3iOBwWkrxbhomjBaWbI9cGwtBNMGtzItHRIHD0sma2Qr3B1oL
vz5AXKT7xDD7/XtsGatafRn8MGgYyZHFjYxFpO8pfGDD8mdx+Fty+vna9YpMdVYNI0CYEJTn32gf
iDxhRBzJsbdYBL29xqSUMvB7cLP+5s1aEs2JzjhfoFCQlYg53io9okT9+7LFNUI+QgRhHwHWBdSv
5TBFDUR4xRyngH6JxDI/CFDA64VGVFGdp/vZYozZshPwL5KODtqxCz3/FWMk563tuiZ+G10Z8lwX
yueoRAvKiK29rgVxp1gAZ63nljpSEh2RT0TeyshIULHHLooLbhJYodqt8SDOZfKzPMmowveB5nEN
BlgSudY0NvP1XmjygDfP2NJi1gh0tDudpuuOyLfdTf3n0CxzsoDqf8JdZKTJHmBPakogn5T/KIfv
KRnaqshdsqJ+abZNWRoXrL51q2Av+woMD4paQU3PeO71EUwVC1i+qPYFyH1P72SXpMdYXIxio7BT
lJ3nw581rbeaHYtqJhl6XDGjP04qWgXf0hnrkJgCdIpGiJSPcnWoDPx9Ck06XuEpI0otEj8em0yN
ti50HR9OibTSwY4KvVgTPmtPprqEwWGOxKBvtN4p21ZXIPyYW/aQqqQMfkqA7T4unH/UcF6C8LXH
mY+GZLA7qCoZaE0L5nmZL+MrKluNucDJVWFJUGUG8/OtWmz5tEzMusMy8wBqrQ+XNcONNwJIZ2B5
Ilr2R97u+H6yuVzNcxfj+gOcJyebpMheAViUbl3QBPPaVFo/8vSLyq5Iru5Th0LwvDJXMvkhviaI
qB3x7rzFtHncoZ1Nx5fbSoEbDZ/X4L+InxBfZv7jEas6TZEcWnY3vou3ZcbZJS8pgVaE3YxKm3rw
fDJ37/zMPHAECpMQd0GktCfHTUJL24edWze89mnPax6eqXxhA/kQrhYrkfhXpp/Um0fAkOc0G4NP
tNZ6A0lysErXIJxL6KI0j7URAoh1tqjpPvAZbKRjGyjji44IO85MwBUkAzoOItHfrPuSKB+eIFCg
dLBc2K/iIr9YljatIZyWoXnz0cliTcZTBZ35XdhPlkHJ57zdUhRpCYU7JwUV5xC0zhtyhHGJ9W0x
7jT+/NtpnZQG/cabVyf5V7nonJO4aclypAg84hXMmVlYkJIbBXnOBiWG7yJpAlX+D7PUqU/HrFuE
gmvf8VCcA5s3W4Xmu+wRKhj031ELv4P4HVH65gDwFDRuV2VVYJEpLN+yiPTwgeIhYqQCBhh15wUL
92c5DmDTkT+/tkL/SZFpCiW+nQXPpOg/o0DRYUTc4htsvFo5mTnOFPENMz+poNw+EpkHPHviQ0xT
Y7mb9E9jZAthAkjtx/uGd66loIukLWvRyWIfkxCPjUPywew7hov0NxbWJaTEquKfmZUUduEl9Mr1
pZXjFJY4X8LblkOHU6soorbm/11/6LZYaBSVqldJLVSEpLKJ6xNFEqesn3Zpbbl8+HoNLEQA60Ur
Uaa5HfNBMZaCkFvMcgYZplqBLCTKLleRyci6xysqKxn6MpoXL+P6ZsbG8ufhQpHI7i9wumFp8Gzq
Dy7e5lj8ctWZ0ljkjnmV8kAZHM2u/wQGbcDdxDBZKOclKE3SuobaNb5CdNBVPqWr1NKN9mJBaHZg
OTxLv5LlERfAGc4DL3+k26rA3OUzSwVHCRJ/Dmfos/DidZUnBeO+adf0R0stPU25SXg1M1ei3r5B
yrcLpUDcpgVT3f+DuNFaLk2WqEJfcA6Sxwh+40HqK90/IhresKoNPmaoVZQ64Q/wiTD2iSsqtXem
WjnNFhExmfhb+Zq+uZoEtGp+wyz8PcRs6rFKUsOOWVaiRAENNzkIW+3I9YABzqIhmuX+rMxl3+oz
TZa3poKYjBs0tC4TlE359YHp2eFunCQUd/BwG6i9XTffqMEtCGIlpwnAuBKf3L349+IImdpZtdxI
AC1qcsOVNUYWj899nIwnA/90Kcvit2nhrFJ1A9WekbygI5iczeUbKd0P7EVnmfDSp0PwjtbYnfMt
AB4UkbbuAhvIYGtYGhBcNt8bQAHwCc+rVzUTLavtQn21TiroHxHONNidd5jDDp3PebsjOLbTDXdt
mAyelHTuEok804eo8U06eftdS38orkiR5qtdSydYra9oTgdWkFoudzYSdbch6u+rIaihKlCTPZI5
GGBIna///05CEbEGCsO/r31sQt+KaDJPlgsVnB17Du+8x8RHK4oxIphbULCa6E7hoAK2ChLf5ePm
Lbtuvc5FY/BhqkZ5bXs48aj+VWwi3w/9pprQnAfoDiasiPmfByzxRZX95geok40RXR75QmPpeXpb
DW9kule+xeML8TO7VcnX0GdWYVHwvLwH2NmwQJ8WYrh1gJL3W+C0Fn8EAb/vmhQRrUa7Mh4wNbHc
766ZIpA6psHiE0P9Rn4V9ZKnbszeBvmhOkCz32CrMq18qOFDRY/kxYLzvJMeXjVJOvk8PY+ymNxR
3+5HnP21oPlmq1JulpG4rugrf6IuZQp5plCsm6VH2oV5Wi1VYImXk0YfNQu7HIftNizuC17dYHvQ
vMY42ZmWoxwSrG2oiaD+xpOdEUJoKUNBznKwTKuV68Xs37I64Ntaxb6NDr5owbjEzD3Pyu+0LUOM
ibgkftjY4navzco9lTG6NOjZE9PONcyI/aQ9/nrNTuUOO70Bx8BH0lOTJRDx5Z8PD7y2eQExPFbt
HUClamr++nwOfoOPb/ouMhxYZlBbHjnk3Kh1900NT5d+r+OuoPcwR6clkpXMcJMFDBS/tXeGulnB
RONTFQG+MwkhwEZdkVdp4CdrdSBCYU4fRhPiSUEagZl8jc1+Hc7KG6sd3pdZ7NOV1+l4K7xjNcIr
6fH82PVqmtDTgdaA21CNZk+P27hYZAS1kU1Zg4TMWBmploG6b1nng3qYRA6wtcOw61W7063VslT6
rkwH5yTDwms+0EFLmv5KMPKCtmZbXx69WIDaOMgNYd0w0CXYoWpxw9qE9w+xcx4HfBEhhxc7Ldxr
LgJc1/FTlaTZSX/+py5+ihYfif9zKaW0/0R+S9Pp2ejgWiDZLMs9rfTm1leeTHQotZargjgNAkyR
zE+f6i4lkABJ2NMgQZwb4rOzpf8dhGEaQaUeUWMSKmfHzlQ8SGH4kgQux0+Amhzh+5VAy+QSNsi7
CJztWj/96J9zJmFScerLWnj6YQquuqzGBzAAIOHjxWc7oMWwwcYJM91e+hsmc1xU1EV+o4QedRj4
Coy4Vp4Ef5zmqx7wepV0ySrABOlm4jP2gSFdPGUrozoscoEezJ6Nv+Cg1+f70BJUfboDRRDW827J
ETeLE9xZqVUvhmWNqK3tIcebgGcz2DxHkIKCeJyocAz5b97zRh9w2ulYWJcW2MKHG+uVxhWQ5exC
CujnMW+uvsnbvwKC5OQpDV6KjW4b6vSWr7loSL/Yvze6jZMuQl2S0I8V3R5Pl/9q1khAh3hUAWR7
+Mhztu4gyHjNO0LYFEHtYIMP+U+3qQMTtmACMa5HYfhbIQtAC/ZZJArgbHNHzPySyAtgDS83QZPq
fOen7ZQH1ErP77DZ2G2Hu9j4t3cquECuv+0Synn7UJYjoMJilZeyiIcp9Uo4mHZ6MoN9hhzDlsTh
PLKHLfrWoSVvK4dAofIxTE3dMmv2xvjlJuIuX7cFkqqp9ptNnj7Gkq82bMyePkTMw2JDlJPmJ0N+
mF8nDDDMsZoI2ieaN/9Xvwq+oQ0bpSYtV+pakF5VlhY901/D/6ykGCuMtmQqxioEhGO31ukhZuuP
C9eFpN/WB8atQj60mGpVo4sEWOjiKwjgzKi6ZnQ1jZOiOvVylTmcvIJBAe9zZBFAnlpOfQ6iKPHe
2vIISg5CZ8s3dEhIqt1NI4fL0HyatDPdqi4k6hOGvnfH752ar8rRzI58+k5DrNKekaCEWFvifXGq
uZjxa9Ih/rhuSG6+YuhzDpsh4Gmwgalhl+K6HxBTTDnL6/yE8wXMgo4WYOyLZLOOeywJ7oqpHlEw
iP/32nvS7fZk+jc+jYIbplW5/sUFo0Kj0ESDDegw4LEATAonCAIaCMsuf8RKxRaxbaaHZw/FlMlH
5lJ8bv+lK/iPTb0TRLqSRVaOB0bJXXW08SpLwwGlnpEYPAJ1FQRRS8qUq5eThpciRHng/EVS13W8
eAeqSEC2jGyUnxh9JbXTMZRixVFKKvZiEZC05++tr6XOvQGxblD2n6TnF4r3WuYaPPX4wckH5vws
Np5WNTcuKjobp3jKMDqOUjPw8y21HsYueRfG8sUrIGmShkh9IQ0kP+gLAVFUwCKZk4kXLHZff7nc
Fy2Wq8Sz66Kp9q+X+QwE63/xnsgWIe0YTVWuFZoZoJQIzUr81YpBpatxX4PJhZCt1Y0TRcpzYynA
oM2AXaJvOBjii6va0qIqcm1U/gHzywGrS1UrS7YJ0LaB/dyjwNHyapYMZFXeIPJ8WR9PQ8umalD4
+zFkAfXXN5epAB3nIHvf6dbszbAI5SSxxkyRvYrxxwNWP/q3f1T9hOHwIt4Fs075NFTuqzuCszWX
o/0YbSviJM0d85iNckQUQiDvfDLEx6ctfg7jD5jKPePJialmyqCLtzt4/VMjBbiMiDcAJ+ouXAEX
PkksI7BH3nRRyVVBbzTL+jLQahupMBIjkBJEkCDJnaK9aqmcWz2jVEUGgcPOhI7DUbkZ3cEDRJ4B
Nh7iKPn0PXmoz30WNe95IB+S+hsFp7Pif5vD+abnbuhyBiUNY8cJqzsgHZWYPOyuQK4zB5RwP0f3
MY+BIL1Ja9xFPmqrx/YCiZho0L7ff+XqoYejhM/IeCNOCWOkUogiRBvElKy29Js1T5Drre9urYQ0
4swfyV6Am1+qyVotU0MT/kQq7F29WMgZyShwQG4tbFv5La0HIkX7C+aXnehq0saI+GZXJQp0xNz1
Xy24JZbqYz8ckNX8eXgBiBzf5YX44vSODt9dsCXMtAHLfHSTZvYJcjQWdRg7onXBcVCPituk15L7
xeZfVXioUJtakuhqiIzGLIn2a0wb9T2diHp/rKnf4ITUbZzkgdhvs1TGjfPHNqULgrRQfRXQpVd0
otFT9rmiGU9PVA6E27AZCzWdMdNZCNer8kimW/UDXZ1JLWkIfqXCT2F2gUsvIcskVtbsZgGLMyku
ElF5vHb0xtc3hlw2YRIo8EPLoFiicXBf8Lt2E9axy4uYJt/IRpHlZjsgnjUk6uJcx7pT7U2Wy5Vm
YSOzHyhg7ZVv7IaDuVWpzHz0HbRHtbqzfT6e8oesKwwG8NZbX/QxKxhWGKVfBNxIsFafst/JIL+x
RG0xqlrfKZrvL8OzPnBdGA/CTTifUa5MvhbK6aA+LmKucVy1kDY5wTxT1tNr49tEtHTTjW9Ysbn+
8NH+ufoiBEALCyqiQ9eiBv8eHVL0LxHUyu23MOTjcIo0Uo5h+kOoT8UMdwNhsVimJrdrfe/EdoLw
awlbtdR++/0QS8Ph1wPZrvJbPFZkpLGOzhiQ5sacg2PVKzowLmdaEpMWID0zC7yzd+YCXudupXAy
+CZlPsKfZhJCOKaUyxYSpJjaPu8zaNUu4ODXRZkrFkxKbl25jSsb2kHZvajZTjmdOAjKD+ZulPQj
pjEkEM1uIvHIKKntE51Ea6Cxo++a/S6yHfE+BRk/JT02aJMLxbL3tnYVDSXUnZ10H4Zk7111DgYU
OkpbsdvFRwY1DvHRn9iB4ikfm0zmHP6sKoWAkUKI3qANaStIqmQov9kQ4cnKChnnwJbdjiIOJO6Y
n8ODfcgK8ybcmvOz8H6t1/GMPLGb3byBn6gqczZNtqzPlDq970zOTFeVps8Qtn3o8Aeu8vHJJ7gv
wBpW9Y8C84nE8ScwXjdLuz0pMfDOeXtQt3ZGeidJgRFBlQcJD0YghRfFBlgwGnweuMnKB+Q9M0Y6
4R3xA0NKoP4rl0WPhIPrlsESGs5foDMrAsprOHwDEFmj7C5wjp8pFn6M1w29m6Ncm+ZzQgnSrFtq
Avm4MiznA1VFx6PY2eUJt/ENZzOHHB8Vy8XTnX7jJZRyEc7c97BSUhMwBAf2N4SwFXZTzCPfsO/c
2OEUnptJBFso56EGOQwdtaT0sG1MqKc8fUNX8ggUsl7DWTCAeQIjHuvIc8rp/ftTXM38vXhEpRxE
91cdUaq9f4ye8OphUeK2KhQ85eubIImvShJdKX45BLHHd9rP7NWcD5vMH/f7BB1GM10NWn9Tqt1K
SO2N3e3XxSiS3GcPzQHVbyQl/S9hJjXVWXt8n459bUXu27qP9/jTiNQkE8OsEqoD2dobBZwCymI6
2CztlVDI1wSIHSIkMcQDez/K/Ur53PYbDa/U5lx1vbmYHVbxpkUStw1mKqXKXxesfV6mPVzXaguO
sK/YBCXpOaAp84jbHmIdt49ttAOyjHkDrfgksLfdmy7hwI3lFZZ8R5KUn+g854E5YhldZw0Olweh
rhZyl/Plojsbu/DIZ3sl39tOmugUt91Y1u5P3hL58lKQsEpbpDU8mU9Etc8knH32eic684iLfJCU
8e/ahtJP0VgJasdqkxnOhDG/mV4y7tYHvamJI8kQo0zBraOkLVKiOBMP2wkzAF5vYYxmxzP9jkXC
UDxDSl4/q6arRq2pM+26ssfi6etI9NalBP7jhdR3Q/iX3KgkjZ/00YOMGJlbko+5sOv8DRMEIWWT
qbzC78UtbW6qpjD3n4/QHbk2jtzKroyVgKzNQcOzkfkyJKedbSJsCYxsukI9dyPyd+QLGVxYUGYY
l4/5EUmZHPOxTtYwG7eq+GsuGNqeVLYvfBcbwCyGHudoj8hUiPgfaOL7wiBbwOl1ZX7Bfl7IUgfW
9zts+jDoYmO/ZguIF4LcwF/dVM0xeoCuXiyt18WXnd6b1WtfcC3IUPNOkmIJTP98APtEuQ/opR81
RoiTgmG+YCXf6E2rVN/I82JxCGys/bg89ZHzZpeVe7jPrINW0+/UsP3XfvVgzPggIo/u7/tNCrtA
CfWbP9pB+5lfLrjtU7Y7yGttaoJmIBd+3No46PEeB+6Aivj70+8PbczYhiyvMqDprIewYF4Y6ckR
v6q8XqdE/XM4ZHK6veBACnvWNa1Raf86zBU6pKMm/U4et/vndAZBqk5vyrF/OTaTzNkHup1YaeCO
BKPdtFcK638BALuS+xceAQMrY4Pk+scUpKDL6w0kp8v3DLwYHRxMnWuvgDF+6dyV3pNjy/4WBMsM
KGuXygriezspgVOu2kjufO88xVEzw9w8frKZtqAHHpvMWx+Df9IPqN5hBQscQL9w+JvorRIlHNdA
FEUWkCLg4cuyIIgFZjs9l30+bjkWxbZ/dPNVKYH2OX3f6MxgaQX1L5+kFi7El0Nlg3ZqpFRAdLRe
7vYBauIaqjv5rqbZCNTwmR+Jz7jB+z2VncVAH5HN7DKsO3lEQ1KmXL3VwirE8AL4gbSzxnP2o0+V
B3hJoq1kcvvnglDpW8PlYxq8y3wTtmrEySIaebanhh/7EvU46QOvBxpEefZHKVzPZVwIjAMflUcK
8TPDlQNQ9p57ew3rUwkstPYZRvFRiSkaChwC9BH2hBiqDtcLVMQpApzKhKeBMzrAbk8Se0p+lMnj
3Pt3Rh20oxwZFAaQX8y4fZ+beVcclXMkBqFc4V3rQ8lYugCH9GRbIBKheHv4/PhdrTzUmDf4/1nX
QTPUI9DNLbTgSHjxFYpG20+VgBBh97NJ01lIzwUTtOLGYde+jJBXCZBm0F+kHFhj33DJ/gOFCEQv
1w+XvxusN6kH1Vm0VS9aR1W8VZTlithUQhWXF4Blb7slmHT/DqSwnHm6xoxoG5MhbpYk4St218zB
o/yZ3tqyl6C7iO41wuDmcWTnxswpZHALhB4fmgtgwo24WAG6YhNQlxCDt0Gm3pXa6hMtB0rDRIF+
lqYdhAwvCU5DbSe2ckIv59DIKQWnqmUujoAOWd8FTC0Rnl0JxByRvmMMXsHAqoz7I7SJ+7VPhwXE
gMgWl2W2dFneus9vyrSs9iThkab8+1ygJPHnZRvNRHlF9EIOPua/0XvJGl18VUqg5nyWJU8qliLK
AAtE5cUN6knVV+8F1NiYnJjTqR1x8Ggfdg9hpn4JQFHnWCG++x/atf4/KivOHWVk2X9fb6WJ1xKQ
H2j7hWhtDgz55CAkaXmyRCch4EtL4hU5NIueV0+OaWNUK0DrJWrlhZlqdNavqnwMZcjIBlivvKjk
cbfV6TiWBNfso02k9KZN5rb98Cbwuz3atTwGE6MeQBsDE4v//OJRAhmu9pQFUpW+M/pCA1xQNEj1
YAFQtMIEj//WNAj8D70u6N+ZGayWFvU8SeQZLHr0KpEkgEr9Oivrb27RKfl2KN2ehdhW/m8596sA
7TRi2UJjz7FTG5zCW0e78d4HwvsWkk1w9UVetWffk7WpbJoN5Kx3ybBgmWws5aubkQfqqJmf+UID
lNAPESNv5TbIZ1nkSdjGYiJ1/F7hGq06kUdn6lBW6lubQKpM68bZpOH1LSzOz7713BS3kih4N/ub
+jCpFj+IHitppmm+bM4837XBtR2StB6KFQErYOkQ+o3UOeSuNxdM17kmncTo98uA3/I+bvuD1cKX
2T8GfvaSMKbXfgzO9WwTnvMl9p0kQUtNcR2da6X9XcACNBSlcBekr1w5h16w4FCX2ifQSDSrxFEK
zSOF/04vQxMJkH4UxCEn14nv9m+JQ12sQF3vizCQFTjaZfKVmFHg0s1ux0kPwyBK63+0WjGxBlnx
aciKh8zI71kNfthblQ6HQCKKy861Ky+xd6Ml8vEPtmQKpn0EkMae64EmQg7QOdHb0So09MmUzNNI
nmhd/GalwENYJg82VfCGvOd+8Wd2YGvJyO/BGZNZkCp8ssKdiznxZt2dIY51wHSCL4nIhZjR/sim
rqZdEQNhiwzmnXbJdmvYcgtH7cTB51Jsi96CCdPzGjasx0jastX7z2wEhtdvqFitCT9r0F5FYe+N
Rjp7n9WgLoPmjiJJ3eRUr4tBGxIqiramnC+xfeQ5xmAq/UHilLYRNSj7MBgeefuY3dqrHHwrr12M
rcVbv1vzeG/dyIPyWBseufz+rLYCLfbZ1Al2sxMndteDpE0SbmF/F6g/UMF2u441ZHCB2v92484f
lpvdcj/7ZA98M+FTAKe3yH4xSsABkJ59tDFIo28A/OdTKFbIh7w+Z8jaIwnP0Ofiy36glqHOAOxH
xRpq6h2mouwOvJrDi1N7CCWSIsZdFqjxnPTONaf72Xf6Ek4w7c5AGd+iQCV7Hq23r7OmVKwnFX52
K3OYRCcCJlrtHUM3X4lxs8Em7EMOKJPjuVwOe20sx1BEMKJcPtzc0VKSO6XrKU48jp/5nqO0UELH
rkRf3sc1HKsU20/rN8hFERDEAW/x6IG/H4Kbjto4Yo2DkT6lSAnXF7yajkAomvabVX0rxCey2PE6
tcNZ1EDsVAagalfAniTk+9Ma3I/n6zWYcHN0rFBhl4tOds/eUsk0vCIeK+VxKSFBZUveM/qwedtr
YcIAPvLERpKSVhsRIGUmkGxP5+Ij3tj8sEhyWw8Fsg6ioFHI3sqpOwwl5vo7pkFu7pOPAGH7/xIX
WvopF00sVRkLymUarqu9pcv+dTijMZO0uaRO+S3KjyqBBjiZQ4XfNXXPm+6icDDiXH+1le4mamNh
nigX9c/+AHP8H22qmdYLai7bCitcgn0MQLDbkxYPAPC9q18yC1gjVldvUPlt1pwJL/Lnw5S5A8Cy
nwsbd/PnVvkOJYEyDjRDisGsfCdX5BLBDF90s7yvH+DBd8VR+73HawStoNHbu7gM0MhhQ/jf+pkQ
BOGfQyYXPGLSxxlolwMtQasipiADHGhO4CLEifPmfuMCAiAZ3hrNP3v38u0wgE8NnzAyJ8NgLSGj
g+lDvHn9QOE3+M1Ky59gAJGFCYBz3CCCHg5RJwhaW8Ue++83zGyFbJtBDRWYATJgnK1kPymYf2fO
k6CiEOh1GxecCNdqQaDYC5RCMuO6S3ISUrCl3XCFeOleL3gQE1IVZICKP3VpPkZfaoRhk06/s78h
mb1VWSEw9fnHxryOOWAelXJeQ4ggQu4Om4lxxH5gLyAddWw1O8zV3CUKf05H1LCvner0MlZTcaim
q1MCUgWA5dZWQGdY4lrYxXmvV0L5rSnJVsO9KLmFzoT8OhWuHp/maflDXqhPwwLKwaTkCC/0SrqR
8sZcywaqMW7lxApp7LtAAxAegIqyn5QAUBRPGu0yoXFqWqK71RaiIm7MA+MUpVGup3ivdGQKVDDj
TSc6AwWT0Nu0LuJg3Qj7DLbWtUW1nxFZKTaJHvNr0uU+pUkpIXEoqxSxycN06cOhf7OigRAvPcXo
G08BWE5T+YngPMXiySQ741HH4o6bHsFJOyE5SzZjwB2rHZemljMqGiNA5TNufCdxcX2n/Qisy35w
opSur3mlho9uYqdQQNbQY0CcL0uQxKZArOFftEgXWx/3AgMcqiomP+vRqquEwtDc86aeHMsMCmTi
GVuBDFRs9+ozzhr77PZkXYd7jqsrDdBzzFk9lKTkGAS7A+71cOdqQJiGlNmvEo2JESbhoKfajEvs
PP41Vf7dJI2LhB7O/7eciB8Rm3SdJt04roB+dLStWXWWUCnO/WhhZ9NDN4cQ1UlXGjC3C/q1LSkv
NTmRntydI1X9bKMbWaxVCIqVsK6Zus7i2NjbC20YIjeyvvgKs/GlC36HDIHBC0TpzAbhn7N9Vtac
/IHamEzIuOW2h+H/jFZOQfKGw/VM9ztcYJEivuwOLM0IktZ7F4CT1w2Y/w0ggqpvltir3ATOCPyw
3qoGHdA/CQifHxJRYGB1jsQmeYN7I68Ors0E4UT2tlD0oCD2zlXpr37Uj5tHK5d8dIS0PUNc/QSJ
gDUC4Fkw0W2+AZ6ZKqXBbGSKgQrDsayCnmezEHsDJaK9ZOFjYiI+uM1+Kjni8uQr2TPDwXtZwtRd
Eties+YMYRhq5nMQSey2z4N3qklID/lHgkiZbtZebgrq3C1RXQFP6224uPB4OVu+umf9WTJQhfMJ
95SQX1M5R3OT1fP2M5G0xITUI3sCZBc3hpYVIzxQiUCUzHYaD1rnCUJOJfE2c62t7jbEmkHxorqp
fLjOrUxDzcydgnie3B26OGzxD4Tg0t2mgXM6n5kDZ6NRPz02bPlg3awxHf2av0BsJjRV9Unj+eEm
+pGO7jvpwK+eOALCdsdM8nI4RZi+NUaunLv/zkU8nmfuh0L/KZjrv+O8SDiJZk05RlHFpOxf1uyZ
IuP15kITK4YxcCOGvuiuUL0WVdRKx6K0OsZI9I8pHloWjBcTFIT2Iux4wK2OyxeUobzZucpTInrz
SPsf8/lDbklGRBOUTKfhRJCs3JGOtlJpbHMJb5Kc16vUO7PNpKfEugAZg2naqPGLlSWawGxoOvDu
CE0h6K/rjygnyq3gLzS467SKQB+ij3X0OPlIbzCjpUA++tQPXvTQr5gTMRcly73tnJne49OlAOSc
4umGE1XsyZ7fXuzFtfNltwhW+Dbb1Wql2/QzPGadK81A+Uj1s5Fh4kLzDQfR5ZSHGxVNB/NkNxMG
nQqKnWfXKwpQzugXcS+6mzTLJ8ynk32Qzak9O4pbkmhfAsZrxu+aRNuzRHEdjUXNGQJUrQbgLs3U
jskN800C1qsUfSaKv/vPW+OHw4E1c4T2rfygjYNv8TTlPt/tzMfeWL8K/2MIdII0Ib/a7DPGXhmG
gV5AGKNrx//yZvwmmIHhFqzu7AMhr8PZOC8/h3zzQYgdzSzlUgg4rNt6bEOx6LbRNzL5ixbzeNZW
nQ7VRTxs0ANjCiQ6WBtSeK32rEkfMO9xgeUYmCJ/ky+wA7tRn7W4FlZfbCNDGE3v3TBxs+dpqSGa
Q5UGoz1QLqOwSuYscU4wKTAUAalVmrCGXZEY3ecrCyd60sfXSi3i44h9KPz4V59IRHu514fW9r5s
ZgjFeiKIPQ+ZPuWonCcrgTP2o6umvjRYK4lmOHVIt4INCgxn19fjq6GshtGLVEHWvfXiLrUUjhPI
z/Y/+tDmsNy5QNtDMG3RIzNoUMpsEmbzcYnHtrWfO2MmLCV3NcoPlTVqmV/3a1D8fzh+5jPvdIOa
sDNxrwOCJQhbxVl8qDKvotoFvPkI+olWZ+JRnwIyDcraN7YRMIfNLyyRFMqf0JS+TjEYs+Tl7Xag
iEKHUbENI/d7Q0UlTpn6xTJfarroN9EICqnb/e6RMiFVXqe1/Xl6uZ5jBr2eRuydU376/Fk5lWl4
KAwjZdmNawYVCMaZE+yRDF/ZA8gqiieOyHcmncyZytQtRp8phP35JbDQoRuCuwL3/owBWlRjK6qE
WKLM9G5SL6wRxnSQC7dHppEs/adZgj3ivIjoAEhZzD3RnH9fTOssUjvs1sACuMXSUnG+RAd7Eovg
pxfZMteMlRIoOciz33dr1tecFndBkiaSactlaFiHYcLDcIlypkL2FGfYFA1TO2ypwAsjVI60Q4GM
zCtEWiNbGyiCEOrbtw4ach6BOy7sCyjBtqUJyRfz3JyXUJIo+ml3uT0zMC15bPziYDY/DxrpvIZc
j6W7VD5Ru5J7q+G4e3Y189ye9D697YfDPDszDaGrgCCYAga/e9+cUcq1hCIHMRCjVg2B6lx5IM17
yEENomxXpF9GP3T4QGt/O7n4nS2cjQ3NqVo1pazh23fQaqQuxwhsodMsUpjAFrFbRkmC5fNJ1N6P
2gGIs4X2C83DsSevHMe5jq7iYaPzcBtXB1EyQNsZzJbmRKkhGnLQtkmqXKxcZBKbkDjzhc3JfmaK
d4qUAWd52uBNAedBmyU4AgQucYBTV/97JXen6gUnTZmf6FCUa2Epmo/pefs5xxP0QC7KYjdfuV2Y
FJg7asWhm+vciHyTskIHVqMpzmONWR6yLPhxgsGvBFamwXCBWd1MZVzQqTIfKnKeo1irp5utedpb
SJh6lLmI438Uqar5/Ogq/DgzTnVubB5157jTZ+taKPWizAS5Fs9+1Qt7q1oGmDaBfBU4UQXyY4dH
igYwSXoZoehs9ebBpZ3Jb00dxwpWSxrxKO9n+bax1lCH6EH0Kt7IYYUfRz1vMtezdl9CNeBng4uu
SvO1cwUSNH+MzXt6Lc+eLanxiaxhjIAPQcuBI9NmWkD+dkhrt0xSC8NU/DP6c57LlL2F4ccdhmC9
sznUkfCGZzcjCHCAU944CXaj1aKtXFJwqAw2tT0yP5S2x/JeOnG7jIgZ8rOhLpg/FpyeO2QMgMdk
5hRsNWU4/6Az8ZMGRgQtWyMXym8G1E24f5zjRqQKLIL9Uo9e5Mn5kOx5NRz6DBnTGB3NXWq5GMQf
2NJqwv9EuWqpqgwtn7qalVYb7YDutdQYK3O9XaxbMx5GLmB6P4N1kscDue+P64dYaY9CvbzJ7TXy
273lRg8xNziO5dvq0o7rT0aKEjus4tYsviYm69QXqwvnJi9J9vt92I2YeGET3yQ9/Nhv1NtuU4ZW
r9zDXtZAbRx2OaAegDxolBXQMDwlfAJSJswkmFoahv1owa89Ti1U1H4LU3ly5CmgJlVDd4P4fPB5
+jknDmTLfHDdxtasaiwHfRG8JZkyz0oW54zei4gBeVm0U0uRcDtpIiYivcfQTjhER5oOnow4fa2k
PDlvPSF7My8BZHWw337FwzJS003tj66PleuByMXHCC83MyGmvyPXPYnI1tvvfdvXTRFOXwoXAZyC
Q+V5RUjagYT80D+6gGief7w1qEM0F64EDNVfeIuZxMoEG0gYsd0Ayy9Wk8TeZUWEep/toJdmq1Pl
oqj4uZhSoLkFk+ImTt+8ftca1xYfQxpasaI5nb59F/fvC+P4DPKjzh2lAKn4LUqBg49PqF9v7Jog
fDB1c6UbpOGk55eSw6eESX0zC+4s/9orZJ2K5dULpz2WLWVm17p0x5fm0/Mc73peX8rpJFyoR/6P
kiffafpu/94fUedG5s0dUUqPduKRZoVyG0VdeHoAmQ1Dm7sLqQDhkSXjCgCbLlO6r03WhorF+rlB
pyL6pIXnu6wHqviLBx7SpOVZFiNa98DR0GWnkkft+9FPZi/RNSTdahZ7YBe8MzB94mlIJQm8pwkS
Oi7jUvk5GHAp39rksASly153Tr7HR2mWVfHbePyvQNGfxr6NhimHdlN5IxvgJHSoNj43KwAcNhnY
tt/PqCh6dK+ysIAJ3jHNNOnOhVKk/iuEf68XSzGhkCN3tx+4jBjC4A9Y+Wbkb7sexDO6oa0yYs0B
cR+wyLrGeRS0It7cSQAEohL9gIPDS/mXO7DjJpfmBZpGKL4kp1iMx+Dmd/SjKNJUgocguTaNATg6
gnu1SGXYLo5MmDC2fXL9ZmHN748kuCcPRdTc/esoOG1Vxln4W0UAh6eVP7B9lvDMUx/MvUxQ7zKY
LZJfE28UuEYs9aR2PE9NiLecxYjnHRaa7Oi5bKWPECymnv5fXTbzAQSd8RENk2T80CX2SmVEeOIk
SINDWy0/xV9Rrno+ox++A64nAKIqJ6YIhQLtAoqpYsDh83WPBHkbED9btWwQ1qr/cgCSj9gVLpZY
3BTgf4lwz73C6ARngObKzEmmhKFq4pZBeKrD4abvxgry9vtTSg+noAQ7CmkI/j6KmHZXo0wNzoBE
O/Y7oifun+Bpr4WnzfWEGw0cU4IY6DBgoyToaImWQsOAULVTuvb1C2djWBmsSwDxA/Kqkgb/Nw3k
j9Scv/R8aeLXb5mhzfRWT4bSyaWNd6etZlwfziI/55Twi7xNlEYZJrOHqPCaS3BCbFRAFdLJASI0
rTAqEAVK1ZrMWiCO7dtwEnReotieu3jg4OMgBSRuO72+z2UxFTjB9V8VL+arszTQ+/i5adstFbbG
72hjB5ab7tK95F4/IJLq5veYf9lHJ4n5OdM1aKI3MmoWNh4WCn1+t83OwS8++bJS/skezEJ4bnIh
jkgBR5WlcO/I0c/NaRYefeu00N2oZAzBZKeGuEnPxsKA0Kf2rHXoim0m+yFkNP9KvYfFZSI68r/H
un62X82CIoIZtn7qo5r9UcGpyEpHHaMQu+sYyFKIVMyYVibT3dvFBwlXv+SU5AEXcWRICU59Zmfs
3dTLNRwz0m9b3ZmbP7KTAaz6VDxLjJ/H67N/Eclhlfi9o4BMuZVOOM3Fwfnfbz+dg+i/HpmrTLZK
iTiOGfyA4+ztqN7k3s/fQjEnZO1xfOtwSnUr3nVKrvJVrJfyXYr8RK1Eq6ldr/1StTYHv1kNJxu1
XSncz55EfZ1qHZoYJxJcg0JiXPOhx74K70MQvggVaCHQ0WbaA8OZGXKFIkPQQTYlU6X/FCig7yzY
3Vb0CtZJsVavtADpFi908w2jRO8fonl24ms2+4EARhkEmGOUEg7XDdHHHLMiSrxzWKqVQNeeNLRN
8N3jxPfLqlgXtE3FLNcc8H9iD90ese9Z3LckK/pNucVPPdpY0YWGQesyaE7w5c6CGSKals5G3qt1
qa8PoT/8DoIFwB5uz8V+jDertuNVCgVFMgLIAQOFP1Od45OFRI2nCtSotK1K5iSlOAGrk2YTaFgb
dVXrOHkIpxOEPYvgVoDztxxDf9nVkwLO16rARLMFeLakXvjvryQyZ4+tMASWcpTaKkKDPndbqVWy
OTUWfJL6hv2UKjEMsnzPBPX/CyHgTd/PIhAQ6V8oF03p9lL7B7az5GA+wxLC+ION3+T+25brxy6i
ZEKXUKBVnkkEQWfBFiKHcCF4AR+wW7RWEpYqBqil1PvBRQNkv27PLPVULomV6E+Fr/j1/iv12oi4
K0DCNKY8Y6X3tivTRLCR2rfzVaT1UdFVgs+9X0v+qG2ch9BgXww1t9FZaxpMbLr3V0TT52L83xwP
FiJsBeCa8tb2U/e1BC1J3ru8jnyJq0HxIDqgdmI7USUmjMBDdbEveIXS1F1yG0v+okqcDluMTCwm
jmRrU6NXzBfLHPk+LufL7A8+u9NIoLVsWUITcMEybt21VeQp02ivzVgXmVCyTeItyjpTQBOWnGvW
38ObBCmSVA0IFr8XC/A+UYDMdiEj6mDcNF8+69Mc36xHCF0lcQ8FUIj2LBRVJwCcL/TVO0AS/mRU
J43ytlMqQX2Uzy5n/TzUp+6K2mSodNJyiJrS6R1d139upBsBo0C4zV76tRmCOWRHekY0szMMfwW0
hKdzjy2utDdzbq3qkI+AvDGtYekWdEr27/KknNDiYg6TAenOFy3vgdmvybeD8aFFowB39uOkXWjy
MiE5MGPotoFtBuIZJ3rtHr7/3IPL7pwFj1FE/pA9XsIJ0dBqCRbZQlCvjcgvyQieon6+LKrIFh8R
r+o6V1ZUm2IKcGnsItvb7ddddIb/4vmXsgodJUJgu1E6S6QSv+LMzWNwIMcmC5lhPMOmV96sPixx
VbLCA65OuHk32yD8tjCMM3/GCQVNfyUUbO7IFtOnTZJEV08NMgFR7FTobMJaUHrSJVF+H34nDIn6
egxm2/Lo+jF+evK0Cd1v/50R9oVvQObrAx4VtFVoWmvCH1Di09KV5JcIx+rxhvpooKCiffFsJ95+
tXR+DmJ1ge+bIAi+KX4oq8C8TkQPsBANksaFiQLYFYRuH35wMssk2ZlScvRZhO4lW0Pr5oan2e0b
aNW6DNdnFDfca4jGHinYt0GFWZqOWnfBy7Px+yYucOLLuSojAsHYYrYkmW/WHU211AwLQ01NsyVF
a5KhQmdxovkLKK+l8IFTCTb8Y3Swnsdu1CnqFBaez43sCPAnop54h256DmGYqO8h7Z6L8ZuP2OHp
hSKk+7BLn/N/vO7sPPl9XykvnsdCsMHVKQtvVv8rs+47BdRf/vU4mX5rviqZeET8ZbJ5c9EXnVqJ
Y+u6oEjR3O/K46+kq+Z2SdgNr78Z3JBstnOPo6QZqFztJ5/sPPeAGTxFGPBARm4Iz5HNEYBvq3y4
XZZ4OzC4RXeKAycPDk6jJ2GvTrOaaa5iJq8GnkB3rYKgac1UakR42VMsReLRb51px25VdzwyGAP4
w/CCzbvwFFU2CuANKBcRt0q4FALGvCZzowellx2h3Xbm6uaOymK4XTldtrPMt1CZEfr9109hplBZ
Qc6nXEw1hSz+sO/HG1gwatiC6Nm2/s7o7BQBpYTDXAzaBspMuZhQQ1K4bR3C2gVXSfKLZVtLFF0K
FhTWMlbwQ5uQ0GOINruz0owzo3QQzv1K+xoWJE1gmlKHxu2RXT99yzhnd2mG/Z8II3XHMxdjeVYi
k5VxU+RWnY5KdFGrTjMYePfCZvcwSKDTobacLz3pK+OXNo1z0ZovN8X6aPlvui1q8SUNvoXzwSvF
OkC8C5ol/P5VHtXVL0x8ZgvNsEYlu4h1OI0ndjS5ChE1c+bgrR6HNly6ZTmBqmwaRf6MrUFVziUI
ULacO34KwLSCUk53qZZLOHBThi9Tx7pkqwlrovAveBGILW5L6LBGj/FnUlq4iACKb3FxNm7Kht+j
xA8Y1phLXc/nmgFgZ888/2yZGCuQ5KWxW5luib9ziigXGafTrAfT586SfFsrgCE2a7+W0bwPChlV
YVsrrrmdGsO6HhonPF1qim/SY2iXdyi7F85JG3//rlcTyp3hj9DqceVGl9FfzlRxXsupu6fwZkHJ
AMFaTfnwxipcpSosJ7zyRLcFix6RBngaXZdztXkFnE4wNndI6JU4kewkB7BDpulU9KYlubmx+8Hn
vqfZMwHVCSk6qVcXEYXpOZAiVXFVfMe0pQyqI53KO+iZVPAmcOtchwudcVMCjntaWi3eNTEoBqNf
kEg79CeiGi4FxsXCmE9PAvhdSC+G8Ribhov9rWs0ENiJkidm73EGWf3F3EBtUVUpG6iHwchxUwrP
wC7Mo2Y1bGpeFDg/wBxcnMxDmIlvumVbKb/ibosGhuFZpVx5gwZYG6W+yX4n3tCdQ4PAqwe0TfwL
Ra43ys5hCzJ9v6kzyGqcAFOefSGZE5Yp0ZYQQ0pLM8GRvmU8iOICpGmssWVEmQc5GkSMvAxG0jhM
jtf9I/MwCWXOnWcjLTsumHVboPezvAmcdhx+qs/vj8EQBdKdHe93OGAYFBJSbE+vsn4v6nA3+hLt
VHz9M3GPaz8at9W/XoxxobQl26H/rLvPulWTnYokpx4yDuEbYzXxOCPsTDdES7Qhqntciba1hUHn
zRDtGtFJmO7CXq7ytRaaSB9fPug50Xi8g/p6vfn5xgPUUCYmOGzX0iaQwPcBAAXkImkfpMDC5WZZ
TC3gRr+kS2i8qS2bfHyPHw1tn2eOAl3tqAvEVjcMMu2qkReygsVVODL/vRfNM7c0s8pQx+fA/McU
fOqufYIFwSfMyztS9hBSMxd4uNpyM5GlO8CI/+ACmpy1qv8Mt+xXwFTpKBGorDLQPl/5/zlL9nDn
DEwazy5mMwnCfkAzt3WdrQd9stBl21/cU4Uw0V1YZ4N6Qo1PztC5pEHWLaA5A6BDuWNyyLaRQQ8g
6Y1mTFSJb732MHSId2y26d/KH3dNNfSTfc0Y+idSBaHmY1DnG9EpnWaqUq1qaGTXFzZ6PDVXfg4s
Ghx+OadQ+O0z3fsv91jCZveHXJkRNv5nhHOz2ppPfdkwNoxQiJ/gzjiGDydgb64OdiVzWWJo7dw7
D3ifeAudJIn3sDfuQZQagMu5tRAdDk4xuI69pCK+vCjqB/bo9BcMyg02faDjon64uLBRoBCbr0Gp
Kzx2J8Q66Pe+WaVco12h5IzPWNcpT8IQe1ua0mccHSWvLbg4cTt6IKPXNK1FIXiD0ycJwlS5XXOl
tkNujvWH/fosuCqMS9hxOPYsHGcx0tGDjxEGICFIH/sgZlMxssSAMRW50iKc9D3FzmiZfZBHwAjR
RyRaRZ13j5qb0ItNz02zHHDfUe86+6cLP9cnxYQmk1ff9HKedk8WyMv9drhZ6/0L5snoNrX0KgMs
KWAFhe1Mg4/Z5Oxc4EFhaB9O/IlDi+XLU2vydTgzFFq9hwu8icvlq2vHLV6y0veWDBL67eU3wSHa
3Z/qY3lNwTaSudHKXEpxXpG9rTwPC2DjddFEXzdQBtsrhgZD9ilIKuTv9T+rZHdvanypbv9yiaKb
Fpy53DxSTE2NhJgZ+9B3/3+eEkRp/NGSfHCoX0feY3gyBtvCLcBUnbfCNwhPdJaHZiMcQx+Q8roB
jAwANp7gDauTI+sj9TbKk4r4UT438nQtqf3kwgsafYPJ6TRPxZQ5BUZO/ZP4S+i1xKENv6VXLB9p
gcZEQM7M/BGuFCjiS2+hrhAFYV5Z50mr7F+1p+MMHiHGZ/MQB276AFApvc386w0c8Zs7/y/7r2YH
iycHBcJyA4TmmvMjQROLZJ1St4G9T5BAqMKJsO9BR+RU4De1Rn2bpMUsBCzsT0zAh8LaxRUpX2XB
qFgIxik56bgjnOqjWIR/9HkXau7/7AVnjV0sthl6SvAYRHgGtPC3NIJrkotC0R1SR0IgPW+5iEwz
8/9fu4Q7UCbNoUfgLEhj8HCzhBmPSv8Dk13OgNr1z2Du/g3p2hw54luAOuTBz5ejozU0I9rlOWiX
qGbUG4pLdKzpuUg7vvnaK6ZsDv3er3kYTx7qM+hsKxeUeCKkgGOd3Sh2mLvqgIeEb4R1txOXaIBa
LsD/0WGtmd/T9pVF3/nfG0eGMxRyz0scBLC/K4PaCaufP/G0wLRSS33fD0sQX5ZZUbk/JUgSN+0V
xz4F+Vz/ozaSKBC0cBHNwVej7t6GtRQChK+lr0aUf70GxfDMPkJvEeZW8aQKQfc8Tz4V6rWjUZ5c
Sdw2PEmaFCwupzB/s6yBaXk9ZJ3wlqdduLcpwW9hPH3yzYtUukQDAz/ul4e8NFCjd+FexJUc5gAU
hasg4lxKCaD4dGH4mKjZqZBQji6OtW1ur+mrpTzqL/4EM79yr/Tb0ajzHOFQZPwLBO13X0kR8Ugs
cguc+c4LTNl3QZDgjKyu/FeHb8k7Mfj+fI1gHb0zT8BYhPb2KzJGpRlLTbgBwgVsTcnoXGM3t19q
k/sJsBVaXzAgtknc4ezyjMxipnjWg9/UapfxGo6Kd1N+GK8J7OzgZtKqvdgkHccOOK9KTQGJz3Z2
w2uNRp0cu/EwGMkf8i8DsP+FPlzdBL3kzSIoMbpIM+3Y7MFgRe6/nnUkB47NWNV/kD0fsW7VQXtR
uFvXLXtCMtApiP15fZSzNonxjJnZUEiVbaqXh2LoJgE+HJzPdXyu/6bb5OjF9Yiw2YZvKIfNbzpb
Kp3QTro8FGdSYUl949NqCj84mAoynKhMoz6wHEk0Z3T/lLdLiMpmysAxEMHTiauSJrKj8M/qbZ9q
6ZFLDycrD9Cw5K5t9LfabBl1AiHbzd8ABvOdhBCCzgZ5ot4qEA3rH5HggzRGQSSQJ890jCjLLNCa
yv9iHXDLhMywmE/vQzNg2R+LE/lzWLeyGlQdlhO4zu2IQ3BZ/fMHGyJWf989LJSoC4qGCJ69qrjx
n988PNce3MSqZu3+yPemgdMm7AcucnXG5Mn9IkpnP3jJQH5F3Ic0Ht1AJppeMGq4e+ILt8ujZ7Os
eXqyaCpU84d9yoSFLGWek8aLtgE0vQrnaFT9o+673ejEGjt9YivUBM2loP/7ar+bbEFw6ttOoWbW
2TakSgKUU1q0ANmoGczvXkSSKRNY/AY5j899RkQiY6c9BxjPPuGvjqaLbfN42GxkFjeCbEo8gexY
bc7lBWybP0h2l0bWpq/nSZeCMw87H9UqQPoKwmmj1Zs8sHDoT6i8UXs6sSxuYNWhTCCwZNcHoCvE
MXkYsxbB29REkHViuFi5PGVFt1orTdxc5iQVRawjOOZlAX01CdtH2vCFe8XeLddUfkg7cbDVBDtp
AI6RSX4l93rvHsAhl21oZmP5jsp3janE32VWA6Ig0FH+iy3fIt39HEvlVuY94pUkNSUMS0pCVyhn
zr7NKQpPOghLo/lUiPovTYT4EQLi/ponQ/UvLNrtwrYIcddK+AeJ4oZVtp+c62RIjd0GpcjQGWdR
uOHvp8lzWsjAuAqvsMeO6StmQv8RotftAHAMOj4SXS8l+EnQ4+7XswJem7V6qDSIBjSRANtnKynd
3QxNZE32JC5gsCrmvHDEHV0zsPs3TC4128SkLYhXGr46nFA2ST0MDGipGPqvL/qqTDx8N0wcVs2N
jDQzJV8P/2ydjH2E3l+I9GmqQEPfQrIBijs79c6gh4nR9K18F775mhdkAxn9PpdfhxAeqEu8W2kq
nETm+JSemjOjset/84DAVlIGVcW7zIQgb9e32zkOsrud1BBHxseU52E76eu1t8YIE4K4XNq91Uq0
iUbepHKs5f5W32XeNk3ygxul3gEABdie+qofayjlFEVrGD9EWx5oY/ls0ArDJ3fuxbj6/h2pGNRK
60Wd8/irIt5IqC3+o8zb3YQITgyAHb+r0qs1EETZWKavtKUVzKK7bxnsUt6PD6BgWTd4fUeJnzHJ
6nvxjLSZLBVL39S7dtBJgIksV8znsu8dh0/Ypyt3q/c3WiwPBcLJ9tnKA+Hb6xm2YzV0e//Q2Y4Y
L/p3haYldT8LUT5uFdwTJRG/s/GsFS6xSF2SuOWC+Awk71pR/itySZMCv5yc1zkyUz3wNMkpsKbJ
9q/mypr1CFkms51rTj8/02M359zjJf+k5DzjC8yl+9yhVdVvpzRKFIVEkq9CXvdrm+khhRHsOJAr
zZom0HUYLlfIcJrEqNrFQ31Ot4+KJDHpa6qg5F0eBn6su5koRVjXL2b6BycW2gmYKqGm3NpLRvgr
TLiS4HcjAV5/GvJ6NBp2DlVvY9zTXkr0zuIWB/MGLl9fMIzpxv+w7MDVqMKWnQav82xP0tR13p8K
Pvx/msfAb+bfUZlaV84asVelpZcvM+Mcu8SNJddtLIvVkbKEd3gq24y2voYP2uF0lunZXEUyGFk5
UrtGZu3yeZScR0bYkWaln+Rihj+6rjjCwFlgT9zlbQmEGupQeBRCUG39tpFTLv/uY5XuDYdar7FK
ql4yDFWx1q3yNnJm+EKLSBwrYZNx0VM8eCEy/Luufe1SmAXKjYJKtIUoszRJkotJVZ0MMoM1HER9
VbCXsrL5wGy7hq5jwA3gNBlf29Qvc6ybc+h+lWx2vzszZ46VpZ6u7B9JEAv8ddx1t8v+J9sr7FJr
X1Wh5ULlelBc8rY8EzqII4ltYOZNEYXJ4SlWggvFzC+/2YviUaB9S/LVqovvlL7t82l3rjYTGzX5
W0qCaNCq8LEqrGClzypmloSlU7mN+5i6bLFJ/P2KBhRHCzIyvEfLO+mxnYVDa5BAo2tcbMEcvd57
KZEs/PFo1iKEfA/KnGdhA3YNaQlhs1mlo2Isdyd7+l55ZLfFFDQlSTzBQsu49v47PXp3fjtfbDl1
FQiSWE5RR7+rJxjC6Gx0m4oECOnGksHqZDludoonGvKXZM8zbTSj7YAQGSjQbYK2xR76/UBrUqoL
GF67CuA+UATl49M4SyvtCaWaqmn2LyDdVg2tUpFXQUJcyMvhDBne+fEKmc9WmOsfd7IKMacOQjVW
/ISfLHCC9XqG/cyYUZjfFAfsJU+sD73Gu5oB5KzmYN+4uIVs0vIFAF1/+WN2tIF2jRJfVx5Saot/
FaN3awnukwJzXlOBw55MaQ3LWeSOXy1Vhjp6RCx9FlHIUHzqrvWTEIJK8fTgJcycjmfUPKuyE3I4
iLOViBvuojSIrw2sbsAGUv8IxzFa3/KJIapioGHMV4jC0Fqshuj6qyVsYovnmWTkEtI1rer4sxPP
5H4ueqRFm2Yb9+DY3nKAm6S2qcwHuqVo4bBLQp9fSQGj0mDIYwl2tWCp05Qop4KWImSYoHiZ8A9l
tH2vty8dlywejQovwPmykxQhryXSs4HaIMMWmE5Cj+uGtAIrzdK5sxVn5nW+wT4KRv44C4G2mDcW
0yqFk/zb6hdzAKlNKw4VcLqF9lPPqCSRCwgY0NMfQ8kXDzbEp2zghQCGoLEp5jHNW12x2zK92Efx
NzngPjIGn8G1M8FsEBCpAYZ/iQPezEV8S8q1Sv5trBa0sHHCNN2crPPY8dt31tmKnw6hEDs5IUHh
pWsdMQ2sqRNiIqGC9jwxlFpASk7B6d/ajXcuP16cMXnddLS++exsUv505LQ7B0i+G3l8jO0wgZXB
7BnjUNgQyqgosWwRQkA0PA4YnZQwz6iVoyMpTCxLL9hwV88mOWzvuga67VUDh/sBZYuxI+uGu4Jo
zckejyrjazyTmP1LlP7mmoD2lguVjXNuEKNdVrz7YedK0tnreCgtoUKyvJkbXheU2Ht9AXuyVCjR
0iYTo/h3ahKm+bCqISCVbu4cXaMaYYJxuVyjXiLfEbCxBOJLSgINTGAOBe3vDnEk7jjgaKpAFfxt
A65NDrm2t7ZPEVNMyjLYjDDU52paJy8KyAwmVxCmEeialnxCbVpIrt+TkO1Hkkar7BzPFNcuBDiQ
w0O0HtG3MXOK7buAYof0bEtZIgx7cgv0cofg9Jp8ZY3FAxZYrUTZaQB60KiEJHGM+tjzpKqX3spP
4We26HKOQmEcl+vQbl99x5FLhLj7HBjg5bUMA18ycdm6AxBeqlaASHnxDzE6r3iz0Fzh2HNITQlP
ov5CQCS1vBCh/wZ0HVimz24sLFHB7odpqVuqr7h4s/Z6wD/XjcI57GHVf1wAXDL4bte3GPPp40lx
Vnx1iBiu3PMTrlltz1wR+RD5JMktCMZsIwxvvSvy06quux41SYhzCQ/ANfeF2EajNa1s6zwXRkd3
CeV1e1K2uPQB5Ianstd2Gp5d4huRhra5lRSkOyPZdvTdOQcOMzfTHHaft+LqdY6zPiCkTjUoPzmN
EBzJ8+finnWDIbKbOAG34vM7ezO+TrQdFcK1BRDT4u8WvWuv08zoDDAUWC/C2He6zKooWeE1zJbK
b3lX0ZBkjAEgRUN017yRWoeTQkpqTqjTpthZbt7zbEh6j0Zxpvmj43bSCrMeteBd4olFgy6ErBKt
gHGrXZjH6L9izaZBbQjmmJHnEuo3IRblmRWEmD2TIJZLvX/O84fUsV00PNcxRph/UwBFO4w3E2SI
C50iT5CtJitbMMhnGxcKm0aXD7K7bz1gaB1+KmhTIoN4G2lrZkHLCS3JZdIpIBDnOEY86r54h8MU
Jc2E1VduB+rkl1S+DLMwuhFzvStcuBlgMNf6kLwPfVo9Xc86VztccNXxRoB4C4AgN/lahWzU1kp6
jwyvxIJuZ1sjM/mVdjV/0n4b4oxn+SyF1lMa5SQHWvW06oGtbCJMVjpG6UqHrgmgsHFv3HU64IJ6
nPs9VHFf+6Cs57BAYuSPtilv4Bhs7Hgp63tw90oS4b5OLxVSjm4E3KvYQe5Aa59lWb/tz2yncyLA
a0fJ4demSKzjnWPnJumxjAS7uXHADkl2z0s/vQ74K1MCHf0vDrsBvAMraXGCZ2Kl9OzQEZnxXhBy
Y8SEEiMAiX8LR1F+Oy7mpWpCvSHjUkCjtj/p2vpuBmlrkxRzeKXPeW7JB+LWtzUVEpG9PXMUyCJu
8JvYcWtJU81xPH9dq7HIrFDu0mY52uyyrnDUfYBp3V7f12TrxyQG8Enf55qCc16mP/0MtgST+9MU
qiv1ogr1gf23AoNVw83T+MZuiXXpBIWH2x3fTADUHoI0c+Mkv2a/5E4abP12to/PylT4+eYtA8Qk
AmFbQkXUWpvR0o09T5yvDFaMl/fOl1z1AL3cr9SL7hUaVjxyaIlYjhmmP/I0EN8ynMYIOwNnrbRG
0Psbi8vxNxy+u0Kfz2mtqsLNQukBkzEI0IhufFY1l0GdoOuIxCDo4WB6hPNpZG+dGe1rztZ+uOng
bs/gz8LRRHabXHJsXNrdR83Bx2VnrtmHa1Gzql96G8szHs91aJ4+gM6Pju7LH5Yk+rTKmCfFxL8U
4ykY1XWpNMYYiKnDG+umwZuv8mZJ73YX7mAV96OkG2wQX5BZ1G/xLPnPTsplBGj/CObY44fq3CsO
KWsLohwxI9uP8BDK6hAfUrLyybTOuQKnajj2EuXxFufr6Vk0xMsF/QciyzMfDTuSu62JBpqM76d8
5qWGcUcNnmHJLd/Hke4fiv0ZsupLeTkMOg3cm+isN1Zo8X6EZGHvJUEuVaLrIlWCLfyEWwZWem/e
x2bdRyfGr6uK/Bsicgjo6uSGFehJzyqnvQCp4XWcWPK+1/J1j3XI3rD3X8NJALVmTbqOgE+v+pDu
GRomm4+BhaG5mCEhLKx00t5+CnpbUh2jPDRHtdlHZ8aHHfvla3Gf3LgLCggeh1mn8ynhUTFDx10e
KsuJD8pLytBesJBa6JuPJcfiJJUqtQ5B3IDHTtsJJfubjoijX08MHUkYbvw7fXzkPfc5ZABVyPBG
NyHLGBY8+CGoNEaWYDk7DCOh8fJuB2ocfoo5JzgL2R1ctHX4A6+jNyo7shskMtVQX+KtI34bY+zd
zRXLbAtJmzkxu8RKs6Js4JRaF9w7gXbQ06magTZYZ+yrwCY9KX1VJ3R/GpvOyDYPQGbrnntQ6keT
aaI99i0k75AlrbDGdwysaE3huppKAAWf2i+kdyGGfIbNxd5vObMdqisnzE/EU3GlULCVf2hv9qyi
jtuuNfpsVZ5GCsg7l6a7qjdaowUokuhhqMoR2FrfVTboAog8oUG8jY7Ji2ZupUWwtKXDQt/l5hLM
jNB96bFJYqKw8aPMUXal9Zuq4XuJJR4BfGy8YzczrlE5g3IHV6ujjNJ1a25acLWN85lHOKM0RbC6
p4pe67GiQ6hvUlaZOjwZB2s3bhJe8g+z45bOZGtLlTTBNDObXJq+aFM9mDieCJjhhCgJIiCydx1I
uPUaoj54wZodDLl86qZsWq7m6iE9yUi+mnN+BqFEccaOayigWngCNY5+RsrtpGY20kRQF7a2kJ36
nFt7+6FhB/Xd3oin/4Toc+pVaoEOTQsd5DAGHE/+nIsDi6aCkyvBs/A0XsFTfcnNHORqGK1CdNsD
fiezsMH3nG5WPN2tcxk4W36ESj9eMQzIruwPmaTQqspVDUQoLVhv+q/+RWkltZI3zFp916Wn3kJu
T+qsD1N20ord0+6GG1VEvEXQfqMcVGNuCQokS3L4t57dQQMUDeIJClECgXRWGZk1RguSKHbJxpGd
iSRWSKjZSofh2BRn51+mDbClJoTgVJBoqCld+8SrBsyDuwxEOR/3ZW+QYwL/HwTLnEWw8tQ3ycO/
ZNK0YQqKD/FMZL6zha7cB7C+eJmGYdq7qSGdGN3gWqJJwdczu8rmHsqGUjEO8B+in/iLjYjFpKnQ
qj/vSGilgZSXeb9A9Is6XWD3tBqWlS/AKbG7Aq6Hx4bqG5tsD4uI6Pdq4cVXCDZXZ6O1c/PAGG85
JXw8iSms8KI5RfGaa0x8T21iuiLBTyA+EC//zWGUV/P5xHzjm6El7Wn48m74iTHfUsySYUY3jqQi
kdvhM5UigWdiHjnqELMtteUzlOnRVR3ufAT0yle/byS2fMOIsmrr9MKbolXTY6vxvSJloBDRqQfw
nBK1JG9oWWjFXuIjcRU1bNP/mmXQLpCJvM6j9wideItiywDg8CvhEw7Si0Rj1nn0O12eNFclO0ak
3RndBiLJZQz446TRqu4LMuO8wjKDY56V5pZ9duqs6EQvmqMH1Q3ewT10Vnl3YTWpLxPCITY1Mr+l
0Lgu99mExwnmZJYxvkIZUjVmRwMCxqIU7fGurJp3By+WnaPs+R4siUULYMMX/ZeDAebAVysyhy3x
UzWAluZb7VHYROt/CGICzMZLqgXs7uSM9jY+ahCq3yyAcaJo82W+ZqQ03H65ye4vMa1cmEziSYqe
ajkU7ab99AaH3EQDSPVBy42cHbIbRNSFcgHGD6faSBY3yWfYYzO9dYFxlcZ+WX2AmnF1oeJvaW+Y
Hc3ysq/FqwKjdWwE8buj1xBaUqm7VmVvzPMASefdPD8cyT7NVx1B9/5tZyFUEjZm8Y546/KUH+yw
lwRtGtZgkt5vBPKQ63SvC+G24hb5QSRw6O/sCCz3SjyV8e7k2hpxqhObC8Pbj9ePDeIdNcP3Mi1s
if2wjL9zRWlig4+p9gMbyQ1v0OSMSk4VOhKjeBzh4oiDeNR6ffRmOFtZjr4AS5jEx+ZMldbVq0IB
44IQeq39yjpXMN2DuVYqeVlMV3sFTFTacjnqVQrZ6B0Eb2Ug1XZSs73qBoonRkHkpZNVtsiMnjwm
9DNU5KxSqzT9umaLkXFB/Rg7wlueZc3ktobJ+KzIBVBs98dfwhrIIR55iBDXRfafNxdqf+TeQxT5
WK3yVSqy4LE4ft0I0/wBB5ZDQyxv+yDQPA8ay0ArFaKtDDrdJpfiY22GI6h41GoxcNKUTcGG/Qo2
ItlKMDKkQXW+X9nzLLMFGOnRh9/fyf5c//KgWdB+Sf9zcb62QCFGtAwcReWJVisq0MxOHADrAmdy
fFX3M6Z5CdBNs4tEvKfHeWfZi93mfoSWPfKr0hKyoBVvUtl/7BK8HNyvNDq3/XnNCsYE47M8GpZy
hKff2250tNkKQnipxIcqBOUixSjCZc/pPkj63O++L7tTvmN0Mqr3Rx0F7JNcUawYocgAquCpEtJ9
0CnWb6nvzHtECA01l7zb34/30HJuF6/NGUuncb1InZyg+9LRZqBGnQPhWNlPTeu17oM7d3pBjqhO
gTndZzQhHlnY+6KTMYcLgnDuzjMBvMBeCQtxIZVr8TMVL2+8G07iiL3244h/eC0802dZSLH3G8VF
Bc1hMvO9ixjf5FHRdD1SraB9mmZ1P67yQJwC/USNll/yEhnajysMJO5Ukm7g4j/VXAARkRWrXPp3
qJWkUT+b4xzgL7SS+V6S+/QiQguKvlFqTAowlPr9hjT4YvEIEiDcTyEZ2gfM0YWAd2/AwgZ9zHSH
/8Gj4gaAsAw/mneQ/QuwvJujTGSlm8WUoYUervaJjhTeAd95Wd6IvHYBnGxgTbJs1Z9nJ1HSV2dY
ahJLTiQMG1g3z0I2vcJBKWnyNKy9X0pVQyUg4jq+W0Mh1K6XZAfP1VfKkQh8hoH6S5E+yDR1hEI0
6q58K+nYxynzoodD/Be6XmAK/AQpt6i/4iPPhRiCciUVuWxhlKPhybONOFWJYWw86v++PSatYhEV
v5jsjC3dsxJ6l3g7Ywoxs1cfrk1b3bZ94rFoTA/aQ+Jv2swefOINS+XrB6ZJUgyM5Q8BAaIyqaXC
Mr4HZlGU26bqxqEjQdrJT9YHOt/wHKkMtR9Dri75yZSfQn7SR8lZ/pqI8OhOSC6rzOVbNCth6Imo
5z20SzgIw5PjNV/+4ELa5JKOoYuFNem6bdUH53NGSNM6A4SKJlOh6VyHvrLKQKwVl7KmKm/jcFAG
4ikW9PbsV2XC42E5LyfQoSOs4PSh3HkLqfNeH/Ji9al+LMh41Mlf7zsZrBC9p5hEjPaqFL1gOEp2
KaegieGD7QiL9iUs3ethX7zKGtMOWTWBCVYuIzxRif8TnBSM9+gxk0hkyORhhoQh/nuHofyGfp5f
Y/uAPyjsd5ldJrEZyrJYulSxYB53m3YIWvxbHmUotkexwRCGb6HMi4seh5m7yixo1V/YC/RTNeB+
pPp26BNHcCNUO/kxCeMj5l0T5KEMYq3Sv1j14c8UsiV+9wZiSI5yvamoN35D5GMz3MABMFvQcZXE
aMFZDq1ou/OqPIC39M8/NN8MNS2wrLliPKfmmdMcdFWNbU/LxZv+Iwx4RYU3Cm7dJipOx91jwW5Q
cVIOT/IOz4kHbYIpWq5fcyrQKYzBMnUNucsTZsEOTE+NUANm7ualkZWhT1VJnYJHL0gNj5dyOlrm
307nc44Y5sdnGSO+IpAnO2TiT7DAhD5bA7mFpkb6fX8m8Li7Kx8k5mUvNPJFCE8XqHe4j/nBSFuO
bPINzFFRLEtWMZn5mbqKwM3BYv+YQjVBopRhI2xM4XQ2KWLjDB+Rf+48PzfKiCPLCeDfUfyPejm5
cJdRkHR3JvyTOjRxFJCudvbsT2/T6I3YJKipLJ3HO13qs0PFUEiSN1bastbVzg1OSBDhXbborDai
w7VafLSshyr/UasSB9LIXGePtOIDIYImWvN+bpZ/0Qg3UtYFaTqCAevBRVSmZ336Jd5QFLY5TJFj
2vnPdaqekfRR/sscw9anfX5QgTdyCuXbRh9PsoAFy2tjodPeXcYDZ1IGS429g5CRoMDoLdAMdMOa
4pPjQffJ8s7jszKEry2SaT9VSl/1iEjk+T61BCgZ+ljpP9ULSory6jbsODfJBVG36IXFo85YZgF/
2/J2VjkLVkNEsgEov6BwAwuDS6kRnvCj1LJH9TnAE6bOntp2RA/WTGtald1mDHxPh1qMFIQfk4CS
ClmFJ9frUkpBqF9UdedwA/x6KlKfjkRO5COXaTwnvztCETDMujQy3GRQ0epJIjHU7zf92zwDiOb3
T5ZauY3dUS2iMNXrHE+Z27IuW5kcXibn8A+/JVvzyXSZ22PzXeNjrUO6qSA2lDg641nWlV/IzK4m
Mi75bv+QC+OAEbaBQgUdU+dLMLHd9RinDi6B8FMLcAm3WsYSJtCVD1bVo6JquxfDq9QWf9Um4Dfo
iKJ+2tSeAllQ1/BzqSuuNVeDUhB2PCFDrnhW5NQpFJRtgb9Ayfzm0jpJA9pDwK1HXcutMKn6VMXm
nFcoSHnfecO+9lupdBoykgVxU3PVJvT1dxRP4V5vwBh/+CrtZ2vZBYE641OaI8J2iSce40HIVrTY
WUGCKKHaSjlAg7/466rV+3dSiTHT3cnZUxDuWXF/bHncpuY/KYd6iniKaS1BwiVlEkF69XZ08Wcd
yZZVhiiDBY4uQjYtGcVH/aoO4W5kpvVwl8bBzOQIN/jg81uJEWE+z6nrPFTUIPxyTb0EhRU9WMwY
P9w20khkjjl2UgkYGrb8rW/m7tTizriazgkhJjTzbFgPGNp6XZZN9XaeSDPphUse3w76siCLRH7s
PC7rXsslSXv/LqvPqcFbBCVb5SjSTLFXhNYgJMcQvNEnnRtBmPG9tU18Qe6949SAhV2R2Mxw5s+7
ve+EjvwSWrlEItbFcT/FoblUqp7aBIcRrmy33H19h9Kpobs+exuQSgn4JqtY+LP+8zksK01J4IIU
CPynV59qTIAAPr2CcGP2srVzKoEc8deHjUsGyLXHOtofpw4SHrLFjtXr1ydEGzi5HtwdTDeR4HgP
4vitjtBjhgQVVjpHg4il1rAw3rUGc7Dfyqqqk/JTeF3yXSflAEbLraSj9ejhH+wZEe7ILhH+K9Og
Sb958cIBt/N0GNvghRYAbxuPUAUG7rAeVjJsxdshQgVupYRppVFwREt4kYCQzx9LM9QzZsODnMe2
oTtxa1zujkDHynRNOTydol1a74g2899Ihuq/shsErExOs5v77qee6fgTQvJnmSiuvNAThZ6YCk54
pGQgb7SQhSMyogX3JzfKhE6OTku0XkKqM3ukVzFvPahaLlOsjXJWwERP3SOvxB6p67PrKdMdhDuV
CfTPa0wP1UQn+m6kpW8HJ4YqgW7Xe492cqPafqFgOCAkSXuhmnOH+ul5Qzfn23rmC294K/XMC8iq
eml24lheidUQ749eDuSFwzCAUOTcC7gApoBH1c2Aj6X0p8+fzszZSafr5m667CNtVv5/tPj8W496
aQtejjkqQA+RWMV2hIYx4PiBOGDADZDf8l3lW92PBnoHMi5v9rvW+GbkMlkFa4S+VTK2U7CqoTGB
CyVvPY/YmtGc/iv1duQnD3j7Dpcx25ZRq+pStpgfGYZUrad+EjZ5KWsMIJfjkX7tM6DVLVhNWnhj
74fFhQV7h3anZMtUBbJG8Cx4Jg9K76jrztop7zMmDgmTXtXzCDw1iY1idMAG4vLfcdDbM0vJIZzR
zNbbi9pI+rXyFaM3f51IHL2iWR+aooqmqdqgcIlDK/37boahpi9TexWaWGVBNslrE7GkyBl2XwM/
vgIzm0q+J0YuQ5k/C4wFv+tPhAp1evojyH94djeO+qj4IKnI73YanKbN15LmjnxD3AAlan1QlBb8
w+uRlwPJJO1d2gVgXU3e0JhNwo9bDaEsgLLD5qF/aA8bkoRi6nxPJMf5ZqzZg+dm2BYzvlbNEm/R
Zrt0rXVltoTd4b9jCKogRVaiBHsX0pe9tyzgz3ezJBakHvcbYjWJq2tFBwnmC2YArhXpN1Kl8cz8
qKCO4IWu2UBNEuBRPnn7E7WWvM4SVN1oPRJfKlQAWWnZWtZMNQ5cYftFiBGxAsip4vkWvQ92VyUV
046Ys4D/vmsXvgekMJQEpcfmAFvhftzAmFt/j8eTZb35dnQt2WhSjbr7Sug5j15+E3W/aqstcw/l
8OrFbwP0YP8e+TuPEtRc3zUW5NdpGfqHdGervy3f9lkT5WejDJhOMsPei28W+iTS8cgx2OJS9guu
PPm/nBMJJhiJKR8appVQ9eqYVEdZ4zd5eSoHLcOVX/ql1EGon62897R5ONERvj0ZOSTpbHph9rT/
6kG4zd8or2ThYKcMPdFChCe5D9Bnpqv6KPvlXS3Gdc6jOwIEEkv6iNn71lVHd0OyngRBbu7oaTlF
t9N5jnJCXieyQ1WgkJW/a5XIhu+wYQGiA4gxPDZxgN8SnZwlruS3aEz6YBm81PJI5UV2U4NAzwOq
8IQb4XU9PiY3rbyvetab59QCOuP2LKTn5hTnYbLFCRT0fArwemm3qnw0Xn0IakU4Vr12d6+7nd87
qeSsNY9ynYh3YtoJPNrkNGEDZhw9iUNdpK0/srySnp810WbLtNJUv7qa2h8Pu7XzBkRUwVsexqxM
JVqt6z5XiMLACgU3SbyuJVjVjUHx/XBhLzxmgNE11x668wrrZBxRMysM2E/xqZkgy/K7zPtJScg3
DXabo5SPzQUwdo0SnTc0V8l5rYsym9eY1WHZeMk5JRdUSNn/l1ZcGIkAa7FtDvobFH8aLMjRY/LY
oorm71Eiwr8iatM5oUqh1xwFXxjWoajV7XlQVhw4c90fwtqqZFCq5enNwDRHqbyXvpYdxemt9grF
PYLuUb0xLIM85bdk+HPwW+yKXaJJLlugsYeqFzw5+8dL2V3nTg3ulHe/48SC3O2PgzgH9dt6+9PZ
mYbcWuPPvhjRE2PGdSihrTzwHFLmMb0U5fdCe9MI7G+pXo8XUcmJHAePuleEzYw+Q9SCRkQdniNu
tZCcyhG5RSaOlUhZvzjnI7lw3MZ1Nceeb4TggB+bY3jGeuHvwZIOn+ObLYteAVwlKAA8eLyjSx/a
Xm9qd6e4mvrw9sMn7rjBJG++/4WPXccZGKxlhMlAozd0/LbgNVqntrSgJijwGcclQ1CpnJl1u2lo
NnBeSiGznjNCvtepPhNwcvFsaNi4qUqtfLv1KyaPsSN6OC8IAysvN5XahKPT/jtRWEoKT+nc88Ix
oW4VLXVw9cOz/MTCT7b9kf1HmGsOisfAJfqokEofB5DVykxZySmoNO/RTPqyQPYTCMH6XAeNCZWX
4EzrDX+KCusBYZkftG7xY885XYV/xlSCIjfcWDhyMfpISW5lVDt3R2S+DfRf0S1TvJo4rF7GvibD
wnFIsX6DqlVB1/VQ8GvZgY1LjsNAEHWWbg4jJUWbnFF2ZsWu4HyC5k1S9K4l+dSuVZXcWnmUKlLA
SqJKJgeZACOYkBSg699TcSbHu7FkFWVtqPZj39WQJgTfNCoQQGfokYInzYQVQECL9Lvay+A0MlXz
i/gH9km0G71ehAYu38v8zxKVDCuPWN18f8S5CcmMlf38J4vG0DBmY6VsfbYonCnW3QNyJ1r4ZxMx
JRtO663sXqpsLicgvFSCXm2J4tvQEFPY+T4qIfyM5PdDyV/xIMzwWhm1VaRJ8CTtYSXG2P8nPEzs
hg8mResoh3yicf6NTba8jmPmt4foN1sN2ZvZ1wSceOFazsph35RM8wCDRHH4+VU8r7mDmHDd0um0
HD80xi93WnuUnYWjlNLR4ypfah6BDmGkxX/HZlhmSCAfwEUEFGaQ+r/E3Ekx8rDlkEi9jARUvapu
xdTloQksx3LG0UVkGAlRe4bmJl26qZTxxw963IlGkBxsem6hxwsZnETpQaB68IxLtp57HoL5LPij
jn49FK4zN+s1d3I62X1N0472/VXKt76uilwI9w+H5gkkzwvfP/+V85P+ooSIGg0hnDSOZL71ZO7t
Wy925G8Nycxom6dwTun+LawFweq+CIxG79c8EgsTtSAD9HW5uyg31xxAaoFoMwuYGnw1jx5iTSmB
hGv7NrxIJHHnxoSWXTQu+5W3kg8GnKMbKxIL5ynBPZ0VO850WaCEbh9EXmR688aXOl4nZRhFr7Ks
eX3gvn2vRtykO6kqW38Yv0LJ/PP2QO9mmWHCT+PWQ2cvyYifvXsqgekUQcwouNWwiLkfwao0wAbB
mLet1oB306nI9tx0HNF4FrbMCYzKTz1IlFys1yfoSS65+DioEJ/n++nsTuHlUnVIwEOsS/cmVtvU
dlXqtbh1l4lgcvTtKvMliPxaCPuDEWiqN4xeRw4syp49I6jYDd+OVvapGGhNjyb/nS3yc4ZncR6i
mU8LUaiF1ctG5TLK9Ttnw3RXCEwPP7t4Uu1XWZM1o15DJsDpEICOpRnyqe2594ggQorVPEQJpxBN
Lf2N+dLifz5QKHcRa/1BSNaGwfCMp3yUVk/+4xmbqRz94+ADtOtl8+VfhbZDfG1tq5UDH79KBWro
eS0tFmd9OrjbstmBzQKyglwfPSV7G8Sh+oLhkf5pmQnACR57GPk11LqnZpG7DZyGoWYVp6QpTxll
t2LT2MNrckNbvAdfaYl2+JOPQWv9JgsmKAhpfjt7dMIaZl9jUTcVM3zYLe2Gi2gM9H3TNQ0h9Q7Q
KZwpF4C0kf8eKc5oQPqH4DwgHy7mpHg+LDEOGbIROAmhuD5tbuEuIBwOE131VJRG8k+Sco3ksyh7
wV+dyXl4opY2FYF9Jem0S7ebu65KuicINFuPC7nK6KlBxoV61mSyzLL3yQ7VLWsUJCPN2Q9M4Ko9
L9xkSRrMpvjOdEWWl3fLKqCdqjwZzQM9qa55kAQrVoduv0/adoJ0/DNnT1UeP2TTOW9MJ7hskxPO
KKsKbQMVGPMIN7rMsVVXvuluU//QXj/msOcm4c0d8qSntYYZdjHTfmCCeAH/raWl+vtUSrFUaHJy
eUBXp8yWIaxc7QLO7egynzl/aFzeCOuyCw3FC/WIfNHPU3To2quzxuVt6JweKHfJ6139LVCiUysQ
EIOwg56wXHgdJ7fcbYZs3j8IpqIxEO2Sd+7d82VLGeFLseV803rYaAfyQfYHaoHr5/05EcYQI5pQ
cyvOm63ClC/Pu0IQVwfFzg7Apflx19z0Oy6VfD7G6csDMNa0rOdvfD8bqyKKzBKYB8V/3lGkLfzw
rl9R84c6a5ju6/fl2i4JGk3Dpr3GCt0yr4iBxOarAhAR71guurlX0q6KXFPBGYhw4whtCjdQs12q
RAdm0BDw03KXIJXMz8tS0YN5vO0WOnLxU35Bfw89STYM2FOdc2Lcu64uGqnIoGuAg4SP+e6qBU7l
ZPdClYj9abEiPfPFH49HBNALK8suE5W+yYUSCcSQlTygfPhwhCeK7jkCXMmH4xj6RAfJ82UQ0NIU
PDzK2F7bpTDQkkX1CKEe3Dl+hBszNRzp5/wT2Wdx4lZhy371I8fPyQxf45y52jT5MzgR+Wq6OS2l
9+Wh5tCnf/tMWRTpDE8/mAGsqxN7sJTT3sWv+82ygx3PSz1BfI+Sr4JCqx2eNOJHb2Z+w8VlFqqI
pkCtY7YwkySAbdR1JoFHXmDyYVOZdNLf5OrLiYKp+xwU6zoXVcVjkzPoeu0YPyLCscbbqiCI7Lbc
uRfO1ordI9EafNJ/y31ww/86+UoIEhxvdLW+dY4mAfO6/+7qlaOMZQ9T1UGHMCfWvPrjnWNxBlKL
3URz1Qbu4cM71AwNm60Bs5AYTw28Wx8e5JV9706r4nvurP9FDMRW808eZ5pJE5a/DZ7ZaNbwOKVu
uLXA715r/s4hzRbLweBpgD4Xg9bgR0wa9LySjUvby3eW7BBMuACwU3chpm7tvWGx4s8B7HT2T38b
Ir2b2na8FXCVRvp4FlSy6Q0ATqA8Mk4D/qPPw5yHaJSl6P2UgcWuAIfBv/eXTEiJUrldav9P6Hl0
xfm3CMxB/yL11vD+okX+BcVVn14wFLgnsbX/Oo2D5LKRTFWl0VuZWo0AYXFpPsoY1CjoNOV0Eq1j
VwAJ+DxdnNAhn6rbvVD13WFJtK5i6IMNX1MiiHLZESXfFl1zsWBUhXG1EbZBOBz7idKvVN3804Fv
4VnOolGD7+GRtj3q4+KW/WucoSepRYdHl7OB9RM7ApqXGjzD1zPACJVDlQWDbhsUKby9ReeS47CT
9vBVj+J1cJVdBya6OLSIl8bPASpjPZcKx/PbiAgMGKH64QU4MfAJE3iU2IZIgeaPke8LRG7DABub
M0AizJn700cfJPKpFgHReOVxbpCKi1d6l01A8MnhWk2okBS36ILHlQeUZRM1Y75EwssmN9jO5kjl
cS2+GFgF+gG8wGE5k/34jJvOqJvY84N+6uF5mqMnqXT0a5la/TaHlYZz5ModGS96c9DsdyLuVBC3
RIeg/JoAIffbhAsGVEIgvfWwPYOQyZngZtDudTav5ZgMVCctTxybg2Z2u0Ou39eYAea8aStgg75Q
YRecfv2UfVYLWEbO6hc47lHPo4FqgB9FCB0ZlfIjHsOUOpgB1t2vWlfPCe/jroyghxxA1AHr8+3/
tud53iQg3Oss70id6P1tHwgU+8gBLQuSsAzbgxT8K1V/5rPz40AN6pv+gSnj4ZJtNU6nlyaStRpw
yTchahHkiruyHwHxAN10/lvw15aw8AEkGPlJ55bYlKLIGzE0oOmIwQWGuWHZlFCS3tYedwQezwFY
4AFB6TlJbkZ2/0xQ1pppjnOGZXBuI/MpIskTZMABVEouuVqj4nJJnIedhfShLH69ta9AfOaT9nWJ
IsXCf4Y+7WtZAuIL+r9kjdNQZUyuXpXp11eGV1WevTo1sGMwxX9Gh5E0nJ6BRrMhQ9QBxr32xUtM
iy0usfyWKSRpguyrTFjvR1HWc5Dw+Wl1KG465WLHjMn0+OkuSA8ztjefU48bF51WkfxyykBdDK4j
kh5YOmxDvchVbBG3Ej/6ZK4lQSDWYDm2YsimzbxVZDlPKcdnK62zMRRpUT9SEr1CTXt0YXtk+kAw
PSU2YE9fI7ai6Dw+rZooZz67yCfRwmmoqrpagBnUqESyqsH3kVhKEo4bIuT/cNUDv5EtOQup8+jN
qAZIcPTBH3A8nWq8ir+YoIcqD9s6fPXaoVFkMvyw0/2JXK0B4c3g3ltBY4iFLW3xXjDZoqieIFYY
ysTcT5UbbnDn+9XvDxy/f2X6sD2/QyQ4R1h4LQVFCLqkFrd1LAX6uutrkCqt+qt0iK6J79pxB0bd
P+PvF0yKzzfidcbVapnNaJ+/yTPLxc09TIaD/222vF+a7sXVOAwm6w8qhwd+2mFM++EvPB5dF5uO
U0GslalnANGgbI37IK4sQEjfx2PsVaBzvW04mRHljLlANmbPBvxwTd7Lu12V10BXAkHbiwaIuw3W
+ejOR0QnvznfJ0VMrzmhQhsQYCRtTwCX70aafzkdU1Gd8hfbH/kAp925MZwRhF5Mcn1FEKduaMmd
qqV1+wL5V/DQxh5TwEv+K+1dWmox/uf7cHUUgXZ1rxZAMKei+w7CEUcpKiS4B2JWaxB1EPzNrel7
w7IFoFsRLAFCCe2zqRXSJeT4mRRu08tgCKCxv2EB5ldd1qH7oxeZu3FXeYjYji0RYeYUIDBrVBSm
9+1YtiXUZ94RR7AoDI/G5k49f3+JRxIMnkeHOgIMZc2+EEwkRXg5PV3F3Q4so9sb6swjX28W1px5
W9RXrFznB/nfozP6JUMGfyJgs2n6sKkiSPk7TQ4lytXXbHdSWavXBhjgJ6RJE5xE3OW5yOpyYPYS
xF5TonvC0563olLhJ+9UQn626GHugJQ7bgmj/Pf8Y1xg411zgLGMEf4U7NeR8GRiAw8IZSqDZX6y
viMxCPGjcvESW9+Yoifg/koXjEBRpcZiqXvjdUAfy+3vVJTVE9wau5GYDjFlub1mjPRfRd0Xd7VU
xsa6lHzClaGhpDRWRoTf7KXtyCDKajDOX7RybDAsFOXzNOImFXYX5NxwmUN/yvYA2+0Bismh1t75
qx2uW1wIzB3tELEqQ9yQswuQgMJrUwqlGzq1TRDBMORD6JhbnftKUMSSGmPt6JZVhbZYYOqS9Pxr
fRyOP7P6ncyzjjT7Pj0tF/n2Nf7wE9JcCN+4UlMNLXQfi/cmirNASZMjrKJYhXU+FpPnUVOIZ/v+
8BkJ21+4ZGXdI+J6yTNTjXQ2EYONM9v4vUhoo8iKaWZbh0hRXwdjswMv8zSQflk74ajOv7n5CzdZ
X98y22sCR7QqJtOUgt/4dIpwdFBZpi66D7nFE3uIjdZmm8kjxOjqNB1A43JIebyjlLachgNGSwge
qNK9htjXJA/ChPV5B64xdV5BGeopbSk+xy02mvbcWOGTCn4R/EvF9tj8iXOihA1lX2tCE3MOsCVT
pIb8pojPZSDU2I8AyiHKT973sbjKy3zmEMSSnmTatkFry9LrbqU1+HGpqIF6271LbuavY5g3S6iu
cvpjsKCjFdqITUhViA7Ha3Ibil+efVQhmGb3EFyuHS2AMBbB7dxtd+C5w5IUUGc2SdweVau5MDfr
rnwiVJfMb26ZFEmiYEKSjXF+KYKTD9Szq11z4cCXHiGHRs5MRvO+xGKjA7QX+OteDlCh2Di5aXV7
f91YxHWiSiFdkKQy5hnD53CEnHonnqIq/Epf6tz7PxJAMmC/p7IS6ZwzDnE6HQpKrUxKjDP2Md3V
XVXRi/Oj25KEHbbObwcQg6k8elG1mKZaCzNB4QgD9hzOstHv5ruawBdgLOCD7uYKomiRCjo9M91o
IzbM/OdXUuPaH7xMi5io/43WiRV0Zhkws6Y4km2Sb8Vpefycai0vqWlV/RLTSxMkkBRio8hBFzmg
/qzR8ZUxam1YkH2Vc1Lv78VATdtJ+s9e6ZiZyyGshAO3JVzYw6SF/dgpAMQtq1Mm0I9OG4eA0u/x
0u3FVYZwpx8Dq/mOSNPdZBEnEtU0+7AugWAO32zPha6YuQwNjNApIpXLHNJpzlA0CWh/ObAZj/eI
rllMiewwmV2VkRFYipDOnQHiVVlLa4b6ygpFHgAGc0Czf5fZLF4AW9Xz813eEyl8v2Q6l8Zt49LA
cyDW2uyg407NeAvPR/6bwlMKOhgsthA/dOccVrVZzazlDJDWsg+5AXCpTWfzVILOzIyZWmIsGtaK
cWr+ykzd/RHY4AqLaPLPuuHC7iIU27yoaZFHGqLWgAYL+4OPrZ67whEmGklFl0bbtXWObh2dP9cS
ds1EyiogDm7zd0ZFwC7h1ctvUXCJau0E79fHwc9UOgv2SjwWMuto/cckrdbmSz6pR10E2Npj7u7u
JtFmexIc33wpqefsjyc5F+Z4D75ZBsuR6j7uGbM9xgN6pG+Tn7kcMsfICM6l9naD665ak/K+M1kL
nN9bcteIs+K6EHC+ut46XbglpskLsCm5Y8idanw0sT93SMLR4NTKAmkzbdWwAnWMkjvRyNMjjjn2
c7MZlFNMuF75uV66qqVLqwWLfvaa+C93iJkfX8AnjhcaWtiL1UY7QtzMCyfmjIsJBaED0u41xdhD
nGOB9S785ag3yCOxVkSBWa0uAZ74g2vBVhIu+w0+TG4GJcgvFS8ileSe7iamkkOp7hGCg9j9veuK
LaKaPVZTdtl7g1F2+i00idCQiS6Iu2bC8k/9In3BLmqawd/sJNxgLV57oBkZI5hqd7obV52UwmR0
E5CCu81j6CfeQjbvqr881Qc8f4CZNVLskP2/T4u99klRjUYX4af/DuFb9EjN8BBP7QiIKuu7elCx
wxpxQLXkiBEoCc0u5SRCPbLOYl8mWDfAS23tt4YjdzIFWc4fzZaaIBXkb21pOcMaSwW6gNZkmuJ5
BQAl3SY/A48h85mQwHPg8fx3gAkN31qneBQhATiRUPJLk6y6hzr16XyVH9Iu2wmmSIdNmG3kR9md
yUfnfhYLZGQrBnSh57dqBPOtWj8ts/SDXKDhWBQ0rkawo5G9gZg72sAmCfEG8hvf0t4o36i1sqaX
mzofwnmzwDRBY5iCzrHGZ2mo00ZRF0xSRyL5xOHSkeYQLDKStqIUm6YLy5CSy5Lk7fqgS+7FWJ7l
fw+2cEb2ZrSqT0vaXH+VhVwrFtFRA7agu1yQpqX5kB/ZIkLv7IVmAiZQXyfkPFvpGONT92qDxlMu
GqluRPm0lJCQ+YONvE4+9ZjQCzRFgnhOZ/+UswJFaXWRqsJ9oVJCPbk4pakm5nTjo9NWeOD+G0GE
BEmHIsqGXpPDlY67auBMA1rb8qzCiO7CiuWq8KPpbGyB8nGMxzQ5NPkSgTW9DI6LwdPYZKhh4aQv
2U/Cd/xmMmsOUKELd9JIhvNvZE6hOqpGcvGrRqLS+Jx5PTRPwxyGzxwdY/LAVJj3hiM2cdZNmXbC
nhVN2EmK/M+5awsxdjiqd/7ePO3Cp/sUrX+3EWoWCeTcuLEvytR0JEvgVAbBwNLt2u79GkuXWUHc
a0rNbaHTU9iRbB8+xF8hQy9hD9vY7PlHXeOr/onSEudS+0d8Uu6+/HPTNbD+7ZkT6TwTwuGyhkT9
fP7NA0Tj2Gsq+xvvgum8KoPgcv2DBFKntJTzeHcmH6jSIB3ouO+31H25my8GTvFxhSv9Avd8addq
wMcSGLWi8O68CRyvGV8xf0OtZMHPM3YSwAOeFm+N7/woSJ5pd91OIiNGST8F8qS/cmmDB85qQsJ8
V8KkQR8B4tOCFXUTP5pTIsJ76HzvdyQ2GO+PSyDFbXy3favLJ9FiGgUCsQpZkYdLK2D2E7DAN9Yk
EsBENWLNmw0QNJKhHL9JzVklioVnrYaU7vE4+xrwZZJ4WkfVZYQNgjHO2lEj2TJ51zArEuYNU52I
bqgtyEhpdFV31dXF9ClxSXQgBY1AUMiaPzSMSyI4kySO0K4hrWToDpPdA6Da3sUPVA7AwVjo06aJ
ynnk5IBzKfmEG9CEHxEmumjOGTYK9Tl3bJEMMras+TPjsdla6HL+ezPb9dCLRc+CUAa2pkX3HSPd
Wp2Ihb7QYtcOkkUFTHiISxNDR+YkTtxGpt8NbNnk5cR7dQBBGH4cZGPcyYO13o+if9XEWGQ1zNrj
GU3c26axWgxyArIFZv2oWSFuTcNpbWGgQfUOmHjEvRpCukDWz74kTIkbwJ0CtGfsOFf/hcMoj72g
B6M+loIXJeLgpGkPIwj/AbDTNJm2jL7ao8Mk/f1nmIMC7p7hIqq3dwYY+H02f6ORbhSVceSkIVIb
KwEgPyjrFwkbLvdO6tRdSk2N7ssnX8CPVZL6RMltjGqxZeF9q1B5AYpL6NVr0/UzM0OYWSOHhwO6
lbHz1HE2MfMb06EF+hk695MZYo+lCB678IqqWDDyAZMCCJkkSTvpDLZAyW7rleeW3966QkXK1Tz1
TF7j0e1UfTC2tA8ZxuMEQB49CUfdcRJWwEkRpOKPR+FGOgitdvcJktaAHRrBaTZdPRHGBCQ3wzPD
VPAg87vtlynwQ5qRpG654iy9chthMEJLC56F2gzaMzcqvr1PRoIjAVR4SgDCLa4QgeTGcRR7gplw
NaPeDrNeMRqB8+Xbm3eDW6kNNERH1kn2mfhZ3ckCu1eype0AinhOMe1ULId/d6tBDCLlZ4Jf9pG/
eTptWvuWiiwb4R6UdbuNPYgIFPipebqYQyE2UqSX61MCOc1UlIL87roRFxFO/nQHtc/5caCdTwTM
YK6v+1RupxwjVvBDsj2u1UB4T3RzmaBx5RlmOahOCDSOZkO2m2BZ4ycJKeISk5l5eDuQTTeP4apq
mnu+lMp3uHCnV00pNbnicbA/nisH6wiO+XnaRRSnLL38wCx4iacGsF1wtltkB7DaVZ/pHKwo7NRf
v6nQu784IqaitnfR1RAHFiHaJpZwf1HN9ph6vxwPm/3bTCbqcdMsNSv8AC8q3A4IwJUP3D+Lr68G
kbSVH9iCCD/vtNqfm3DdvmpbK7BWOA6uChzO5PQOVBkwfecbNIGtGVn0ixzG0PXI85tgzm7UeonV
20Mgbbpw3a0W7nskhMIhrO905OEhjiZx/hdeHSasMY/BHy+G7IHCoAHsgDyZmCg5vjQpRBbq7hJq
dD+mYoMw+m0fiyAPsRQvG2G74oUNVVB5dUUTbMBdyOMxf88qfFksQFJX5MvGMThGXAsvXnmmaTzd
mlRIBi/IIpOacbnbK751zWrRrlmSpgGcedI/3KjIiTr6nZ4sF8VzywYtDUCklzsZQjIRgG0seQvx
uz8spZcnBSiFT8xK0rzNYp59A722qjkTFzXgx4v6d20KMrHxK5d8U9DiSKOnECBNoickLDhIb8L5
3nEIWRNiS2BQjjxgQYXxI6WlfErypSUYmmsj+qCCk2cTsqvYTAUqsuEJwlcPmgeeL8l+uhc4ZiSd
Zpd7BiU6aWIrc0QILt17rkguYfVsL2+bC7kToIeOV0g+FGQj0U12pEw+35+TStWJVMFSjJsZwk+5
HRUvmBAAXUz29gofn6AE19HansolV9XzMRoRBq80gq9NKuBekpusRXeXCkDsNyEpw9bDxn3JeY37
FfdOlXhhJ0v21EYPqwjug82+vU+K+djTXS5wT4jybvzeTYXR5r96Y2FPktFvZz8zCDz+PzEpLo0e
dBYdd1FbnEyADxwY9N7N8ZHy1tdbva12/TvgpW8mgT9mxZDIuqcETEWwQVFuy98RVJECwNBR1IBJ
ynAI+gb8ZRsg2i52j3HbHLoiD+F6CmghE2/h29M0vNp1hGYq9gTXcIxRUJTGewT13G09nzjrrHdS
40Jo5Hdwj6M+po8dkQj44Gqxobx/KsTpQFwvYQbW9itd6y9v8AjWX9dxNrLAn+Z0ZhdBFoMV6Wyo
mJcYS2dbB6lvMuLf7PkAKrids9rU5rIvIO6Vn6JtZBrlyAHLLMEmStkJxpN6/Nlm4Kt7m5qiEHjw
VneRtygHWnch4/2bS3oFUJVPetIDkg+0uTj8+0y1LAJFI4KtBAsBSWH8d+NXD5pFAOZ5g9yAxPoj
FN7n0607HglQqzIljdWDRVWaXJlMTF1G1i04au5re43PQZPu9uNdntECun4Hifn/4fRAoUl14Ild
EwUihjXpocmyYSJWVTSpr8euO6o44hDwowJh95VYrQUCcO//uD+PkLrtsOAcFgadHi6MqSE5LKc/
k2cpdQHYhsk+pQGgXZNB2FMbkUkxSTTyGF+WW3taNrDrQKdIM4+fu3x6uWBRX9JgtSuN9zrVpNzy
FcQeaugdVgd6llph6rZut44Av0SgLDzU6THxgsucSv/5VNQW+IMg3BvlZ9d9jPKEz8CBCiK7rAQ8
PvCpYER7FC0JR6TUEYiD9yxOu2d1S9x6Xo85jcECw5ssUfl7Ujgt3b2eWxx6zygsjhXyZEPKhU2p
FsSPQZxA0BJWE2BPtkUhu057G2qxdoq/YbKLcUESWpvXygeMo2M0j6nx1K5DDA7sjLkSx2xuk6xG
nhwQb+cpATZLBbUN0eRF5CvKczxuTZapq5FSdBARempEpE4ccSvnpM9BTBAgR8TJ8pHA2sLN5X6u
JXxxYtkbrJ8oZifMFB8lSJjdXmIy0z+Sh0yPRmeQKNXAwc/soy/K9dJsE5637Oj/G85scvRfnJf3
/kiToQZ8/L7v56yYOB4tEJr9hUjw+5HaCbeBg81SYZVeHHgTL/z6HGyIShhDqTXRCRDFI66OWm8I
lLkaoQ2yAEeg0ay6HurAl6zXEP5cv2VsJbiFgdhH/X1+3cpzZc0X+pRq3myPhP0bhzc3lvbBxD8g
kjpf4lm89aCeIia9/n87c3JBTn8XHXAJ1Pbz1k7yTdtSPuDRlZ5gfhXomuMfxl4h/rDFn3bY2HI+
GaTwFEDvnR1GpQf60GclTmY4b1yHrRo8WSdCvFxv+j9/mg5LUa7GVIYC2IrnfQ1mheE+K9uU2edB
Nn5iAJZS3tU+W1yLCxZzYI0eO6NqlfNrQyN7DygT8ZMgOjP8hFK1il7I4FaO8U/fJOdSouz9pK6A
+uwf0GaUwHMuVO0ouaPMNlxi13sL3ESobq0V6YlsBc1jJIMu+hFZcmajY+kj/sok7sd7TeWMTIwv
x5+lXzgPlNndtnZDA44htuv3OvX9UTJfoxzPpRyUa7gw8YPR+zF9U05KlQZrXEDJEPEX7RAIej4x
YBvG56B5/KD7tqBcpETH7XaS1MeUYRAz5xg+kuudEYm+ZREDFLxiHwrBDwNLj5UZpIGYg0nTpSnf
j9EC7JyvXd1iBAj+ZeXuSqCR6NhmUyEQaPFCE6JrLKWRENsKyvTJuxIkqMC3G1YfjFDxegmJiIMa
pZko6iP6emnmZFGYdMDHRtioyGnMua0051vK35YpYf18t5geCyWlbxVDtf1nFLc+9Ca7pqJ7HlsD
89Ncf1ZsFcfrFn7EMtp9OG/hwccJ+r0ltVhW4TO7fcSUcA1SS/PrkV/KFNfE3jhZ0W7UoNcN2n7I
jufXD/9WIgUmsW+EWKXUdln6Lc3y8n4YBaWMneAbkg/uxtpZGrok6buRsjedu2LhBOLyLSoTFC5O
MuMa3emDbf58BKQdwUJmY5+9dt7o7NNJNSjhJJeE93WCjWNnmdC643a55VfLavnqsStAoWQIUjoj
E7TS/PY/UuWdWbvAF9IBMuqA5fq+LeRPRxxtBe4rOqbzJTZyDrW2i+h+rQ6qg+tPSiobzFh+dSBj
DOwn5JmFQ9tLhxwbg9n312pZXzmDlNatFonwMBLbxD6a9GZ7LKjFjbiBqjvVF5ZZ74fNsHayImTR
a0XixpB+9VXQta31+l7TXW+dAnV+TV6zFUDMV+6kK5X89kwsrpfBf3QbMiml1j8sKNsvioYRZT1K
ENYwXU/upZeoAOugPYlyK4g6NWSA8ysTv1ynq464NmqUHGVaS9L42QteZkGUgyQlTibVsJ+Q63ml
OVJScUGg+QQqlckGaQNhX9L1o3xmCco+VMeHY9bGjBs9Z5xBk1zBWg01Y9vErYSAb/fyodKE6nQo
pF7+kwVnL3Vz51Y1t65QE8P7Gc7VX+dOkSWVeZLUra3UVBJaAbDgD/Wn4TrK5nr+MowWsSy5V2cY
9Jo5zyhjJHlzp5nXHsuOzP9knFOmaW1X4psmI70R8NcQ3b148EbVUxldvlV4LhK0oHmAnOrDHDHI
k2u+VwUXwxeauh3i5eQvv205sVfqgwf1SG37YzgA/N5Tixkh6lRqI4Nh+he5pcG5R9eSaJUw4atX
6iObZ2F5bkz5wezrb2pFbLEWmEP0wIJ8iGKapD64U7FJ+OmH606uSWBhpGei9FcUTjIMP7FQ+m7e
4VYJvpwmK094IlxTF4AD7Hp6banfCjFw4/ZVf0NZG3XmA2/vOmyhlmw3Rdro5rcChKYeuslkPgcz
OO9X4quNjkihYIwk6a0S50rGgzqCzU0oYbjx7S7VSEKPN4iYIVaIVP1qAEkEllV7l1bFgvEiuRx0
orI7hIvy7sI4m8IHT1UA3OB+2Ecbg2LoUeTGNU5MIRUq++co0/TRNFwOLnfPiotMSTiMQEA9sORp
qemh6Fm0QVjZ0d+iS48w4qPp9ZuH7qH4xHGoI90MuuOVyGxlxi1XlCBSl+N8mcKmqQofx59ISIc+
yUqK8DTEQrcDQlE7ypgSjG6/fN0nkfnDbi9EqUo/3BqUig93Dps5YMzhv7aXAqvYWju4KD0LPcOF
Mp2Dggcirg0hc8TUr/D1F2wgOWiswgUXWdkh7gH6qkv2mfU8a2B4HPqx+fPAjDHJtdIFdBuPxd/0
QucPbU3DQ02cADwGqM2AAP8gW7JgD/7NMbbDZmOumNgKk+l/LCrjFyeMGxbxOCPSch6YnIkg+BUI
TOYEG+kloRKCGUMYIO29NLgieFkgCbXutn5oFjaBiQkqQDKpMPCBHv+3T2rlkx6zb6RHQFKC10j1
E3DZr5UyLEueiQRO8jErx1zgZuhhBwsxCfEAuXh+DcPA+PrOXq8kkpxklT8J7pTsbNgyIXVnDxTL
rLzBo+A7oBWWVp0rrGojTFxybxUdLoQ2BEVMMwuBLJkEVm8J8hDjM/tXhU3+6CPpc9iQcmhF1HfC
7i2PQksof8ikwm0VQBn7JDhn1oPitB5283qS53Jun9ahrQStOWtKvQ7yRdRGVAZx1CFtFApU9JZ1
qgbnD7brXuRitNBYayrQA5+jJgHd68RGGhBr5JCvTy5W8/eIdCiHbHuWDFZYKPNNvFkeJCsXLHHl
puqoQjUOwStS+J5SXrggJFlMsZjvzg+n8ftR3Y7Fn6jZiTWByHRF2K6ZSndxBaYYsluk09Qqb2zM
bPkVTdjS20D1XDCdBSU3ekzomJwsT2mdcfaUMIEI+YaQ/xENkPbhWI5GGO4fCZCYcFt4tNaQen2a
JDIJ6fWP2G9NsOh9MSwy0Alu9DdSkeaQGTVPHT8Cf8RGdLkSWFirDKaRKkBjWjhg2EHfD5XvLjM9
R1qzp96w35qIIxbrvb9N6C6j2l7WFT5woRwOOp/WIMbJNOgyOKD/YeWpf18mL/WYn0UZfSjPqbUl
efR0RNo6x5p8hu9q1K6SFX67xwlfnfoemgPTlnKUivZmTdjqgILLo9gjytj3FndMduqRcb++ZqMe
xMhLI3hqPLnDVEVUTVnGSlRE+VJBvbMJY0plJCqKQnbPkHCfL1rXX8z3oUla1koyZnbqvFw+lTbN
pMrYfHhQgsH/7TO1Nd9oFVlH+xWoTN5PEawBjLhHX1b1B/FbO1xqhH/0iJLUy/bWVJguYaXW6Ixf
d5zQmLoyf8Tg5YajyhtmlEzZ5MqbvprCiHv+V/3T691NHlcw7vJlVXZXfiEtU0C1akClDNqmhNoK
A6S+f3K/PtrDuC3MEigw5irzeH9rsDBcs+5g/2TjVsEFWIty40lxJQ4TZnA8XUiXm1TWTR16CfSP
gsiUspZabKE557N+zOHJMa9nxb06Ld00MECsrppVQWY6uykpnqjs983vWZs7T7EnKiJJVyghKHqn
DmJYj77frLozOtnPRSSl4kZohLuAlJg5nijRJumExaUZdbIzviDC3ef1yRzPEs5DfL1mbqUS1Yau
9KbTSCt0Cb4tdJ5u10onfQNqGhkTEOdjmBMUg3q0+TqosVtGQW4R5OoSPs2Vpx+1qjqwU+qWwZQY
dB0Nt9leUOccWRP/Kz1pXFtNQ6h0bXeLEAWL+NCfM83xaES20BCOC0QAoVguay4OON7REo/t0ISi
fPCnwcb55boMyZw2kc34aiKGBQOcicrCizCTDRyXBb17TNABkdH4QZcwMPHKYd99nfTG7Wcbszug
C15K6qt/bHXW3CLf2NyNGA+BpuPrS9uV0yCGXTg0D5DI/nQMS7tr/wFFzWncD5+c847DVtSULYHj
TEtvNMwBVSmkNmlRZDGI91vY8m9WWHtpzpctVwOj9p3qXIq2Rh76Zcmngl0eVQ3kwd+7hBVl06Ge
k5hh63OWOxBE6pem1qft6/92jvyDgxeOeJK9n6qWmY7zulIU6ACsFulHjLD+urNT+2WYrBeuwfsn
mASJqm1nEO+odOeJPeAkqBF4UTtfHwFnbHhqtGxsqkJQwW+WtJl8CRmwmH5ofJ2h0+wGiAFnSWd/
zLVqFNDIretCQ2JsbMeRWonxFzON+CJmz4hGodfD+9vtWBvtQdLB3GCk8rfiM4NZJoD0kM79PM1g
HxdowF7p53z2TA1KumdDKGWtdzFrofmVrIy6NWvsmk+19FxQ1btYbdGmuUWJnG01fKZqnepKWGUe
PQLHUvh0oCJkjSuw2F3Y4ElI229hcN15qyuQ9gZYM6Yw3o8IEU/UNMtxCDKgizwDE2ofuGKaxhPw
BA1UG9DXJ7m33WT9gfJEm/dfs3zT2qoBYKg9aY0YOYd6cT8d6+q8DseS+GEx8TUOTRrvIAd3Tjx4
pTw8WyVh/pErjxaJ5KodcU0Oj2KaZsWYlqAILbT+ZFeJtRjjT5mkzn1pO5QiNDxvJyaxm+f8heEs
R9eYAp9vC5YUruKsJta60kDIG+e9a8ep6OsjiJgIGHEuXyA8pA2Wgpf1lRrRnZ3QnmVaT5TJEoWz
jQTvYSsfNBgHz3k8E+EytZsoExrE2vWhss0qY7vmIH2dSBE/0zIu92kLF7zeQdUmBMJ0RWvMC7gu
E5MW2ci8PIqktYHXH2V+NOeEd5I/eoTqP0w5O7UO+MkkzS0oBEv76sf/QQ94hifyXjMBe8lj/XXW
mSAnIcvVDz3NT7hHdy6igmU2eI+o4Tc/YBgMVpZDwa5WhrW7kkWO1P/0AP2zwt1cNR78Avyz5Ojw
zHNMHB4eIzoZw9fgY1r0pBYxhILJ3L6RoGv/c5t6+H2g1g2Waqwge8vVo64GAM7C7BbH/fF3xuEJ
vRcKK/OiDS+pBm5KIhcE1OeykpZgn1j08LEA0nGzQi4Q5W/Hdy8dkGWiMlz1dCq0qfTJ01vRjdoi
107NIPOS56Jz7oS8EumGheporrOctEe+VWza+eGoXv+SAhRd2IVENPjL0iUAJ/pUAgwPQ9FbCJGt
6vL7Tt5079Gs6SudSbtgrvNdjJA5VPBqJjyMtENxpLgJjbusTaxeKTxtU5RxzCSq/MTy9ohBfaUt
XDXLV0MG7iCQUYPtOGLigfCSelmpWhY3dHwaRWEsP1A2UWkv/P57lRvx1A94fuA1TR2maWgMkQ99
fEeKaF30W6sPgdkr7RS/zRTLXdwehleEf1/yFHBNLdsCf3XbgMf9YUtgOGstV1ZpO1lkm881KFC8
A8C4o2PNg+bBbwe34bu5HEZbzVNmAWcP0XK24pGw2jUMSJ1lxKFu98o5t5IixhI0GFpPJDJAMFr2
I0pjnikLDL4IQpLcWhV1i6Mz9EFyV75+pcw086Q+bz/Yynqg0EJtxTQShPbRJExW6V3vUZSd3qD/
muvQVPdDg0I0pszGrZAiEjhlzJj3kWLf8CUF8OQzkKf09Lqd3oyOOypBfj7LWpsAS2QOxb8EBXcA
EvaY/dlm28HTtLLE5PV/KlzLYx91XyLkDFLWCzbDd5QFBWeJIn013GUsgg7pRKd4gu+buu3DivQu
mTHV5ZWj0+eo7NlqW7oDy+jp7caXB64wvrMy9o9ROuobX6GvfOUSiqjQtzKT1YMGta5QeqH3Yp8q
Z9kVKDDiTVVNMfbWua7JZ9277P0nfsdJFoBUIj8qjSKqyj7s1qClmbaMStnZRlRc5fbzwiNjH/HV
gU7to9MYzVOqJsGCusJOCzTsFVR9ZDI958W3caN6QYFuA2Dc6Yaibw8vgYmjE5C0lOeOWhGjMw+4
bW0yaBvWVKSXfOzQWWXD5B/KEpOWxcG9b/rEbjIe9j8tqz2ZV83zWVVyPjvY40cC4b9eFDichGMU
K8a9n6rFZAk0Zq7m/rbDthyMdpPTp94ZbZcyUQt5QW6wao2NiqIRCle/jlMJf9/HrYSmDHxkn2AH
R7O5ZIu+V/yCfAx/D9ehSQstpVLG5+SqZlw/TcxpFoDaL84su13Z5vEQK27cV5ZNW1HhbHeqDFLJ
di0cA8q+E0pWIVsz1tyKgTA9YDKRJy7+kKIlkvH/apKSQSrDTG+rBoTOtvQ9VRd+Icf/wYI5QYU3
YgE7lurvbu+YbT4r+gM4TZgbQibmILaKSia5XHBdtEDiPQSgPT0GGMfs1BWYxHu1db+4k9U3Zqf6
hyjFto4NNVtPfmRRPxkHd2Slu+ptuQ5ACSU534/NdEIXHE+gLDAYHDdne0cpwIBRs6w3tt/4p/sE
GN0dEpXG0qP21KJu12Hks25JstVF2N6ffyhNGU1JRhPl/u8kUeyNPmQNlrJsUK8/zm0EyBkBF1V+
NwSFbJRVASs6L3FQnLJU+21Zm0noOWipeo8dYH/LPPElk+1+k4pJu4kt7yfdWShsUum56IPayLYn
7DAgD1HD5isvyaKQU84d+sRDSow6pP2q8HBnd+5wwCwiaOVUhG+cqsKA/NqX/QEM+3g+1Wu/2MnF
7D4EU3LzT4FuIPqYY05A5MoQ2viSlryg9iVkHNpAJTwieWNgoVSvFjUPEALszBT4+LSkcDDPO0Ow
0Sq2lBoFAVXZOFI6nfhuvHWudlDWZkGJc5LkbZ6c89ubBr+dVRqnrJjNWoA5kI3DK2ycNH8Yyiap
zrcOf0iSU2X4uD6+4IrlfI/pNvQgtjWOmSHWWRtKM6iWXiMCs7tiYoD3uKgpomk1zBRQQOWlNuV1
HR5w7drVnrMFxlzeyrG1xZde5yi35jwEE2rbtn71+OZG3IolCLNQ9gU2oFdpaGYCfx10UBQhP/7s
6fnG9DEJJOO4cz7sqTiMINEo/mRfEKlOl76EsKuDNlO4qoz2ucXjREX+Hdd2ua/bci3JRvbYCz+E
NUf2VlKbUShvL5YUkif4Oy7SdXWGSqQKnZ7spOvKcfzfHDSOBFipagyDoXFNbS5njovmfjKYFTTm
IrReJLXHsz1Cpryi/YMVRsSpNtRLhQ4BrY0RN39zeHwOLMENzT/DFUacNWMYCVf5pXaNyy4UE7Xl
LVj4XgwMzKAivTr9dItGe9TAjEjxZlxaG4JNFwlRGVmFGNjndDPd1lgJO+w8bJW5ovbToErO6Ay7
Qgwt6soIGUgvNbDy4HuIBWbk4ujsiNYMKXTPCPgaMbKzHDLUgmRDZP4cVCEQvXXkDvx/XNSKBT1r
NvemTJCD/RtP9A4C2i2lP5z2FZuGU/JhUfHcpaOaUlFykCl+KnXTMNytDIQ8eND4J2RJaC1g4hnW
pg/Y9Z3ZhVQe8b4xSu3HhaDJltNOyTl3Ocb1znQJXUQFqKoqjG15hzK064t62+g9F/uBvAfgIV4N
LdaCqibFk4yHJlTWyLqU08Cdl2ftPurFpZxfgv7C6UbuVE+GNqpuFFxREfC/0aQW53wTVYLjSg8L
WywL8TPg1EsKuZAfSMl3dN2vZVfXfEGg2/dgrpbv+Dvrz28mQ08RxSPbQEnJDRkAhcCX1NPtLJhe
6cZXnqV84RnAGPsGAFzUtIcvLL4ZwBWnKva2TO3SY0rSYg0rZJBXf61iX/kLQHa38mXTQ+vF9Jvg
veXrbB4Ku7gZR16P+TuXZn/LgxzsxJm5f5tCV3LYkQ0McGw0x4XkDVqlBlA9hAj+nLp30cFIDFBN
3NszKPIIJbomJDeH0halyDVjYIdmGB3zuvHVbQuUIAkvZymeKGgo1tYLIJ37sWv1bqW8BOeZL8SK
1Bdnzrz7RsDHk49sG1L2NG8gb47SF6T1WYjA31fB95oYsuZyOkbxiP4CMBmAcnE+wtNb3zpwMAsn
XG8D8RCOGBpTBiPFsOtcawb031GAYxeLW6DFejrjqlp6GGO6vHmn0QMXchz97JeU+RPOnFsuMxxv
8VX4V+z8YuccTYbV6PB2GoQ4FSwO2wtLnL3xcErHogzLCUCfcvCtssjPY0STj7wSRyjsLwuzyPgy
sa9pdc5dfxV9ERtoLwBh1RQHiB9iYoBrxU9Z+I1j7jZO7EicpKylfFXRDikk8CFZ3FniLJcK4Lvh
zZxACi9ZiqKBX8u+F5kFcFkygKgGVYiFrN39qrYJxw5dHiRA/0g4XQgTjDaG205sxEFbZTHFJO2v
CtuaBSrbsaoh18qiK/sqHXqtr5RgZIjTOq+snq0fQpgCcwbnsXef4+us4Pb8HoTRBamb2pDY1Tj1
9uBdFSgqV+R/omZMRNp4HXHfuzR3qKImJApFOclEG+9KiUuOk4elTDFrms9d8g0YfYm+geEXTcsR
/BzR01MCoivzvbIOR7Rnd5ezFf0VufvZyZ9/3WmRNtXIdV3gig1QDhBOzp5yUUqcJp/TkWneURvC
La/m2WBz0kJMYW90r3Mrgoxd+c4oXMiHZF5JV1bPsmWSHdtsOFiENbsjbPl0SD+pvBbelOyfsaor
tV3Hc9GoiBDO9Ve2+P8Y5HU4p/LEXzxxpDMffA6UPOoVSk1kD00nLq4gGCmluE7TInn9rpui39Op
6OyKydZsyyC1EX6L/IOfqKAEXgFhdGtfdGFh6620SstEqjpBf0JyDfrja8bn9ZwYGbgV5k70hG9u
osRVaN+zCbosc/TqTnxYNk+jKmBgilNsCpupC3LimyNbsI5RqpIIHssMzGtALRIkvMpWOqvCwnzb
2imXhJuEv4J8KARS1+tzjQqE0m/3WQuPFGHFQlWbrCSMfXfhgDg9rFfNG2qkWVVBqnH1KbiocUTG
NNnl5A/P2z+R3Jh8qb/X5ld0FqyzB2qiHTYCzleQ+1fGpdgAXcsbJ+coILMprtMkV0ydf/4m9vbE
lX/vk7ztE2JlFQR0ttLt2pxGenGq7tvKOGS/c3zMae+Rc32w98xYy/o9hOF/SPeDcoJfVIoWFZL7
ICDidYjZf0I3Np6bkYl6MMGsnBalLK+4NAdfsbCIpHbhAQIJTX8apKrSgLhhmCJdLFHwUb3lf1Td
qIFP4Er6Myj3rQC5LZCAvnMEfvIkJPI/tiwC7n/WkDjkOUtKPWskDM9tW25r9Hp7j2pKIyBbbv4g
FTTP6jo7ZiGxwwz1611ZpkINT05ZOUJsybu+WW1Fk4RYC2c9BYK06Zcg+CdSQ8mril1IwrWVySQG
OFxRrufA/9Wc951AF5VigiCiSnWd3oT/oljvei+0sZsVNYkpF29HDSg1hC9iGj4U8ywDq4H+dX3x
ZCnXL1yHQUGJy5PwO10KMzrXIlqMMs+91R2IkuUsANC1GqMpfkzzvr8XnxqtB/Ij29KupLjRZrv9
AY3+xrXA1WK6eXyK7DPEDULpzUDQ7NGYPC+lwqKr6u5eICpW6aNALFOqSkPMR5mpSipdubDP4cNE
JttatL5PM85m7LwruoeRZ+LQoRqP7Udz4aIIxe/ygDbP9AMkxl5DSZZV4zAjkLyuCZG6rEJn0gUf
mARELc8lklyLTzhccYuEgRlpiZ/CbhpNBoY60dxxZsOH6apO6i6QcESyORyyKWvnrGv+JjfPj/38
xeE8jVY0nk3z0+vJPtSHV1f6NUjaOQgT87Gb+1grLg3UdU3IrobcquXUqLpMAfj5qKuf0t7Jg0j/
Jkb1cYagyqzjHMfg9hyKpE4NSLdCEbuPruI9Lpw5X9URlKRbaQEtxRfkblpeBMoeg9GQa4upmld1
qAGuZyuKXlET7qlue6JwRVJuM5wHFMQWDlTqysr9sLpoPchTpUhC2a4Dz6forXf3Ps6mZSFJbJjp
P2tTwuT+U3XbT9TjuYZcGLIozTFNCEXdfEdAlxfkWbN65T0VCWxXVlaR07MQoDdAW7tgvUAfrRxG
ZaXu35VLxLFINQiagY3YzThe8ZIAOaHmSDB4uABo+K9oP8/ByPaXtnxS/1JveCCKRLQWiRExrNG0
eHmsXBocZCUTTueRgjVt9aOnfjOxLseBDOgBgqq2leoGDEa6vr76X0Cw6bKzm78Qq28tHIgRZXYq
ld1eFRp5/H127o2KpbKUHB+AQOTDaQc9aFKLH5ctp0jlel73QNCes7NJeqZryWLJvHiHnmZy3HaJ
TqdXBKQ/+Reopw0hNecTLkQZ+oCq/41J1iRcJJUn305CPQLHtD/Ktx3UkBSLhvaCP3h3O0Id7Sgx
f4ZeIEZyzRE/5L9R0TseLhhn27DMmL0kZUO8rMK44OlFsZa9iCVONcfBuNIvxcL8x5zaorXQnZUz
3pFtx4JEo1dUJkQJ46YUXmk1z5rmQ/d93bh7dZEhn0ecGlxRVJIlfC93q+wbB+hpduqTy+GhEmPk
7qQYryiEc7q6i0ZR6J1rbg8SNU/WxC1yIHeM5uPqEqu4sNrg0NXPCJDm+nxGXyBrinspijgF0ls4
Lek/LWuzQNfOGe+XzCkC0lBMve62i5goocJcduyzN2P6DLZBugVJAWWq7lIB9eKc4fDYc2ZCvgPO
eYaHmX7fEetORX4D0mnm18S89NA6Hu5QQZrF29gvLL70biZm4EuzoITbhM26atpMGAuQqQVydI0e
9eWUIn80X0P9h4rDjIGXEDqqdV88h2d8AR+2n2HGJAIJyLkantaJnbEFjCndNifiO0pDV2Ax32F+
K790TNdPv6fq6mFGJcMScHy5s3RntO3QSX6ASfZBCK75aezKDWTGuIp+PUl6IAxzs7hnPLmrC6iT
MDvmDPSxrKFWRHi/C+UULkJ8+6t4O4eQtRhTiPI9Cn29MHihJf+EGpsrDNMxNaqCzQeYEMwMmIvz
KYVRjvQd7Ob9ul+BaDD18Qa5w5hCvU4n/snxjSqYztC0gM9cYNBfDRvcq31j6CSBOxz5Mffc7yr8
hks/jbWxdQnQamAkgkXhX4YY7urzcaEO3Ktb5sqdd7OHRK4ylS4FiX7BPOzKN9KONA8z/CvaJWib
nZ8pFtsr2Woq1yBrVcBwuOYDg8QmodWjH+FF6gajmUz6Y4KXZPAr3pr1W9l2kNl4COdYS95Wnqjq
6t3L0zeWgWOKv8aXBkcecq7VDNXTqg6HlH0ulfEbI4LN04Vcwr+WGJsKSnMX+ST5YrO6mULrWKOX
wGh3qkCG2DvLm7zvEuK+fE+aZb+YJMM2aXTxfPhKT6x7/UIb3xFGAlX94+fF8Rp9BGsabiDdvW35
639PfWroNjUQy/O+mVnD4b9O1tuRrUgG3IYyNBlHLEzIb26q0gS1da9m3lxOyQf9ECVN2ssO5slf
2e1vr5WMoOtzeZk+YCGooYslytSAYnoxu0SBdfvjjs+WbP5OFZ17f9WUTlAG7NILxWK0Qth+UQO6
o2W5QOn5kCfBruQCrMt3rYvDjzA993+4MGRzjD3x/CiTLYHM+GEbUAA9VPwNRYBagLta2Gm4wOTd
+W2oDram1XDUg/JN1kdiivtMbfzHk3VxIpYLNHChOC7JtiiF9u0cuBnjsJVfaYpvRlWSBYMKRwx2
yENI29qXk3K7q7zsIKbSi/344RACacHpyBNVzDz96MPFO1dCqBoVyYkvIYftctFzw5VNWn8+76Z/
5AdNjjz6jJrugPf/8Woj4ac1aFC0dH/3oRXGlmnH9Rf8IP99ZRKUI+hENixvIwlKgDdf3w7tnkFt
xkfRRluML3Htkae/B88DEoo/1K5C7wpD/TxsVE4rhp8hiGAXmMKVi02tpQMnXPyWiSZzijaCsMGa
0N3C2NHd7z4auvRBxbIUgdmhowOvBGARw8nGCrMGYuKWZLtAQGmDFqI/D8hASVJmNCQhkl7nLjyS
Aq4xX+w6UzBSSQ+/ERObgvbx9eYZV6/pRv9vhd56RdSlWIYMgO/bBvVRZtfdBOiF+2DN2Xex5lg+
BcnBD5mzxQpl8n79/sVeSpoyx4dO1GS1ArKhPmILoEltY2HTx89sv2kMbK75djMQMOIfdME2hgn2
gdstC5SLg2ZWpu0191DVxET1Zy+h2v6QhckF0NoK+FiKT1m/bPBVRaO6l5x39PpZVNN6FRr2oPym
3h9k3uimwOTLhtTXwUpwS9CknYt/ghkugQD0QK8oGYhv0NWjzGGAEoThiK5zii3sYudrCzJQ9nHX
mN63+5v4IKBQeztOlFraHJOJ40TJ4VgmMuIzODU+aNHw/7U5BHdKvwStN4KJHFAk4AcZ9L+A7lDW
uV9HfdCI5N5mkQXATy7BrDWNIUsrioNqBYt8iQOOKsrimmYPZXhfiaoOqQ83xifPW5NUtwfZjc+x
x3bf/cjev++CghAD2eDKZYUkwxufDnT8AcxoZK0pNWbIaKveGQtNZqdwFVaWqjARx4USfWD9UF0T
+2MgloMpu20h7aRgEwzV9oTQbROEqDQrABvd12ESis4fuEHmptDA+Na2PpHuWxFdscH8dhxvITQ0
fW78CPzcdO90xd33j61xqzrZw7g5ftXxG3fz+XZEtMDHcECpilssOjZFL6C2oPAnuPTPvqbnpVzM
gaD4viC+jgWPY4SWpmL9QbCwHVzaQIrd4vsZ8Mvl7J1DfCMqvW5949oZU3CTONaHKOh2ejgUhoVw
720RVbDDcEejVDyD0Q1oPdvBosfzpmYK8VgE43nyZXUm29f07A0ZNo7nvEOyZbDttYAod73wRpu6
/JsYCkEhkKbGIz1Yu+vc2/qV16nvdr/NuGEP5/6wcRPcqkRXEAob74GcnQCvfIURcxhdPd/IIrBO
apgaabUKyUCgNpH8jlVouCwwxqPu4VPqUqTLSKiYoVp60gvXRP2xCz70s/fkd3rzRrZxjkdKwLXT
k7v49H3P+QzFQAhLDW1VVkrEVtd5yXQs0Ui/3bQjS2xRHdGgIWDGNgdJdOgZrVBUqxXsoxn4jmqw
eXQQkqLaWRMCItzA+cHYPSlP7X8zSmu982qGzo3z/U4U5SwbCsrCmrTps/eV5UpAjF1OIVwa+eQg
80IHfzTLsCVRSakyJl/vfGPbaccdOT4x0YpHkhbO47bxbz90u8pI8sZIN/bVPV2rNx+54bKSCXSE
GfHCoMjSAwEO/+Ot3QYWuwes6S/5YmFdeehZotxyHYxa+Q8ZI805VSUOTiQyLFDh18PkzKzxwMiH
XCgofcsfuVHUY2VfZH4ORLE3mV7ui4Bgf3sT/goNXFfBQgWRkCLFSkCUtmpDXp5LRf3/O7DW5LE+
fvSVYY4326biFe+cZp0LSYRIJ1XKvfndiLN/jRvIAp1k2R4HULNJeUxxpNjkoGfZdjulderPVteO
4NuLTQq4eF2Wq4oQH0/kIqRmcP3q89waddDlUjeN324FkCGUPbHk8apYJxWHl/t+v8OtYYaQMH8L
ebnYNT5NBmuJJfb+PCH+6qqjlslHMi1sQ2/1mldqRS2eni8qXuQyoGy9W703xfxMHgYPmEC/HU2Y
ITymeWKudwZX2DTFIOTTkwb/BicPCJalnrm6gbFgsNu/bVvG56d98xXiHZe+S9ICHg+w/3/ojFNT
xQEyO6wbSeWYJgRajpGQt+IQWwqyQqiUdx1tfnPQbCMySMOzC6Bx+WSCKu5TPEw+mgykkFTj5x6q
gLCwACmIQQJSe9cWjQGfWc7S8riDMi6SOeZ2iFebxTIobDgkyPXxenir+ccbBTkm+Fi4Iy2oGa34
p7BiVibJ6ORX5Bf8ZjE9C2v2vvAuhLK6FwLFmQBI6farjHDMXgdosswRyYDfHVidpcH5/FfgJN9k
r6KxleBCMl2bDgp74miYEPbmkltp2Hi34G/sUcG3ozw4b92MOiTxTv1izFucDkRfbWmAGiY6Xdeg
gGd7y33YnsDVDe8+GBhapx09+wjg9jBxCYJcNUhD3aS52fQAJG4rL1kDF/jKXvYHAK+3udrxLdo2
GrwZJTRuXLse367oKiGPKZixiIpvXpj/aSZZl5qIHzccZkKYAx85TZmEbW75Y3YtrlyW5UjkF2e2
h4AHEeuFnje97jY+deYZEqtgU3l9yEovQmmpFJVnx22r+hLzBqP1xjg5qGc10ixwKDi9tErIrPm7
7G8cprhymfC1ewH4DXn38SDRSFGo5uL79i+hn5rW60jr2hHyOPaycvmJ1E4bVruPO+xcI0iGJoW2
b8Janehw0i9zSWDnu0ZHruwcEfocZrwv3ZVJhvFdTnliRnUKqs4uS9X6wtJQ4XBMnHYB26S853uf
XX4wn488B56g91KWzVwhR7o8PuliSLWLGlEuM1xdAmTrYp+hyhiGY3pNIIVZevz8yP+WIx/tcA5u
Cc0VRWHDLCThCabee9PhVGZWa3R0Mjsg4rqLq+uLyo+QZHAgenCwdDQXVlazzV5C2CUjL/Z+dnBf
ITLQREc79uiDPBztBAyJJS8qFLdTs7rhjKp1srqW1bGyBdeEg0nrAOyHlAjsnrx3SklJAQ+1yriO
kwVEoWLT3AyUMNHXzDeNi140wkHTa2uaWT0Dv639gF5W1XTst+yiqWuCoveYdOlKMxTBr5aX/0NA
ZLMIJ4qENOxIT4sLa6r1Gn7ayLI3rGFCGCuBG6FhbDXTcRTypOiTgvwPAaauPRmJeQ5r1e4HafCF
L8lnrjDQCDes9UfKUE/Xn/L6WnaX0UaK4O5/nPs5dFhvX6C4jreMmiQwCOqDZnisQeQF1OQYOPsn
im0eql6teM4h968a4/6fn+4vP3P7IjhqhtpHFm1LrLY92iEdsRzr1rJeOyRzcR0SWnDLvRajASOX
xBL3WJhYc8Wlrj4izITyxABI6sIzkLcYqDBQNERPkFry1A4TOl8b9gOWYgDTMrxBlVB4nWgBhIyc
heQFXMKSSov+ivMLUNNRMBj4P8FXRHmYdbQnsin/L3T2MS+Aj22G243SfgHjuKVL7dlI5ZyFDNwA
+3Ec7INGMAXBFZi9ddeMsxLZjEEl2PEumSvLdLcQ8kUlIn40Rl7Ck0Q+PQU/yRGJnB5lPgYq9F0b
HJ2P0wQPFb+6kwDLvUM13uled0WNd9jPW+wMTCpDWYnTCsnYWGj7XFUX+XlOtwheB/gbFonJuQfF
HBITvyx52wXYe4O41KvdFd4chaLAhrSD7xa8ApVWl3l2sNkQf86Ik8eN6tbFlqC76tlmLrddZ8Ry
yN5lrgiL6BzkFuzbf+zGgmeo4iQysW3ALP18R9aXT50fy7AAGtO19cyjHOXylzswJtHT7s7/YqTq
3OFQ2n+a83jfjht33EzitRy4OSYvu2CYf8ctN1grMqF9Gkul41/T0+Q23/sqFoa0uF3oF238S9O9
lJPRezj+cBgbNVomyqwmZzz0tZEPR5H2gnEERljFwPFFHN/nlf4lFiA08xizfUEULS8saxXYb6R7
twKW1+7AMkUynoC3/dT8hm49Bj8YKl8CVppTNCvCZuZ6+wX2pb3TMvKggxzGkheXnw+FNZaOeVRT
3SgqXkDHvXinl7u3CXhPPQR37ZPXRCAh7VgMSvV1nFyedE0TBHXGGBZwz2nci8+pwa4PaQochxzK
vOl3jvcS8OtF/4/n8QlELycJrQRcapXUUtP9tFHSe+rotDPVe7T/v+OkoocsfSjSRuCY3T0jzkX9
wHncu9XB1tQJMKNJUJKyrw/ypFrpNMgFIA997e3qOX8yc9OugXQIhcoqRQqbUm672G9WTeEcqpmb
ijUX3svoRKUZy/TkTZy2lrV7FNMY/WHAoznGOV5z7ctFGCCiyMVZVeKAAp01WSbKB4p8KGr4xfud
vwzzXRUZiCmzL4elgyiXkaFm2AgMVp7m9qRMCFiAf54Rtoxfhcaxa8oiON+4II8HvP8AJAcRm4n5
KzqWnFNDtLp0NO3UHj7PXXgXJR5n48RVa23g0pFGOACCt3jvW0cbGhYxSQvRAQ03is0h1G7ykK3l
n/Zw1jwEEmqS1m38uWdEn1lYXGQzP0HL+vhJm5MooG2e5b4RfAsyVCemNYf+6nU57rz/wIWNqUya
yiMFmRNOs6mzy6Uhn+aJHjmMIAnKeeJscPsmkCxD8B2Ncdjv/UurUecb6Za/idAxUufzyWiRfURd
urPLn/PVgUi3CMJvRhNDZtsB/7cTaRV6a1On51v7Za59l0T//mxOmajp1WFGrgyRa7YZRv3P76B1
fQmcumpT5WLKcCFgKs1hU66LPaKQMORuGUkVKyACWwI3kQ87en5xquk1I6kdHzSWgk7e2LkNfRKW
MXEkNF6ydFU/Bnk0/PcZ+oODcCq2FruVN6vdnPpzSYjwouw+Lh3FpCxNuYIOWRXAtx8NBvG8bDKw
zdMEWIbNxBmI2rxy4HBcAFhD/QOriOrckfeZdv1dcmdpRjAPnWn13idhO1CaZ6LxPbhgO/Q+QV8a
bEDNrwizWSnqDdfmI04jwzn6um4yUmiCPPKF/S31PgAhdxEPNIbtoTNitwhmk5scrGfv0yUMPtF/
z9GrmdmJ3iv19w356EgWsVehBoKjxYmoDKe58j/t6uvZLHRgjaQI+vRpdYwbXhlPuXVdNHvWSl7r
0OwuE1itC/fUGhfGLwgVRm2ymFe+qj0sbUf2IgP8z6OPgkT2BXoQ2yHyVHQb+MtAhya1Tl1LfJh4
TLUnt8C+Oe1aczCx09qVdhdA1mUe9IDGRW68pwz0QshttDW4+mKB56XRp6dPxh4cX3l4gpCG7Dwh
W4HDpdCkc+p+G3WDzSsMLpAKHyLYd2mpHAOKFaXanll9/5PfdR5Q1v/Vgk4BJbAoLbRbpB5BWlnH
LLZJq8hWHddFh8h/UBGOrS9uu0lg8zjNRibgsZRHMQAvQBd0zxJjOY6vf6203ViLSgUAkTUAxAFV
eYHvF42LL1bnaJBalXzvrqnbZ1hQpZFRCswI55ADDt7+Ygx8J1MArkmLBplu6IA52tSsM8CpK40X
PdjovwUwfEDUAV9uK4y/5cnPFzsEybvPX0lRYc8MySpBI5JUHd7lUIMbPpdYvUhfHag1SxeF3KTu
+eXKh9o7+aby7lMrT6UsTiwslYTq31cMldHu2nUzh4s3hpeUnFrYjzju5z1Cf2/3Z79ixOjs2ryq
QGKpB8aWBM/64uTgTHka+ospJLdweH5NpPfmHwaxJv4qt3+OOrvxA6o2+TYnIPBt9pPt5cYv8kfb
Vz1fCLbRRG272B/w0k/oyUyccQ8WddCRmsRRhGk6pPnFraZzikfa4ZEsF4soJIioPK/z2S/rHu9i
MuEzz0t/Bc6Jk8fGayTwkJd01C8hvCHcAUgXVvRwUgezMKQTtolGRbaj4YFMpM81ghMnAubAjf3r
PhNWczsKjB6fSuBklkG6pC7+pagU9a0o9mAkP9NxFwPwBxq2PVxhIz+sc2LBjQJi2DvCCuVwOo3T
p8SOzm+rSDCsuNDxdBiBNoBwjUtxtvyOY9ibGDE9Vc6CjXEqNdqHpgcIgDd05+kne9E2OfElf+gD
cDwFboh/oksL74Ra/cboz1Ky8cyP5J4Ib0SoeNaz7X3Tj+BvXTTyJTx222PvfZImAc4yUC9JUZLs
lkV9YA3LXPxD673W/EfDKdJMMooZu1v5RmDR4emeJYFBMdZtDmQY38SIgx8woXHOSbXQUbD8e67q
a/sX4wubBOCt3z2+QOpHW/dyru7ZJBTIUQaWqBMsrHft7WuJKy34QPCp1GReTcAvG9+woZIOVfqc
OfHuUJZ9mIYoSWQ1M1yxxv6fCqKwzsB4LEOzw/OZPEwSQT8Z+nvzPSe2YMTmVyCIA6qfollZY1Ga
dIDxKZV3oMZRmyrEge7TmPhGu9Eu3UH1O1dMTZZGpuNfFPVBjzULoX8FavLq08wDcc/uczkrETDa
Ac6O/6n6yxXTkFTpipsGWwfMkmi3mBME6N/r/CuyeyANp7xBcTOOyNJy5auSEZ7z00eXV77tgK76
YKrRcHRysGn5a/v3XpSBapBq7M/Ft68NIpXZkg1rxR010TKc0kIlanqqkXc6hfKAxaF+1ITpKfK+
SrB/BaPyI/odELLTCDs4zVPi07u3ZMpRkCat5H5iGt0/LcjSWq+SwNgG/+Lb8f/5f9C2ziJ6iuKv
8TXQ7trpC5VmycNFuetemNA0hLXHFoXUj+7qe7c+lGMDNlopUzZkDmDaEHPeGGHe1/6uINiFsEBw
qfM/F0wEksbEUIIhi6erKJXXWCehjFMMOtl6/s3MuEClpZZ/n/jAUnj0/vmA5qiN6CMK33KzpDwx
k1HEZTRtIda+Z22D24bgyn1FVGjJ7k7rzhqQYG8yakW/9djK/5vPZ88ELYac1zjWGtf5QW6wRm2g
SKkVrtavB8yAi8kKEsJfnzez+PO4ntXywvsyucWFTbVLccTKY3zON5M8RXAdFhfcXfFp5mkrvURO
20dh8CiwyXyESevw/YJORimtLvTRBniaTHB6VEwqHaZ6cY9Ud1BvBTEIB4KQPI6vtKCvLP/60Bfc
r0ueEZqzqnJyxIYiLLCZAig70+S79dT9LsCO7C6sFTReVD5zg7fACj0/7BGQFPH4xfxurNB+XcAF
Whe80a05G4OHZa37u3GNJXPlvUNz9U0bAwqVQ0ToIWPeggGaPT8fLY1mGULpwmfHZ0Zb9f+FCPL8
l4agi79V8b+mKEsHVoS6mW8rWebipZCh8Yyqbvg712DZc66uOlDcSLYbqLIOhpjOfrtGKvSxjQMT
vAp5P/JDiEgqXxNTtqCtPebsyXghynX7ph9SryKwClgKi1DEtYto97oDHERf6BXtbjaQt/LJPk+9
yBK22kijNrtNib68eOTT3lfLPfFpgFhRVYC3mz8kfZSIZif2sDXqWzvHBCnwOgR99iyEydlv80a2
1W+JdrgbZXqyIBo11a99LBTocEIv/uPVCj9ng5uXSbti5XL8bg3fSzvC9laep2PzAyJFlm9qKZZi
tcfZcOVgvm5Azi4fn6vtpOHnAkflZ9XIJHXQdjhHsnYs556r9i1IwfII9eehm5WAYCBtb6rndTr4
+r49DKQyCMz76A7zqz3SEnx/c/HsWhPrMOX3TR5D0X+gbSZFu+zaOSxFDNujQAlhUmycJz290jgo
GcplNyUaA5lR49UPmAhhlufJxagpnVq4t0nHihw7Jfqcs3qBmhOjUz9Tf12cHfMo2xl+IeYc20KQ
Vn4F93rcl7WFMdy16lLO0OFEVwhNKYK7VaERds5MHbdrQQZaEjnA7mvC8IAZOIcpMhlkSwommVkC
YDNR8BpRh6WyybwcZBpKC8zasbJ7RJHg+CCMycoSFvkSXfmBxWZ+nRnFN4Dc4Vb2OPas0eCcBUto
M11MTK+VV0nBm9FS6huFlL/Hj+7SqQpcC+3Xw1EOLkK0goE12uvwbiVWgZdG4qTT81WtCHscUyIH
KVnDF8JxH76R7FAu9WqjXp2Sv6vSy+529vIZ4yV5sLI+A1I8rT5TGO/kXo9yQEBU92+2KoQXqSUL
I4rcz/L/g7JsQgjHRWYkkw8ZGxqY7/Zo/398L5aX/cCI1TgFzBIpxirRUFGXbfhq9MZyyLWtF+S1
OkeKyBDK61StT4OflHh9G7avua8RoY9+DSB7GwXESYZZzU4MWir+rLK353pR4k1xvC0ooAhcXlUX
+MeQsJUesGvZSY2BlYw7dxQXII/Wp5zzgPGuE6vlIUAFa5YnxfG9ktXzUciiq2NWccB+G4hbhiE2
2K4BMN6nhy/UUv1aH3req/zNi2HbfSD3DydZxPgmpC4xS7SbQ5ibHlMSFLoEt5KIY/6X9qPnv71O
FqLUMUrFKKPSBalRty4pqqeHsMjB1kPTXqseeX8+J4wlp6X3f27VzEWKErtN2ZYH2akK2V2Oospk
yR+pWfu1s/IqKBKjaqtugLrhR/uwVoq7zChHukB6e7tMZdvZPGbFJ5VADj26pn9VJUQB6q4rptUP
557llbS+hM7i5iHb424BiGQUpRyEf19CWaUyFfM7BIYSbTfZpcgoe96l+OHnbgl/VhDE/0cM/Qhj
R25tnBUr7KyulYfeyYtBMVkMsjqzIJFRcrv0g3JSNIKc+lNg+hSKvqhcWn/rIPFUHQZYyUiy4nbJ
1k9M26caLDjy9sl9i8CpmC4hAHPmVm2XpUPQuR8fdwnv/4jDqWjcIsu8av76oDTwD0iUDLJUNP4M
8CXytG2xsFeAjjX7mldSotvnJBubx1YRFLTvX00Mi2hHf8Q5OUiusWCn+5uz1lMS/gMtfdhvu79b
C6/JV88Bvw1ZcUYDYZ8zj/exhCEmto94zLV3nTAD3ibFhOLpaQE17SjqPiO+QONa7DFykdK2Qq9n
/JwD1dsbfguzFBmTu00R6CAEGOkdjJtguO2d+Lq30geHRh+2WrAl+IFilFSpwCIss0TmX3tUN5XG
SFQi4LOVjEMHi2dKIKOwObgnBoybFq+nQK82U+Ts8w1XAr83qTluw81YZi3jRlnI+bSO25Xmfn/5
UL+Rf0OvgVO5jRNh7J1N0ktWUstV09JnQu8Z0iN8cumRs6D4VmXmRa4GjnhK7rRfd3pRa5GfUkCN
v39jAu3+Hfw2C4ni3zOrrsjNm8af0c35/n52npTX01+B93I0v5dHH92u8hDmzv7DDz5ixtMFvwGy
ZQLqbQuttBeHKEQQe1lwUxVw63tKFtO9ACW24+cv5NYj5GwYzcH7gPdNxLAqQaj3AUqN2YUkBKbf
EMnGe/+hUw0pWXfNJvo3tSoVaeSzOVBWlsNQG1W0aPQVS4Au8RM5b1su1A1GqpcJzIbR3Y5KlOmX
XEa0CuCKb3yh1FzrF8Ugu+tvBgm4LQAL2mWQmopycRDFEYfT2RLchy9bxptd+ASByapu6GwjzPYx
Z5I+UbdVpXBTUQXN40FaUNiagYqqHmUpgZo+1mGMCcNwQIy+1g+niB0anENNnJ++XcbxjLqP7VuL
YGGP05WLjyryIAzh+zMvt6puKSxyQyiB7cscm4lM3YhpYYz18A5LXUkfoJCuHzl38mIjkktMsTCz
D73W+H875LkxSJ4UdZeBMidFPciDnWhZFImUP3SY3ctVXRHamKqkF12n75cxvP8owr/5A2N8CLpb
uTBFpcf4UK/Ag4hr10s+K3gKZV/ynS6BQ5RSPRAayfHSELF3J1xJL6hWQGqCh3kMsqgDnq5HzC9n
kGwjAJ1ba9evssCDyEp++JO30HtmZH3qG/H8scscdojL7ViuiTN3dly7ozOyzZ3Sx7kbHIJAh3eU
bIZVkgWcDBXLkFZMT5eiPRyQVlv6f4sPFwa+ZLPHygiqos6J0cG1VVIpTI2lPtPM4xYfn7xSDbE+
7O2rHQl82Y8MLwPgHefDgXUtXs7c+QQ8GMf4BJewbryqbsOV78T5Y0HDZ4pdA9fO+pwCh8t2Y9Ut
l/CTf5pYvU9PCxz8iJ9UnjQldbJtTnIl+qKkDiHLJrM6rDq8Ong0o4G4W1Zu4VrFmKz1pJdwo0a5
pQ4jYv25ziud+WNQieCzqSXwzkycDsw25oUr7QkkIRwztJd2Rsl00DfjLuDAzV4DbokM6/fnrHVG
vsUispc7JzpoId96y22Wa4SYUAwH8HdIetks5DIsH+4tpAXcT9c7Fdon665h1Q3dAx8jxkBBgKX6
IcmQ+ipuhSClPqSh1OAZry6sR0hi2LqgMEVuZeNVGFNUL3NKS97PVcZkVOJnnoMZuzq71yIR31zj
105Ypd0LZ9IeKr44SAkVKXrypTE/OQBw+bnTM8KGXPZEsGggi1fuL+W9txHMhorq/C4FTtN/BdHz
E3zX89i5DFP51bscB1nM0/Pa9/H5k4amDnTQQJU7eKjKDTmN6rRznqqtrwKdZgMSI7IkJL6EvqGO
3hFWTCoAd4SW/WW2I6VveHH4Hsxgbr2nmxDH6PhDprHzg2uZajMLlAvLbL2Vf0hIH5ZUeoCPWrVk
hdZuyTwFIavW42WnwbYtkyMasbCWp2Bk3QT9jqc6c7G3p2Yx5MsuSXebDKuDM8TgZMH2IO0CXg2y
4i+tNjXnkwaCbrp+xR9MdDspvryWsVToFCM5ONWtFRxgFyvRJT5CIdCdmsZ1fovDktBqIDAekmfV
7xE24ec2Mmw7B9iXwYS9cYH90E2BDAdgOZPlfPR7W9CqP9fn0ot96zpww/UtcUbbTEBWMCZFCLw0
9s6cIWuzXyvJ2LNWGJ/hZTcdM+EeIeT70RBLblHBxHx8kd9wKSS0KjzaTN+NZAUg3z6vfrdx0ygC
n6Ss065YRITlVtetW/A8szlocJT62l8+gBcRd+stlQIZOE3bN9UHHdd4FQ/cORwlnagEgRI6ADNu
Jlt2tGHyU4kJCG05VBrmc3yqz6o3u2O55qwTR775Jycp3BuCEaJ8wA3ua4eqrJ4zTMia/FYqqbIc
bLcfLaURXO/9qpMpXHOIEavUQ1Rhd/TD8R4p/J5z5DXSQy6kwzRQ+Sf4qWxzj/vvdtQBbqtlQLx/
hVOuvUyal8CIMpsr4rhcRMI/wCSdRs18L6+4Eesns9pVoWq2rNTR4QJAEk0Av165+ZK/UUoaGDJl
CE78x6ablZu4VTEsk4wFvWlgVrG4Ge1Mi7YETH93eG/q/MOtaNoItHhdyElmEG/CAByGiG7lhI6T
g+cBeNFyyBtOItavOStJrnphxDS9+aaV0Q3wU0/Pr8dyST99Nb4VzmpthUFeaHrTqj/Sw4H0kfzq
KfkdtS3B6dqpu1/VF3JQ9CmzfajcTTpQp7dW5JAKHV/bqtMP5va22Q9XXTcWZpWAJN3pdfCPDdtJ
u50l1c3K4NxXN9OpONTrXh+Zg9xlrumWIRPLwOMJ8TqTK8hYQKeEFKtB26u0MKPCthy9tbiZrREv
7JFst2xw8clcTA+bALSEYlJb3iNiJaCL8jRbldNXrq7lonEJozKrC9Cuu9OkpMfdzsBZwFIv5/IX
9WKsfQLlhNiUFomUzZUP4zIPQmJWmNJMX+IJz9NZvBcUbxb5e/B3OcJqkrHKOBK2zdg43hYSskBW
p6B8lDwodEwjIYPe98J/wseN4fRohR7s5zoUe+hxCZhv8YSrMY1tyiMJZVXcnLCjgg8mFQBHcQ6x
nxLnoJut5KzeX94BTzIzP7qmrrL48TZeqUaqQnsdzC6b5WLbNei1b+W3kdnvlg3ASRFPg/PyNhJT
IxfcH7Vu+Pz/aVsT2n7cLkSkErxxrLHNwDFm2cvNc9Ura3yXcTwLNOw4Hmug6DsrWhLBCHKECC0d
hmVryQzAeq+TL5oZ8WfWCov0INJyyjJ2l8aacI8t3SRM5QLnO0WI2CpZ80Wt+JuNRiD7ztOdJSSr
svPx5LnQTNd/62MWE+xUmLeZgkTPhqlLWOcfpEgywrlm55aMWxr8W7PKJUnsMVftLiJVMH6Qp7LT
9gu4IFK+NlT62hyOwf/udDRxfO+7dxjo2KGgLxtTVYr5Yqjd02bGy5fWPzWBkkhwnygrvbQ1caxD
3Diwi8HkwgNCoQGgRib5UeNFuhMounMZoXEKph8zlxzcBVHyL9mwVt9i5+gOji0V/cAxiN3eWkPo
LOOvFUT4+xiKZGW8hGKs8qA7wMrQ63vaYhyZLQDe/R4EWETmokgQFTni3ENSEDQOrAkORaXpiKpC
8w3wPKFET44BK7GScx20iWwpIcsShW4tcwGo8BMnVwWKizCMh5d5kn0ObJi53fzgTvYjR1bqQ/1L
337KwUviK0IYVOxgWmKApxWpTpgnZla80NscIwxzqmlaEp4b659DYAhT3r753wOBZcA0ANvBAP6R
qhYyrUk5Wx817u7irtZrff5bptt8CoJex7472ARSGXkTNZO9JvZIDhjjx0GcmCpi4AYXphx0AM45
20NPFZ5n7cvZ9ezi6+Rhaw5JH/6mk+6oS/mIw0ISDVRlMnpT6+G4D4Nlo59WcfD9/VwWiOSfQlbT
UCLmjQlnq5UMDXDAqt6L5+fZ5Tg4frE/kZZgm5UQ/ETACG1GCJxhRKqoKi+PQ22vI4XP/lFWQ8o1
arr5/RTaWPOiz9CrsXpTIYh71r20hp0jF1S2GrUNhti+ij4TDkR+PKrjTfVrlJJJEl1lFDUm4J0m
T7hT8evKsIxOD8cEqPCX3q4Nnp0A9yOnWNxsF5jbNtCCMr4v5UQ8RuNJjBJRk7Qv/vya+kOSUlFA
wKmL4IGrVBmbIGIYFce2XyxoxeqHYvrRTfYloEvIQQxGrnqwcmbPy/pVOdjuqmrahAziitRVTJgg
rLSxNKqf+JnOYI44GtbM/f9CCzXx4vVmleJ2EHt2owZNKU7SZngew9PgQ32hpLYyoeE4PYkz4U8z
ky9Zh1KSgR+OTfT+RENBDly26VfM9NZiprF1wDSSxoFG+6RUTcQcqHNIvq2nj7GejgNjx+Jt4kdu
q4FBgNGjBSq4an1wDfZ2fOL+Wkk4ZE6G5eH6djYnUeb05opZLhY5IqhWTv3y608BdyrOjNXLPKcU
u2t/Z1LxaXgrtJ6t1Z5BvBgH8zBSJA8HCg+//aObo/ina6LlyFTIFEJo9Ut/4pRElDFbJ11Inxqq
Y77Dwhfq/oJOG8und3uIhc5bNZ+rDx6Yxvz7m6AH3zweHTGijAx1MIQlNnnFwbeGpLeUlrpDjuzj
Lipyx3YRLSfUSpMRHA9qF0gAU7nCjd36bT09JuPjNIZERFdPFhF3X1anokedDOI8OQatgXBwF+UO
TsG1zj7U/C0vku4W3bkITp8K+5pI9iKZr0EX0X5hwIBa5LW+W8BrzMJJsHV18hBq+118YMef5sVW
I+WOZrG4+HoBn9Ww+AxUQFOFwQS0tN+/JvjdId8yi79KO7Prxa/eaHAcoLhiVtyzwihQxCDl9/AQ
ubvN30U8OkFQKilaneWWgYzNpBjiNS4DUdSP4fJ4873QIEzEhgMktrtfkJi/TzJClu78sXHsUCBW
vWrHEBU8rsRG8w//5dBQMESloQycvzRjzQjM4J9FL5Qtg5kWuuyjy7QdS2lmzIk59iSydYi8wQOJ
XmmPgnY0ieVEKPm3NG8FngaEDAsvIfWmElK/yjKFlsGFCqilaDRKr+w5NAJdxVIRgGil5Jw7UGjI
Fw+5KlFeCxO0ozSNHyZuv1Qj2XdhArkWP7gcjdDu+LmuhFELDw5FQ8tNzB0dD33JZ8upH2j/TNwv
mIy2EvRRQCRtMrbSE/m3AyMmKC7hfOaNYn5Vi/7sijodqfhtE7fM5IrzieNl7m9nNsTqmM7Xe7bq
437TfHPpKU9KfKunprsFQAGkzlD2zMRMhTB36wXX32VQXrbNTKcwpJSoyYhrHsVryCVFL9WVXxh6
XwEHAbyauNOVVXet7FFNpKAWYHN4ypLCyVY6NYQPPdLq8QsNf3YOq2rMJLIfOnsQ+4d0gDZzmCGl
BpbMWugP/xthaI8Yg70z/iqrviKPacSbHHEY1h5pPQycmhf3J23KZMzoP2np+nEr+Tzs11dGnZBZ
2qDmk+DD9Joj7WpaF78vCAZlwV/mbz6yYrFeM9Z8vCr5+qP7bCVS89TtraamIz9wZrMQMw/OwAio
8PbIuVGuhQLcJrcgNlDQB+k3ZbCKLTXI3rDK9RrhSbG03dzy96I82a7HpQcHEycF+gMWdUpL4gDX
bKjcTO21SKq/lNEoo1lM/cRZWvYp+TQogZBxBzdc/jYvQPVi+uAcMeRKMBwh9gZhObaNHB3EtKQB
OnCQpe8GVeZeNc8WplY61TaZIMDXlAp9dDvuNG/0AN7x4rPC1giqo5w0VuBWclKfposh4mXKGf8j
9g9gugSgFxi584fe03CCngU0Mst8NEb/LTtMiBk4KsVz3ucnpQ8Q0y3c1PzApnorS0D36n+z7uOK
Lfj43mCPcjIUJZL5e+s1xmpETxkSoDY0qWBhp8TmkS7OlW67eefAYysCRY/OT2ewEGTulEHNs0rk
TKVU1mkIaGN7U0ZbrkcOG+PiiX3KkwqZcW9fP0GfW881qECIR9knyxT81oVsvsAs9JQZXfIrloCL
F4jF4CAVigkz2ZbOdQM2cpy+yJlS9vZL74oIx+BVW5qO10huPqz5dZJu5pn+RkujbVBfcyMnnTIn
dL7Zcy8fC2xK+kk2vF2LkRzq2DYoR6eARgGH1+NBi4HFuqYFOYvG5VxDyYlVdGMeNPAkjFYCs/+d
ZEYyEpghKu/1+dXaBUrWxeLmH6GRQ/SiLWVs+BFQJncYdk5aJPQNfO7kNKG8mzhlFPZTNQDgebmO
P5/dhEINh30traONtJNtqIAxQsR3hRos9GKNBwrjPfYYprk7Pg7bYKMnE9NIQf4oeELxSUhelrU7
fGY1B/N5f3k8woTfNo1HKWTsijViP/1QVHk8YwFKpTMRYulLZTDZPZpHaTH85ldK0wnoN699Z997
9Iem79zho5ebWbcef5JR64q3acUI5nyOJScHmZN8JMutr3B1Ds+3U8/xSrF5AFOW7ROyb+VzIMbm
mOP1OMpmmsgnMJfrg1ygoLvdYIix5wamAjDG+NuTrLfrjk+U3HtU4HXSgtGhwqknsMfP+FdZbpK5
wtZJVU/0trWLzy2QPCP+5DyiGwPTizGF9w31PJKut1aN07F1U/emhiMYHCz3kr82AbQnZZGGL/oQ
Sf9eta3TlmvC3lJtkNFWIS+FGv67Bu0VO52bogBH556Be7NzOksrkW8q3Av7O/p7fTcUB2+cTXPR
5H4mZcC8VnPJBbGv8eOFqPjHOz7oFlLIIzVLGGieD9Q7WB9HtvSATXmKzNFssyRLJkAieiGCnUMW
ynOPzcId9xKdRK3GylQku1Dg80j5xTRmZ8IP/fpnk8rOXIUwpuTK0g8JR0vRh1CxLo6PIzupemTZ
EVrth71QLjK2gT5MVTqIAn+L0ikUMArIh26NiTNWjViJL99EHJxlbQKPGuy6hYu1VjyBQsWsAs7g
XC/z3s9w/t7srhMO2v5ZoCQCWxRwR6YskUavEN7+QNWIliEMP/+OLBFzn3JbVeeFVd0EumPR4Go3
kuuN+1bcyzrmQmWFmcm/spv40e6WoLzaMmo6u1tRGYZG9NLFKuXvcSBHgx/5QhQbpEbOlEqCLEKt
gv8mDaJ/NuP/DD2pvQuhHqcSe2iXwuvZG4Vk8A2vXA3HngorSm+TfsaIfbsLjcf23YKPZbFbaFCV
r7o9HlvQSFIxvxRgiqtWRLb9o5vCWb6ek1kkVjbeSFOFTvUMTYFvPy9D7rx/y2csLZgH7r3xBeoc
8aG1G1OQu70XoKBsYJ/B6Ls2ryk0QfKryn8xsZ6h1nNSrElXnmPlVY1ZmFIAPygsMTV+kA/MP6uR
fPTJ1w2JXqI5jtOSagV/oOr41MOwV71qw5iJ92zWo/03AqrBFQjZGGAdJtFePhoI6gDMqDOpYZu5
8snJx3gGycDehUSB2RR+JOWYWXAtdN2APL2+H9aJYMAxR1RbwIhI2ohkEQhuq2kz7jY13ZJmGfDa
JuWwmyev5kVj6kUnBtIl1rCHY6NNfxI8wtcFTRSCwCDdnDU3INK45rMFfQvYIfDOsl3g8DafyPQG
RHu6hD6vj4m4ei6MqYAdW4Twp7pbyJlxH28A0cnrRNuTsMqeQfborbaCtzW1Xn1Y8UKUhlrjrrHo
KEyyRK1DHrBv0sqHsz4GjNeAut8YChlI/7eAmaeJcowjFleaZov/WMnzo3gTDAxlIMIktel2VDV/
w8p6mC0WqMpP5LTtzbJnrfz6j4m8sfjn4KScpLlohdVpnyLofaD9KqR6JV+R9w9x94DMoFAibnh/
FDXwv65gFuTLINl2H4SBer/B0BcXAMwlCuvaBgDkqKnWN92+D8pGs0WbUljS1sh7Gj1jrnq1q5r9
dd9JX9a6qUtytslAMtSKVZgEbYbvUoZqk4QlPq4yEMiTuVYjzWQF97AN2L5NVmBJavxNtWARs0sz
xra1RYIudJjWdiaFzWBPMjtNOrEPk9qiMYgbOny0Z99y9PWoGi0x7zvuNVUDu7SeXDzLjXN5Xhix
K97WY7aIkMl9429gAyg7MjZ9f7LOgqP5VgowGR1WIydve33M5oOQwvLwLv3kPudTWwU764q2c+Gg
aQVSCXCNIAAIz+MbDBAlIY8yOtJi8B4esceNj6ffDxIKS2bbFc5m5MXRoLAWcr1aafRz/EeZBgUD
VuuLeVFXikvRrDGMj7Zk3IegA9gkGNtm9Ohqcpzrv8oOtnSis4abFT46HhITDmDPGEoI/HK1wAc4
B+DGK+gNAvhulgQ0jXCfMXcNRn2pjyaJE/z5HZWzXGHfH4WR2YBPEPeZTrqyKZVvwGCqI9NchSPu
JNM8HNfPDLkYfHraC8eyO9nIFRMbPFjMxXel1gizq9b6SSTs5ig+wL2HfAq9ZmGOWGHbUEYtFxVY
9UFzD2VLB1PL7fkiiUnpqsAG02C1CDH9+NTIgKfASQ+CpUP7pAKUYf9q3cX46SnJnudC/2K9jzwp
mQeoc6TEF8IaCyX1OIgdQl7VCrsGxL4YsgDIa6DlmA9HvBZ++mrLNbJ0IsjVwusFzCpscysbhTE+
+t5Dhd5IrJdroeW/w4CjwbtDw+gSyah7uD2dXcOTERElkvJMRINCDYSdRwkGDW0mKj9kSyzeOJLG
LnmsRWGcOofu1TinBM73LP9+DPu0zdKIIM++/boai7sye0WSPTYMfN6OyHTyuj7tm0QynyTP2iRG
vS+BZpuhquOzmgXWHu6JN6Y32VVIZRuPPsmelIWeYinyUp2GVS90PwY0JW/SSTmixw+SEOy5dNSD
fXbFtjwQ3sFNxUeLxLa6fst2NZgsFzxAdH8jZOprCs2udENbDXIH8XUrxZ73orx2p2VxfdXWhJKE
i28cwWzWeVzmv1HeF6PfCTnwmlOqVwPBbq/hdDEMN+akfmvASebzTWEO6VUV47kjpIDu48ESvyLS
SyW6RVPUErwEY/LryqTJbsJSRTaCmAxtKh1YiOOimnImoo9I0RZ56zxPmHKn6+80TicqGm9o7hgN
RK5O0j3CrQts5xKhzJM6AgcMkQLYH2+om0uFbr4MY09rJKNPoW2LaFdtwmxqQUI098Ith9/4E8Mr
SbnpWU2XU5F5bF6gmbnPn7j+kI88XLrdKTN7/RX7X6k3l3q51yxKNY3GvfghaBmqUl1fBQPyniFP
O2XmPZQOrzZt+xfAVoWtZvjPfo/kSnqr0jscAhBgT6eBGaQG3zRa6Q+mfK3kzv0q7J9pdjL9Q0tv
kZjUEST0jIG6mJSClZyQLL8LUxUswGojTiG7j7f02XnodlgWAdnC5FqJZA35cFSWyaF23T92s9Ps
8Ek1snaWus1EisCjkyDtmdIb+wkAJA/200EuqeIRz24YwtUHV+U3NznIPyz/MP8E7S+R4YP1jouQ
UWFfLZeN24+YQw8E5TwzWyLjiTuJ7FtSQs7wXYptuSX/94F0JtZAxR5aNenUezDd8xcmH4viXN5M
0CWMl7IXFlaFaM+8zDnWbxm7b+cRbx7eOeDeolcSIuv2w62QsQDKY/vFxU0nVMfgN0LFo11Tc8Ci
6LPV0chH2oJZnaGad6GsH4LiajYP6J3SD+2f4BlEsphhQQEN5g+Fd96uitObXcPWFU20Ao1agYnP
zNsJmZNqxX2IZPCWQzyx7YBXjqQSPWMQiOBvvBnNOQD2+QAxLJpn1BOt+sJo1+8+cVEqD8oBYwiQ
bU8fElKHQsNaJBODxT5mFRwPqE89DNdTJI3WiGxMc2cc6UJ8Us73eXdVZB4GAFytV00kdqjGxI36
JJXljFCQWa/jGhBFQFYn3cPv8CJ3hujQFwn4LWodKadgW4g4eZD2dOoAotvxRbqoy+WHVLSMti2Y
h+Uf/UPTzuTjvjINsknyA31PqL7wb6DlGXRewDR7rC6FG0cFoS/GeqVRtIwcATj/P94dCIN/aRZs
T+znRz3mR04ZRMnqplBVhpCCZ5I9O27Yfb7X8vERgx7fa026hIYUk1nE25fogYSR+K8ApfjOD8G4
PUZQbkzQ2h6EMIkSJEWjE65VOUAFsuEVKIos8dPN1yu/KVr2UY8Usygu0x3fEMYWhEXbZT6KH7kw
7NaaZEbcmDj2JJKp/l//UiCgchgisNR/uPRNmqRvnKwtABYMW5LpZNuHCjLhsaYEzySCMOvLecdJ
AXq4h7rYqeXLNChGCkBnQf/S2gL/mk+W0Uq7pDOoKzR/jGTxmhHyV6tmd1quHgKmNkuNa9fqqceG
l2Jj5YGFfAHuJPJ471qdVn7TkN72GzBZ92m+nDa/w86yyYX/6wsYc31b2msbwHUhQElE+1lsOIRl
7LOiQuN/OuZGsIW8qfFLZ4eQty2e1Hz3g7jucIuwnJ+e3XpDwMLDc2OhuPyndNZXs6PaLRn1ms6N
54z5YPOVQ1U/UL6l6rc+v7nZD/C3myJv+yHWmrqhZ1i2y4wIo4UV/actyelJYXGwLVhUE/0zzNVK
qVFrVvPuLSWMvIEGWJ9W4Tuc9RcW02RaKM+l1NO+vdvsExgs182YlYq7ZrXG4XF2SOlcEi7bmLaD
OVHd7Ru5QdfU3pWtlWLCutU7h3jNVuj/28UQPewgRvVFW+DlGPvqSTT3CghlT1U86EU1ybLFy2SK
RRjeYOmr1Ywlw3n/QTnJ2WMFikJZ7YoKGCN2bxTuIwvUoOoH0UfkS5EbCDXeFiGrAM9Nq2K3JBwI
jI86D5pt44IpHa3nYTrdyAn4zyTN+LRiwol2bC0RmhfH3OiYmgR6gt5tWiqqMc5yDP9rvLqYbrsf
nb5b4MGSrMKIs4dF/1rF8762lUepPPsnhc8kWUyIqmrj51PBt+1BqTeu74WyKlUH14aHCr77QDRa
GNQ+3G2ehEwZp7ilWWl+efRQ1B9imMzOhGZpx4Fzdzc5hm8LTWYyiqIedVNGfbhtY7b+5iWZv/B5
J03Se6BrZ7qpe2x0nzlpSop5TzifJNWhTP2FD7ZYoQxQaLE7sBEhLkScIGt8G561VudDfkfoBQgI
PN3FNfJJzgQdjGulbiqYzui2fD9/Y1WESPg0G425eXDFebaBfwElykLI0dQpKeYHmP/SK0tAzGO+
Gqkl7x8UBvIdqKxY/waqEJhubXanAuLFUyzGnEfRa/dcX5uNfbc7vOggU8i0M1Ex2VbdKBxuOrhJ
7S3HpgWxmZFyIodrB/05+16CMO/xFCDhkzMjAq1SxknhHNCyNk3N+9xlDtjD3cB6cUPRblCjrpAv
0RzZMDlVuTwNwNn29Hhb15IW8h0CiBEfWRgvzrWUJT1NesK67xW4beMow4cBZfsqUIEfbDdNuQjB
sdM7x1CwbzolIHYyvEQRsl/TMA3nUpmVz91sAgiqFrShZ6PmwIU5C69iTfWuisU/mvj2rxWeHRIq
Kdq7nQjZI/f2iHsh9xXj1wQE+8RI+0kI/Pv+lU5JTHgyqDzkqW0kyDjgmgVxXOFOQqV8LJrtZxTZ
AfAU8muPI1XWNjSzQqlc/Drb1aXkYE4X1LzYDQmWlxpDXqx8rGfPhP0Sfc8kiEwmcFa+qf6Bgs6E
BZpuGvlPsD4PcIOf8D/U8isvVgyMWU0UlwhzOJgFAU+iFlgQIrED1e5oyU72+cBiyLwnBS3VD7ty
4//zRKH2J+zi3NBhCWHDGaMlCeMDbBCPX0t/7Rgay+RB0UG+BR5LBxx8v650OLtcIXOgO6fYqDgw
I8pqCMr2RQ9vA1R/kZ36xX837g+kG47srHO6JTLi61PumePbx54fYpnL3N+ONJrjk+IbMGfTMU2c
KLZIVGaJTDeosomaSS/UKep2ixRchUUHBq3UeDEDLceYy5lpRYbUTEQ6Sa90sWqrkvHY4Xd6xwQw
m6rOUruT5d5dgwbA63uhfaz/DPRxDxQTCXOL2H5txfvX/CD6g5tmoQXZLvH2DAPxnMh6jC+27gyn
G/RAOq11FEZA3HvtZ+FJc2UD/tugBhZO73/GnAaxSpIot+MKJY2iMjhk/EFtoxaBraUBMa+oatGC
hL7VjUy1BCAb41fni15wg4ltam5qaQiAFx7FgH/szP5xRhYrWBDGMFhquoetv6Imnj+OUdoPXKml
bP6/4Q1SHDm0MKEAj3rKtSXHu3Ie//U5kMSGJ7f6NIst5ZDYIjIGf41BN7+VmAUUurUy8UtJPTER
wMS5+c96yzUfIGEMGA7ODZQX0IxjfSAWiI2rFwVtshoSDWkltoGytDOJRsQhKg+kmLQ1pfXurC4J
VQbysSSGF7OnuW4Q6i3a6P5trxXh0s0a2M7TQxTQAuCIcP1mlpV5kYk3BhaNGCStb4bhixuRQraE
hrwkmF786RWCjRKMV5bQkLGcbG77JK1HypLm3JtR/HAz5hyDxhSwMf2GmZI/f34X/j531zoNalUa
iaLb0gZzikFAoIA1MzE/RLGTZJd/Rld9Ut5RdjnsBQpqAatStBNS+m3igBdDcahg7hv+myI5VOrI
IQSyysUJYgYsDN44epuTUu5SSoOS0TEFQKwWi0K6uDj1DZMLfHUqA5hTtTvErGNb+ZwSVKDHhT+6
o2GaIVDDFZ6Q7WOs9pNADu7aUD7b+PLK1PQnf/MFg7Sz6/cTNXIYeApL4aRcTr2TVmydpUCnCrt7
8ceFTkhGExfgX4g5uUh+NyPwR8EZKYVL88+0DLaTo4L6yuGkiS1CN4lQNclXh+OuRuf0ee1fYldp
jysepeKfezQMIxtPRX+Rf5AiKtCVhbB0zFuWcQJojupArQBSqjB4MGjBxVgcDuLfPBVCTQslxHmC
7xM4nPIDZHsWInHlTF6YG9EZpUbRjZE1oZ2yktIIxdTczsfU/sHzoAxtMTQI6VgShz+fIvoiWNFC
kGtv90nIjOKydXOGsphqGDOAlS8l8gYxIHAd+RDygJM+7l0StP/bXNwfs2rsMdYSHbBN/b1WvU9D
qnxTEW91QMtl9cCMmun56OqLn5amBWmNk9z7S7Os8gdlFEFYoIk3VhWLNjSpMyG3QmREYYGJGQ/j
BSGm67XUsGlYPGAOR08JokMiDZwTNi4R6zdP7xJjksxqCxCa4iSHpHaSEbJdxe37bBv2byy6Jm1l
+tMMRjC6d1lGhQ11MBoPnF3vDhXyIzT2SGlhusyylYoi+mz7+N8HLUi99fFwm+7shfjs3cGXEi8T
5o+pIz5V6904vtqZWXv47f/EvMVEbj/qJRflaoH/meK1trG8a7r+WPQQPokqCwrlZ7YMUxml050K
1VKubIaNGCMhSxgEYs5nSmwOcccak+V7+KwM8QB24NSmA9D8jAPUCi9TtLRdJZDgzT+cnsBkjdPC
2HwIi1haj3xueFK5z5huCommqnRviQwv9pxkaiZ79itSyl1NZtoolgQhYfcO79KPwejvSIdzWGBZ
EAVncxFQKYTdtJkzaj8PrUBEFwnl6o8lDEGwdXCMxkkkDZj0gP44OUotJkq34X3eYcwg2PlfBxNd
BVa8O2p4UHa0d/e9Hhj2gzSE2WLxixaFTQLpLuzprgWAlWvoNv989pbx7iEIyleWQMkAHyBUcy4I
7iEUoBj5yn9ZT4Y+Vat+zWsU9KOiChZW9acNH2n/VwOsqlolrNlfmuR5KF163HPAxQKIjg7gRwAO
umf4vSPNVHWiTz+18zfZ2x/MexCjgCzInPMvmrC8VjKcoQlB4NnFPpvgKQ9bFIUZhd1J0Wh7n2Hv
Un9KOJpXd9V2XPW11+S60bkTItkDbRIqAN4pnzd4HuMiSq6uBBEFMpeFZBaOIGIvIrgG1UTRXWU5
ueiRP6FsZVh6gKAxVXddBpHDzuRNdLalFzViXzCZIGbjK0g5ZPZ/gfHBQKVGkZoukBSYJa4q/X2J
0ymPO62Afv98RXAWshav4vXYFWNMZLxZVAWwKmiHU3MPaUD3ksy/beE5aaSyhdP/8/+JYom7Pbi0
mxjK5ndQfhTt8SoFpI3yjGj7TRlGCUdkqslTE7blU7czqiqk3lhJecbmBOkHY141579DbaKo14lq
uvP0KiswCdvs3lowmzudvVg8LAkH9LATjcJPP9vQoKMwg2z27O+hu+Ax0+SbOnJnldtX77TtUir6
TRalkiOldDkrrweVFJp90ItWWyZkBj2LwjthT6wE2K1UiMYWu3Lib2F2pC1X/oVdUegNo+WdfXyC
YdM5NQvlPO2XFOESSanJ93AksGrfIb1h+V0RWncIzBUlv2qO4hHkrAzW+wbulXNzUWda+zlWFlsD
PCi1i+Y6FgwupRUCkyXcUgZ7cL9Zm83iZik125IUs10iDObHZwsv0sBWniAH3cqkQEFByi+zvTwJ
dRM7nxn55p/FQ7W21UbmKVuwfcgcsg4DUnAlElXAURzWKEFaerJZ/GozVAkJvq7o9cNvJlDZdOTC
uHMIFOja83dq7OsiRkKiDNBkH2I7w3smh+mjY+aAQ9mbka3Pn7XDyjkNpCv+Fok0YXD22G7/YMgS
yFVVM3ddiYTajOIowa74mfrGdByV7QM4ZtNvN4TyryevN4wXsA5qz+eF+LUH4vdmfbyiqFP9tapX
Gg8d3ajAqHTTD1G6ycxyg4Pwk7yMyIG1w3gz9mwyjBKEvwWHyc3p72C0rLTj46Xk1/kzXQF8JeBQ
HkpPm+7uC+7FEhbZi2RCZOhTmilpcJhDG/6YKc9njenpvicC+MNSQvW8tCdmAHtwQM+yDsNzb7e9
3izKRKT29ji+tzxSVGf92J7rv+1I88DpxpbZ/rKOHP10F+/lx0W4wq8MZaqFXpLQRCcTnCRECraU
NJM/qMWRDnUD4oIyZ8TywHeiNHnkUpQixixF2axIcPfrqhHyNSzmidMtfbYEH2vBtDHvQDnnffKo
Te5iH+B0X9UIB/xSLI3xvk29QZfpzIN9l4RxOpMPttZjgPk+iEWNl4gU0PLE2TM4lULPqmNZKsbk
wqp+jR5EN2tN/tCuqKCqF6JVzh51Gklw6kgbzqE9j0mrtYB0QO9AqFslLKyN/k+B6ZPQo9AbYPCb
WrY5R45rRIhHjj8UiVweYaa26uefnqO29StJFii0UHlg4kmKfUCi9/WP6ZjeFJndVV/j+PKb8hEp
j9K+IqUb+UUgqLB5/1EIBECkPeX0erLHOPl6AvAU9Lsv8Wq0auLjCc1bQ8qQY0KEsZWVJEnWyAIk
9X0aI0o2YsrPl5KA2nHrzMqEdyPSnn4tFK5xa5YE84Dd6zzORpI8+942ZuhaVcKZhWCM26bsrw9E
5G/xknCMInbBmtaFy7j9xZm/oJSSWj8vPzNdaTof0Pi5WkUForpHCRyaPxlExIJgbg6PYcb1t/kA
07dN3UfbnDOguQhYRpysugQCnievghVdGWidG2lhzJwzdLtXjq+e2lgDYc2nV1+iRZqETo53PzdO
tuJhNwDaoCdQok+6L/n1TYMMtF62IgEsKDGPeBZHLT5B3ArsXeEDCCfEKCwlsJrdbtfAhTTxpO08
KSuGrAihdcJ7Q8bAhUlf5IRb90rmPEKmeuOEgx8QfKViqK2bSOpkuuYr706hmKIEsSK4oi3OoI94
STQTuN9+dzOvIRdptYwz/uWGPIqXXpHcmb5GR3rB64hEFxCwfzwbi7sBP3xKN2GZNv5Wp7sU7tzF
fkmpIgYLcpJ9adrX1W+LRWzzpfhcDxbsxxmTX2ZfseXqa79oZA5vDSvy978MBS9Mr0ByNSsQ8CU2
SzzGwBsvYxE6MKZHxk/edFDl190v6SWRxhLVNBWpqdWfT7XbxM3Os5RivnUtEdGHNRlVhiG0ReHW
KkXMKUUOvdv08m1rGt5Jk+SMqYAcwJ6j6OuyebB70fuPdVANjAQat2WKNgtAsEjI73jZoUJ1tzqc
kxNl3vz8oSJ3n+WPiSy0FGly4+87X4aX4q8LQcDueHCHL3IZ1x1bPqsjBYDpwxKnODAYKxOcxZ2u
Aa4xgZOi9L3c4SnqBPQIhiDpNM3/KCT11A1lEiHyPg6ZZty0usY3VBm4TTVpsjEtwOoHWygP+fhK
CJrEOrWMA+OExYmoCS29SVcPTspvYRkqugJZutsK+M8mYFY6Q7yZJr2uhqYCEvKzmmEErWwprhXt
Vtckc/h018Z14CwqhJYNhAXSRebOrEDTB5wOzGTcp3RIMXNvv8gCdREr6VBl5SXYQBpeHl/oXdLY
lJ+T9w7hh07rdkITqdg2wvvIS+NNuKn+5dOlL80sKXMyS95AOs184pE2JY5BixXjfcZ2b+Awu0Wx
kme99zB1hOxMtgxmzHfmMUc4LoUyX8PC7e/12ciO+nHDvOet8PtaxkKl+AqUKpQ6PexyJxCh4oMr
1a7r8IkOAXLszboTF37s/i8Y9rNoJT/jTbZrVG+NafIeGI7HITM874I7YLKEhzylxMOHAMbqevWF
rOpSJOK+OdZK3GyNatg92U5nwrNDgFQM3p1GHXR1t7RqWzRjaItvImU2LSMh/GifB0nPmBCI6QxH
mDv0+SbbIELjQY5x4APElmQmXnYpbyz7NihFXTz5D5ZY6Fhuz9wDSYzORdN1/znvGn1ZFTNpO5cC
dLAHzaii0oaALnXc74+l5dcVdiraKyncdZ1TctVKry0Et9tHZvylw20zrGPbLsD8eCEECfGmiFII
WCdYUYJZcpyymvBx2Jv9sX7uMQuWfZd1O2HHzSr4MRvCeo00XfFHovpbyKm3Ijlvk89QMMk1dCfC
wRZNqfAAnlx5zRupbPTnEzv7MQchvHIu5ZDTq2hthjyD3/mBNdAlASAwGPqFLZBub8dV/K6IpELe
niN8zUZ26KUYjpmTOLCsYstgq2Cn9LO6ZzYU3y4lqujF1SppJrScZtdyGCaT8t+rJ9op17hLjRmh
RJTQu/ZZezdtQI0q4XYtUe3MwEEZd5Yh0fJeFryS1BTSdh//Brrh4OqYlzI2W8iqRuD1IlTTfNaK
MDqptT8hNC8QJ85Gj/K2D0vU/E2vAft+IQu8qxL9EX13ea4CEAYJs2JQlFErLs0whhqPmW+Pz9Y9
MM62fcBs1uLDJqHjS7ixid3PAUBTW8D/xwzcV6dN4eD8Z7yuOqn0gUn/Zm/YxOFXw7dJIHX1ATgh
23H8GAKbnyQJx0atIDyxHa83CRo8PXg78s2WOfZqxjFdNOuVZHRfhbhORWzq/Q/zYQPy09sVN+Zo
odNb3eb1+c1Aj7nOvP1AyLYxZsonPNGa9ZJm6V+GT6YUse7XQJwHo0QM4Su0HWIR+oUoDrUBDu1H
Xt8Ijrr/VlHab8uYQw9NA/CmRCRsd+h1We+wtwFiUxqSQImizcxMkM772zjYk1HTaX/wx7Sl2q1F
YhZQ1y99m4bATd4UcnN/5D/M8Rd1x62sWu/K1iDhXbZLQqmGlEqrEpifANpjjUUPMXHu56xE1kPF
S4i3lEe6GUwyQNgq/6S6/+v9wErCipvKMqsdl5hTZUfF/9dFG3ZyW4JsderuouWGGgzwCwkLCSGM
dPubcVDJbwvHaiymlWEyddBnyivdZ2l+29JxFtCJ7WKu2ezMJUdu/70vxieo7PYpqPzlpSq0c1mO
2RuVEbnKIZOkgItWiYsbmi+vFZVPTG7iN6OmE4Q1eXAd/wa3+PNQRVdiBXonuTBwYCJrvwdyku2/
O5CFQqkZ5LenkCQgDQITG+60BZfzXN7iL84OMWBf9aSZS7OREJMb+DYRrItyZiBlqPV+jc+Grl/b
4LxEqZLCOnkrFa1C2VXxoV8SJdb4x4tRN5RT7aWlLZMqE2gM5hGC5XYMxsHIOCP+5UTQrnyJ2c4c
qsrQStQSddklzSZcc6AJadnEdoVqTsCkO+6XNXYIIFFny+4Xh4X5xwt9dLSfd8TZTRShF97vVEHH
Iwft2tFK0xAoonAv9nWws8cM0KGIhFhuO2q5vA1M4KaGtONW9Zukj7hP6B6fYgtsavo/BBdhXlv1
sqXz2cte1YyOX6DwBkTLCzckUqJQ6K5KLhAuBxrQQHlenzlAJxTKsJc8NdgDAllwZIJ0icoOnrSl
12+ygzaJ5yogcc4lSdZajkN53ohcA/mykluf8J4DBePR/ns6jnlXbUGKSRh0CUN016WVhMI1QV2S
AKJkRqCvOAAiE+xFlFPLGvNHexmcPz+SRXMGEEfja0a2HLGgMa2/zuYXblYymaN7wX0lUJSHlzsX
w/QZe4DjeSaWYQrS2CIB3wTPX3GvW2ES4s0w/lwnGfeMigsQ1yJSlpFuWf9X7+HfbqNnC6yTWUF5
tSHfVLgtbWSCo/9cEZ1kT7jX7hCfBOnITR8TZ5lY2BdAAPcrG1qHRHEjbcN4YOc6QLdOf8kUuknf
3smrIS0xNBFfVp7ULiP9YtgZcmqSkY2MuFsGn+PB3z64TrNmvNms2t1MO3wMecSoUu+56y8j0soZ
dcvj4anA7Cp7ewkYe5Wah8kXBgY8/mRWbrc8rnrwIDwVI5S5EsLJdiuWx0cvt44l448sjkDKYlhY
wJrBqxjc7Gzuwx7gRIa9/lFLaAtLIeP8Sg4V+LnTdjD+9jenMNRBZtvqAe1nGTDbApze2PyzoWt8
rhjlR1wGLFSjsZe3z64MZwh/EePZCpsF4Kzt2UpgZuSSOX86d4sgSSJJYOwaB+Zj/dOKjhDppUmk
+fSM8PKOIctBK7mIqf3GuhrqrC3RI2142soxWkEpPnbhLgNbu2+ZeVO25qXhA+lbdjWO5tkYGck3
OfFhXDH72sPqnoDj3looxwRQiTjWULZS/BoesQ9BTOvgoljkndcDuSTsFPgpuxB12mcrq1lhxHZ8
I72jriBWtiSLOn3OnjQLILnLZXWecpuqKjqzXtdjLt2ofth7n7dZGHKxkvt8JNfA7V2tIcsUzMEp
4dtm2hc416KrX85h6aNpUfxrqrNh4oOYbIU4OxjqA5UAuTzhMDOxW+o1dYOSfNd5gbuOOcXX8NWH
zNo7VVaigfmyhFZN3fNk7aYNXsgFOofENxr+2wn33dd5TXMU8iNb6h3cnDmuyAWpK/YXdaWBPaTS
LCu0xWWa2wKWXg9ep9C1F2IdJX2XLZpyBbPiYNIiVpSwqYbccfdV/IaJ0jDp4i6jpUXt7Ze7FMuG
IlOaahEztOr0FA+A9zQYBdECUrze1ER1aMEPvWE3Drha76UIVsAFoM/ubEG840YoCx1fjN4JiQqp
b3VVDCkoZebVZJ4PhByw2JuNy1P9Ko81hd0KI8n3C+kLOiOQfv8ydTjcB4eYSTuk8Xvsv1afJHoU
2YK+q2bESmlyfofV2U1K9FI6aOyOzXCXxpuMGhP3CXsdXsMquj4mBP+5gGCvHi5ElZ8pB4CiikFL
542vexEQq98EkZPHlthRGY94LCsfHTiNgc/rzSp6nNAk3eaxwc6Vdlh1MfzkSBRd8yt/XrXz29ez
VyQdTgrRB/bOPN+jAODMlEvX5f/UZ81LPiKZYgY2OeHsabDvlJPFnufpaW96warYhEPJZE5WpfOj
Uxzc7HX+EY+6HCZpe/yj/1kzl6+XKu1SODWnB5kYzige84w2ZJ1cYw1z/ldEOumdwdAF1TIk6PpE
BX7EjYVdPzCF0gsL1/ZO6MiNTFHuBfJ2q9H/siaQJ8n2Q6FWDm0w8oOn4V+aYZ96cLPpCVVTR/+O
9lOvOUCuQM1KDoR1Z4sEt5Iywd8Uq40RQ9ZvgIuRTirsM8Xp0YMSkgMghj9pEfddPE6eyjdpwZEd
cjYtdzmwAfaasmHoXn43HzKoOlVGdO8/U9j83MXkdUlNVzlazGhKr9jA14Zkpq52buyZIzv6LJX8
zwshlG/TWVm09w/NHv3pTBIxF1X/rHuE3pO+mFXGR4biYl4HAdNKR4HRme3e6vvkcZyRHk0RCgqW
z8Gdvvij/+C1D2e7AdI7a/w3KvLGOzkV3rdkGTaXMLYRRGUthgvMYex5njMspinRkpWug3xWGhQ9
xHv9Xs76jNfB3ImXhWhwmESn5cTNKxmEsUYGMU1EjX+TgMn4thCIpetIogy0GzgaxfD6BpX3tQqT
/XkMryCb7Tn+31XfMw0XSIU4c/eBwez9G8G4DayRxM5eZOFtt53+Xpho77dBPfqhhXe2nShRGYjw
vdMJeENnjfjE5GgkWl3ALr1EvqSkfPkkMO5Oi3IMtFK0AIL+qaGHvROTW42f1X3bLyu0XE1Qub2j
+PDu8SjUJ2nP/NkXI5qj9Np/o1OYZZ/WEmZE8sQ2jf7Mts/YbzGDni25jmugVuPvoh5390tHRA+L
gCcu1dLyj5iWIWgx32xkr94ri8bzAYk3hxAqf9oMhVm3ZWjfB/tg8T3/eJ1/GCwwUOZdsVCOvSqI
9AkuaR7Sz/LfpqMx5E0GVEONVZ9A3pB/XNpJYAI0hAjUqGrSzfTM6m3tvZeUD8tow5FsYX0EsHNm
1Z1FwB/+TGPJPo3HVN31aHpwjFBhuovcM43KvJG2LWbDqZLmCwQ9/LWoWDc884yfSD2KxAVQsm8m
anF0eN5gxgNfZ4GEYMA1WbQ6bbAMftKS3saVgs4AjXXR6Gh2g0IG75osWn5OG/0rQQAs58Cmgt6e
BvQt/A3yu99zKMpt7zICmPScwM7pZ3dZ4eib0zXy4/NAxOD+LbUJ4QQfnLYXoNrorOsNgaD/nrIG
SJsY5e6JFdR8EvihM6gMYY/vlnBNXOrKHfGxpEfc48Nd3ii5Ac3zve9Z2xT94odzOEfedfn/4929
KqrA0Pmm6Oq/zdwL+iK29owr1DWD8t4Yg1TVRwN5JP6+831g8whCbE5IWNb4M6BkFZOmuhvw6klm
ZzDvNhmlMtZyONFWO+mDgvsxTK9v33EBjoLH2XrtBo4S0xgG7DOpyL1Qn4HOPAclPPFYE8eAb2vZ
lUYl+r4KdlO8B98tRUFiqD4w1YDjtzC5D8WumgFbNOYbRjGRoz5/ldPCLbU5S08dDKAesX/zImcV
kCCNc0679RiW11ng0qZanMfCUzM8U+9ufq34ChA70LWe6540JX6zorN+IDElpylSBM+fdITrnxBx
0sHqnd77DQI3keUrwTw2fij0chwrejigBctaxcf851SZ4qnNgbfaJe23kaus5zFFfhUleC3kGvMN
xyHiG4k7nKtevmgVjdwvaoOrxXC19tjKAeCGjyWox83PaBZC0rdK+nS4bq/q90iWq8PWh7DFveRd
I7Yq7BjucpMo6w93FrxZIwO1lnrr8X8l5vVoL7uR4X3tvkGVdeduSR+LVJLwUtKV0hOck+G9DbeF
lpFbRjQEimayx1XNtSiUAxW5zchPcFI46ROZ4ohShxp3T7tX1AwQvhg41w9Q/dc/R5A8TDhvUe7U
RZbsuHpT0+xY/7Db6NbStZdwtnzLe639LNHIwkag90cWK+BOEm+x/N/tqt+WoHNKJP8Zswl5cHPB
RLVUqePDLvAMzp4CepI+vPLKy2kth4NTYAmYQp8e+gpOpxqba4+G/2at0k4MoG5cKthhQ1VsxSS9
+4mPFUF6WOWkNNVIwBG5aGtSU+hzXig4GiK4+M8P1c6N2lFc7bOHGSpbg1aoDZBge2soYu2RFkz8
JrX814lDcgDhYGAb4vc8Vkq5FypIQ6wkPNYrqZNA6gZsk7U7gtTDTHAHmO72bVidvi3N6V3EObu+
wD49WAK582Y2fKEFBDs/ftkoea1lUwLtCuNf76dTQyTlK0yHWwIj9r1sQwrzFxaOJNTEiZB7++kS
2YE8YkX3yYRwoGhnKZRW0GVfch1LzJThvidsGZHUTYjNeQksj/VlXvJT5/qP0KiSswy5AEbEB4eE
MUlDMGcjEp8UdS2GIeTbqNOGjBRdvpFQ+Brsx6bTvNUg0btGqEvPICZb9s45PSEvENgVaGViDFc5
B/athOZMuw5VHS7+JTnwlHrdC6B3aPJ94M1rrcj6ueYCn0ackyNVneWMxnsfJK7d4RIiJP9BabWl
TpL34nfcMVwDKWw5Awr/26zFs8XELCWypdmrbRP7pQ3rEqpzAV5rtJLMSCxE8fsVnFcXWbmlKPfK
5MENGgnO3vhVPhlLZA+DHpaGYKBUpVVdr0vf3ArYjqe/e2MMjYC2UJ4WteN3UT3c0YM9VChH8YK5
8hxAlZGLi//EhgWTjG+9ArmbiIHL6XCSdYJo/QDVXopsr/zT+ThqQjpTSYYKVqh6ku6jJGh2RZbT
YydlJJxWI5jaGBbaZqdfK4aQ3Sh/LoMZX1jGpwlZQBh4NGyosHKxem+Qq30Ps/L2MPNm2gWFeI57
RpuPIJujDaYxO936FzXe5JD0FaTtOHDreFTUqNmtbgNCupO83vqQl9NeahOAfKKjAB0gKwOHdR+Y
QCu/HNCsG1Tb5Y4rDfVsWPxZGlsNV21j+MUH+dbKexwqy+6nR39Kz9FsPx5STKl+//P0UrRiyJ3m
Vh67LeXPLNdb5biq43haWlf7XmM7LU03OuF3jBytDz8uDz+lbSU4lpc8hckOfQjhS2E5S01eYIXu
c2qvch479e4uZpx7M84J7MdiTQA+Ync5efK/CIPk3ccD5LIos6Js0FbErZW1m7aiW6ASI5kWJjCM
HUKisk1NUjxrrxQpx1lIqmiOCFLiZMrZP54x7Wg/st3kCyrzaZeN9ckXZZYs4mJDiH9ZxWhewqK0
3tbaJqRI4BNTTkjDtCaMYbynZgz1/XAQ5dcbV+IDAx0FgE17yjfK7gO4cFqVcI5bKZeNgvrN1KN0
7ABsalH4Ubuca1TK0MptOibnmlYbreBJUWse4/H8hJ+rOEUsH1KwCG9EnuejHKCAZsx9dQOWoASz
V1E94XG5xX1CUOBb45isxXnxWvTLLAdM44BvVE/cs/XNnYSC0OjlU2dTrj/yzDVV3BbrfdmaufVW
ADhKxRy2Z6wzoQoLWzlt4ogbrINjhzqZZy2dOXUeyOFE/MJtrBokbaNR9gpvsokdlS1wkIqLfs1n
REWT+Ty+DtWUUcJrLNgCKq3lKQ3C4cwoDApoyuebESGcH3JqtBKc4+IUiyYMs3FGfE0E42rW3Q7g
xPULrOkQjZ8xzrfHckAnGrDXvoEXN99b52ovulyI+DAnrSKxYJ5qphS9quY80snw38e3z/eTM6sm
/C08a+upSvgWmjkg5We0eR485VotnqCczuXGnpeDBH+obQmsx5wwz1d+j+eoitwHzEITzHQi4Em7
WDOX870ygSoiV9aA/IC3w8OhiEClU0nLZCpaI/wKfervTV9E5nydYO6p4ah63w7bGFD7VISCIlJt
fVkbfd+zn8jGh5jZLPnO2c2+qeoQAReFI6lMAGi6gT7tA15ur7ynCN3uZOvjMbXeYnrb76+rKGaV
uoU7NjwYVjMGtl0gt1betxQ9RkllumpOmdjzWC9/1QjSRKdR7GXQZ2cHbxVRpEpld7CMKIv5qpK/
vLRzIIeEPamrHYRHc/z8yaFKhSWm/HdowM3xOPz3P3ekNoDygMFrAbOB+4hYRaTYEGlf5+/0XJM/
XjGRX5DIDomM9Kt+hDp5jK3gT8JrMvbcoPWVqQ/IFEwuU04IO2e+6Orx7XVGwtdqalqiII9Aif/L
3Tcr7cJx8VBoy+Ikr9pLiK/mgV/2kWOyHeNmFVeSyyHdoLgVxWTmHvTKQDh4hPebVz8pv6aMLFuV
Ex9aMbp3g00AKIxxi6QwYdlNea2kETvaFaaFb9WEbzo0OJOOJt3Tzg4zWyB9qN7Y5vWU2ecGODcd
AIhbTec/qiSubqgPN2T2tjhKF2yTkyXwMarDscNb8FbXW4OdSMB0SqVr5xegHikKUAkidz3WTqkn
qGaMfo+OXIwydNNKMCftqANA+tex6CFZ+EjZhEq7o1FS/JcyJn/MgQSxXE9a4FjWFqB7jh0UMPWE
+GNzH0IwZpdcNkapzsdm/WPx1Gt57Y3F9jAhzlCAgjqaaBcEgga5ARrgzGre9bK7yZrQkVgYdEdV
Moz247avWT/VoNYedZlhUaTb1nOA+2yrbJ2qTlqfYvIy8wM1MPvsmj/dDh2qH7bi0dNY4ennHYZR
61FnW8fbB8D5XFiA570R+Tff5mRkBbajTljISN/QkUJhHaY907WWrz7QNkljU3JX5s2WWHO3uJdq
qjCWt4D6zCgcZOqXTtS/xtLcc2G1qp+B7gcfRpadDqO2qU6XxMRoVYDO0HPIIZgO/x4pdj2Tmpfs
kk09cY3NiHX7sUldVa1TbKAOujVIHCsXgtieeMVqVd0TNGICedETvHKUnTN9vaz4kHbrz9cn9kau
cuaVtxs/s3thhxbn+O5Jg0wIynbo3f1XCg70H4yfjfm73Fb3oINKsJ8YyY8FuOzWlufDVTVnbjSI
nBnlW1n0R3dTzoG1sH+Nl+QYOSo1rrxt2BB3cqLh+RK5HYvxsYW3Ksz12clArOd86YLwh6XV+MpF
nko6zvYAOzBUG1B3D+bYvB4CWiAT79Cw8gZe07L0LNOzQwbJhD7upcz/CgPxx/VGcMzyZk2k8csC
M8KfAr9U8NOGymkLqsupPdZ7Teuch1AH7Euj3bPi1HbG6Q1WqYb4Dd5l4G+pvenMyb3g/sWZbmhS
30LLZCeX5UpuEhH19YlR0j83Hl+b9PisxwdSHph2dbUVR8b/nomkJdA9wMrPCnwoHhFgBHyow/0n
sSCLU8wtEJ7kjUDaBGN3ZngMUVjkJW37kJ0oMBYBm71OY/dnid/YU1QsmXQiwxkTrh/JZqrZvko9
B55eNkHNbuSBWzrgJESRiIT0tfyY9F9ZZ4rMptva0aTxsqZ5gu5AyNrLgGpU23SMM8TTxjFmqBHQ
kvbhlRmUitO05qaFUemPP0TfIYFjPkXkrtdigw+Im3LwjAqLu8OsslFQOI37HOgDIOuorO3rCEcI
0Tq5HJ7tdV1Vgr2i887KsE/ghDCe+SAKHpWWOwn8Yx4MHVyIhQQKzrO9uAYnOQzvg/SgVwUesgOy
EprQiKXn9oBXi91fbhD2dA/Z8EjMzghOXhQGgM192jRjyUp2uIorkI71rwCxPemSpUJqLspcX7U+
zKROZRlwDlilDBZbd6VFOQaVt0TjlvMaKcuKdvF6VGNCJDNRhZj/f9KnTzoHdNy3L7yu7tqk4czM
D2eTLUBvwHwS1ZsNO1tTiSjWLCc2AbgHBwv1sW6ZWz93/l45tfqQpk3n1nCASLGUhB9Hm0Lb1MQY
PKcWeFzDd5IW53zgsSJaPzph3jaQ6Vppar6Xaapz5rCTKSVRL+MUd3jaVYabXq1NHFjGGeKTa6m3
bncgEWRVI+mUlraKF8KipxFF1GaHIcrLPLqr/u50QvRGTIqf5NKVliiG3YlWK0ZORV9nyRyc8G2I
Svpr9U38ICNt0NpHt7g5vgyhgXbsG6NW9MlCwgfUzqd5xDX4oHtsS6J7jRLVi11HIFWfYKvOYNNl
mpnEN3Ewq4J85Ion7A3VDwPRt51PKM1J8jGPqcusBq/9pgcd4wws+qIEpNyBu2OgLVsc44M9W9cK
UTSTH/Y5css/+1cbUcqJ8wOK3I203Eh+bFamZo1xCrz8Uii2P2bvs0pYRP5V8Y63iNkwPbt6hjgA
YM8ELPnXvJOs0njyGpg9cq+PRLtjEXEQRxk8iE/IIHDTIIG8qJRWnt6Its6hsp61LGnzLZV/GkFc
LPwXrfyW+CfUpK6kL7M5fg1SpFp8/iBS1qotQ2keRabJO8GhtuS76MhDdB0HEDcW28Z6A215Cjbz
afuRTFif2g90uRpjDaw7vdMqLmcV+LkhxNz6pt93maNck+1wyrt++FB4zmkJWb3jAeIebKltBw9Q
M2ysW/zToW6hoI/kbqrmWYP5g2sYV9bIaUf9lMUzsBRJ71y+bMVflx5TGyn56BeOVoSWynJbFTD7
BAcvvU1M3X3kUtGlrilddO9liy8GmL7g9Wpwv8j9YDPM9quSbKjoI3sll9JWSoIEsmZvO6NGSz6g
tQIyiuEvj9TzsG22mDFYRQhyysr0ToMKnJpc3p0Vv6iGtPl7VatRzT9dgv9L1pg0dje9XYKWxLoS
U8txVyDbup9KFg913eqMJtDmXcCvgO1Lqe3GAFs9JlMrLAZfqMkMHiSmmUWXeCJZzB5gkYTdrMoz
gBXRwy0RNeaWlrUEFCJK4zdmsn2KgMVdZY5im+DbbxpWnbd4YUXvijhYvP28ObPSE0tZRI0E5e6A
++tWfCqecrY+TSnMYNg//UNW6PAn/ITYNyu8aACZlK5VYypvdh5enxtah0RE0I7Zki48cfgUx+7Z
8BU7x00u3lL2GNqkaAWGtJb9/oYzCDWt66LgoX7mf67nvD8GdlxLgxtanj6KYZPxyrv0fSFGrphi
ats7zgkaJiiurSQ6Av6s5dG8h1tLRo5bmA2A3Hi+026QDrdC6ts8npICQLAbjo4+VvCT2zA7Jobc
zgF6yqpTF+YxEA/CrQBaIwTDvj1z4cZQrNaqYKRoqerh30Gv40pvJRWCNOEZZbVL77BvwFov26f1
/xjQzC4jfHervelrmPrDA0iMCDAP38LaGpyezNgcGWOhB8atifEMsBpuUACD6sGxuYN0ZQtU0sln
WJ/UudAOIrSOGh9wWiDlGlK9sHDfFbVoPckTgHV7+nFPGdt7HG7gTjb0o+ny1eGgYnxPVI/wwlB5
Kn9p464hNBkzy3OlHTXIryZwkS48cRqyWbYVhRGUaj8vUElLoKBhK3RgOYWsEPdw2HupRNz9RG41
nWXinXBuAlJsxukeDi38KtIfC8TmSgy/CAOSSfrq86fQ1tp7yhyinpQRPwZRjEelXxyMYUdIjrkO
BqgYz87IIUGY+EJtbpqq9E5Yya6FINuzrikzqgrJLtRbGV1tOmBAKUnnZy60mt/Ckftkc5nTI4Ez
xePhVDsDYhq8JRCBsUv7NQLhfCIPxKEWL2dM82Ry2o/OfM8RBqFhfzAWvyZJ1e1X5ucitDFQXirM
mHTj388wuLzGzsEb/2iRlMrDdwKxc2JdU+i0rJOYFJhCiZxdLmywXd4HQpCfuZTMdXme6VuHDTgc
tFtd5fhuTs6QoSWsDrCB+jSxIZ28SsAjP3EefUyPzlWs/HAd1MhllWME0wksNdGHEDeDctm1oSuB
WyOzx/EAnV+FdDpS8B8muONGQQmGgzitH1a7rif3JQxGdqRTeQw439mYNizqQxxr8ML11PnWQLJS
RyLa+hDEOQY+N/9GNxxIhtsOtZpUi04udqOMQM8wmo/Bv6uZjeX/L680Q+0byInI6Q+kExo115Cj
dI3aNCrOG2y0S/sZKfCVi+AuCCmUO07Nw6/kS/vri1EmqkOxkRB3B/8SR/DrOeAF5EwONcFEvDhs
iN1LVbW7+RBR9f07e2iwYoo+7Ff902jr2d0P92tsMPcrc6eTvtQe9ALRkBOeb9d1F+AUtqR5ww/I
xLgW0BMxCdlfn6kL8A/HNL3IW1V9Ua1F50YWZwJg/KPm6a03cCUQRmm242tgoA70mJgj6yfiEolu
yLPIJKU25pOzLWgEnG+fOM2/Ucs6yZaVjXaghLyKMogazSONIJxLjUz6B05IqGQ0DdswA6WRxyDZ
sMM3iM6L8/xjNj6o6NfE1ukUx1vrTKitlRYPnMJX7J2QjMcSdt0NsDqXnw2rM7z1ZJbWIH20mFQW
mehIB+tRy6hx/TBCFJQI9WW/lGuu+Wl0I2/dc1E/1I/7yrxbnAC5Wny/XvsuyEDavxglwkFogzpp
FYmaOgK4IaoYwzwQquoLbi8hywJUbMsNFFCdyNtlK+uvfB3ghSE0ODXf30PJo2BvN1WrCqZy4+bA
s7s2De/p/vrs92/teqPla4gETFz4RaMlfj7oCQD2Ki+ksV+rN7oBq3DbR37mLYM35aRbQ27ByFRG
8SpBofw4aJpf0XDTCPTj8MSnZYEndylM4nDFtT82IRcAd0QhBGBqHwSzNFoEvjK1Aw+4ml238IjY
y4rBoPVqK5EMHaZVmufoLQLc8FfpA6bQ4vFYxpFgfxs3mQQOy5+8gldummSUyKbCXCzyeGYCDEmj
XgvHPBPdDGnFLcFTx0BGTAibskLJVGuWQWcQ+mn67PLaRl3lNCzG9fuVIBV0f3Vu1HcT/7YhanBW
oBMe6cjnGvmu0l/KyedMIvqgLOVK0wmIpQHysXUUiVRJjHCr/bfn9z8w2gJtVtfGgA4vklcbatIq
y02NPtCM4PqoqRsqzNx6Tt7MCDfkJU4Q7L7v1UUnvcJcWlSLmvp8QoV2Uai39fEdynJ+kRVBiriw
SNnryfvu/ZilzTCI5cbDtkuITz9SwN1uXDGXdXiej2hGpnsesr4yLZZyqamraNvhdfX//zES2f6N
TieAuHgxALlysJy86k7G8LRFpQvrL+NaGKLkLa8ML88/mflvW6Lt4DdjnyUx9PjGL4mOfmlulCXC
7DZ0wsWjzbfeX/xvtk0j2UonFGjOkH29ojXbbeEtX+JkWKFUT1yyLLLPzCG2z1tXt/KlizIb9d9G
mBs3gGIX4Nlh/OQwJU6GgSkPxLabq6hzMSXQUSqrUgeGUZAkl8vKxANBwTfSdpQYtnxX2UBYVXJm
l2+W7pi95lGhhBg5+mmn1p/GtJntCNChZSAzcFxX7cD+dC+p0vkP6J0KpH64pfDLMvFtdyF3XYZ6
/2jRO8Za8/IUh+i9puDkjCMLfgdgvsVBzUaRcPcOiApGfIKmqrFdS7fny7mcxhm2SG/3ui/WwRbk
Kp+J2n9tleRRJKuqC48XmwqGvTym8YJh0nR8TbfPsdMBVsEjd3TRvz26DAnCZNcClM5X13fjK22w
o72KhsoB65VUjsPSs3UUEauy52/13Mbpv1CsAZUKqo9kdpqtgVfuJIo920rwNBM5iK9nibnWtuHh
coo/wdew6m9Pz4gB92CjFp9Nxno4lc7p6GE61eUFnnNlqp1BKJd848y1R9BVSlGtbLBm8jR1yP+O
XbwfPhEJe7ViIcQYaUpQkHAhAoo7H0JuQqc8n92Nek/ZDQ8gi9zQcU/Jh0/FK8bna7n/oCabVcSc
rol5UsUNxJ6XkMPp/ytQly3HknZUxRMqrIOfcXFDQMUT80LLdHJ/yDmTHmZXOT5pukWS/AcOLvis
7cQLDdMnngZ3j4Qyyfbgd0b7fP9MKRfa1A/BJYZVKrvxDFkSN6G2JIllTAgAmjlmEeM7CmxIwFQ8
McmnZLm5yW9X1xMbzv/Xc1xRpqtSFs3nyLNcTcIjdMZ/Ib4k7NCRN4op6YmUAX+OCNt0XxzfZDK2
5SDefFqDqe5j771Zl+fSmr2PdLzq859aomBq9hPLZpw87V4Sy+PvbfA4Dcs6DN3f+KmRQWVHotAL
a0asAQl6/kXDVYfmPEDprIkWOxDxN1ZdoH6tU8C/mnK2BBMJTTU1ZkeiRDQlfltIgdyNirOjGgQz
9xbtzHB+N/2txLR7Wt0oZKfp2wY/XRF1p78WATEpfLizdP16gsMk7ZrilG0wPWlx4IgUJsghKAsK
HSkwrg/ggtqPUQtSL2+c7/jzy+2X1ZEdHtCqreRgKu5VwtwUr5c+nHUH8g8HyPwhNyiWXEyDGTzG
PqDdxtk4OVol01rTGB1zAzvXA0xf33xZAuRUS3DpOlsJuAgYWpjFMsK3aw0nzLfFOYLDOIqyotUv
yst+iEqI7Obq0y1Db4wv0YB8NbqipthLvvmg1uDS7sm84rasHGmg2kVTCIJOndLk5Tj3aWEaPI61
t+FmMUx89sUN3+gdQtUmDNLbZP7N2g8hA03xXPOR4IClaW8/0gg/DF7Mi5qzcTisj43ulj01U77w
pctpgYwlPacx00Yc0sBTgPiXM6ekgeTk0Rylw5k2kR8Oy107lSkrLGEUbVac9NJiB6W6MSyVN/Su
mXdYQ3RVZMG2nn8lq7O2jeCgypeytkG3AnyfsFSgs1qUkshEbqCKUL010sYnejTaH2NrPxtBvaf8
MSxwseHpfTCv1vxgy9zYfcQ8yLdrHZf+dQW6pwUnSvfUeIwrIS5pq5T2urHFEeh3wCj2NqTFsmlc
tPckRdYTahfO0YyZ+7/fC4yN1Z7tzw7hc+ROKuLJVetdzHiKo0aV+rLya10sTDB1t95qm1PpADPP
XeRt7nUsqKDEMsFggr+gGXRabXY4GUZ2A8O8oKXj0BTFfW814X9EvcTV8pyWpI6Ab2she5CZKaHp
noxTNqESffZbKlt7tBGgjUNOpND1BRhJxOoToeFsqvs0H2lWB1lGmAuyGaqzDN1g3hqE/e+ry7CJ
+4AbywYyCq6iPo1evazF/GhEt8h1tU8O84+1dmQ0J09YpX8z+dZIrlUBncU0cyqNLcE/2SOr7wJF
6JUwWrL+GKjAALEBIIoqcvDdoeTnjmNrVmvi+Jo1zuFO/OXOh2RNjWVkO6ifB8pL9iCzGUzjf0Gz
4leQM7+nOlv24lsGWvoSqYjAVYrrMzr4HwTjv6lzB1WHsFssp9yk8iGfI9wh/jW8vAPIQfg/HEyy
RDzzl9M2NSR7OI42NhEzx8aYFq0iVTss74S5yBE43lu1r2PBz42pWTO4D/rYZA+WVf6l8kKuh62Q
6xUW5oPvvPeomZz1t3uM26RL954VlaXahT390aPctiF4dKkYHVm54PQyO2YEx9ZV8hkcnj0h04GX
qECUob4TUgAXVqCB5Q0KFvDwmqDi+bR0TKs/ENhA+SC/mfz0xCB4jewe2iAHvGzOZEQ1Y2g04bLe
glGAjJ1suKrmcLpe9ugv7BSbO6E44i/tAlzJjdbQqQuH0XiA3FrgVOqfa3+hTu0N3gDggLJI1j9c
Q+tuGxl7lA0FhPo4B+TlIeJSov3iTo6m8TPapsdioip+J47Gn52P4tYvoDX4rtmVetmvJHriGrgQ
VCq17tpyQMyS2wgzs+HglUaJXfwFjwM0ZjJjpYG98yNj2iibccK+DjEBqyFCHNFwN5sRWJESkMFA
hud9N8+cChLG5rCcRJ8Iacyubjs5lU//fhov6f0Z0/8Ui1Ln0OaNJNh3G3qbjbBtU5ZPrUv+ezE7
W+sOtiPzs432F5J+P7gGb9uJc3nq05Y0G8nx1AFBgJggijPHVHbtHxfflZKQFuhbfObTLBYACOVR
cWCYocwPRXQXHvIon03AXrsohrOOzUcDOM4BL+EfriIOi4t7EE0WKv1kSQcChu95uersso84+NOl
eZggSOSNE4d7nFkPsnhrGZPImcaEHhmfn7A418qr+JA73JoWlrMmN+V+K1me3qTrQ9ndz0S4FJK/
FgKozYh0xXBcc2dJFB3n+FPju6Q1qc3K8VjZ3aGC9oFQmaJ9EaWxX0WazJsG01gYr8dfB7XIyxuk
WEbMoerPvNNKIwvqomHTOhqjJg34aZsNVVz8W7CVwZzgpLGmAu7pcP+1Nhr6biHi4u/GSUHCqPwi
X8RPkM0RQEMNJv3lwy9edEtY+xwkrKrD+yrrRnnKxjYJC3+XGx3uig3MVaoXPN56xfuSYxZxPD0L
CLc9RyhYk+aMUgOXtKPDRrqbyDPDUM51kIvJUiCriTCMi/8QlkAvhDraVlgILILm+JObvjA4KH+i
kG10EITIfBmQRVyre7m3T2Uub/m0YLwRyg4QBMCZbBcoZ5EsHPiBy4JNy5Hy1nAil0DbuDjvNW6v
gqc9nCbf/XxRgZRHgOcCw0ylzYCiBykarXcVAiRTjv2z1sG1Ygk5DRW8P5DQZQcRT0mAKGgiT8I2
J16k5Kk0l5WL0hvKoUX0QcF/kpmyDRKKvnc3e+1uYyonrVuOhHhfpGwycaOhErBuRYMPbjC85JOf
sr0Xx0rPVOyQ0hvxhwdc2SVurWb1NQn3UjOVLhGQg5CyadbrOSMELijaeJiIJX2tW+LP4xI5ABCZ
ptN8RN5psgPYoCmoii9tSn7B+00Zq38R474M4FB8yIGMndU8ItGb/kj3pe42WUj+Pw2elgyQFPFG
yF9jdt0ZXQzRgCltCyAGW7M0k9o1/mWCLmELGXg9MBNDXrgHSoF5S8+VvA/hgN88OXovLjW/aIpN
0LKWegmHWUQ75/KOGL6QcyTdhFM8A9bH3ArLjWhEVglASIzdQWuu/sQQXDUc+uD1AahmlDdayIHu
2Lp3Vht06qEk2TKgt/QfIyUxJebLxkCaBLedwIdBV75YEv/FQ5kO33FG7ww2LtnGLtV0UUxCelEE
wJ9fSTl1jxnuXcr4PVZCZy/dpRuSzI/C5CQdgQIWyRvTxJ3JFeKSXDlFXAyzWA/Pq2ourEsZwWZx
77WnULcVW3JoB5osG3fPV/Xg5trrLHgB9IHJ6+GLHEXHEkaS6qml4bui1Gd1xot7aBxwOsJx8NzZ
C/COxIoN2h01YpDFIlH4EPUAFrDDwR0EQ8UKDKTAbEibrxNG65Hkpd7Mdlw5R18Mzzh7la+vA6sb
RMCL2l15gaC2Vk38O9Z7CnYHWSQOthQUy4nsNbhCNYuo7dSHOe2Jrhm7CYcbJCIEP83cUNsGTNAM
rcxBxB1ScJ2i9V62zJdoFT1yiUQRaFk7eZiDPvz/jnwGHO4OwGiNxR8sBHbyvW69FBq4FQ+ExOf7
xxew2nsVVPNPDFzq5YUv428QPeIEjVywsl5syxNjst9/jXo227tShiRozIF0g6EDIKWMi6bWN0H9
CHk0B4//jCXARqwfWLvScDZU8RNn0moIQwfS7gqT0Qu5WKJk3U2lPRP9aj4b/pOZif/WDVlLlj69
J0oCQLTvMm0i00cU1qyM9gaWuOh4DitpjRTDUuR3Wk+mx0ctXPSOxSJgFi+M/9EArLbaIO70hMq0
GfIO4lt0lBY4nwmwKap3Er2fjgkCrA4Oqdp8A7ZCu5SvSHqQS1xFC32Qg9GL/wyna0ZSZnF0ylnY
A6A6A6/DDXaQJmLHceklyHNd/BfknxpaltU3NPPXUV2Cep8sNITenXKYH8DK9oPGGm0w7+bGGozv
xiusKuJtZh3dHhkrMmVe5TPiGh7KMjwd+wP7QiQSS5cl79+Y6/dRqT8W8bjDUFIUAXIHfNBiPO0M
nQcTNpusXf+jnnyZ1DsbRwBcZZ1NFpjGJMO9Xfqz5NNHvg2CLdpZ6/SzqbDGBJmyveeF39F87PEI
1n2nLNKFBrHTyHTwW20LMmy6lZhe+AATYBLZy7pAzLIm59i/l7+HfGjTvz0R7aqIVhYUNoRPyJ3I
6Yfwnm3T1wh8+Y9cE/8brpU6wCBZKCpybMl2yPMucxC1Aez24pVom6stEwPQxTbgm/EJdbd+BWk5
1ZIEkUmQLBc1p+FZ6PbSQJjA8wRNbsGyaBFaERGIcuq+ekYyMEoF7a3OiqsXi61+ZmT/Nfu96qjf
v5MGov6LBW/dJQcmZtj8HBjq2wdtPIVl4rHLY1Hk32KsE6GcKPaHngGew4a2hMKZ2AH4PIsE6zWD
sruLycdxN37ikGqUoiFdq2SxpMYkVWSaxY5rsi7gVWkhNU9RARuWQSLeMLKT2iVQI0+OAwNPOKCo
b+g4aIugxdNhnArWC9UuD5NGEGR/GX46uUYR9+so8aOuVs/8fMsPO9miIakWjc1K6O50sTYlBsS9
cd/4yqKWIg2C5EOaqcZYN667kIhIxAUMiCIqAl6BoLm82js9/DruakUK4Tkk7Lfhm/VYzjrKdFv6
quY/c9HR2KFm8/V27nb9OgTIn1ufwhrokN8+MM9sXA889C2uB8kF0ruBspff21NBvR2dWlTaMlWz
eh5FTFz39YV3b55yWZw9j+shF+IBiXnnRzUebOcFiwHIdED1Ny7FNGDBpRlylbdzZ4vziifltoyd
C25q/wA7FVpzGig4DhI+nkr5NIOR3OyCa+cIH3QlT1A3p09CO3Ioszy+t2lXorcz0xfm/ktY3WXx
82u7eIRlMU4tBfr1r729ZNnh9Lm0vRJCZ4aBEeUnrlIGKuGCPFlohmgl84XDkCChTCQX6uz7s521
88M5z2gg89pUxBtJV5KBSa1tt3bTZ+vkC/P0Yx8CMhVxUdZnZ3wJerR5rCsl+0dKN6fm5j1XilZS
I3xwrXSiZK70OLowtXpfVTX33OXz2ibGWluT7MllknjkfHeqqoYqp2l1CBx2zikNMTTEc9mzI2S5
aMvqfwoSIDQyuEe7GvQzJA+kb08dmCy8vtMKsbYRFM5v4AIp44CzcDQWI59y+7lCIv3UP5N5CrSA
Xx6GaBky7ICZMjl4aSF0EZBVmOLDgiQ/VcRLaUxYJHNyiY5eAgf3Ms1puP57JBFDSvkZ93Ul/HEL
NGhN/0TIgkcSDOOTvFlGI7c6QCgTYMsj38eS3jDIhvYHLhB5kGdwO5s7WpcO3P5bdXdzi7uSg/CA
qVJpWBgW4hmQWg/tIK+FMwFnmdbgjYEqu3Th/3rv42153K9yGw553+e+iAJcuw5Zg3CLIOHRQfN1
ZChgyW5iqBQXriGL142x+4edZBx8Uf/miKCeA44bv5ooev/eo2FDRLdBDwCGlW35ofYC8doxIypj
RndoDo1L1UVBf+/gx04MyYoYZdfW7ECPAdYfgqe7h5OKFatbP4f/FWniPSDZKGSTgtivCfHD4kj7
Ubv91idyJv17HV49tLZnSOERJyj9LTqjzsm9Bfk6ggJ7jYaBnCOWZt9q1NUVA2ZRS8pvrviWEkAt
4g8m4y+9/TfoVW16uqgTShT6gkd2kNYrd/5wm2K8SlPw/YKF98UQadD+351aH8313/lpYvZRBjQj
MhJbXUJHfTFVXLjrpjDidzLO7H4p+ylYmTwtJMPh7exbMtQDyaBj9PsQGurJjOikpG/0IDe8hqHj
Kre6KRM3jvY7Ue5jdcToqkpjBjKm57L06MV+N2M8s87P6T9gjNztAv84GDVpF1wLMlEUNty8IIGZ
zLum8Cc0T7qhnQWWHkfliIoNREVR+SiK7bLQudTR2hFu/DPVXmFWA9Wk8lxHl9fhqZl2hutjRy+j
n/Hqp0+7+/IQLSiYORGcptJxda3PR57WseIt9vk/mhF9/vlMkve+j8s5KCA7sUWcXAyB8I2kdTtv
w5cFsmeavJy0T8Xr0yOJM9o9qpz6YWqONgiLPtz6EX5GuAUTRFy4RDJqkaHTsolrrPy9EZvmiaLN
Nv7Nc42VFx2gyKgLL6EyIfvmB29me+T1i0Q5tCJC6BR+6kCkePkovKk2ai10C8aGj12q7QzC08E8
bFa5XFvUZ81AHTGdKXpEOI/yXUPREle2QSY/1yJjxyaKMAdyOOkDuDbLA7IduRQ8/2UlzkCopu6q
pswju7uDgJkKtTzw3iRZW/wsErIFdbgXH/427bytRikzGAOltye3M+zVBA1mLtLJHR7xtGm+Wkm4
xOnIvbYzPrMUIpqXjsXbzYZ1ER7mKK/q+YxIf9xSHFVsU1OIzgx2bRZDV3ov3NeNTnpvph8rk/Tk
aGtKzfiM80VH3n3Juu974bOYOhpBRQBH638WfPXKR+NNLKSNs2dLU5bjx+huAGIbLBKf/pcCcx9I
XN3e+wfK0n5RkqUZnPRtVzV2aMumhZkgZe5NicAvk82WxXBuYQ5tzI9R803Ip+91VRIZgWitHprM
VB3IxG7j6kCKzR/gLp5r0wiJiJmLefaku43gLi0DdzgOOAbSbVzwsVOMd1AtHcdv4HlVs68QU+Wp
CObNCzfPgYhjtEegs/zuMNGm9gnvVyz3U2ef/jQMw1QZWEjxx6x7xtfX/Pl7dx485ZZyUcp/s6Uq
mMhDf+89rnaaXJ/6svg9u1wKpc08/UyUDhPsuLMZL5pmmzOv464zCKIYenzVrMv4QvfO5Pg46XNZ
1b0Pah8Bf1WSWw6M4GFaOto4kOLiIwZbZJqgaRdN0GohOB7e7hxIAVI59p3QG8jz6GK6IfW8rJXu
3/l1e2hDpiNz1EEfzM5lyWPXY1aTmefslKTxuerlZ2hRl0D3h7iYlDURFK3hemXAjRRWK7O6+Ag4
fl+hoZbz/dT+ke+gzebHlf/Hug+AKQrTB89W95swd0E41osQy5FD6b/e8FHS01OIKlw0cVxZyib8
xgUW0nwYYEW4D4DrYTBPi2eAzFNzufWe44s8HUKKTUJH8MzlSuGVXCnDAqvSLRKogO4NTohTm0hw
XBM5DLXciQhz0b/DAmsG57UBJJT1ygaotw1pnCM0imX6A8p2tKQIlSmUwjvSNUiCKreLNjRdf49n
oWEwjyOHXXcVEfPec2dlpH02yR2sWKzQmYUDq0oeQ1izriu/DglsoJz+FJ9RmahIatOnU8LRd7Ib
pjoyUaJbaErDNW8NazEdhqd+8lZPUt9SR4TKo6Rxsf+TczrAmEU7gl1/Or02y83pkI/HnRVdVRu0
QMuT/T5F7GI+fwfTDKxVsHSHUeGl8oqN3x0mBElyYav4/uKYCv/XtYcO2PDn1VxqSiR4vnKwFZye
y1gY2PgU3v83r+aZMvxsMmoXvqb8vwD2hEUaJQVv1+6YXwbDBveXq8RWpw+WBpI41Ss+hlHNlRPX
vOImXbTY3OPmeDfhNOJXnmPIfMcv8Kcor1nDyFLk3We12lIPhCc9yQb1nMLi0TBbWlsSq3cnq7Du
2eY+077cbORsbVwOJZlHdg4J+ZCviHfaAwunxfZVDmUNLE+h4B7PDM+kQGnVgCGo7muqSPoAouM0
6HIhFN4W8DGHZF1+Ji3fiDNLQoWTIz6WFgJfherrcM1r6nvQeVe6v+Yzt7/+x7omAS5GBWLKEZOb
30xykrND1x0Q2yrSUkqYKKYZVKlS2uo8DDvinlf2C/wGX9xt0HdS60p1HFbOaxmi5AbRb2x3RF0a
j/mUpHSEKsX/Quq0Jz1JWh6loFmbZhsa1opN0DvzV2ED5uiLGqUKwCfr/7kphSWMD9YOViYxj0hi
o2v2tPMlS22VvgtaF+y1de4rQSvK4Q5wB/+bbBkQnoPBGlz5BlHv2vMMLniRG8ohhiYg1R5qaqsY
L5lUshZzyQ5NjCUZCQUMzIxuV7THBAV6WbEC4RUymN/m8qirN0UYU3i+H2GnWcjTf4ZpWu8m+m7k
C3dALobHh+rHqwIIch+UqSQBLRfYS7IU88oJ8yLxypszmQ4eFI0+FvonVwH0+dJX1b4+c8XAbOPi
FNjzIyXYG1r5Ucy0evrmTBHtlrWsmM0vQGZMDfh+Iv6Ak4WVvcpGYNm87NcvcC70H8SJ8NBNgEl0
fjrLPvKLAy6yzhTicfLnwE7exCVHIKkLF2JO2yBMRz9j6kscOpMAQ8HD26oLo2a6i4Weddn37n5G
p5kdOb4lHzwMbGwbU0ievFQwfhy6kIvbIsbynw/OQX4T+HszgoO2ZBkAZ5FtkwszcCWmKLYP9WEt
IEITiMJpg6YhqD3V5Cw0E9l8tIdplOopiajIGibOeks5Ik0EvS1rN9ltRnlHpuqis7Li6E7wgDYY
3KlkLs24vVWbEa3SKgoveqw2E4Ykg4WyevJtEyUhS6omoWQLMn0pRLFerCr4J+w48976l2V/QZbm
62Uz9a8PnqS9JBO/XHGVe3hmatOnkYLNreaF5G4rSxwAQNUS5rt8I4wI8ePq/4V/Um6XZRV7xi0x
4m0xhdezuWBE5IU2yHNTTMky1UIBmoHpUMC8BwKXKn1HqvDu8SgWP3M5MDTeVDOOFL+hsaDZu5Tl
zyAPZS4TvgPsEiAGpvS8evw88Ny9Oti9aVLGyXQVK4JAY/3IpqoFRNR1/lYvG+E5MBve6QFeOjkz
pw7ffVeEhP9WjLEX0qABFms65+sZUSBflOmDLt3wknIvZjABjcamnW0biDLpauiVgzgNQsSo8xHG
xSeJvAR6HK2Htxk3PXVif2n3Ivp9JxXQjHLAgY4ZnKMJwMMH1E/Fn+A2wUQw6bVNMATHIJatE8is
6rXNLHz+6MhbFlNgGSiRjYVfr7uNMnV6eURUJ7fetepn4M/pzavxb1jnZKoj5qM9Sf/0B7GvwdEi
TgPNet7Wy8gHz7QgQ+0NfZ7H/2G//7nGdjX/OBHht+yAxjAaTXWkurXtbtOvstn0aztznLlLaZpx
4PBBMsheT/zFURymlEeoIdMwYdz/o9jb/zb0ydhf8k2NNoCL4s98B5PLtt76onCCDwHDu2O3VRxj
2m4eESJeJ7G4OgS1pNjsx4NxD0KXXF+tyez9u9tCIp7o/FezuV15JAIQ2QpTTqFEzAylumPkMaE6
EtI748FBTrdLrcT25rF+z4wEL92ow2AcAUXh1jj1dLnd55nTXTAYVSjyifUyIqkEgjks7ZxQwod3
ysBix4Ha3wLu81lKiLyQwhdo1c5ynEvvyuuKj0MyZWAfAngYxNu9HUi/LEK4Bi10nJDbUkyZtj1J
W3t9OTFjLVatwid4agBYYr2BzFs21UN/2kvIc56rPiJk++MOFw/0C7JkyA/jBKzSeA3gPYO76VRT
iGXKxjxcmu3NTNjJT6oKnwkTsn8kfrnExN6qmcW5H+vdTTyXcv1gkV2km5PTJhKh3Jy/XY1Ebsbw
qMY7AKpTbZWB4KVuCvjkQpTsHjxb7NpySGR+6jOpSq4SKMVut3JCG404x76j1jJYWwAmKW+cGW5i
UNXSipE/7fL7oPbx2Nz3qjdTDMR1D9/58av1bgEFAy2JEUi/c3glRye/0SD0bnfCLrsVL1Q+ipS8
NYotZX0h4v9TrhlRAwzavXqNNvv3XG7mub8I+ZZdkDN+/FAEfwHYeziMKU7IZJ/PyuBfQTbu0m1s
W45Eg/8VLOIREaN33S1jlmeEY8n8B+eDjUU4ia3Ru1bNMWgei/MfYZm2WxiRfG4GgmzJKlr5CXlc
c1qUqtgEdwiNTcdsag1I4gJRwr79MN+Rpshdo2FNlakcrKCtWKl5TjsajGs9DXzpuUfNn4noIvPd
fZ74ogHiBN6zV6/CHk5JkcMTc649FAd5ns3+OnKKM0AcYJ2vgJbxgyBSGQuoueSrFPP4+RstJUFv
OwG8sRgtqeW6y9xqME6s1TowlNnQIBXuas1TQ+iI8Yl0csjdvtfkyzc+C1LLTuwBOtM94Jv3iwj7
mjrLKOWtHVlYNcrMrSrSdwxHQe0kcdHBF9f2PI/8O0c6lA9TOJ9/wS9KSPRdJ5ju0JLmgQF1t8Rg
vIuPRBqhW6SFT5gfq3oKKOW0Wspfznp840hosa2KLxldrkNK5uQt/AUD8++Gtop8KVcVtWewkkah
/rG41pYiZm7SJe2QDp21xVWVFEcb+R3Wi9f2vjEPCEdpeyA0JIN3cDXDDfOVSsOKm36zoS18up53
IEdJp6FU9tEDVMGdpXavlqE0vUoFhMjlcrjs0c6TQKj0HL+/JB/9gMBVm4CuBQEF5tl2Bfu1rFDJ
/WzUEMvDsOmS91xhaqprqnhkTd+KE3JxLdmg2pULWuXg+5oqBfp92AJ7Y7fv5LockOYZjtC9VzbL
lA8m41SbYPCkhKO46zE7LbkIYMWXhPwlpJd5IFDd/hcdqgr3YfU3M2U6TbwyeZKqJ5AySMa6rGep
NeKS0rgatwrcK0H8r90eCPbKHAzSDW4dyojT4cxHi1TrH8pRlvjvzUK8yggZIdZDT962N8usoky6
tkyxqQ6zSbuMUo1skfiRHIcbhx/qVthEYLpRL3xd8QH9AmUGreh8WBr8BBXlaASy4J98KsVfKJw4
dyYI2N+mpy09zctaTlvTqdWDnk90HRbmVe2Rl0uVdp7ht1K5SmioL9dxd967QE+t3U+hX3gvZfFQ
Bq8Z6UXTuMIDq0YLdKy1i1fSz5vcoHsxWvpso5f9wglDdxuSB9KMwWaJ2QOuEgTbZWmsW/uG51eX
ac9FV6ZQlIZLnfvXRg9i6FL27nrO8PRUmeowmbNB/glzqUlN4ZwSGjK09XYmD3gDBRYKk8t2U1HC
J4ROtfXwPaj63Yb0BAvzJ/dxdWNBFhMp6notacGn/gyq737EjzIoLOtFyYuk0ye0Ux6pPyhrpQiW
5iwkV17CLE1NgZJHyJDdnWflDsJ7IaalZGhr9rInjiOcBxOVQN9S/G1kCE4zvDnlEvcJWXSpa0AJ
ipi4HqT94SgFjKHlf3xhCBqiERxT8s2lMqSflYNTqRXjKs0IOc61H52McM/6DgGwkJAP3JoYm9QN
f+T4T+MWu7BtLoEp8Rh3z0v9WV7ziaiDDWNvsTcvgKSHhJBgiVWTbxxpGm4Zf2EUNMN44o4YwK0i
vxI1TKGIA09XPjxKwj72hBCISeMYXhkRPALSklNRdaL3rOY9xGPzFRUtqXm/xeoQyhbnCAJkO9Rd
BmdOqUn8QM6K3Z1Unvlf4BbrSMaEUNjtQVOWYv5V4beNWt/JJx9Mn698dnyqr3K0CLolVKM/DyRu
A15LyHWVrC5dlemXuM/55yoW8oC5FFYgCKLN4HClSoU6IFPMroEI3KgUynkXIiS9QEMyyeVU1rIz
U58ItriivUhAyUQuGNTptRIhK3pVpK511ERamwpjvrMBkT29L6sXY4pyptU3sU/kMRADkcjxJcx4
KfwRPUn4MIALP/i41Np7IJGcfG7Whl/g4ao3B1NYngYHBf3BmDqQNpVv/C/ZPQDizNjOXiyjoZLK
2LHKw+AiLOBkipMVVeY1KPy5PDnKX98BKNAERXTxsdfcmFEvocS8xRVMUqjjmm2fajwxGurIFrTt
vB7BnQv8wvsA+TD5c0GhxYA+98rapty5BvfHp1h25/etTFxKir2jvrMmGEvJVPJdqd3uRCFgsPm4
rJJCQnIocHU5gIW7ba9gdw2VEU4MtVIBekNYdFEu2EBxROfCK7rS8EuO8lihKiRsUcuejASwdJF3
B+XtsNCE2oaYFoWLGQ8StMTrYT6rRhPhoUCt4aBBq20oWOc3SIhiLA+3n0pVO5WvYhW4KwCHLb1p
CnqRFs0OwWLd1zXA7iQ7at79Y7VJDTuPgf5AY+rIySOG326TK47vBsnGg0oT4YEZfzQ32PdwbQuv
vRvE0xDHlyyluWJEE8Job72qG1I3UrSitg6CANBUkg8OLSYnYqGm7XLXkUEuGGzTEkn/J5xj/g2q
w4bjnR9FSh2nuG4KUd0uR0TSiXJeMxNV60b211/hqYiKwcySJsaixepC63S4b3LGS7B2+WwhxGrR
yuKtg9p+IVhB+vaw98reltJt8ekdsIF1i8C8J0M9gI7wsLPM8feA3sSGdyo3vOdvSlF9QAus+4BS
uqgz7p9slM0LNABlUAtT8Opy9gP2RmAbLL7ZJINBpLHRCgbHjmQyOOp+9SnGBIUTL9X3fCmkHxeE
DeXUj1AHyDwHan46jxNKh4jiBpCvRg62GZpkvUqbhbCc3B3DhJaLDOsvToXe2uo+GqRIAVEoLCwj
h9+U4PiJrRzIvNN92f/8PBHKYzJSK/jXtFbLqSq9Va59/9x6bNCMj59fG/7qXGYOPveUxi7uJswv
8tp6WjEysCPIiNnWULDQ7hysEzFTTMeaLfc2rB3V6ONYftmEjyiuVUwANouju6xZ8pmE5zsJZcG+
IeobEAznRcF9lvLkU2KjIYTtdCMk8o4S+JblJKP5YVu2odBDLwODxSzmVn/iU/dPJWxo1jRSuavu
SfmBExaSjsQIe88u+rJmb1Tix/gcxsPYulrzxeGCLeYUgUcXhUCd0EYEmKhpv2frxee6UzZfEwho
GXQorgSW8MmkiFpdsWo+gE7LlnM7lrX86LST5NZPthZ8DTBlHr9AFQgpwcUoIHLwNIcsnkPWUijs
HX4+5veyPmVqC0/UOoX/3BJJTHvMGOBjj3ahfYlGq1U3goKAPxpdQ5jl/N9TaA9qNB5Sa9zW8G/3
U9U2xa8LcF8/9GgP+axuFH43KutXXFZ5BFGkEw1XINtvYZa5nDNm1erN1BlTUYEC0D+W0F7LtVee
2BkgNcSVXQFoO8pilRkhXBP04JYkRzdz2qPLMFyJGQ+kJdCy+9mlZeyUwX+5n2YcCUssRMUWLNaf
TI8iCAhMgeYFX7NG72faJe4gT90DQ4zZN1rwcDLqe6iC1aEN66p0eFLR+BGcdeHB1I36h+sEmVt3
HKARy6dq51zpgzqTQOQtmYLcSKGjns33cr0l16NORjbFVpYzzHaSUIsSK8iSZv5WalEDTgzuPApc
npMgQoAtFYItE+5oUk1fxewPr4yxLWge61NyccqnCAKxujI065h/wb0fPuY+c1kd+v7DP6hb+uWQ
Pu9gYsUm98tFJJr0R9vqFJW8Rt9n2DEMS/RHPtQ1ZcMjl3fnOws8w4BMcXlbDbqZpa9uGmReEqhN
Z9ruCKLteWXm/AfRv0V6IhwS1d7wnjqYumnloIEf6/5+R976CzIImp7aJW1gSXgAczobxCTDr92J
Xufu2jbsSF6WsHX8VnwSH7dymLZ6Mahk+lT0uYlXcRXr25WpvYhrJ8khA3Mn1jKu4ZNQF8eGBi80
jKUXXYhZhv9Jrppo3Rl6ToVEt4WI4TSliJh2UW13YpJt2sT1kDBZJMOkxpEHHT5GJNu7N35kLO72
xOU6IIuST1jyT8+t9Vk1MRFHjgs0Hq7I/QGqLnUHIxsT3fjZjciygb5QJHrggkW5I0ZXkudlL0+V
EEsr5h7uO4aBwHeGttYoMWD97NymVhYl2HSTYZTWBQBQShuXTGki31rTqk5mTKoS80PBjY5iOC+p
TGOK2jrDVfacx4q8fCm9xu0GPfQFWnZaxvHLo6F/GyVrB83g8/x01PsQ5SzMFabjoolxejI3ulxK
H/CxiZPIYakjMCDISCZQSwsc7DQwuzPOUPuIRl+se1N4hffqSUqfJD56+Qs3ZUV4meb3swF5oSJg
sivoE1sTHjU/06bJJv2oQAJqFqL39ZBQNSbHSi3Rmp8C+8vKA2lK1W5smeUpLbOzn3X5SquhcDHX
xsdEJ4OQArIhbw8TfeAiX3uZ/LX+uzX2VZ/c5b/uleA/188MPd425f+MoYSN7x71NoFZ0JGshze6
ibGd4qTjgUD7hrpHtTcQeMdD60MSqXkNeq7BO9sRN1p6R+T+LuBChA1imtdztjHobI0Cnup30Z4f
RKRudQgXoN9b31MZ03PU4zq7KdS0M1Qn8bIBN0AB65OEJM/ihlbUvb59kQSAjamdIULQLYi7R3tm
cPwChlQ8PcR4kgVSrrp5lRg7HeBCPWn6R+RCrK5kaFvfohUIfqQp9RxKGYSjAUXkCPETUbz5nLOx
dMezUrAWZVli38yNXqCwu6UgQqlX0BujGooTVEJ+guk5qVKbGLR2Gm0bpwYWir0qlTbQWwzdPeZU
Hd5F0tK8vi1Rdn6vgZCaJLkihgVOD1hWSSug93VH7MhMkk+Uv2AGGbn1hBQr0TWA6D0a2bieDNMS
pQHE+ZTeZDRt9Dalh0j4inPrKYnForo5B8YtuR4cqeQ6PMCtBHgNmg+g2ydzNA1JLv6Qwt3sOp98
hrqsjYMM7SCV2laF0H4Fg+xDTbPE5jThzKhQcCc9mIR0fEh7mPh9JPcTb85MG7ZaUYhE8oSzz2pr
WsewC+YGvDWL/MVS1usYJgmc5af7mv2aFuAAJN0X43/SlevLDHCFMYBm51WD7FZgs4kJfGGJeVWq
ksdeCqHo+0l6HsK5Kiq69bbPO/HGopX+rFvdu4qgGFFo4JVgMlIQ+jC4aLszazVraFwd9vgoAgcB
rAsMxJUfTj0f0tIdSkhuTbMOYu3qeaY8d/abeds8wWkFaITYBK5YaMPrhvQAb0IGhRtpYeElhhsU
tHLa2b34tedTEENaE8Qi8ncwYKFD8aLl1pXil1HfI8c9ujjdZP1s4j3v7P6FsHp3HQSSUhxHSp6p
qGa9HXYh2UwJlgSoGJOwrBCMxKLiEQT7Grb1tX0lpCh5etZGA+Nc81t83FzcXP2/bsYHcn3q5Tm3
LB02TKt0v+0zZb4Sr4T9yhom3JYPL7h/Ec0De7l6gGn7VbqonBvFyoDrxLsto9cRHZOcukO7JZYk
QjIEYv27btgQ/hRJDmMnJdU9tJ3Tiutmkd1wSXyRXXNBdFPyY7EL9WVqWI3WND55lbX9AXHjQh0F
BOT43rFNxzwE+S67Xo3UznW/LxCnLUyqH0hBRVcA0M5phVwWjnKLbVO540+iubOC9FdpT//xwXzm
Vj1/aQgGKyQBSwVEfVzxHVeki5s+YriN3EaLznt8f5o0FInIJ9OpTVfKzu2tbaQ7Wyg1AJ43FoIx
NXfq43Rts5KtxeezfZqsIJWT2CwX+0kPiHDvheLuammgd4gL+Wf5GXgHoS+IRHZhKIiLaYPDCGkx
Zl3hczF3sQ162VzZadYHjmKtv68Xsb0HjLaHwK7J6gHn8IZnisd9OTscLUDDE8xyFy/GXkcDpFID
vp5jiXHLK8+H1l9e5QcF6Py58bEU5JyAwD3BYyBXscE2M0uCepjAlNuB5h/zYPHGhS2nZ54fB8aR
O28j2HjcEs8Uiq3I4pQ6RqMSENleWUWjPjQRH/FasjDbnv9wB2hYA4Lf418DYCoqD+m9/diV8VJo
zW9kF3UWYipX4UNnDd4BrTSASdobMec1dXheoQaQPvi91vldJMPcvqR54f3YqNtKmxY+pWNfeH4M
7TRTjLnlCBPo8o/S9NrxSIFQz7SHw952t2mp5izZNk/SaqV6i207xkSExU2XGWRof7UN7vNFbTAR
EqB5vRlCTirNozeEd2s7iKGnVupA90pU6FWNGrVS//3SHjQ0nuR76OJBRThxk7CC91fJEul7/+8b
H+R+KY4NwO8Rx02CTm0LqEx8w/llNnG4XJFcnDxlI66Ty+x28rmxQOVsygMWS7cJo143VjG2UnUV
Tf909YnC448FDx5wf/ali9o77bvK1uylZ98FYMQBF+CwqVRF9YooavfIJBuN8xtLxrC6VtAP0Uam
9lhsP369wbs6rmoY04oZpU7bwaDINsbtnXQKXxb62SuuyJKp1AcWVVcRlJxLyhWfQY4qAVsCdw1h
otf3kVUFMqfFfab/tK7gaXzhu88cddSdhHGiepzMSSiJOD+4cYKJonUVRkfmHx2taZvY041ZsGaG
L2tIL0m8c8R3XutfoOgIpNho4oxQ47nUQZeLC+VK94AqpIAPloUTBjMHjmNnmPrHHpvraOVx9c1/
+1stumrPiO9qWe3ZqgE7AhBQXioZrskFhPVfnZXf+ODD9EhCGxZ1yJtznJKCNZZC4LBMQv0bcWOH
vmufflW9R8U+sJ5ZKUl9HwdMo9N3W0voWiCCH37XqXSvtm7BV9KAR0BRJUfEVCyUtIl4RExV2NXd
/Fk9fFfZpR/9nGwdm28/F/HYS2lqXUmcCbIchxSZFSCCj+h9xvYnhfp/gyv/4xvQ6AJLNUWyVmVH
FIMNWepbvPdooQQvBah5W0/vzRa8CMuJVhLmfE5G1evduoS0PTGvM8p3V2a6zOMz5Ui0RQibOZ+I
PdHKYyJgr2ckivMVbdu19m9MgB8uEda1LLA76roOJ9IvnaOh5XXquHTtLE8VrOjS+08/Ozr+hUab
dQRviS59WstARHij3yPWcsOIcanvslavCtqn7VMloXsGfLs8P/Q1+cSHgIlCM7ehwH+CWqq6+Ehk
711g+LensMVSizpi3mRfwgQJcskfT5DTEvjzoC2kuPmOBcIldHSvKnlhSuoR47LwcBXZbbU5JnSx
3cx3SyazWssM+jnLIgn78sF/PYZM5odJeeeLOFEo+EgmYRB4mSu4qddrxkNbLzCVUWVMH3jWYnDN
aWgiCs3EUXckNKYnFzXXOydPSa7lFS6S+nNzV5HRsSx+hsOdDJTPUHH7dary66bQbc9/p4hCQETV
mPFZV416XWsLWT65mlL6geiVCCJgAulKfgRWkQUSvEtpStue65SrfGP2MMdagDiEAiYRjlbDo1J3
G94slhgmXnn7dE74yqDzUNh4i94L51wXIv1TbI6U/vH1JGfXIEq0jfkrLYalIhDzDW3t3WInr7Vd
vF59dRgqUnb8cEl2Uf6NfmAI71iajMHsMmCqUySmPjGCpJhePEfUD80ab4FqPbpi8aSTaaRKMzsa
8N95El4VxRcTt8CIf4qhh4XFpSRc//xBQRa5t5X//7Cn4VKgpsK+QiIuJPN7AvKqMzUppvYwJ4Oo
dVQHdnRRgsdJSk6274rf8LDkMxJ0mC8p6l+XzfROr29iePCEna/slT7/69mj74NWq+cnwbP/yDW6
xrEs/6aoWUNZriViTPHzACQELYW5VkkcIvd+LGBn2NQJIOA0R//x7ey86X7g470+I1yWXH0oyS6s
T8wlckysEDI3Z+r5tCW0MaVNwON2EQTrxvRxUgG8SCtOR0UYF5gcWHUYxW1lLyx29OSfSPbeRV9T
CDqIgJL+pdXZ6bkYViNNwhF38qcMHaCJB4iUORVNWpMjMQV07eFolDZXi9cjz/d4sDO+UGDVwZ5k
hvO0tpyqnAETxzgr5hlil7jX1gLB734u5B67PcJ9IgKO0YpD5BxSpWead6YJFuJD+RiWAjheCbg4
G5wlMRsQzML9WPYp2CcarQasBOAVZGlGKtRytJ+YDJVjmjfaIuhzHKmXQcOeSk2qzprp1+uJ5S8Q
egF2equweC0j87+ANSn1pRuWT+te21X2vqMu+Rz1sc4GpqmSkAo8oae6cYSeweEfGUAM6M79V/5G
t7TM0TmAjRt5CzDlblvb4R7Ge3cVvTHuwXUaJft0Fe/xCsy3f4CPLbnbeZ8aMyQLCOOB0c00w1Co
gL+oSD6f9sVB8mbNQrePtImRv6oGEctJtgtO1KEsm9ejeg7rB1luJmhxW1ndAz0M8jeivssYj6Dl
QOHfuS0s6h66nF/uVtCBC2onmE196mRXuOdYMfMOQBZZeqIbDM5iQQy19GSfNsMxi8zdzHasksyq
vYIT+Sw58AX1gIxbvSmXL8FteNySI8Bj8eMyAWkAiWQdPAMTyqc+a01ZWxYjhMFiI7oZoKpILW2X
59zma+BuGlw+A+p2tHblBhdnlvi01zAtUH2axxFIIVxEeyz6lbj78kN0DmZlENY4C84aTJZD+mDd
VQB9gQlXKxlfu7UeH3sxdlWI32aDXt0PoMP/Q3o6WsiMK/a2Tj2aPOXRWqCP35RmgM/4BdRO/d4/
/TKWefUDz+kL+s61HMNmI4oJFbXSNz7rT+AZr6OD4+uVobR05gsm/I/50TxCJoL9GVu13i0mqZXe
yGcyv9/kIcgWE04cUSxAB0o9irFYBOjkb8QyJgUZF2R8HeuyGlbNzWomPIbMQZsoI/nXBURf65Vr
sumVqlfWbZqOUd99Br9+GwP/fdd0AHjga3j07qdBbsAQE8pJDASfNCfoDYVc6e5Php342MHqPt5T
fX9Ov1v7ZpKAp1MD3GkXS4d/CLlv+wAamDAy6rRqRz9dAR9RrIJZ/qlUUmEeGOdE3QMnWxfLV8vD
T1FUDdKu3K36CczSs4OJqr5a5HlYzqeF1FTKNXrda6NKJSQgJEH39TOWbO+YwWCnPaPMcuMz3Ny7
aJ6NjUbsqvzKwC1lgRPheEXCMNkcVIYjwiTow2J7dJnqHBwqnlCFo7FPMlBqiReoGLSEYNbk20p+
Rt37Zg0rT/JjkzYlMMdwW830T1HRqWsHNsiHiGwbbiR+jlDNeoKTg3ZV79XCHzxR229SUOXTN9Nd
OvNrl8PXbZSGDYnbSGo/a5wwhY17MKDXpmiCeGyeun2DIiGfm/L0BOkOh+UUG2X5nh7YVPgS0h+g
yCg6Xqw1G4wjfUK4x9vW9JWzSVZvW6ZuHVbANVqogyc7vLhoAE8U36L1AjOPLz48FWpGi+Egj/3c
jEaaSxclXubAVkRn3oQ3HQwgpDZ5tIret4QshyAdKP9tbNtwVWJtD4KgZOEIL5Cn3STv0aEcV51r
6Q3iv8MdP9vuRxko9AavzDtaYVxlcMK48MUubO8z+IYNiJi1WYNpPWPniGtdocwjMGULLXsalwKQ
8C0cHBCDfc4b/n2PuwFIlmxggwFp6VQvqEKwUQMYu9Qmf/21PBiYZzrUsoIhcvgFVKe11F9SUh+U
ZHNTgY/ej53HIjPGDu8TQTJY2mxJ/85GdLw507+jsErJl5rdXJv86lxDA5SGpOiLrNrFtlZHclh1
ZhteKC7nFl42pkl6MLMUXoSNMccp1HO0O3Lkvgty3doJBeEvnjY1ARfEfOQ0BcxFddNmlk4wwmnm
SNcnRZXXcpg3jut8ExoqbXMANHujbEzjwvEQC2AFXu5RAGcYioFsQFXCW1bF90s7aiD+KWOJNw2T
6q5esFGh0p9gFBknzzxxTKL0dfZvDdpLrVtCQ8W+lZ9mmOST65r+zrcGYkkl/WINcimcO3b3QuV4
KG7zuE+BWWRbBXyY3o3nsLhc4btPsQtdLD7uC5p+4/JlGMhBubwI3otiCAYNbiG5CWYzVxzm+neF
0+d6sQPhZ03EG1OV7O54EQzyPGrJcGjJU5bpzflVj/jw4k2k4xUo5rDJ7VeHsjDQFVkAWljsZSS4
39iRLnpjdhXgzzUACVQF+rSl9rJYgL8b8slEXh74tyZDjJeUUmnB/D4NPrfMeRTBR/gZhYh80aeS
HTsKgzoinc7GYgT6gRTsDqpG6J+1llTVXEnvC4sFd82lxNi/EIB0N1oE+RUX0jLL+VuH+uhKuI3o
JTEN4WHtrAM/tR9R4z5YRTLg5ZBBU9F3Ec0+6yCuN7xpRUxFwCFUVKd6T5Bd2z87YDuW14eBTPeK
wJWtRXzjfBQizuaxLOkY2QRZIn1MO1vBvmVEou2kJM+5+v/ZL28lRoVfZjwxqGPMppJTLNjmYPO6
a5/DiO+ApmRXTTU48BFnT0OQygE8WDVgSrOGr4DUp3XnL997rrocGr3yl8HYSFLg5lx4aVnxI4db
revgsT9QXnbV+lQEs99vidoSqJrMAn1S0QwTUvpNnPWWnXA/ZSE2jToYfTnEdGzZNgOF4XEH8Ee8
JockONWuDIp7slW+liRVCNdLKiAWH8451PrEoIYonECsJmZ2ZjzLoBJOPQKdaQWPsVa3mDxJjl5Z
xDikV71adh8tTOs3pe3+fBSvZInIv/dg+kUwA7ZINw9eAnSVpM32/gA7x6WJ7y23K+XN55Ogb4wH
p+hPNDj9xIMj+ucfZZyRhu3um9sSZFs/RVusrKW1918EkqqOnBSEXeDm4AMPEzIFMyAWiPCzf5o3
+V1jY7Abh2uJYsyd5ycbJT1cRmhJA84E5bvAwnpIAva4na6JTmjAhhIjeT0+LzBDdrdJq2/lpVTm
Rl/yJqAz5r+6yIxhvevEUstEnMW8q3yrK2foesnsjvFguGvk7LB9nK/1kr1nUuOIDSelZuDeOD3/
QB0R7NIHyoEemBOu1yYAt6052ODtyDE9WkkFGledrt6wLA4pBqqIHFKXzSn5VSrF3IB6xRZ1KWWi
jDipLDI/fgxJ7GbUuQBwA6HMgnJlqvYLyxkinsBHrfj6WXgkBMHx9G85raHq0zR0sgYLSnplALO+
pfa3xDgKErS9+guVs8n6PwDYpjYnTS26r6GH67aGOTyDV7GnOlrFotLxKabrYq+QiVdKPOCrC8sC
gApHinKnSn3jaKkZRlOpWIQyn7UqmSk+gPU051YreEdNwSuQUTbVzub+0YYCtyG7GlIIfXJ3haxC
BOglgnxXB3lAcaCAZV95UInUtQBupdUVcA2qxSentg7zlO7/GJsVRdv3AtTxVXlakPEiw1RWzCX1
vm+gwp5KoQJyoHU40EIL0KYfuA6Rojlj8dI81+UnKNEc2UFF1ypvIuqALvXPgGWkIVH2zOWIAfli
yL8YNrNKJZKI2v7nq+FVEo/GyFiLwwWdG5LZ8QXSubwnjysBS6JYugE8dLCR8OBrhS72P8q7KC+Z
cjnRQKqaoQxt9KI9B1x4odCLxCTJ7Q32zyrvmkRlkNjHO2hQ4qX9xONaSrKzaeBzBjOfEdJAKQQZ
WkMKrGgJKlna78XsP7CSHecyqjZn6iIerk+ewJLBDSmWDQMAVyPbbs4Ti8HvX68Nj3PKJsiJTCNp
clvg/rgMs5rxISZhdFnVzeX8jC0gLdn4v3X1rHxE0hCDD070K4Ohjoy1PqqFakLqApKD4BkHGxjl
MH6TJzAU0O7zaTjqvi+NrpOAVmXFkIrbPT+7sMr7yCYO5ZnnzE5scOu9E7A4P8IChcN5lwUvwHc0
V8MGGNv9gO7lo3cOdnDElelBFc8v4Xj7tYsLpXmTEGWVn+JQjcsqQ1G5hdH3thW2geYk75wgGdkm
cK1EoiWweHTXux8s5kS68/gToXoXiyMal+j20m8BH5UT8yGA4s/q1oIXI48lUffTFxPYDEyfs/Hx
ac5AWw8WPf5r66xjcn1I00GoABdQ343A3zt4cADCjrh+YyxdeM9bTkttYPTT3TMaz/sFtNm30NDf
Z7T26iyxO43y1iHnckcfBknn59+WyO3+6pYgGK8Ns3Pi0iNAvdRbwaQeqJppbfHVFVN9fSImB8hV
lnFHEdmllGLxbWcvLGzfhZstdVnJmFCBeO1HR2QB503HZdLvU8ErYAgLmSapXw920ZSFZjMy7jmK
ii9wI4DRuDSDRjT7k4jdT6M9CMiTEOtSaayz5Qjw/Wn3W7Sw92yew2fVr7Bk6D/x/BsAtApfDsBv
t0l7vumd9nWdJXQR5vrlMNMitFp84b0tLqZ+EqxEnZwgksj74P6NJEJIka5gFOYP3vle1aMCjhej
V6tv31kVPJmWTGyCHkE4mSIR9rFZh9vyeFKAxuAfq6etxzYvJgYj3aEsSkp2A87uKpJRYe3FVFMj
qg2uA4LfmQjYD+i95bVXWefQmCHDcXgs1NwYfeM9iOePfuBGoIzCE3k5POjgwz94/TgVpb2qzl6m
D4rxPw2SA+w+E72o3d1+D1bQ842rDK94FxAbEk8AK96ucDFOrXgwenBkHWQ4bQxvSiBo4BtDhnbS
OxzjTpSysrXxldP15AhB/gMAC9HShvTlq1op2qdNjk80Rojg6Vyfcivuq003Xpbnr6cSYJ0/j/GS
bh9R3No0UNAOzPh3S3QvjrpJfZ/5jkkTrN9rk4SFOifY58B+aotD3TEuUHqcmT5YEwgrziN4y89z
yTS1wIYtx6OXM0rj0uEwBamXoVUIBMBOzIXJNEOxz3xJ8OeBEwdQZxLLGOqVW+Jv5vUVaZiE83+Y
lEqOdeAXirsoGQKmgnTWFWYS8ADQGxdLVh0fs8DZpnqpe3Zi6+PXvCD9M/5CDZfOclvRWeyQzLw6
dmY06sMlroR0Qsc3dFih478vrDd217yNBR33uo73i3GsbU6vJ3jB+YHggx2DnKjgm7huoGluN6QO
SbOBOJjTgCuz72fZdCAeL1/392pFJXO+NYWCHIfS3/pEXuIvOcUTe2iq7MKcCGqEYU2kBsYO7Vzu
tN/zk0rTd9SGj5a+DZn1HRIgwh5Kau7HA32jN75JVh9G2gSzrI1QKhV8OC837jSzxo7ugw760NA4
NNtQl+1susq2XXlpvh6FFi8efj5n+hV/A4RiiGs7f6l0nCb5G3QWhrXbbLce+5oe/BQutUqRIJ6V
MQm5t4KeVrqv14wmlqBfAfqokesRFvrEjPEiDMk0NLX0AeG0FaiEVAXTBX8q3iaEnHIiTQRZWijm
coM8W8Xm6opxJqaIYaKn5FBO1TquLsyNwKHp0wHcqR9eHr00pp4o4TMtWI46xbKaFcV6gnk+Cx41
GcGRPXtXLufzfyGcip9NSDa6o5jfUygoeWhmupLrP0WUFxIwocvfgZjMVNdiLO29Vk4dh7QHIQu2
V/5XNhSi0XOViX/DO/3dHYKZKO6ldQFjNyPwPceQ9S+rW9/UgaxN2k61lCOxJVtabZHUmVo6P42t
8Vl0rqZNr1SoJOae6jkcpVFMGKekjjNVaxGEoY5VNkpYhRoEVfVs1aaJB2F1qrZ/Oby+Gv8lS1Ja
VabrPsiZ048VDfE7dE6EdX6AMro2kyAePwnqeBAJ8A5v9Z+tAC6vpROqOtYaoqMJNfLpdYiyFCaX
m7AXmsdwq5aJxm0fy9i0xPK3uZepDejIhptOhbz4t/2IxZ43fPR7V0/rBGClo3qz1o6sMEcj3HWU
Vg4iqk/nKb/oiiT9cZwk/lm+GFFCRamp2w6eUAUVP+/Tn4b3hXTYm03ZZMs6EGjO7ST8E2lb3tQn
JNoBHlCRIlo2EmdxF5ZEkZUHrXswClMbRvM3InKDa/9liQXzYjfIXZMHlxp3ArzNoGVwBMN8TE15
5iWFalCUeac6+QWZAK4RKmWwGgWcjM3GNr/ZBwbfBhPPN8KOTjhy69eYId2zUdHcq5Pwt9NGxD77
kSR8Hic8mK1kEoWxEAramXmor7IObY8h0+sOutDzIzCCfj+yIo7TRK1+bRccQb9Q4PTRyJm/KmKe
I72Xc4uZj0OAOeQFOOFjjAplDr5h6tcocnGi8X2AMQzAH6EB9IM46j0/JJGt1d4Br9lFNSXUvqxw
I42SZGjrfYtLBG0TYhm7yBshiuQWfrbZIMToIGgDIa4JwRAIOCQck4RTfg/eEu0rXXMDuOr/eWmB
y5h6tbf/MJK0hMQDoL+R00ncrRiKPiKqefkyAqgJe5zBolK+nZOVaAtfPLaFR6S5W+e07W290D7u
v91DkOVR11kc+vuDcmdMvliA35wLgFxN8Jhryhcdg7YGWSDHhfEMBG3jEuL6gCK6ik4U9hnsepo7
D4H2lhLI5i/4JXwG7bOXWEbzFCvJV6jJ8kpFTu1eDl2s0u88Wxszy6uRIZnarhw0MBN4F4aAJyRM
eMeqR6SBcrAhhnMQ6dDfbWoq+ON5qcbpzYc4Xp0Npsuh/ImCsRiJcS+QMOtcbeV2j+XWPM+s8sXK
Q/WKwZzmA0iQhw6NjPiN44wvyaEpkOC3jMh5AvZFPX9R97/oDA95XRALWRxHaS/Uk0CglT7mrnZO
vMmRufLcmXqX00Cb5+QCJF/VSXTEWtGuc2rjIxGPqFV3IXVv2djXVWJxL7YjUHjXP6gbYN/ncaFj
yEoaePAyAhCVY56SY7EGS68RH1Uz4zEaGdnv1mYruUQY48zP1tnncOLQspmja7nenjhxK3nQvZsA
Rv3ammspVesOrJwvr6dqZoeIv8qfDxE7B1otmndhh3DPJx7pd31+Eg/v7JPHls2kXP6QiuSwo8/d
ZawidbeLVTh4mQRprPEoLfM+9VwKK2ReslkbCjqNLQ3A113nBbANi1g+7Uw2SWdpMvF74V3zf3PZ
N/c/R0P3CisH30cFJm0yx1Vn4YbWZk2lfDafq/iVpiexZBvSvriRwrqQJyDL3U3yJ6X9cs/WkDbP
vCS52Qcj0XLr2Q6oaRJfZQl6tyPgMbk2AsMQzVlfURsVpiwDb6otGtBRvyABsyROzbphbMFMcAhl
8Kw8JyMdNbdP8LJ0pazDD/azFgAP+qC9RewFZHUeku+PBkiobd9GJP3szax1UkJcJVkK/HWz4oLG
2wEhgjThK1I5ijPBbCIITeENGP6xMxVg6ytYoOrVVWOTsYiQDCMKIzhIl97jlF+lWrGcLVEsdNMR
1VHhWY2q/DNtrinaH1O7MUcD5YfKNClxfZF/DFxTVHPoUIA7NyickJJoLWo9PaZY86vgIUtMTrU+
Y8lREL2TeJxN0j/TQpVjjGm93i/Z6Z0vzTD4Pg7pq6NczuZlBt1i2ac4fIVjnL0dg4jwfqk7VQ1t
lOuLnLlAD5THzhDlrQFTLgHCWNuy2hCH6UhxgVNmvmwhNb08/kLaJKpRI0JOCOFhEgSz6rEwQwpf
6/xObR8bUucpTyKyAV1E7kATOBmVn7mr1fS4dYkWyUABqkQcd6O9ZV3dyGXP6vrBJIOLPrU60rzz
RhLP4KRMovTMbboirThYBt47BjQyyagoMUQ1wcldCSID5nQHlkLmm83QFHlybEnmfAqojjXaZIB9
+iORywTsP/WZQXnIYiboaeFsy3EU2GZJRm5N4qfVOnGXFCgvcHsAKX9NfNnU0QcEqVKvnjLD+Sod
hJEqVa3yXtFIb9TuFq1BS3pWZ44Du98VuXy6869VI4QyqsZyb8g2tm60FLDtgfPGbqQYuLZccghd
qEzebmcBYXttOfTZvDMt+G8SF+GsVHyeco/A21wolU9hQgsjDEaySuH9js/4HvpgpBd6MhUPeKjw
tpBnSdc0h6DCLvDzLm4chmW87C1nsexMFs2nkU44MmA52JVF9gfu71LuuiOC0LQWWK9NuZu3h4X7
Ohot5jvEkPu+zEc+yIbMm7CSgKT/J8KyucX8mjc9E6X3evUUP50uK5Hr/yNE/GVGn9ByPxjUqH+b
x2aJAFdiiHoDTulABBc/rFcS3nLRiJ8fk5zUIis44yRSfvWt3Sf1cchUP1GZyu9inIS9sDJsi+3+
kgX9/nT7JUKNe/lGyGXCcYTNB5cJAYmWkUeJY6MG9n8C/4dGFdY1mbStCMTcvSENlVwJ3NLTGGO1
zj2C90W+Qh8cTXxMTxojt+MF5GISSZOX6Wc+8RKMxXjcWqFqpv0MVagDNjFaCRz5Wf38ZgZRgsuh
DZN/D/24NIM26UpVeq/yvUEqQ+otmg0XHlbK38x69zXwVONAx9GRZQz0WKF42XLWTPLOS3rtQoc3
s1tjDDGj9Znk3Pc225AOWvgWBigXF01s4daowkq3ecaxcRnryNS8tpnlvGMyv31BKE9Jsd0s/DzP
yVOdMSHDrf0qYBMlsuAI32tLqSQ1IIojhjfWEEe6PLFSkyTYZNXazYisDWsAC1mw6SJc0196ls3f
0ow1O0cvKN+Y0QgGD4q6EU8s4yQajzPNzbjwC6W9dgPUWWI3UJLa4K4RsL60dkuHRFQYndOVpHy7
ePGBnssx/aOWRuCWzt7+JvcrVUku/Xiy9mxVlQRp7myfarWniwK6ZnTreM00pVI5e0R3KhVaSajC
AirfxwtW8UrQoqe58xTMRkBk4PD8CagA9iFmeUAETCIZpVebFUboUVy9GcSSV0GjwfeHY7rHcRiS
bFu8hgqzqUSFDZfAlEwA44fvNoPL/xJakeHEsV2H1/jyBHXwnYT6O7vGTwXzVKNRTbm1tRdRAeuI
95GjTa0vzL0cE0y1DyNgL5JtJ4US8lo49kn27iAGD4tAGz8EACGLMLAIMvfjsW4GPoYDixyH8MOn
8uDdHnDJkQNtItcujPgT3QvH5a9gY93hemFPrOfvWKYewUoLzdYpAumqnGgs8xTq9X5b/DW31wsq
RroMseUPMeS90fY4VBuvaq2TjuT4KfTPBa6qJHZ7eZtVkjyUKBH0nSS7Fht7NsPuHdKIjNPXqvMO
vQXCzmy4YX3a064myMFFw71MPmLy4CvGUeFlmQkahAdKXVepFXQYanjzoge/EEmKmJA2hWlzoGfp
+AGWhVGBkM7bIo01miL95QMKhIBdNZvx4wNr7v4o8OsJjjt4kgbHCtgAdY63r1SDlEMfHfeFvskO
W8Bq5oGmnv6mOC7F238+6+puHRN2WH5UT0zBoV8GvGAzpbsSuq+rgftdApTOnn8Tl0LGhr8PtE97
lL0j0F6xmX439Yg4W0ADhd4c9XefRBbsE0TJK69oBcwOYlCdbFrN+kfwuDc535KxYrIl+2wsie6u
jC5mitZoBuWvl8Pz/MvrsJEhD+EsCd9LyaO+zG1l55ltKXUHsIpKKn+l3liv7HTaQ1K5J0ubKISA
ulu0hvazl/tz+lm3tGWY2f9fWfWisUrp+7AKKcfidx+ecvR6RjvD3h1WHyElJKSQDABXlWy4Ru5w
R7ataar44GmWNvhV9PzJVHo6EVAefVKL30oHBIPh0FtVGGZAnxw00YPUtnffpX/6tY72VpxxBbg5
hz35C+w4FVLDaB5V0OupGYPTqIe2O+/UQTeJobyn2oeLz0WXKhwnhxLzxY86fPhQsc48ZtuOVqEz
RyQwy5GiuDiKc8YYa4zWJq9zUcHrQQUNLHpBZjcc0f+c0V/6HOSRFkYShcCUWU3ZtreTQbIjit6d
ZfzdHN/aI4JsITGPHE4/SRAU5JX+rWxc+7Hke2+IqKniBDXKoenumbFagp2rrAVhpavzb0yQtBFA
HZgexgZryvgnVkDqAl27XIKS3KZfzQWmIkhShlzd0mr8/vQmpUEh2NMBL8XIhe4xtIh369pxY4tu
XvxPKNAYNjUhzZ9746MV+DlyRANcv54M8KFqUlQ2xP+gdlL0tOpNrBkBaewaNOQNDilUvJCkriq1
jv9dv0VZTa4qzhrxHDqiiEh1WE0GeNUFQXu/mjKu5ESgQRJUzRs6EGfmKg6ZJ3prf4LQINZoajEc
JlTcWrzv7Oi6QjKFcYC5KqBO1fXH6z0XwPEEVRizZ7EEXQBomVhyZAbqSgtVRIoxZVDU81qiqTWL
hkkqn+ho3aEBohqD65oPbJl40zKDo940gxsu06C76Gyl4LBuQ2oJx0chC17+/4ySTsDEYcYugIKV
xCH6NQZF6RO9i96e/AP1WNfpcwjM3rDuvCDXxASM+GQw1fHNfrLP2ae9wPjNTMfSeLk6sNLvYEMs
T4xSV8xrh89amPCb20GSPR3n7634G4DX7b/z9IWvPxwRWZz1X4NMysbpeGIvkVWo76H270a/4iRW
IDU78Yzs3+2wB7jJpyPjDoUJSi0HrEt0zU3WV3dh+QQmw6DFHPfyGv6Dzk1dppgdd2SsAa4aI32g
JsPNLGG7U95ND+lqz2kZX9mtzg2v6gGx60My80sZPR89sthLhiLj4ZBlX+4A6uoCh+p3ntPJFo6g
A/Xa0wLUT8SrECG5ktJapDS93CVlWp6fuR4yuIHzaMHDMSQZMEH0AYo1OQUKrhc3UW+NNLhcXbUT
mY3AjTONHRQ+X/fvmarzRlTsndoQdWO6Nap3K7Qrnwk6AZSOOjWsgo3lodZqV7IdNUhWkpveMIEl
2V/Y0hZ1ekBHZ8Ixd1NUaenagPc+DnyQoyKXbMEbYrqLJXIgZYgvysUb8gpOaB2ZxjmhFPrJAIAK
FG6cjdhpkdXSKPWJRHKiOwEv0laBKQ0Ny31LznVGG+0kb9y1v0ZPPj3b2lsggLTgCLdrECOPpVrk
y1Xxd7HwBYBXxiWT6jknmVLY97FQ87VEf46iF9VzaF7ANUWXQtTLollQH6AICaOT2RFXIyc1I0c9
CblKKAofyyrv+4R6TEAXkGwd07Hbw63RRfOwUSLcGNLiXV7byUVXctfbEu3049SaeKEX4SVFaHjv
8lhfA0W00oWoSPjcp/ARpuQdMBA6VyUgafKShpmoc2jL++KAQ5/3miyhCKXYyL/4AIo/gIQXjxMb
/LOf+fIjbVofNV5nSMzgizJgdaoC/B/jNkfEUP5itEWJYL/F+b3qlEt1tKzsKLVKodJdf0DHB/7l
bLuIRzX4OhBAiYu0baPCDqIDLGiLFPgodhFjtfYWbF88MeqGG1Pz4EPreCQrxmW64tg0OoiPoyDp
yftoDP8SaSvpZ/MDPFQAyIx7vFAV6un/RYgs6PU8wzYy+f+W7xIVCw/XcTijA03eXMMpFiGruhIG
+ym5UQgdgyD/tyoMWYE05010TBERIuLbCNtUTqi/BBGznaxoczJqDzuZn3MD1HxuCoYPmSaCZW9x
/B+p6M58ZD1LEeU2zm4gNwOzNCmHNdDj2ncrTIeERSIrqPl/qdJyXORdwBACUvOdfrq8AozeKWpf
UHkMOcbYIsJmHysXnsVI+LU0FwFrEIm6jrcb2RU3uYMf8EBLmiR7Reb0RgzPpq6e7oyhaIJ9hmbm
sG6dGqtIcXZ/NWDzKZQEugqATmoQoiBg4rLB0YDmWEY4jOnw0BbrkcymUUxRb59uS19Toco7qQ4q
12TZ4WTl35e9DpHFv3GmlPuogn831xgDdDL9Y11tY5Ma1YFtgrTEXH7lCKySLUEpc5IeAOle2y0Z
Ruonj7X1CmrVCMS0bn9ai9PhgsUx2hf2avBhsiiTW/7EeLyep2rxKZzelxv5Ztfb3J4+Bg7Ivq9w
NWVPw5nqG7lzG9MbeVbqgPT2rucRX4dOfSke6e9nuyK4ALYUST4rhoERhomknrfJviYCelqJitM9
e0+l09O2G3drhfhpEgXudPKtLowgOlYvUnHim4XtNGny1kk7gvLwwpDaRCTiv1YmjVcVWnOo5pkT
ZhNssIuJLm/mJvaCZqXfNAQuWbp337GCBkCOJ9r/T4nMA7HZJb6s5ltf/xWo6P9eanNNCyhP2zvv
QaGZYw/sYqgmvHFKKz4g6psdsXy6IMHU+6Q/qqzedQ/D1NRrLfN5OJ4F6NXVDk8HdR2ChJK6hk4m
cqs9qqkZdYYAxGJLDwoKyle1v+qJf3IG7tBEW8MGlniGghvmxZlM4LpuHTwR8xjQUAgMUDdEfHiv
y+cTefSv3lw+BnJ95vXgKlEwWZQZ/rjRDSJSj9mHgyMEFzI4tN1I/IlesWMhddaopRGqb314nlGf
9L7ZKAVTfEVSijZdCUFGohLiGl0Xo39ZKDvetYmZzN+VANwfQOYYZH/voKoM/LhKLy1WhHjK/HV7
HoiWTcLHVoz9sZbMlrbMMt9navbbY0AZ2O8z+2mkZs0YI8ilyL7CSI49FxAEypqyeiPJDaWSJTnY
YhCh86B5SGk/zhyIbnY9wWtw7dDe9m/g5LdfMmbJSEazOHfZr8Uh2KKr1xfd62iaD0eMMzE5WGVC
fe3rRkxK+FAPfDpZelX1ql+JScHBDQG1+WYtVXo9CnxzGQbWZ/eieqScwGKrWtNfZ5oVMyW8Q8MI
3L/HLePEiVsnpCLcmhJdToHmkG8ymNBO3Ob4ZBa25aYLw02IXznfCpauEVVixvyNz6o5didAVufv
dpNsKISJe+/BzvPRgnP2fJn3U7KyK9MjBzBj3NfhN2egycrxglcsthHWLxqzbTLq+GtGO5VXqjvt
wYuitkPAsi2cggxF/bsnSDB7/wDuUx30ooaxVIwXgffQiizhPHdgECCNWvl7/26IGb3QtRFXKT5R
TqW/tF19MR92fDk3ZTb/hzPV5p039VpZleRxainCycYbTssXO4o5UOq4UJ94QLnWaAYTi2djHhSF
5hJ77hs8zC4iOA52s+2GvpeoSagFT0J4xQsk31wm26OWbT+BTr9dKVfMEzswAneBypAgjfJyGjdd
5hqUoqrdYYixDkFJotvNPXmuEMSF0BagUdzWYfrtG2c51wz8PEdOgUd3iaXLLGYMadovg83Qp+Gq
ME3OKcb7wrdU/+s0DzJvaUOz9dcb0mJOCpCMQqN7r0YAilOi/QwtOZtsAK6aeUWjC/dFAoKWa3/p
zOsJhcvWh5PScvryFCMwOn1qZhvE4YPb+NuUoOd1TLi5qEwAYj5C2Z3eN84VGeoffPTuUjf55kAl
3716OhCony7BXd/ycI2ZyKRK5WkfWUAXcC80PsowP2oGTLJoT7ypHH/m2i/yRJkVdiIk6NbXDofY
pqh1r7MiEiWRjhRif6tVIIiamb89U17+1P5UjMYG49o35ozWOCvJJVffGWcY7RGV1IR47xj2Ya+a
rfksPn9T48TOg1wEzqXgTWTuH+Qg5xvrt3D/w542c9EygUoSdmXtMjBtXi1O7Egv3TuTuj0dWoXD
f2KrPYMYMs2o1InWEKJloe/KgDMquM+XAPwq4MiYpT244j4QLfsfsMS5EfjtxmcJnXwxB3uo57ed
ZKi7nMU20D9HdCxLVY8u+Z3SOQbpE2xD6OI2CXF5TN6hgpRger6t/uyScuqH9JomBk4dbY2GYTip
e1AzDQ/dceKaW6gZ0YFnD+YxOIvsKt5EdPgN6rqH/eSpd1bXrtnaAAj8ntvEE3n6sPTOqes07eqH
TuWPvQfJUr54XizROjMmDORhUL3il2NihI/Yl2htrklKmvTyQ/zmfevgI0xaVPmXoEGjX2H7SAm9
hFqNzqtVE8KTwEyTgcQFBglKxmy35+WpgwXYOpLqItxPLgxKst00ozP9MFpeKeVigM3/Tm110Bqd
xZjhYYzxiWiX30BoHfpYgpqudJL2pbFMZodJulzdKbjI9i5KkKA+a4e/em3RJEBtLlpC2TsklRkX
dUv5yoNSUUZYi//PF1iZVUWHYICd/vWxfVa6GPAvinJgdWwpFEgBhbn7Jnu3GvJB4Tah8CprpN9m
mUjJghGHVpRsv+hw5Q7gs4xcrmLkTNecGe06GMVHrPTWvHI6QgYBbrZdGADjdn6YR7QZtlNCJluC
lrepuivWKvsnih1foPpPojcTLFRNQzvFL4QNky82ZP0sLcFHjHqn1c/5ggtWHWzp0Y8myKvWwN8+
gr8z4Y0BIp456wf2b77Esi6+DjTCKN8PY0zYSp38SzxlgbqPC+1GLdfZ1zKQXbYwYMwi2zBo7kTf
Xr1JMlcvAVHTfI9gWD+u6a0fqGZbBjb5/yDeLmg1FWWJtGepret9YXlgbeHhHuZLkD80JQ5rSERW
I13D3NO3Gu5DONTLKX2y7VFSlGfXUn9/2CjMpauwFXWfTyE+5zg3EfbRiTfKtrs4B1l3K42Ctmjh
4cDpxe2uKgrwAISBmnypJuIEFdFIyGI78rP9ABHPthb/1YqVtsLwmeVGpLWtVag2h3bQEszPe7Ch
Fli3+tFcCosDUUj+oHdRmIQY1VNEZcSDDq8+GS2dRCWpTUFcR6pLvWdBKKGmPtVLdA/d1xdoNjG5
AK6dEDkTlHCBL3KGwzR75MmbFabPINaSjlfQjQjH7kWKue7Y5XvN6Jl6/CtiWHZPdkGLbiNEbuVe
oh6IYr1iSuA/KIVQ0uDRWQRXdWYUqqeGutPlvQyorD4vza849wc0ZqciGIlNCIgecMDEcgZzarXY
XNfDxccjj4vLPB69qte3pqbJjXgwY/2B45f5IfB7Ok8obBzb5kNOvxOIC92MrVHXKefBRon7AhWx
3Xipz6k2Ui9Ip1VaG6OF8N+7OvkIfAogymGYqWo5GA1jEc4/68kgutasjbu5ry7FXJ3RMhEI+xRG
5U87U6O8olL6O7QU50++x/36CRCwrEJSckQuVQl74S4aHHWoZCTy272CnLuqlBox9FhBSyhQNNyk
h1xbr9PO/h+0e7wK6bI9ti79M625CxOAKtj7T2oIHBBSS0Br42JmIZwyKhuh6efeWLB+pd8ay1jq
L3C3VxxF6eli7U16qblwW5FpAAU7M0ktHroyss9AaxSMDQLygs5qk8P0m6RmYa3uSz2rW+IkIT+L
q9Ha9YYmTr9pFAFhAA2KDhnfkAa9IQB4sHe+lHMozku+Kape2EvcZT6FurOpNJDl5kmrHg2N3yXr
vBZrYV0rDsG0EEfh/B/E5f+KETVImgnWiiFuvIGaxAXxoUdN8nPCGKfME1DwVAd7Ysi32F6IoSg5
ipXhxluvTmBrYO7fNlECVCOKRdFh2ue8Soh8k6ZAAR709LlqDxlrLK2qmBJi9xqiM/NiVBqnl2fN
5NBUcVblfr1bpW5W1I3IxBePWhDK4FIWqqvXaRk/7iOgoclk4V3Pw8vFdtrwdbgbfUTMVhSUIJ2g
R0fARXXsa1+n9sXtcsXb7KhUyF6piEKfcOBG9tIKVfjUTCBIDFgaX2dD3hR5yNXzcimalJpcXay3
OkNd9gEihhk/Q0K2M+Pa+zEDd9LPti4lGRyjMeyWh8EMsEi7RbUM7m8r0XLXENfUUWUBtlAGpVal
xLXPtIsYy5KKwnHtN1B5yXn6aTSv4WzA100fLLb97/FehxiwilswIAPgOITuuRQg3PpNmPoJzRAp
U55DaQky0gp72PZn4Cqej/ap/YmL5wMUivMu5gRO/HThj1WlVFLCat4rkAa5odJvUUF7dLrUMnxG
wV0jRkrnPMn40aYr4QboLeFtZk8NJ+g9AS9H2+6/nuVUbbSjFtX8ws4hdnJq68V/FshD3o0xxSAz
Qv+mwPNZg5FLPjBCdx+eR/n4t9k2Ueaj1R2mS/MM8GGTH9L4nZlgCLpwKGrEiSMFL2vakCqIG5MC
A2y5/GjE5DA77MxDBNn14NA2ZXCZSd0geHfUqj6W8FSleqMK/aPoEblkR08dlb5FReQP+4tdiym6
P96pSp8LKSARAi7EayREIMRZvfJe//oPCKMaq9cjxvBN70HvFgGbE4y4KInIkPMgObsxRQcosYGD
PMS4RW/J9Fq7Z66Bmi8+W3ENeVQjvrACB1c0kHphZZ9+6z+cuSjKnUbLDBtdFZlL0coICNty8iAc
/flLawurBsDCPC5iE/30PR+/IMGFdaVAFeyOIctX+QWYnhlbi0y+O8bxWKmWEegT2eGOMrHhXR0m
ibr3SpPpJFJCkPPqeh9IUpaw2lyC4Ebpu5gb0m5qdu/PvLQfnfyw0nvlwpGkvGUL35i3a3/1Za24
BvTeIXnGkqFFrN8yYmabWLgDxuFq9+zdCVlYjUUO2+f561vEYsOoMQT9e8+6edgEWRWpll8Gj3sS
xyg+wCtRgxJ/Hss2EAaBzQ85l7phTlfFDax//MZ8DfC/AJhe4nwDlDoY4hV5CaCtdKetwqPP2osv
q0QY6YwXEuLKe7dF2ak3AGzTcGMcrcJIuzcCccueBabbvrOlBd6zLAoC7AwQBB8/kc6z2rPCRWp7
IJ1NyFzMGkCW1xYMrXA4usEcesEX5zJ4ylDGpv3MxLrsAWHfJY89tfHOm0Lxrf10J5X6jZXtQJQ1
LXA3gotCFuF22Hzx3MjyIP0z7aKsGMhXiiaiG0WBqw3kyRNQKtf3ohHB0iHrBGIbX47xpIxUcihy
dVL5uKo4D7xPZYZWd+AMsppNFPHqC7asbW0Uus2qv0U29TKl43NCPXCmo/p0HChsSw6WgeFY3Oi8
U07obIvZbbbScdVc+TZmUq7XCgutnjBlteKjVtvhOGrXX4JU6fQ8qw8hMn+T4hvp4Dh8+PHpRpJM
UVB1GcTAl1eLdq3nbEW96y9aaxb1p/tf/Cq7VxPMUK5pc9lTfQ8S2k2KCnaAH/hEw4xH8dz5baIb
Ob7BwDdtHCOfON/LWuqOLPolpv6tvvkToj8NsvehjZeVtyN4ES5D0s2IjIeB3gwtgUdlZEgIK1nZ
Xa/NSmBQmdB0mf3Qn9BOtmXiS5MJyIxkV6TrWJ4/0Ym4bmNpYj3A1D+154aNEYHRZcE5NqnMAIcJ
OLfLgu9ckbM5UxUU86NuhRZSxDJhzS+Is10l28bILaQO8DgnFToyxR0Y+XNd/Hj4WWr2Nc1/3Zku
2Vpn9tKRLALTv0McYmjMFX6Tk0XqDj/Adu0/k/tzIAsoQSfn/ly/YzXRfxZyeRfwNjzbd6AkrHfa
qQCf7x0ICzgG6ijepLoZ+zti4U+V8wXZp9stAQ6AE2V7svTE1z7Vvh6wQms31xJtizXk4J7Vkt0o
Kpx78+QboOJzgP9tTJvz0t1wEH+hNszxSB1aN8CKqrJtxOA/AaooNjuJlKvYWt+3V3epmYaFYM++
+Tf09WBbOjfumHHNhwbEwnpIWIl/JhcDD+1mU6Z+2TqkzbX+Vi+fuvgz7kj7o8JlzJasWrZeZDF3
+94XPxnCD6dqYjtqNvt9KT5Pmz8K+jUAY6ekqMgJHCLb7I0je/p98KvGyezpcn5rllwF6/b3pV6w
XlGRlflHU/8OTBoZg26dkLVburVUavdeE2c3b0Jchy5vm6v09NVXy6kadMS9UInTQ9YFUH0FCUAX
j1zrPNBnyo3ZY5+xQFxOdmKpxVjhwNfb/mD+yr0gHtWqkQM07FB22zhmKsYjGL4pNZ6TH98V/xWC
xz2z5DMR16Eceu1CsjMtHcThTesSW50bRH91tdDxjWXa5yqFlfsSvoWUKeR+kQrLnlw/JdfTpwov
vnjsJaiip3zdXY+Nk58rYBSTpJS3BRtiOtXDtfVJOLYF1pj2SONnb1KzwczxSfT9CM0PBiJuPfAA
Olkjtc6XgKeMbAqhNYtFzy8u+QaorFsUpWJ/jKMIkCadf70pi9M6hDGYCrLglYlP3bjZt5vapWDM
IsRXRSpeUNuqz7PznbIJ5kZaaeZsNBG/AWsRyXyzw7lGqz74fInWPcJbV5QHKiKdHZTeUbwp4dw+
MtKwgLq0sj1vrhW1CYksvVdeeeoulj9X9C/yEtbMQzkWnM1aKnVEvRIsF9AGSXUIjwt8AsK/bV/W
aVmZEzyC8Ga2N53DDPRmFLokyoRCWMQqbBu7Vo+3LsrjlHBs/zP0n/5cUWJ1llPpe5vf/Dj88T2i
wtNFoCfSLd5+xZkW/51UW6adxbFDVDIyLX/G4mssMWAunXaVglf048KMss5EDnEJ5/4koaAGyjiz
ZW3DMi3QvTwWZQbBT8DM8TTfo2hglS8VpDy2OAP6FugTKQRhtv77JvwUMbJRAxkp6ELSCdgPhxXE
sPinq0toQsTMO2ib1I9sqVU4SVYAwQu+kb7I0ENzLFA5yykx5ipJeRkQW1uMqRiFdX49Tp8CgCt+
mhFlfxrcYmCJCyjcyu8NeuoJgpgDA1u7zaNMVxDSFOz2DBpNhCZDK8YUN/qLtkGcoQk4T2PsPlWx
Tjz0Kj4762u9njJ3gMr4YVD0NtRd18yR+NUG9lzdBhP7UROu5nVy/ecvQqPw9GTW5JivbPp+0jHQ
k9XCDtLQDdAepEhVeoOmaO6k6X/wifrSv8pGTSM8eh7fEcgpvc7ZaxsNcVXlr0LiG3CQcPFUy2mH
0IVp3e7FzsqopVFxJkACibZlLqImxj/JWgOEL1iSe9KfgKaJtoWxrKiYMaW6s0mrKaBi58jTjFvE
ROd/H5DhTjOcr4XVBsaHg1Jwjh6x4rtRRW0i53hRVArpcqkSbPnB8EO8gvosx7eivJShi/Zw2ZZ0
kqAH8fLjlNgiH+bZO6IluifMKRlu9JDquE1x6o3tzsdlBZ/esouO5AkEgpzmoWcI3b0IMHYvu2B6
1ygCYM+x0wS5LhoW98L22201ug6wJ1xJvGvyM3ndUZ2LpmnYPc2b0+hmqARlOGyhCK66Qonss0Ej
5L/B4XPM+Kkptn9cXsoo/S27laiBEDwrxMbYGjAc4CKnuJM6d2xM3K15iwBxV+r1MonODPkLJKVB
AnQgqVn49NTcs0dA8cfYSB6vM2ytJqxSlWZIqR5/1JsTsYhmyQdieowmacOiARQs/xBwVMr1cPeb
KPc5ELN0/vSd8WxC1g6Z9xBleApwFQ/p5Xfg4jmiG+RYgROPIpX+EeA9Wbz2WmCe06juLshqxd3F
I0GALVh3iXMH83m7Ho3CWluByDLQ6NnjpV4jOxkN1F29QtuZc71BQrgv8WiWqNe/yXlinD/GFJqP
3d6qGKidJEG8XpjVUXUOSJIrYK6YHomeHaaJ1+sA1fA60B6/IzvpwBemxrOjPkoxUTYmDhB0ULaE
JrQhLMs/onbArAYYsDD+pw+Iigbx7GSj5VYR8COdEvxnerw5aSbPZDaP/J7XzlDPsMD5/ja4+tQR
93ftDj1RS7XqR7Q61U+glgzc1VOXGAqVc+bfzUsg8b0H+6arE7Jaad/9D/8W7wnqIK/XZaANfIYg
65NlliKTOvr0unV7lRfXxo8OgRdUnxQvnTeorhXILhO9wxbYHGiISbczoZHCOD6WgfRcgRXECihA
/BpblSQoy0u3nu9bYNMTU1Aos66CjPwMAADEISfzwGxfcZhIB10wTgoY6q4NdrYgYh6qrruYK5ie
zUTqRg/ZQClnySZHywOAh7X9mwy9/D/iZhEcpQUsaL+sU78vOTPc43xf7JhkyHDb2vuP83Hl7idf
aqnd4kgS8jVS/S4JfvRLpYksywcFevtI37s62bcgtrP1Cl7eInVdv39Qq/DORvhHKfJG/r4BsIY2
RMU2f7gzBIkzRsLVN+ynCTCJuSv5Syqekf0SWfzAgeoTQz6IAAR48qGfxERYDByO4dsYEVrbOwAm
K0Y/agwwRI8xjw44HV4lRoAJOXyDfbmJAcKK/L2ty+kxAN6YHZr/O9hGAxRBCIQwnoclHqL2OI9f
O/xdHynjW5rdbKi8g+Whr4GAUmyguSm+alAMchtjK5bgb9/eOmSYLsZCbSpxh3xf8dQ8xX2rJzXF
ZVXm/lnwaxkBQ1vOfeqd0MHniFfRY5u4/st968N3XXF8VFEikQ4hUdsxmRgaxNgcNWhvKGAxGZnD
6pyAGi/ojkDhe4s/7z8nOypuYsj7jKajvlRpoKvLDBjvU4vEeJvvKPjj6CEtX1GwMAxtims5liTs
WBJs+eqLov1R0sTZ27HG4M+g38f6qZIVsKsknMjp9jlBRgRawKO+8YFAHZus1oOXSiSXcCqUJJMv
RMlZPzzm8JTKVgea33CtPIWbo+T2gRQshb/RI2cNftrmTKP9asUW0TXwAZ/h4juL4JmfPJLOum20
xhLuKXMtedew+Ay400dhzSm5fJ+YQ6nXK4dJXKx6WulADehNB8Eaff4JxMC1ca7/w+NyYxa6OeCS
VcEBKSWGw1bGRlJ0Q99750cnX0It9raS35cPVB6+HMjmoqHeAnRTWnl38d82hzIojnw3VZD7d211
ecL1mw42hL683bzIWV1rYb4JdU3kVqSGU3LuawJDVudg6tDnugYmmaWb6kZkOtWQpbYjtiQd8N4l
uf2C+cm8EGf1JGZjFdV4B5NwDaZCET/9O3EHnv5det9sp2teYqzNKljNWc5/1iPlkWoGk2SCld5l
anTz8RGyocDv0gIv3jE3LU9ealIpoj39VHYd4TpV0fA707E4cFM520iQsSYV0FP/ytGOx4G2+EZL
/qLZJUqfkz9BscYzLlgWTUgETvytrkAtdndpSCyXzQI7cuTbx5ocPqvtT9wuodXO1aprTauLO5De
qpObmD26OMVaS8WuoiNzuui6GqoS0LIg9pSWfee4zXz7a035xpYRi5wZ0bDhEtVFMz9KodJQo4f3
8hzCAIwYfUdclTn1XLezjopKH0bU9irjg+bX2ozpx2jHzPu/UtjjGtUuYYr2qfFBSpdEfzAGQiA6
uZkhovDx5VhglvBjo4Tb2tS/VozlhaSYsYAskiIQzFHDxZfemV/fCZoNLkkDwj0tsmvqHlmD/s4X
HYIHYoPmj0NSNzv9twxoJzgtRBbwEXzo7kZFXOcjoIjG825mgY2Ylmt1d8ob10gXc/uipRIiUXGo
H8JOjAgQn0+WkO55gCAmyNs3u5qTHhR0GOr9HpDEqkcXlcoUVDn7yyX/M/LTkDg6ImsbM92zczqG
K+ZE/W4RaqBP2Onzu61e//HEmgmRo/aipNXuJKL1PIBPcMgi1Js6Vv79Vg4XJSUHHpC2V3hEI6UT
Q3vBaPBLUQkmwvckBprxvUxtLiLFA2vAY/RTZ4+A9Bd0Jg5nu6OhdDUbfUb5vevgNvbvvlAngvGo
HLDbQLYMj/gMtJtC/GiEpvepvEYZ8TOU2KfyrxFjCzUt+njx1FvKxvwAI4Lntkx7A8kOvULVFbjJ
L0aOVCxF7hyJ6F5aQ+3EqaParUUQbIP1eE1Y4w33lsZizdfR8rNxGGOqs8cinyiWQfqytwshkmTO
GHdOraLCO/pBKqnlIkY1nO4u+bTkrHl3BQrpvZvxmZmLdVMHYkigrY3V6WdKSI+5lKLpTH6l7rOU
YeQ25/ozqv6rLaDa/RqGYR+a+oNQ5tjoa6JuG77wbJR60Xs+cHWzZX5GfzXoezsJ/grjRheT8DYt
pMTNtuV6YtEmB7q/67ypYIsBZSm98z9/YbSHUYVkMqO1vLRs/+oEx7D74RzY0Qq1k2Wxk1gNs3yV
hrCN40js1yuXouDjdJgFFbUTWiA5WNfNcNvYTyHcC0hk5RlD4JhXEQl5c1/giPt4di1zOk25plwH
e7cBruZvtY/lZydMZ6zqApxrMS36rcXsmf73K5UFlQUIznlPbLnwc0jqDsiLjMNe+wmsqPCSbYRU
4IpHptOHup79hJthWomXCoFGQoph4TilclGn2kwygW+5d0nn8mhfHG0TnXhcOWE2xIMnNkRsqXK0
aLdC3Zqa2oFssNg71gqA0L9ClUlMQm0tYjdIaQox5OkkLGldMyYZX0tnXCPFho4ZCalRLPOrPwD/
dh5QwfN5gZyo0kUxw4UQp0kh25tTSj7b24YAD8OXA2fsTtuAoCYKwGgb4ncgZ51026OOEUkn6QB/
86+Xwd5oYY7JP5InpNJqNVgieHi08du/siFIcHqwhyi+J8ZkbW5KwHZUEpcQDraBLJ+SOSRKW3dw
wEzKDCqskLdvW0LTGco7PMvFjHxPvTSeJFFJVVAISwqlGGm6VGg2H/D1ZfqUuuCj9j9k/kZM1Z7j
+jwXjI9lMwEzdjXMqLV4PCoFCdfFTXQ++SMz4Qikj0gqkTgfUJ5MqNeVcuR25S5+JUd68EUnL92p
C3PldZEfyZOro9IdiaRPOqum5HTOMuYY5P2A9l+yjNop+JFgGcWcR/G/7acvKQtsXY0FbiOPexPO
Xd/CcDdGy4RuswB/Yr9CUoj0fRZr+9PZSqiZSYE9UEJM8WURcfMmyEW6vSQPyF88VQM3bXvd0au8
kHioBBnCT6qrxe3mQqkuVWOqAg8nglIYYm3fUAwAM0qSCEZ7d9GECjeuOmKdP8SSSactQKhZyEWP
l4RjefdrHUM/x7B2NoxHxkBf2Zt5xz5zCyD4u312XYKxJrR2VQ/4df4Fh1hwCWy/87myoYDLTuZO
1+hnUZjp+W4tRDGw29jNgYK5IYEdYIAwmzvgdZnY2MvDWezHU2JJ68oIdOEdYfjxlKo7O4ewY9GN
8AeJ1rBZJxtN+eMbt9LApGsibZrn+hGswztkuMsDp38zkJoQWFvX+La/qyTD0at7ee6jLrp7RtHG
SS5XqkisBXfsufd3w/fhD46rGL340N0/V8NCGuhA80nGESl9Acq0vACboph3eUjdXpmn+MZVPJLL
f3DI8smKYdT6Y7Gud7+0v9envXA9J71p01My3qWzxXNa2KN9cj+3c1UiKPtUgxtN4D3R39c2qeO1
f9RJHTNgZOORzHJAnymrrFcaaaTYMaRv5seuWeAp21nKEO8bKE7mNB9IJ6LT/ZGOKoiOHTe0xEkf
7gUPQJLW097CgNfq5EK3zhvxZfCjA48FjILjxJBmaa1Bt7toVpwGr6hkqoEVr868sHMDTNTpc25/
hzljMUo9yDpUYOW7FWG8zA8FOrlq/sfJB/vtodaigHtOFDxPImVUCRoJt1+q3Gj1/Mwh3Bsp2qal
Zs99+h2EQXlrFdywtKHo7BX7rO1iuvpyXUmCtkZ0x2+fQ21pg3WSCoURzYGM5tDJMEQChaRVK8L5
q0jXvBG1kz9/ebqTnNRWKD7wButi7asmBVA+i7CIq9Y/2dPg3UDJB2E/xydvDu3RLu8/ggJhjgax
N7VGHkBwXYIUb5gtG1g6mFMGl7IX/kt6AWpl2s7Yo0cz2EW8c5NFMRR5UyPAwSTG8C+BL0g2spwJ
4u/k/GY26FB9GqA4e12qMDFeIigxT/cM9lNGv0T0OYAf6MDH+y4Z25PkgoEp1JqTMqDSU3U5kk5p
a2FBCJU3kQdMy2/JWTUxR9uDVV1i6sO+gT2k7CHca6mgovNfb/G7Hsnkupa2qKd6DlQuBRLT+UZR
Fr++8DWChZyKgl0MRZd8HPi/7OmsVyglHzQ5qm7aThAYzNVR5xVDdNdu+7TEXumY89Y42I5I90BF
KFsAs4WJ7zyVeuQY5Jo231dOoYGj4NIl4OZ020Xo6KKJyAFX5c7WANVaE4cDwVba521i5ldYiZ+S
ZZV6gs2S+spsMT4kD6clRlNNZjPHnrnbYsRc3MlSMgXVd37U/8cltDc/Ge/RkOswqb9aGQO+ojU4
pTonNuWQqZb1qlnTh6VAZuM/dDUZwzVV9mL9ALUEM6ozsK+AHJw6AT23IwnI8j936BeF6Nt4dl61
CELiZ0slIiCcydNw/pJVkNQrxdmtW6fKC5erbhh2jo5MHb4QgJlLbkDStgKNIJjr1ijbxduqir/B
itozzy4Oje/BX0NjLk2Ty+VZJDEOujv+alL+YOP7XdG4GeW/HuclWQiSN/d0VBLrQ+J+AB0M/yz8
oDk1ugtux/L9Dha6Xn1H30m6GQ15eCAitHlnoJ5pVCUA1e+M/hyW9uiyZLny9aH2G8xvB8dXKKK9
vFIE8YPu++FwtG6caUyaG68Tj2pOAx9c4rHPEaO4Vlg0QG6PNYZQb+VRzc0okMCcH/B9Fk1eUa+b
qx8kEtZKRC1Zc/ZUCN+Rhi+/0ufh4j3qae8uqtFBS4KgbP1yewKdNFKqmcdgAJmT0WzORcXwExl9
3WpBhTbeM+/MJgATJfpQjDph4aRVRb3Sqk1rQxeOwM61qVncq08US+B18U0vsgQ5DGpo6V5Sno5r
oRBSUsZ+ElHOuaERUho9jejr133h42awG5yJQu/Ab+UrveHRbJLQ3kHs44uq3vItTtpOSlqilvJT
ujbK/kTVd9YxuxJFxMcRQ++Z4ajqFStW2Wb8qxmVOM4EZJAiKqd52+OMZu+sfp9JMZLWc1wC9iVg
YRSx5Hj37kpVID5SXShzGS/Jd/snfnd0w4/LZ0catouBKbTsLs/lnRVsULdmJb/DwVrVkTDHZjoP
V0Vj4CQ667DYYc0nuNd4G3sCngwT1cum78LXJ9a7DIIBf0Pbkhg3VHtaMlQRAGEbsP5pF1E/0CkZ
GzfyiZn1ARo6ZV+DYCobUJDsbjkzx2po30jw/KAvRoRDnA1J2rCNh6XETYEj0ufWbW4LPlY2Gch7
fMtjTU2ahyZ15jQqcXD2sWpz/qCr6avytNOpFlT5CJ57s25GLRsmt2CwHOJSJCIs3S0Po8zWDk+a
w1uASrtbY+ffkKUgwygeiLarnbKacQxVskzDT9AJmAtXUkfDvnWi28omN105QfhfomylaTQA92rT
PrvcD2Vz+EOcncjap7n7uQsNQSx/Nw3ME07BFG+mbJ9QbB9KzK5t4rw9+Bdo54QRCI4xrD3+uyP2
dCjCpB/I53MegdNU5y566KOTCdg0KfeN184FAmfU0Q69J2wS21Udar4Fmjurza8oROqSUuRsEgtj
EjPJNvVBiGlK/I98JjVkdkEl/faMyU9VieoHipFWsyOS4sjR7hRN0ubkZaWhnz/YlObqf1eDZVVx
lggrqye2XzORuSjEOashNDZT7C3JRVHhax0R6JP3CvO3Jc2pRJ3vOrHVED+AaPlN+RwsajV5lY4r
5JV/Li9YySy8h/udviY5oT8UV8Ov0CatRn4lvMDKnaTZl6awZjXvRRw8Aj56p9RJxv1S0PZRyVUW
ZhxKq7NJ6wZwCWTDV3BRsi3LY98oqx9/qd0p95U6dxDGXQhYS0jptk4XaSM3pws9IUox8MIeP9Pc
e/9n06x3n9ZmcNGzLEwYIa58gE5OjkV3jjc+f+GgWWDaVAIL4DDbyp8VDuMsVkLVxEAFadx3HCmx
9Hkml2QPo+zjWU24u8uVBASsqqLLZ9seex09Sd6xemLqXmzu7tFTH4YHgWhtcOruLUmzfqekyeMk
yUgrhEHezRsoQnN4LAvPm/4CFzdCk/WroiJt1uCrWCczQBKqbFW2se/ZiFLEnPxoZRUdvJLXzurc
p11KdlZy67nvnc5ttihiIql95fOa6pzAp1RQDD0HqO/RJo+14Na5Tcag+2V9kmlWblJ22wxrdJQh
IEgAZ+TwoE5UVeecKvvsgct8i8/e/7qPPnWt7f6lDbRblI613HCDfix+TndpSqE2dN/1/kbswAQu
Af0cmUe1H2VAGZaRgtWFhBwB144/WzFH+nTf5wTEIO0pCR9jTzoCAi4Kl/Nc1TVAJlzk9Xou/PqG
JrVG7YbOhIrNydz2gVRA5vS00rkb9BWp6C0tUlg04+8s3+GezpwxjRuorWbCH6HLLHIJsaU4wNwO
8r66XSZe5wPvbtRJBBrlUKlz7kcgUBZaaFBMT+WE9Pyo3TJ5oTYgrjUkPRKmFV/oOFLzP6QAEfNU
JLHjvL++2kpb7rOnLlgxwS/2TjZzPucoXvgya1G4gvnbbpLFES431afsrfpQNromKlqnggYDyRgI
yN/v/RpF/dFIhUsyVYnU95mfuUVSHAYXn2P+iLcWtRrBQW+HB67L3ylNzz8Ti7qYRCNcxGfY47UU
5eIS42uyVMUKRfomzaksH9cGBfUVOY11OxLQkTUHO4atOkrD8le4BoZeKC94EhPMpG9UEbAySpOB
98Hf3imqr4FON5Mhc3wkPShZT53IfMBndQ+NoHjqMq5iAzTJGSYYNVnUucMmngX3UPWm66lljgOt
2KbGx3elvg39PnEKH4Fkj6iq8r10pD8GJWUaOmQvj5Xcrk9afymz9YVIWwHzWyzSdJzUdLCTcrXd
T9vT8/07pgTD9J6+Hw0P9MsmqE9h2XA8K3vJEwx18kAhAfj1ozp03g5f5mOz90499TZ9469mp1x6
I2Derme8bo8j6MUhZoVERFWooDxi5bO5lpW8B2b6nJGdGtm96PIvVZnXN2kbCE/N/yUYcja1ry6x
GcJ4O55hp8UKXRrAgurrjrBDE24NC3TeInVMX78rkC4FlK9a4NTUU2IdqM81IY6bEeXmMRbvMfYO
xI8O6KU6RxQXmkaMASWyEOqPiimFuN/YUC6fBQ75GBVLdjcpFgIrDFsZnO6NVrLy1Nb1LX6W0LWt
cU5kSOGOyNmN1VNpuob9RetWm0OgBcUZCAiIFLb+cShpoNbE+BrvKhynFJaWZ5jeQSOSmw4BD9iB
O4qOirKoiKeFVyrfxDa7GMHQ6mN6LA4nqRm/0JuXgLQ/rDhV7vCpYWQnZCOQz40Emb2YmhYSbNJR
fRb1R3ehb1jzoRuLTzq6U3RpZt2ZY9wPVM8MEBTegmX4I+bTPDQu4rm5pT0epy5WeBgs8JWOG51Y
fWqQzFNx+0eROz7xmcP+/nzJTzp+g1PlCHaRCBV82FElpSGueEswkOL+bfk8vv3P7AfLVk4gpR5z
p30SiiQbgeox4oZh0wyncUoTx3SWSbxnIRMbfUis+fakaiBppTHTSpDHpgCZJBU3XEay9aKUgpKt
vXgRE50Xkh3/sC0MwyqJkcsCdNmu+frxI938eCBTG1CW+YqVCtq/FvvwzIS8/snI03fdh+zawOF6
ha7R1rMJtCYEMZA3aqTEhd13G0tlpk9yNrQFIYWruxZR0K9Dw2rVVeQRsjvhCzuOFGt8cRRbnkAZ
Bf5bZFP6H98/2sAldTu6DtIExd3mrsrgNtdfMgtgQ2NCv0Uoxn1JYOI4Mi1ZkrvaHWdUL+0fdvOu
KaVpvvi2WI14h84cU9A9foxJ/U35DWqIGkVxzzGnty3HpX1iLt1DLg8/M+vN1sSI1Vwq6FfIVpE9
tBoEXHy+XCC7HKr1HUnyGqXcSoJ6JTXBpZENmbDk5IpBLYjwXm1C2JtPgJkHHTFHOoRVmsSFlFSj
m9VbKqyQE01v8ipewsy9ueo/HeaIIwOx9OFs2/O1+3fv17plvhl35Gu1WrbG3BDN4R/ZDzLfweo0
FPjKEpenX3I8oAAdjyLoonWk+Pro9axAReKKBGvbFIU4HO6mleIDy61spyHWydNCLZriq6YbOINh
Cj/HPMjke/T5h6OstEO2gGmv/hfkNNPsxrmu5BBesFvHFLh+cYOmG2YfvMwarHcbZFVWdmwoJU6E
67fgDk9pHKs2ExLKpn01v/xkBjxFw4M/k9q81zEOG6fm9+XvXyeQ4EyqGG/7FxNVS4uHlSnRDzaT
jIer+oIvrw3Q2vNPC6NrB8jBWnwHpZRqXdfw2xmh3iaSkIB5yyAV/VO4ZcHjxlLcT8u6W3cNr87M
HjcWQUZU6koKJxq1Ekl+mWnpsjrO0Y9HrwTjfBIwR4X7r+xDSA3Le8dLEPejVuFhXGhlqZJCK9Kh
FYVizh6x1syAMLI9DtdexpKq4zPxlUgzSl8q6EsOvjevmdFOR8EDpcDPjx0X8k42ejXfw/1SENex
atJCFtt+o7xQWKZAKh0qRbSFgRnMcnrs7EI1V3q3MXIB4T9l9kVxaaQemYxEmJV2Xo8DeEmfTTSC
PovT3FN6cpivpRq/M2IOKYGitYYbj7JkVamllYJ+m+Z+dAlmR90JNLdeLAe4BlLMOCnxXT+Iro/A
DDikq8JGaGuBZjZCs0cwb8JnBjP7mw4SUn/jKvKPmw08X44L9oMypCATm5eYtLIP2iBXSUsUu9d0
k72vsmm7hgTDt0wYQvKpvPVJiO1XFBNRu0EXoArv04Yr1QelUJn0azAQiEwE4w7Rh0h/WrWJjXUt
rNEhOwOLofa1gqT+ADe6XEMV7E7C3/hJnBxNKhf29zJhcx54W3W+2wp5U9lwbQcW3P5ixg1Nn/Ii
4D9CqI3tOWfVXK2/ALhZ07IIHVC+VyOXLstLPRp31W4Byj7he2RN+pPYwHNvsd6Gl4Al3KHtONus
5cFnUAgEj4I6SCUFH8cEpe3wDA3QNKhonhkOVmaOyURm8bb68IkVbEGgAQwLUh6ttW+OhHjZ3n4T
V2OGol+hVp/cSlMIOXestOeoQy70d7jFn0yMoPhxg1awjR3iCPHZjDSK+h9uTURXhVsMmRPvfNsQ
C6jzCEJKYMcGzKikw8Jn0N+7vZEZEmTijLb7/qXnIP3HIFNRP+TcTarIbAo7GcWPo67aiyle+YSi
7JbgqPiGgUrSX6wt6L/ufVjajU/K9FuaXwaJeGTCqBcWC2EIrpIIL+YNivK253fElVDpr94yrCy9
OabL0Ic8+0XSfLLvbqL2az26EZkn75bXrHuTmKHiI2PH9pbxDismhVftXrS/7tpNT4bN3PHnweAW
5ulyBrvrdVKLrVi12cPFcqQKoEfDxx/8jdILFSYzEg6+1nc1qeZ61gWJ2pIAn6c3mcuuu+q+juqk
5XSZaLRJNh9RZPRA+g2eRkRsbgAZ6cAtgo7Qmu6uqvy77H+51hosQ3uvinFUkWIEJ/ndb8mN6Gj7
ce7DKSrNJnktpzagiaDe9XRiVn8/3iECTqetM+p+KGI47wfdhBsDXsK3LJs0BuHlnFhEqKvW+37f
p/pRpsHKlMfsduTnA9EHpRBXFEI9137GiALmnZQwTe5+GulbD8GHk3Lt4YYw1kEX2ert8TXvb2Xo
+tkkDERsz8YP+9wPdZjmxUoIfg7cznJIEpOu5AbFvp8N/Vv2pt0LWtv/YSdnzTfKPRsaMKTql5UI
+TbraVcFYTwyiNYkH1fB9H0Rm2H+57McGU5BedTS72oqyYzLirCwX+0YQ8xUwXgMOPSL7bo1O0an
u0ptfKkSGB9IwFo1riL4dagXFDGltOzjfOhGgY+a09thbxsfM7goSnH3vuLpDUIw9uP8XvqFHHd0
NRpx9itkCzAooJ4MMT+wqfesfp2D2kXTSVanpYVzu6a48n3lDO69vbRZfDT+b99psZQd3eP69BgN
nhGMGGlB0LtaA/YCYpjZSM/ayHla2qD1cYJ1TMq7WCoLW7rc8x6bLCfcYlXoyDx8ql95YIEMijC9
JCd+8PQEy5k8SvoNbfpCnuqYeIm0R35yU5IhCEu79TF2KkqmqsStNGxWK0goTIoKMDwmhl0CfNZQ
mnmmoKTmEgMqwhP8h5SEsR1JBbRG01sjEvTJhuCT95zLgR8iU/0V++7KB7Q0uTt8ZCks3OHoAyGg
5Rp7YyqNB/SaqOJPB/HAXQltxcAw46h9Hok7xCB6jxa/O6d0kIv8rZ4yVEMDgh0//yiXNTkZ6BjY
OZkQp6c5cGu3Ktm0oqtcDCh1mxV2ahU0R/bHf3rRPKLoDP1U6FY+WapLfd46LNQM/SbFUaLcP/Ty
TO3oMEHSkg5bYJWBaOZZuUWMQM0LuVzXu7TxrG2x3i5zhfxLLfr2PX3G7pUcPFbIBCI7W4XFdS8h
TEdTbh8/UZSxYSuGxdjMadygx7Ie29NVlfq6AUSeJvHD32P0zCXcDexzpN4FJFPhbEXJX50WWQj5
HN3nq+ulSb7EwMcwXVefFeaCL15YUqTBNQo015Y6QQmXwhe18fqTQFSr/KRco3foEAvA164v/UDT
UkGQZFEf1PPP/RZqpG5PbLGcFQaDbu5PBUzj412wu0PyNHR6KsmlX2NkggbWc6t3xxamcvW9LBdT
LJVOw8id9saWBQGOTwNJfW8xvinVJ41n+iOZuxwbt6nGvOjwwu+QBXRYh2G8IIdZ3mHFCMKX7OCU
0eTDoIm6BJsxP7dy6pGmfyWVIS+FGWQ7MATY/TIkB2Ok0+I82Y8we+ZxjJs/0VS9dQv3FRci5WE0
B/dSWCwGlmxi9qhugdgfkGz3Nn8tEubWrVbfQSbrfz1HNPR9AMlbv2REbMWl7YBi8QIeyuRR9k7J
9UlYnouWz0BtdE9+FQJfFPCvkOnTjXlGGj/Vy2dQg+9Rc4sjChUPMAYJ4nsnNaIHY9WqF66tQ5aa
mSzuElQtL344RNVAqe5/h6AMil5GAY50M+cZpf8okGTRuucMBip2QH3KRW8KHiRP4YbvbwwOU2Vp
bIkLHCyZwLACE2K33l1cl9WmAO57Eqk2Xc7rYSox8Zj/SqzQWBwpDSHCpx2tv5GDN9RViInDSIz7
RLkZmuX23koJQ9DhXCK6WGEFqWheKZka7ONknsW+FTEQnAakMSKDi0MpfHCqfMuBkYGP+5lEnsUc
MxbZ/oZo/Ixs8z0Jl0ycCamzI58Nwa7cj/cQtfjg90kRXe23FmgRcypWMfj8VUlMOH4wjAeW97+y
vFAlCggxiWnLeoY6dIG15StFfBhaQotDiOXfQO/ax7E/zKGSvBtuURVt+UaZXwldFFNLyRC8SoKu
Nv62YFWBsOVeV+t2PoycH9QUEotyW+LL8SqYLCC/8QfEgOW8iplyv4GVwziHcXeusUCGTV448IFw
k/ouJWX/xt4ZW2HQNz5gEEMPFy+8gS2bEJyRQYVBJkcCFJPF7YipxTAwEZpLOa8QXaB0dDgKxXLB
RVMR7KzQHNFEeelg/fgBzPWVfwCMiPtIVXdTubfwNgAJGh2WU5oq1Jl5IhmiAtEDlLnsFBG0hwQ+
+ewoB0Dlh6q2VfO0An/OVg1C0DZ9+tOzsI1iP2O6MvZXeffQYD4Qny3jHImR8/HUCv0NaduU1V+8
UVr4Bnb+ZRQHycspB8qzQf2ArK6y+R6hLH6I30HwlQgIokiFVN3YyRQj9M8149aJc9jYJ+g4LRym
UavLz+a1Bi0Luj1QgOYb4IoIfK0DOuKwI4VAcblbmVPrGfZU14E52Lg9yTsnK+DT6sAFLIgmJlNK
XtEEPld0aP7mwTVoK8/na5LiCdSY/3DYYXF02GTjR0STx6PcF0gu49l04+IEMcC7qxbtz4YPpcD5
MeXuxeqccN15XXAcKpz9+S889rY9FNC9oJOXOEYMCzUoh/av5e/GEb0S1jMQUoAHDOrxrTEcO9/a
Ojmncb8UsvRzY6pHc2oPbhvdGztFnTQx7VpWHcouDtkXpVPDEqK9V/OmlZGI/pJr0lXJ9D1UJSud
h52VpOvp3YLL0KkVkJ9DaxEGSnasLQBYf6rNh4eE0yBex7gM8dnr2NNgWJLmKZ2XKMQ+ZSWdxfuG
YDgYsMKnK0ViRHd9c9TZ9VoKXdfYQoyGPVuxYwggwA2maEoNlqOj0a4i3PiGsVS/R15zUEEfUuMl
qRZPZWc6x/3Ub2AoHg6oVErr9E4YxFr1hLGJnurVm6xROoUzHAa9LyByV9gbSags2vjYPFJ1w9vo
BLtFpu4MP9CKgFLYOWiexgbMZMV5PylgYu/Z5Rr0S5c8YWct+R2lnz6dLw9CBSq0yTO89aauqP2T
5L7/3pwBRSJdD5DstvwBe48mY1NKq+6mcggqk0XC3WFrB7jRc2UkhBwl+X/BIEOo5VmzF2S+fvr2
6UUQ9UrQyS2V0XKmmuLvyuz3GXOBM53WR+ItlIwOIrypjjfVQ9693eKY+vQkmOkacZrf9IAsrORZ
f2RWf8H8Uhwzdg2o2vEUmJzv27S1wU4bwNTFD71XcYjg5/Wd26C+hRVe1/vmKFHQREzqHokMiL0K
MfJDb9CFmkFl74MMcGshma4hGFS4PQWLladdAO/qUePlbNm6YXi5DthZtqsq85/caaojBKe5Jjt7
rNfUZceezRFx47WU/mXBpUVc+YTocmn5nVz/BZ+HVtg8fqqScXbuGpNoOV9pFQ/cyO2LolL+c8b9
8z2qD1u9uYuHze7VQ53yJdMY3wulZnaso7OQX8xAmQleJT+h2267tgopItV4tQAWDy+pNY7aaGii
uhS01RhE81PWTF2irW44nsWELtmtntSZpgUNwRZKX2tvPiaUUH4jFCNdJSIYGOQYEa3xJfapWVYq
HofTzBNhA96QFYkiXgnMsR84TBUVI8VTH3wSH9QYBe3/LUW+cWXtUGbm4FIcfx618RvgRe/8N6qk
59HVqm483ogC5g8Cp1r2RsnS3Z3NwLjPPylQ37rlSk6DcStVo5tXVCTToMFY4uCr3uJCQorowI9a
moS73Gm01EKq4EPW6xnd2GfsGJHKun3W1c2J3OQDFyk9pC4FpT/l/fbKAb/nZWcmOLgSRofpfnfL
/UzS4q7ioOkUUt6T2Grp694eb4Pjo2wyoiyw2/vkjD2CWD39e36X4f1UbR3EjH6zheiWsRclsrhw
I0YBergMdj4b4t+hVLDHHN5NMxl/leHPtoVY3JheJQJNEJutoPOtigx53VcRwdMwuPLgPsVZpVkE
UyXyJrJlxWwp9J2Axe6vrHjuRpWRjwmIHsbG08xsFdrAO1rO7UrxusFa2sYcQshHFBIcg5pWMwU4
uVLeI48gFv9HRggma2w7sbzpr5jw0xbfU3DQy69KhKCQV/ZHCe9legnf2HMovmMk+mdsvXOyOB5l
74rFWDXfVorsTCpqIoXQDTobBRISCSXWsCfIJYnziXs7hBnn6xx1J3Bqw9mymoHmsYu/jseene4x
7qXbzoAAIX+YIhDJ1H8Pd5q9ZegjA/7S8b7hxbsXPhaT9oMuilnkp+a93PiFF00213h0N5jhwbg/
UkvESAkbhIcXRLAxzcGuehNVcBJS4uWUeTPgVEBuJlVook9Yp6u9oHf7ireJjNujZctn0r8qwUTG
ov5aIbVFZB+BWblxaDrncADEyPZ2nwpGLOT5gVwJ8xtWNitJ2GDz2YL3OAqY60ceN0uAH+qqEyJ8
2i4nW4LLalxmr+z6Zf9zXQB8WsnlSMp7gpXzD7yzsRKebGtSgt8NYcuHF5O0vBZTfGMwek+tXlHq
ZSqPQYix+ErUYuMN7cNVg5cbVUft6n/J7/9b2KCFURZjgEZqusI9ooDwqDU8LfS0vuFaIEB3YAev
oe758W70SxCXTB+MjbrmMq/NXo7Ma9fTvKGjYe1UB/P/PYJvYKbAkfsOejkFuTSpTLipJVcj4Ad1
l5KH2bIvGAEBIxbUKzPeDba5hw+czwKlxOYciLBIgOIkEewD9qITwVwsNGT/1Nd0btZBqRiSZTew
iO6SYb0kpzkRPXAxKY9ZU9KVxbhirYH2wCK2IEQ4Ch2hxUqA6ntGjcuZHZEusbfjXW9n3+t7fbFo
bzflVsk2cEhjYdzO1UazlmYkk5cHp5i66QRb1ef1Nb4lh2MvHZi54jQOCilHocBZprLXK/lucKg4
KFJdznZD17yU2azgM7A8/VMU2YzT3c89CzE9HK6y6Gsct+6G/LnPwOnFyhtXlR/O93Fin8PrEMJX
2y0DdSbyydMjPw2chB8pHo9RFyLH+0hxzv9KATYoEGhovCqXXbwzoqRjuqYByJ/oeaYK+SotaFld
uJN3xpmO1Y8cu0AxmCXzBHH9JGUEOavXxgcGDfHnO6e3fBULUekAJJWTGfhS2vgUHi8ysGaJ4frD
Oan6GrPfBk7qGSELrBjF9wT1GIvMXjpus49SoDZPA5G5iyS6lPRr++f4Sm0VzxUG0wJAMYzYSris
b3szjEWfvX8Y8NGn3pZgfiXbqZAt7TLFUsTsdvvI5d610v2RPeBPnxYcwcbpcXpoFw2CkPnQrO2o
9GaDwWkbtVYLRvmlywlMUytCOUdJ1Wjfovpz/xUxCR51Bpc+RXDCT5DczeiBuUQJAtgMazW3OBlj
ksNx7w23IJzi6DvLuAzYmLoREzN3/v/DUpqFLE6Fxn8+nBdtlcWboDDJFKHnp46LaGpO92vZ2yd2
VrQylLDGYeHzsqkphpqHrXqry8UQDg0Y7wLtj1+j28tIP0mIvcu++5pX2Z25uAdgLlCutj+WSFud
3HABquzVCgK41URvX1E/q0DRll0ut5LUEfPF8p8S4Lboz9GFEBy+n9qxkbbFX3FZUulS3LocT1pK
j9NNpN9W9amAJQqsGO5bEPB570YosTesdEJdYKJ1nt5hpvu3MR1W5FUX9qhjlGS1n3sDzzc5FRhy
ht3wvjgmljv3ZI/VUO0MTMSQCT8h+teHeg/bt5MaoDhmYAtipGRXog74vTzntQK2CLyV7quKQeAI
5v4CuTYexRXF6YFBUjXNmVe6emD37xZmklfKMdqX6+w4hcdiKy17KZrdbAiP0kzGZYyV1b96bg4S
fXalq5eNDENYHx69VmlKvi7gSZj3Kw3Z/rSP14htQbpfikKVkOxgNQ6YUTXC4kS0uZMn03eG8TO+
yuqXYqqVNJJCkxf+4R40D2PxtflPXGjRjjkhZUV0sWGWbYmK+ok8ePzs2UBYKhL/7YEuVvvIQCwZ
E8fAHpOSw/orB3O2wCcbh+5MRlYHe/mVi+Je5OU2/TajUw0pDWlpm69KI9TUpSTusCl54IEfoers
+jBhGDGsNsOnzgFcOWY5epZ4QP4UNqo8IGUeemqXkrpOXrSjJL5B71Pb4Hv+8bUxWBTnyss7MwbE
8p8fPkeoaSkK6agv7RhFQF+ORIhfh2ppYmymXRKaFHXkLNqYZ440/odZdGQqYKY+8IX8QzVH5Bm4
wRAlEVWpVSo2w3PqTF3QZRs4IH3ENH+ZJ91/L0VvccVZZC4h4pYMc1Ol8Fh6S+gMq+rZb8Gdheqg
hSwOwkmUOQm7t+ksOwhZogeEZWuz3hLks10Y30p9ksygdQM1BBiesociFfA5RDyX/YckHTzulz7U
FmRpJy+tj5sbSh5/LcpUGkgqywU7ix5Kmdh8wrDjGrqkIHsJiKdK2I2hZuFwvcBak1bR/73KwhaZ
qCRNXl9kScSO7NLvIKzAw88ja9X6o5gFTX/sxa5WVr6MwAM3Otg2hWCEDDWzYwLuwfs+4bQ9Jqiq
f2hNAHCI9JBCHxq4bWjlxA5/sRwt2B2v5AkwsK8IAePITesMRg6wVAV9rgBdhMDSxTh99MS8WZ6W
s7CVem2JTn7b7HZRlnw1MbqbtaqspUB/MvqNXcpaRvRosW6No4+UGVr6KY4Y6xLJdpCqcJKgA/p6
1wGcKkvZzok+WCYXlFN92T0u4tSiQ1ne3osjcONruqLolCdSaqIJda0mZHM3yA7d87HnJjUHTUc1
xaME16o5QCqd8+PhSBJZhvswRcrl+O9cLi/raR0DFqe4sEUkfgcDt2N/f39UJlxtJO7sV7+2q6g9
iA0uI9am3XStixtuFKkw1NNZcfGdO+L34VnCY6i1Xv6NwgKl76j4mVk7kpFTupdvRcAtSebBOATr
+fdaabkrydZ96gaFITR37VTsv9xN3EtiBHQa++Z9E3U4D5XZmNAPUPPWfcQBTyvosipVgTQSHqON
eQ0PwEVgFbtQOIDUxlMsi+1KYnfRJx94G10rymfPsD0ecrdxf9csFyjHR5F7wEahahHSe8MnQokG
wnP44ae3nQCPvG8WsBvyOtli15Cn/H+ctGYmuDQRQRgdCH+jirSsJuom7IUjQ48oqlpdE/XDUsLa
Y7ZfOeL3LWBnaWld4E+MJdzbYoY7o47xHxmWa6Mh2YNycSxIRXvINJRpRiHVQd0RnKfQDrYet/BU
DoYbXIkMDHY9YEbPbgpsbmNIBi8rLwhBf89GEP5ZSpC9NeDJqvFinnvTx28cPMBijgCBRcjfpHZ6
k99QbclSOwfSooKjvfjCgk7RmlPTnCvDUe9k1C42f8in+1+MqS9Fqr5a6LtG/0DjCs521TqdW1VT
N7ePmGdFrLZppwZluTH3O5x3AHlXFlYKdAH0OCNN0MbVQniB89snadrbqUm3NOxFg93VW3eFh2Rr
FWm1EGNaE4XD3pgPdkQydlx0qVzecxl9MyDsCd6kwdWVtuBvjspygHUHKppA5G4q5DNgLJbzGwcM
JvYJYmXvCuUGMcPtAEVY/PvZuFc3jyoiqPl6S8+FMeUslumY/9cI8Y7gxwjxOmG2MVZbrjYG+H/U
nDGwuWV3/fgA2WsxVuOta8AZTbGI8DV7DZ76U4n630NXC4EMlOX7ZjzswyIp6jVv44nVauMDaTBf
Sb5Cwn+E4F6FDX2bY/nKmubvd3MAlX1T419u+4Yqpfd6erAQzMg9lSJG8Q9SMuQXjJo3Hh+U+YxN
5yYCu7kGQaxYcnw8or+PnRzA14aezeCFHwZiDO+4DfQSg8l1u+lxDxBb1COvj6zYjkchqxL5BSY8
SYlvfXb7omQlhn8AehTXwcaQfYjYF4jg38MxykJhXaToWlxATMzcqXZZFu3lPCi3JdmcSrgSSCKn
zIb5jVxN0Ak5bdPvjMgsYGID+9ORvy/JEQJT+Z2J92N3Ei2ZU9i8JCRIqWViumUPXs3v5ghJxMOE
HPwzKmGDid9/X8tupailQTA4btZJELOc6onfeRuHfvJWuxVLqp93TajxXUQMcWWtsDR3BknGJ5AY
8owTv83gH3vmCmzkQP6ZyYvg3wRt6HWoyJUM/ZQk2TRrJl+c9j7yCF1MetJS51/t7EO19E8/vENA
b8cNZnTfdxOlkFT3HJ31BD1vKTf5eycNtEuElWyuIEEhR831YeaiozDo1s9RMBRe4Az/dVeMIofw
e07nMFZAWno/tqn8/wiTy1pDi6rE7056o/3opvtlstF/segNlIWFLqof4WYeXwDvofJJLhOTiV5J
a9sijtW4DXyyhMueZBeQekM+6Wor/faPz+M1jEK7st8cKzIj1+1dJM9853xV4XIDv3xHsV4MtQ4v
pT6wU79IAkNETKqX2ZcVvPjLpxfhfza+LMVPrd3A+b0mL4JYS1G2fzMTDShDdHU8suXila7vZHzq
muFFBtg6NN2Y5pjcMd/p7WVnty60issxTo8oamgordDCc7NnRLoMNZGXLAjijz1eJ83tY6KM3iT7
omXoJQSZrGer9lnQI1+s0FPFbrko+vc1if7sJPuxF9eMLTrdsbbZxR4lU1enXEw44qOmWGSf4J0d
QXpHZHRgoQ/Mm/rxzbr6sMzmFG3UZZ0pIxhJTHjLIhmJWoqmHYDxmjHairc3zhcy2ZBs7GsP8n/A
wX3DHBSFiV0vAuCLorRICoH+Poig7rtDLOTdPH3zEafdfiKS2F1w1VoSwmI4F7tFcPdNZs1OcECL
5S0a1Tuj6vEcCbiqW7ffPKT+3M4zTbkm22yYtSxS1tpQ4+NYq6J00SAYMDa0qAaHjs3PPxy65o3o
PU7WBmGv0YFjl3boB8tvVsARXsiRvI2JrHa2AJWmoKlhccGbCJ91NqOypfiOmWcRrjjC1SHUbVi7
qsuy8XZ0gCqFobMDsfwyCMDoSBbY/KJ5ykGZOcmu1RYjJnbUTaiKSzDUhQJTAEOauk/fw5i8MBt2
KAllCl+uj+2X42NbbGlNyAXt2/P0B5Kvg61Uj2ZIdk2pFnwE4u01LnLfMRTVH99RfJCZwoqGUEx8
YqknSmgpV4SB3rKqoLH3+SZQ6Xcjf++PQbCVaTq+8v0Qg1Fer/NhOnA7LPONP6Bm9y+OCsjMhE+v
YutVOW5u2Khd8dUF/a9yH9h+IRsqKNdBPKIYpsqn1Ptl5YDj6XBvEFUs8WaFwu4OtlyxVpNZo379
wJXIwpb165IWJoZeukJhhTD04WWrJ4yGddpkKaK7tuCJaIpXT3EduEDm0Bf0WjmBhiyzHVdSe2+Q
IAtTZpvTE00pikLtp9va8rX/IgQzDMWEuts6pIRgmMb1yLfdrQwQKxbn+rMxFKqmrhGND8Nj3NyP
TNhBVPOwEoCPfQrGVezCGJac00liEf5bZ4w6pfL+HTH+nFGtOXupD5ZWDgqYHnV8M3cxm9w84Ong
Lh4IvLOrY7tfYUjNZAXHbnSoY5X7ig9zABtNSyWXfzBQJVO5ymbGlPgOZhjYMKGb0fb+QRt07gNW
Nf7PFg4cn3hdpmsOW6XFC3gBeFxJa1RG6b6UgBXpdRmXrEMvmDneNFaXRLf1bIJTmqhKEREvZ00f
y4PEQME3m6WRM5TaBrtFtN6ffEg2XIviFgot4tWslnas7AYJBkfLp6O5RVjaklRg+vbr3dLEhOyw
GLZA81hCoxjbdDRHcbB5WH5ecY3mq38nprhoM3+UwInBS//Pkc6NRPWgFMb4BGtA7czcKrzLocVQ
wzbfHxZB4qSb/Qxoj5ikVCOQ4bSwBIucJP96hqVRQxREuXzmNqGrU8YEwFE75dxhQ0Vg2liVqvCN
RFgXXNg/VMZxPyvfFaMAcpHCRTx7mxb064Wqm4d8sjvU0TWHGLqlUPdWiDkkoTZTmMyl9nOW1dRN
9IOFzsJj1ncvb37mcptiv6HQnjrRzVUqhEGLkJcYvW5lwDYy7gkj4xBdUhc0axuOe3Sm1elOHoDS
+uAAGmKqs9YaceIltKue1j9aPTC90NKpPwn2LqicfZFGVmZKx5XHodNdEjN1q4l75dPD4rX8nCmk
GNCVnmX1/YWRVyUEJUKNWXzilxComNOQslVsOMGV8wXHX2qOWBi2FvPAbqHLn29p/dl98uyQVAVS
OqHdQCh1TIjTqfISUoCzeHHJFIdY3SY6zl2mcV/BUJjC4YBYrFF+5Bj5sNJVLeCpJDAenyFKo8J9
Tuz/qDctw1Hbec3ofqoyGMn4ZMKU8qEuFePA33oNrFthY9rU/hkImkTeSL8EdDKfLJHzX/6Om8ad
A/p35QzlX6wzM5EAO0VI0invlfjBDnF+Tti01+0HpbU1A7xPOc1LflG21JCs5nyDQVmK2qAhRV2A
qFNxnkYgBmLKHchdo6136RdUt6Kd+s2CMZcN9tZogEr08HjxszrQQp0+Qm04awpd9ErD9LOBo1LO
iSezjdTKtDouKRBYnjPwKmOZJflLHxbjMOQ8fSsah+LoAg31+wNBkEj/pb+NZLegUWj9OOqA4mx+
hmQ9cnn904fAj0y8rnk8GijuaZsy7yTGECnfLH8ZC3BAjLQAOwZUq1rCSarqlBt1vezC/qtZ8n8w
IGmHQ01uwHVyKwt+1MphtAe1TJU+QgRs19Q3PRbT9brA8Z06v2GXEXbKH1NkA1bsANDmlZ3hXKlW
OOf0Ol8Q5LNExv7QyZnDY257QXXzBfn191WC6By3fnNWBPYPPngaAVkOdWrJYOXE8f50bpp3Ydhg
0k9cNgCBZQAwpjEqNtWddEsWOfPvgXYOxCb3C7lmfl6zLIrZrdPYkScQB5lwGvdFLPGH0/JJrTuF
mQE6HNgwSStB9DqDOqp5+fscDkVPf8FOcetoI52g5ubD6Tou0uOTBdKdcKQOXqcLljkO6mJESCQr
nXETIiNmsbgG5R+QCjuSxXJSEq8AI9lfGA30dbLYtvqB0sHW0Q9Eba6qkkTD6FgeO4wzH1UHZ7AE
qjCbAAm0xsg0Epbq0/RzA0lvYDvMR1LTaPqLo/z4PS3dTC8WDX5djv/a3tzDEK0UE4YPrlaH/tNp
3/PVbIXcYsM4MaNc1Nyb9UN4IJhlCurE6PMYy9twOokp66jweeVX99lG5BxvvO+zCKCbDnK1PG2X
151u1XB92P3BklNhbhdtar/WYR6471fa50LDeifjuhWeJLiHdClQ+0hEJum7Uh3gbRp6wqCHpjUe
Y2GGxjwtFWfVMXJSRTimNUo+eFwRqC9I/LR9L0Hw85L8OkzKCaUf7BUnN7YHy7UF8VLF2fGL95vi
6a/OVEJoDFbh9BbVeG2wrhltHsEVNbaCIE7coFJNd9bOcbPdsul9t4v6FN9lXr/ZUfXxhR+q3tcU
dLUdiH/3SXpwuEbk26/EKrb4iIILXDqWY9CvbHBbEI87qCMB49fYXErPPpOq1emTeoss19f3Bgmf
g5tEAGS54r0lAtRSKyzOQKSf6AfF9WRTc8FRov0LIffl/jmhUTDdQbydT0kLejm7vaA6iJx9UHLd
1V+PGDbA/UbSyFOO0CasrMqq9pqzaArk/qLLj3fFSCqzZ4rMM2mhSwtyM4jYwWcov8SVb57gbNJ8
ZETyxz828HbLEBGRuAwYYTHwkji55c81Y93yPCmyHht4uwTKYg4gOTKCkNe3QWnvRXeTiYpUC7fZ
V+lRhdahMuDwM1NVq+0kgVADtPumVy9odtez5djinNRrZ1aAZAA2L6AAwejgXvJJCTomPcqNRAqP
EUIjOgbNyJvJ2UM7CC5GLRIgKr3VjCuycf6Vavmh9Sdyhdeizv5nEMQQeZj3LQ99lHGBWUkxVuej
phS1g75TLb3VtrfcvjOFIbtAAfy1BdjSOVS1qhIv2gr5vaCRZKisWtX/cAsRTg16MKeG8AOL0K7+
pEZi2cjRedyofucPduLHCwlGhx8HuF9VpXt16yr04yMDQjxx4Hf2ZBV+3enQzKxLREwgkl0ppjSH
bJd1GlxcCY0E6tM1a1+eVjigMlBqCOShO+AYSTawqn0Cd8PQeYxBO/GuA4TtLM0WUo9svyNMvMUj
3qenrrc7esKcnhx7MWt4N206CA9PvuqBocEEmhsyGE4YM4jGRc5gMgbEoKuxGMAlTxO5HdLRgmbo
v9XTPJP5cPzWYOLQSwgLKFQmb2z82IL4FXqBb3G8zJBLBUVxjafUVMhIsyBRM21fcLFyjW2yvZVx
8DvfGl5tin7EJvFZgxlODjaoF8AOjOAUd0SUx5NmaZxIPCQTyVw6e2JznaJzqTeUkSfHz5UCo4ts
oDoEIu87fL59XRM06sj9WaEB8sAAlMRxMBrHD4/5Um6Aee5SlxYmBKGVWmRJVpfERD2rh1KDJWrd
U3RYpBSFqqglQWsbEGbFRToycYJNGxrnElqkkbOxNMV3glWKYFSONLanAfs/hgvslKYU9vhSz8RU
1xpbPFXqv31ftONpglyQKrZOJaTwMMi3GgETayorCApK0f0Hvu5Quo5TnTVulxuJFdTPjdatSb81
hoNeOvXfPUWpC8yo/NRwwjrhIwmhh/XzDdnD19jkqISIWkFCGQBl9L/fT0P3fpTKSf8FM5iMh7DO
NOVdbcG4NEfZuYuwbCdf9dfWimqOFRd8HZzr6wJonxn7mfU1M+EwHIlVVMC8BDvAt9yHjqTE5WZB
0Bhew0ZxlpE6DItlG2TXPxjUSYfVbqxriap6NWQE2FSjaLys+YjrabrcuDvIeAULMzAV+OlYZ+2E
oZv1PR6nY5I3q3SxM529plPTLEoa7T5zQrY+gneQfYlmhzcXpSn8ns778Cg7PFDl5QdBE9ZeO6M+
rnnZu0Q/H7nfkO0hanm+JHuzkfkHRjcKlL9hJxx5w+5nhhnzxLwuViKraY2vndUX6rWxiZgzD/Il
Zn7wE3w8K6GxphZeMhK/2y3uJGRd/kTXtzxiy8arN6Hnw0VpLRyIJ6vPJoqm4jcuZEBmJUTJRbPk
+V6zK07+8pzP21ncuFEZ72gE7vWcRKC1l0FrnNC1806drTwiAS5NcCCU9QlBDrveptpkJR4PioG9
/ZB8tNGHX/6q9s9j6VyeeOFaVZYKI/Y4P9v+NDu5KtHG1m101aoF1bs6TiJTdceaOLrv0mihihPv
4oLNmrxyyqID6saYCsHif3WWOSRqLIeQW2Skf1rVREqTTlH6EZ+C2wm5d3yvvz5NGpGLpOS3Kszp
UDBKSv2DJHhAVWgWjSBwOfiVARAkPL31Bt9RdrmROUK+5lsrByMlCyX5lOukW7G0Uf5F6BsBe+7Y
nlMYYlx8oXzOqI2vKwhtP4JBrekLsmau7IkTj/vHj7SJQHBYcAqQpJdnxBBjWQeEslFBC7QjHQAq
FJfD/cq69UdxrYRIkUTHVBmN+cEyCLo2FfCiNrabapllahBe6+qlHPtPXJRVFkIjX0ju9s1YygMP
qbvjxC4ID0oLrzptgDCvjI15WVUTCOAb4w9yozmrYsZinZGJPItCmvBeOfTgf2B3K2+VA9MwOXY/
Z567rf9A7e0QLhhiNBmwCsJ2SXtvyvzyues5YG5zuFwGOmavW/2V967XAwOHTM/6fPkWikRrWzEB
xC/QA9Gggl5Keop9ZAyVPTJLEGHAW2MxVoxzpO5zHA4bDvtupohqM69+xoplXfmgJlfrbbh2lCEO
fp48TzZVTmdY5TVyzd8ksIDgr/0Jag+ZABpzF3dWO0ipY0zWVL1cTTOABfkrcGPpzc+c3W0iyo0O
ax5xmtTvt9y9Sd+zpjTgctofJkQA75Lb5yzUwj7Maz8iFUgl22cJlAwoJI3AiAt/apkZwyp07MZv
8aTTg7O1Vt6nPQM6tPxN2fiiACnVYocvxiN5fpOliTfYhkkQWRD2/SI/oHKuD3gAIhelkvlYyg0S
+ED5lUUz1P/rYU7jO4988CuXKsajQENV218Dr4Q4kWBl33UFoPD+slk1fKW1da+8NyPoL80KKHc5
FQOhBk+pCUUOA1vXv9XVYirWk81SyiJVCuJAscec6GG+oj47aWf2039xPmoWruI/ZqRDkatbZUI4
edH9IBp349unCDsicabuFKxFJLHdxqp8A7WF8OyFAyB+KUaMJ+6aW1npQ/67qVpUhgEp/2E7KaD5
5uxZVfajlr/m6jj3HrdHLqf/v/eAmxaBJV7oUKz5cOWFMnOJ/tCf9Lc9npx72n49Ay5nIX3kxS18
hja6m81HAahNGr9rYvU+NiYf8aOQAJ/FIU+qXyr7EPdp+vJLGhygWWUlPjb7JrEWXV3vFyawUK30
I80xPqoQNmVxyvAVdlb+4hZsU1QrHQRlmMVquZWUnTDbo4mtU0PqbYToBvTiOKNuLjiJj6PsWBrB
azojhM6MBEesgQhcSQduakHki9wwIxgcQ70PLMFE2RD84VOmEbh+/iHPTB+y5p6smXjZ2sWU8fKx
QtNR56+6yPjJ7GzO1wxKCdePyAnnq9FDCJ9PK1d0MjxtUjsNcP5jGl3XM3QtAtlEM+8ZUnaC2VDg
/A0L4pl/RnhAvoL0L9PW9O1nm9nsMBAnjQmb4Hce9F4DKfEU9V/RAQERqjhx7IYjL2Q1jk4GrCZW
G754fnVTtJkE8G6ox45blKXtKOcCvRafycFbXMwOlyo0etL3ev4VtwhSN7jPKKhdm3KWlQKnhQH1
k5uAjzcAt/CqYgzOe7mb0Ey+bZcG/jpQDutTMro7o9z2hPPGUU/HgHmz55QM/FBpXrqTrlraSRjH
5nXpOV5zI7LaK2ReaySKVTXhWFEkJ8AgeUgGdrDKzVb2tRzjle99MayntyUsmPDs0+yFF3wUV2NO
2tojZPomDtzN1W4nEDtpot/FfPKIjeM9QZy2Vig2tuIQP1rBP4+lb2KmDPoO3+XLtRY/hsNlghus
hqHxAT9GNUZmW0wjMk62p7PVrhpdqwJ6+mvYqBSCO2RHMKpl1T/SMggqTHK6J7dvIneFpoKknY+g
Rj251Sn2rrCamtIeGUnMkHeTsEqMhjAuNDYutbsuwszCNC0YY2uDqt+XOzE/FUupBEDi4lrB+tl6
uIGwM/nOX563GCT6m3aEz9ZKUzKVtiH4YfffK9FGLVctlbmxesUrOt/w35GLxpj1BCxJSJKYgs75
7yOUhonYHbdUcX/+qnkNzRnAYn89aRbZrzjn+dvJWnvRK5dLaqyawo77BkwSBjEK4qBWDD3qwbei
aC0s4ptt3DMwyiYXsXpe6cdV7Wvv0qLbv8qFwjLz10mHmFJhb/FwvLf5tXbYX+8AVP56uMFR70sk
3sz/Tm6wGFrnpewZPWZ9eUOl4rRgjY9bO2UJ0xz9sQYj6cKXkdZQgOtEkmjjTv+DE5sNZT6SvCds
Sj/u1DXfqscLHhIU2PowHYDap+wJpvRyKu4KhbBtgEsiO4UmcnqhNArPfmzVYYTvMdBssylkYsxt
mwTj95/Q5QytYQyV6eSskVF69DMq7BAp3ZABz1IAORBP8JISbJAZtJNb3ooxygnnrDRny9+8YIHJ
z5f/oUybcODwKlqRnoA4SrA2VFfaLVPZZYtWzO9MN3i2BwCqfBnxCwuGfHk+8pTu1M6X13T1ya0j
ooaJI7dwzVE8aKqp6oUTR1UPVgo1j68mAJGiOTmcD85/Rn24LMKQTC0QuQajvrPEaQvC9C42Pl2Q
2jIuHZgS1W0Y6rVggDCKn1u9HNK0KeLkNoFCYQ/KNU2ka5XXTRLBeOgFGc+ieTH930Upek3s5hy5
NYc0kItYfTcvc0j4iU74KAmBbZQPGGk/nEmQZ3Et7pzt0xn0coRFN+1St97UPzLPxNpp/Cxf8kkv
V1U/ONMoYj3hYyaG31P9Wm4L4rK3rQqe8NQUkpZYxGMiTBuB5J5vVgpQzG8gnrGeZYdd4Gw8lejO
kOicr6foNVwNYJDM1ewJEK5+7ic1LxYJwvGZ5X6v6Ir7QIJCeYwUAsyTQoqQjjoDaEljJJ4qfety
+GjGE61mAsYFRt7Kv2uW0XlIGC9ZC/k8PpmdRoMWewdDyrckYJ3S3FH8vaAlXX1YKiWRflmNiO3h
2m7nA+Ti1ec3shkN03Nr/HpYdNVQdO8/qz3PO9cYVlZECR8+EZit1igkjHXMXFj/UkDvr3bvGRxk
0P5PMihBewFLmSQ4cfpKJ+xSmbiMSq5OPw5w0ghlwnwlzSLgUCXV4O6xDO1XrGEKLbzxv1D0In4f
0NY+m7np8gFFPYDFcCBQwEw14lgJcAVM5xWoVDV78khgSexPCk8Qu3AnISpLQDE/ViIjPcKldnez
yuHQLqMO0vo1vqemouXof2ZPPofhYB6JbWLV5Jsow7i+GK59JnhP6Y43FcF3HT5aEAMEBlRP8cv/
3eNH7e+GFUgtqXc3F7O0H/wQvwewYaplgSvM2f4r6vCWjxfOyRCUM30vYxn9BCx/lRszvBV7clLD
GqAcCbvtoAz7aCTfIOtXnZnAmOvczQS+yVZNdlhyX9VVTICswpj/kU+S60VUF8k7mcuG9XniTw7f
1+rW02LSjm0euBetKpCnRXKHNnSoGB3gafFqIMieZ3Be/dMKpu7q17n5xR3H28aDvw4rHTDrn5UM
7euCcY/dyZwBohvD3CAMcMuMx7DPHIvkViai0q1inKAI2xwS6IaPyt6lYgVypa4wljykHnF6tfvk
h1h89lmSK/qqtrR2MDJNOasFDgqxPgSqkWXDHPB8vKe2Zu7+NjSEas83Z1UFZUYQE95GOhGe5qxi
iZ7ZKDL/PG4ddTumWr75vhr1t0oj08k3/ol0xviak8z0TyMMeEu8FGUx7kf7gLY67nRo3F1jwRuQ
PtoithGnJgVTnnlZEpnk0fq9gQz2HIce3cbsaH3CwPBzqLtx41OeWWGI6XT56atzDvi9J776PlA6
CTEwfl0kLcCYuCJBfloYIxRXCKQANTrZhpnemp6CR0ImcLo9FadJ46dri0CfUcWLcci+41Eossz3
8HR6jSgaW7GPVTMXjX0AaYWi356gda5XVz+xOUDU6gH+kbY2wb+PSrHBv41ZvCAvyXlzvq72eNNi
Gl3W0kwN+wiJeQVi50aOAwXO5WL5KJ4UNxCjNsgU1x2YS+n7YmivYQ776l7f9V8CS7j4zegl+XNh
l9gC6/80POTrQcoU/ILBYvrWLXDdjSVd2tpQ0IXM8j+sOd56hsG21IlhQM7Lv81BjR1r9H3NSP5x
S/bj5b8+6O4MDVLLXqnK9x/w6ANmg6zYFUWF4S/1EuS3lvUL/e6CulX5Qh405UnYzEOhFN0knDIz
Hn59Z+cKluBp6BO516zFtHQ4NOi05wFXKyFLkbMYYdHsz38PRgMhaCgO8NZOlaluut/tNF8Fs14X
N6AyD0V+UVSLZTV9H/LJzPGsd1XDoNi7BQvKATAbbjuj1707NQ7IJKJPh9oe/GK2HLfToJTfZUaP
TEgByhRMYLkxnsmW/H/ICuWiXGclBEEInrN+xXZL2pOzOBKcHRfhNzv5NfNPCh8Y60sVBD2e1AhU
tYnn+yUHQkDEmKI7BRd5u2e5xLj8pEGHIb6TTrbRvRIdv0b9v8mjkNS2tzHBvO5vB2DYxGgHg1c0
L0qKlLlrNf4HFrkLpWUr3wRBJjlnydmxeK3bHeWmmx/3UNuc+v9aOp0tZlW+DWbbe1krt97lJ4Ai
ValCR7Cw02KIJjxJv8eSCjlHOCsZLWwCUTYzARPuS5UvhUqjSf4GxqsmqU3T/FIVmJKM60Bp4jo5
YwKc3eMjp+geaJKqzNgFDEbPYUuPGsjJlpDu9M2BUbHMz1exUgVbgXtDiUUTCuka3QFAiVoIZ5Fu
sM0JOud8bBBBPPuFh07qltMaXiLsm3ewub1hnH7GevZtjinPsDvKYQrr/IZsbAXQVha4sDJCT61A
ITzwPGCMFllkkBB0668UjejXA/mmp0DYIkWHinFNrWVVC3e5uhccurpfs169BIlAmNhwAYi9Cx75
E/UtwFAh41A/TWY52dOIVQaUMg4wBbulWY7EX+Xv18MRVpFC/Pwu14Tr0MgpFr13DyKtha/yP8Mm
+w5POUWY0579828VG/LMzFbzBxgT2lFsimpzqbpJW7OpkCcg259WuV1iZrqqByipIZWWWxiaXKNl
usArYkjDOQPM2HxPK8VvjfsNzVSDI5a2PUzuk/NEiOF4xihFqvKp+LqQ8kKMWPI7TU+D4JYaeUgv
n72pyFPzqR0MgHWjBR1Yv4BnPLdY2gLdM64DUHtf7TE50ad/NRCn+2XwC/lUjGRi6Y9fZwWvLJwE
B/hyhg1LA7zAuU5GCcXOEsUYjUEnaK0SUiLPMmp4LmxJLdh36wxrqcOlIU+aBzhqOhpUXrXdKnLa
jlxPuHlb6Bp05srOw0zbfVomdWSpYf8+Rn25Pb0ripd75XLXy/XOsWx37d55T0t5R1PIBQuT7oPf
PmUt8pnuMlq2VhfcUhc+SBFIFmE9fY5Q2f3YkUk9kYhr8CbrSG6xj97+Ct3xvxKXV7/elwLT7ZAP
jZqhVFgUTIj0Ye2V1wJGZMQEK9Ft+5QtLEvkcl4gsQ+3j1RHRPZ+WtTIZFlFQl6vSk8xuqhLGpQm
1hkUFdASj+Ha8qXU4DbX856zIcfsp8u8Eh1KjIkYLMU+7UfhGhSIOmCTXaTQp1NDUJ0H+ZWA9CEj
H88kUn9l3qwJKf237hwKGU3+6MAgL/1PZdTXfWb3SlvqcgpIMA9RF8nomSkfjfh+UVo8GoPlBpvw
NJeYHZSig9mMAH5MectSsaAbEbfPGxNh5Lgtto4GCrn8Iost8XrykUqBGNxtSYm2XzjSNXVE7Xrx
WIYHEE8YlbtLvxzGdnrKDtMkocmK9yqDsQiu8qBqYLK2eu/Mq5RVrQZFCSDo0NVi00wAR2scS3oQ
oRJFE3Wx+Kqr+RwzVI1p8V/GegWR3r1U5xKqMYMusdOUltngFjyQ3xzxvyZLC6UTlFcImwgdgUgD
5UGCLsgduzjq3CFmnRbX4SSEB90ALn+USYu/axcdRsj/P6NnPfEqpHNP2bouN0e5DFCuhVTKSro4
t6CsIHDDzIIw5RhnH0CR2GIwKOpyFm+m16xJRrsrG99Ty2V/7QFIalXG4drjNYpd2kfXSD5InLBz
LhkhVOUVE+WTXP52ZCXd+/qY5v7v4v8c+lAgbFwCRY3rjViBKYCQQRc5+A7pKdjbLXTNgEyJ/vsS
U0iJwqd7cqHnHdvF0+Rl7FX0flINiK2DLQtk5+jpMwasD/nRp0X7gZewAoHVnWyCAcdwq2BmbvGm
BRiwIzxJ34WpOEMHBjjhzK8R4Yb6rjj25/QXBb2KDcFQg7mLnU8eleZ2wZlTFfIIsUofeDgFWRbz
6JixWUxRXwVyq35uVMHHxhC2Bu6mXK7E2+0492e+cu++eiqQb6KMCIqSfrynjriGOSBruFbJ7GeN
A4f+MiXBG6t+kJQcByjp7tKfRp0crloh0dTUk8aDJM4V75BUANyrLx82yCYLKzc6hou0HGxJzUhU
0aa1PtpEgIQh0qKizreZKUf0PsOTjaOBZEFIXdzkrE//QVxZ1V39cFKtj75pGQ0X2lmEyl3FdnaR
mVx64ueZ/GQUyjMrsrioNQ2fW/9cT3MIgoDWDuNHCeSsJtdDJLtR7ETErU0S1cbjWfsQvyD48AbA
iQwk6e3ZhD9MeH8ABeBNJ18GXdFtuNeZPK7ZMZiQLL40DFEjPvdBo8vzbxu+AZX764G6lySrLTMh
sESDzt0VXC6T0XF+eXaK5cgi+nUGjpo8dXVF6NV1GyWZ02s2+is1PzZwu1336+zAvgi4Nk2JmWBh
24LPRCS+Gzi+vMdB6Abo2LaN88LZIB2Uy97oznSWGJlsohj5AfMAw8OeogS0O8uYgm5yCvgRjrKg
u4HxW7s0+sbCT8CrkCfvij65ma1iv7qdFp0lKjlLc9wjkcNUu34VAw0D4vTS9H7bfbuARp5QkDru
SjoTht1KXjPNZcL3daV73mqQk0XvGBsRpzUC+8kg/t/r3eUBW0YrvoNPsPctAWvVAsm3d7QBuoIe
jLvG5CnAmjP0qRYtaLQITS20qClBPHwXCtmvbcahVZcGyzmukgkjOZeHMJVxvXCtHyffRD+qCLhw
rBMwI9k/7A2bssbNo8zcDVibfa+d+UGKO1aIdGV9SvYsuesu8n5jDt5v+Qk7H+M6MW/6WTxjUSVn
3IXfdWrOEHAo6llyrSzwC05m9XPeVhZmpr4yiYiPS6q2X6wQMulYzGx3EQG2XGPxBmGLdlLGHSEF
0QC3fh+t5f3Ccvy94TESreetoP4bLu9U226x4eGjIBnWTBhTRrv3qDq7udUtxqD8MKmDujg87zCb
KpOmhCQSd6OglrNpj36DkZAG0WINFsS8Uy+FYUrZ0HE+yGhIn5HUUkXwYJVHhRi/M+GgpsLBHGv/
vyoUHn32wtujQxywYk3mb3RGZXyUnl3NF2OAUd3iqIvW18j5AzOTzsshVptmVoLA/ci+ksZluhld
cC5f6fbKH30GkNYLzBjRMXgEOpy9J4256A3bwd84bNDvj3jX+6SZbWjyVOSBWN92KLDf7J+LcL+Y
Nd33PPQJxNI7GIj4HkibXwROnuyuCrEm7MKJib13v9+WnraODSozH+jefolMJthH+EY4h5nHVBVR
K0sPh+g9sMB5dI4HWurLek3ommgSrlilo8zSHOLUj37JBfJJX8fcSdsoZwCmb+8AJZJRto8jbucW
B5hdJKvSKRs5XWotq4pcYOSk9r7fXyYpax0Q+2tmgnW8UxY1AEk4xI+TWHKAe1TTaFmEA0JKJxdn
WLkiAVlyT50u4cnakcYboSRfPS6Re65szcNl83UmKo2tC3wpcFtqmMrkMHFCqDhSg28DeDubRd5E
KcAJAvGFjVVOlJ6khN5OPYo+JjNyatWipw0GVU2yMHJqckXZie3iEUTgNrJlCygUXsy3XXN0TiTR
3iUi4UGxm3ve1AMTfEnsHCu+vXE/st3wNY/KdhLll97Tr3hIKJRtxrzgaHvihfdMJlKckS8HhruV
vD8BFYvy5FH+++M23yl49Fd5aNyNiiYkrrVIfa50GdFfGZAaBOL0etJ3p8NX0bYqogcjHpE7blWb
Fcm6Gx2j/+p9RWFgyxGqiJ3x5YXWiFWg00sjC8fAac6xyJRtyoe/x96WNlM2y3xq91HiYn53CE1H
jWx6LNzVOsLHQO70wQ5ByGz0B6CoRH7XBJX/dBbTv2mfs5AMZRJGokZ13F7g3+ZtomcK0VkFuILZ
bhpdKIrzBZ0RLdVGka4AzOzca+I6/FHBjLFE6VdoCbNQeZsqFjiieDkoLMeAhNlak2EmEGzB4jEo
LdB6VJI5CRfUESRCQS4iDSEJwylKFVjw0yl8MV/tWXcup6mi7rpbNTFmPfegcEq53lI3rf8ZeFBL
dTbg5UL1vu+PK5rJ/eeXvImJIBRZjAuHY6VJ/gMqMCLOiq4dsz1WvJt1wpysqBod3LRcaTYmavvl
SBmt+UYpb17hP1dI+2P+je3GR5NDXshc0cMCqSDbj7d/B6SKMTN/BZ4+5ioXLMBT8q/AeqGR7D88
KcBJQ51RcZBjUe2dx8E52GqtAnAAv8LAKWgiyvesBdfZybluJDe2PX8shxqCZcyx57ssz83E6jd5
o1jnxCQildBfLd0AOV8Etqo/KJV/r6p50WpFx7DJrIvTqqA6ztgu5/owDlHyAN1Q1LQhCdLsNyIj
OgK7i6oFrAVNSPT0mAv+CMPhBE4/6W30Wqmlfo/TK9eFbU2bPv6rjHJdd8t3Ec4S+uju/AFfdLxN
X1vFzOLEEB0js4kvRqrFX2Pyy6Ej8Rrm0fmAz9MmL6ekJ9wmnm9GxsIrHQDYToT9PjgbCcYV2qVa
O16GtLd0gLDsLodXwusg72veH+5IbVbK6VZiBBPWdsqhfUuq9jn6YrtRyW01DJhtNxD30ojdJYyR
Gdax0qgryjdJx2pKYc+lpjPOKUJVhNkUvYm60cy0fioANIS8R4eIdDz0N/6GmzqUQK3BhVzy0tM3
5P9zWbgsW6Yax8rTfG2PIF/lSTmK/Y0tfxfqp9u/hkADae+Gbg2jgEpxjAvipWxomzyq6JM38Jtt
DWsLTIraXkldjJgNYqapmTJnia9jJZ6LKXP5wafRFI4ZTJoQkA5PewkdMl9T5DO+RuSR4Hthjch+
3Wow9WPw1XSTuldNcMKqDrPxHlrDExND4TJpbXYLyxIlFkcnLtkXnLTLV7Z76SZufHIlYSRhYcBt
2+EZIz7qfPRmMqXBWxjEP1aNt0HQgjgpdjM6anksMBGoVMSPnkUcpkjo259s3oa16P4SnK+JAZ0l
V3n9l6+0P699s7zzDhTooEXN0Kxf/wVFo1YB7wDSGzUArxWM4ZX2WaVfvJ10ehuIALv4Qi1LTdmP
Y9uq0ml1f6l7vqhwLcng1+LfId4cMrm8gViMalu0FsftJodlgphuXR7OTbd1iP5HsUoaEKyM9sQO
GCCcJublqDLdt+TlsweCvpawZa+PuE60Dz62QX5whA/cMXFoLpaF/csJHYCNwfzUm4aZItC/bN9m
jS2DlvrP9Q9mjjmps+WQVZrwniOtbGg+AlkRwCYClvFD/gYwwGwx0Jk6uxXUwvkPigkrB8gImS3e
EdHC8/xSjG+DecYTK4qUg3pdgeCPqR+H4O8y3TBtWE66MK9o2SfXfLEdNb2/Hp3Os8hrX1eHGXnR
+4R9guRs1gDqacGFD+eiLr5Y6Jq6NsYSX9ivbaI0OlLQcsmkJFO+O9Pa7B0DZ6UqB8c+wAYgqUAb
xEsibVeTh4qUsFWhsBYyPTjleCG0jvUx4PIlsnoODSvJRAukgumvvKODfHiZZsXRfX7HepYmSx6I
sYPWUcpS4PYewzrArhtX7AeR+yfiht4MjuDUM/lERH2wwu2//0JpbOgv2SLCN7kLqc5djESU/J40
vzvTpwnqLDOkf5D9g/gR0M7ppqNRrt8+AcbQiAQF6mhtGtdpbn1/1fXRdtOmnueCXJXaw3GhkRdZ
lT5qRAOUJzC+YYzrFod4vHdm+jb/SGHAjAsI2lreUhhuCUqMN0kwPnWUU/p+rOReETbnpaMAVHaT
G02V1lW0UCziT2vnrypBVR9K1pqcdc9aYhejC5aDsXc9GbHI69zw74EI8sI3KkpCixRBQJ2kde6Z
xTpFlhEEPgltQso6b+Kta46yGSgjFQsHg02X9xk9/rR6YwttwWB8cYthXrq7fkNDty9nKxqlKfCW
sez2h3XK1schG9sdjERKr6XT4okEi94qKvM5LSomOxWH5tvlwQl3uzA9Wf3vrNDXWEZU6YTFBzul
DSmuu2R4Tm+cBKx+rHh4UzvNyIzq6C+XiEo/3j4ECfOZyl25bwr3o44+0aZfWaLgbqT4Ukxv5cIA
rmkxDDaIsVCaTWaJeOrQr1EI/Dir9RUIECOy/U7hDTGtrJ0kRUq3EByC4XITl4X8GLwUTeHuazRP
UYHUFjXVcCJH7nxZ9t3mMu19Sy9Ouu+1wGrVH6c9oFzzOcIkcuQvzRXXFi9tk4DxkegdUbRop0vv
f+kXyqO26J5RS6DW3GLcev7sMwz7/HsZSGVx0dMR0NeX68a9pc7GaBxupGGb/K/6DqB2WJHNaRdS
kBiJhra+9l81cUTQbbds99ReP5ZupgwWk6csj/MGL1jfwHfGFe6e/6fgRlL5uLMwc713RrWk09PH
MuME/Vt/7bEho2+DhCStfwKpOCuTe3HS8tDA4Gnk6ycZKKk6WVkw6w1X21HtfWlILUxDthKTiwJU
Sp3yST8FEIO/VuKbC4qtlpDvtA2z6qWRfeIsVi09szxGTkySAX8JktOzkXzXSYfro1/7ZmpXQmiV
N74uV6ZKtPzZSferjb/yAy6SjWuz3v+Ti35Lhbn4RA10K+nt2YKBBykeuwlO1MBjzq/jeKA5YzJ/
eKb9aITGiowqsZNhfVFP41Dyn5M7eLs27yUeq5hEuLtOcZFI03E2aVyOS+3tW8AwE6Qq07BFdyio
KVRKn5bl519PGTceqb5fNTBz8gwo75vo5zdRDQIYmAvjhXCnCwnl7Hw2UJmKtaZGRXD85Gnancsg
E3/AbVk+fchkEs9h1BNtk5NexQv1urbI3wgsXmdjmCcBIBbkk44h7gvtUTBbKKDps2/IP3xONKh/
Ettx1FowlmBVynBQhxdhnSZgsgWBpIo50wnXlBeY27CLXkj0m7UJZHl/RxLj0ZtLEkzbufQZ8jZy
FrqnvuJyfMrgnEziuKWhfq4r1AImI3PdDsf0GY4eoytcjvZb0KVSOv7gSFkjLQzpUDISTL6gpcBW
Hwh/XAy39/CQ+9b8kuWw4vB3ia1MLp/VTA4sNKwopEaprKvyfWjagxUff3kUVs9HlCqkRG4iaDC5
at466w0FRKaiNfHM4DtH5R5UmqB5C2wE9lGyjurXhJYw9jXo+/fRVjAeWA2V66LQm47hPRiObEiE
swIxLvhdJxiIw/3+m1IAnZ4zlxEJiHJ2BsxDlCiQJqCdEomvenxSf5Opsuqmps/TxXUg/V/a4bBK
KEE6oDRaGQ9iIgffph8jF+2aBMeoNaPzlrp9EXgzfsO1yzBtUQgWT4qx+ZXoaMuCNgLdVo0TU2Nc
dSOvCKn4HekAE3cy2ej/fCEkD+b+0vAhHyEEMgOHPIy7MyqyYP88evj9fv5HweAe1xjuENOuIAUN
JzCK2cF8ifioGlU2X88g/dx2OPI7Rs3V49aKx3ZG9QviaHATCS/AlzAtoet6GYORQlrEa2IX9I4o
JNaPhMiEzWYutSDA8yHjbG67wbv3xntmxANSrKdUF3ORtiqQgFeMWOjWaEjZsFOVBQG2QqkI8QJv
8rY1XUPd9S+OeBsjnyVa9DlPU5cuTe5yQ6TI3weWFLIsUE/swF4JQJ/56pN6vE/AzjhadaSVJ2eG
WwmUlG2+LIXlMgkEyGDwosMuwfKsCaucX5l7T8cHMlHGLPkY0SrqQa/s6SJMQoZimDG3mmo8J94V
MifGQmAcEu2PkRajk+hCjyaIJ7NpCeooo7fp9UEOLxTlV2gEjMlZgx9jy0ZQtUbk1WLiwSWfZdHV
Tqf+e63ANgCFAM3Mc11+cz03MXqk7qWkUiPZqWLYRWfBE/zCWAk6AmYiFSU5DZ1lGEUlSEEssYeU
Kb2q61SvEeZKHHXgAHv7y4ZOrjM8fbyO8C5Rz7F/PtDAYT6+u1nmYXFoMslHuFQzIkHVWeT1xtNu
ERcFfOTviG3J4FIBDCo17BlntNV6n3oDiqAVHgxwhNne67Y6fTIi0hCMwx6QntX6YASt4ho7yhOn
cq8QOy4rfISb7KNLJZuI+SSfR9L3lN5MRnREqE8wFaIVLJhUOtv1D8LKHl7S2OjpuHKWIB0ZsgnV
yfKN9irbCVlJCJImvYXztebKN+MncV6E3Q5j+tJ5hr3j5GeHzun2cD4eoXTIU2cArMBr/UDxb40n
MIcM4/jaIYgUjcgUK1tdmcq6Q6Byod+FHib2HI0vUuOSgWNFgSTcRNZvHB/7sbkyK7rXTjoqaKHH
NYuktc9dlDz7oVcunz3plwt4dHjvwYF0UiB1vj0RsKabukcNbs0vMsrw+RVkJBj760VmRDHGU2Oz
vi27u/s1kzVcdtWLeXzMQlSvVEeAdjy1H/qbHd818wUnYYbGqnsy8a5LFFKGNI5HT2uMcK5X/TyO
CWXqRzMHdtnHadYdLX5NVomKBU2Tr3zYerMZ4R+RyH1KoWz8opUZDkQjZw1wJLS0EWXtJP+mNUVJ
tpKwAiUifbrqZ4IK3AzZHm8JKW7L2qjlJF8p8Y2ed6NuwgYriUbtUq3Eo7ePZkg3uw2mnm7fCLYX
y6Wu47w+tfFXXB9pONp5OTQpZjVbuUwF9z8Upo2qiQuaoSFS+Kg2aXrJdLzchs0C//oYjK4NSsZW
ynlievceJDG/hqoLO/1zGk9qWIESBE9BDhtS8yE1JFTveCF+3DBjJ+5EVO+m39baX6qwHnLO7dLd
q67F6dhYG3MfOnyFuRK+W/ubLkeLT820yG0lywsLMgW0kYYYBUObltciQNIm1u2ufW5T1m/Q2SHv
8bdTTXSUfvssouOkLadlG3qb8/7qhLwOX2/h3BzACcJjXIWhzDsrO/Z+GpcgqJStVhrgWO2HHR8k
FjCOw1v+RYOgVXkAWBTTdf8b6B74VkldciFyoBYyGpExZhx4Kz1JTfrVxtB4pu1VZiZY8HRzPlUR
9OzCDMZvpAnwlm1rUFB33Vw6e/umDwk+RyCqdMR2qv4vyro/q77UeVgxUjpsKWg8aez1ocLqq3lX
+J1Md5DGGoSEhe+mxm8uBOZBjeTc6yk+4N2wt+JiCRKO1I26P6FiSSnVdT8RHV+q/q0KsYEU4IOc
P0usvbMO6uPCZlZ4okfjf8rwkTySj0aVuOt0CCsIFhmGSE3PZDl8GIOOjl+uUrVHfeBkheIgLMFe
18XT4CNt9UDmy9waWN42rB102dJiNigHWdvYLicSFdApULy81e1KBp8W/iVQM2LFb0EjKK+KbRu3
0Z2S5R8xl2qOn91iaY0E4ktifN71r1DVse5OLualgp66g3p4vyb+dZT+f+I2Zu+sofYtobxkLp2M
j+dLUdcbF7byr5hWn03lEeFODeESjJiRDHoC2cxvHMZD1wTJKpfwxcZa+0JFDFH55t+5U2AAYoWA
gxXcGxaOrOr5DaiSTTx2CF5jCKcCbi3V+ssRI2XN4EDoDTnBjSB8nmrKRco0CJ5sBOWD0iPQ3Clj
RTZQfegvFXJJg7hVo5wWnKuEnjMMiHctEDuBlc0xZovysTFrt2aR5WngkZ+NRT8R/j33G6+rpoa2
/kysBFTAE0lqHxN6Oq0QXpsiIG3/Nbujcsnuuk0AEDPcpiX/nFlgmQgDHEVHmLlZvcwCoMS97M26
nWYGRxF1yn4bZnyui+SwfoBb3rjq6ot9L2YjdX1d+xwGewgo/UR7PGDhdraqpK1ar9ylqUmNyhzH
2YQuEmQz4CT4wpFUxlYYL85Q8dD2abj8DVIMHn2vb9sevLjjE/4tY4k+vVdjurc5cLE/d8iVkbUU
UKkb03mea46HSImmc+Wc2QXTsoMOQXwIbs8164I3us9Ywbc1POd3RfyG8/DjEruc2JXnLO6QvPiq
ZDEOdSpPY1kpL2yyibHH/9PggrvGAVkFBl+ubtFthAw/1w5z1fSBBz30XD9KzGr1N24wBEXfh0Ra
JoWD8ncY+zuRzppxhtzZ2W45jHDUE5+3twFLmvk3Fp1xQ3r2ngwgMSlEORNViM78P8GEIYqY6nRX
VPNQ+JVulxZR1UmB6FT8ITR5an+TZnjohO6VQKXqWev10IHUnJyP8VKF2/XwVWi8WVp/Yteh7ewy
gVOpyKeWoIcKWUqmXfMcmAZdXdsDL2TVjWcL0FgQWTiD97IvUvl6VaeYU3JyE5TBW9PELXYf+SGO
SasizknIiIf8SlBltesP9V8xszKmAuTubft+maDt2d0oON95rGszcaxUdU3vFw0EPs5kV9xIQ/62
Oe1D2DvkfG+TL04yDMoSvd0JvnDRVLgEtWnwyPGEcRLbrtF+NOmtetklbk1PseATxHgNDqH4S36Y
JkYVvlkFd3iYPbrsoWX/RBV8JPfLnReKVAHRljRzYCpBgQklM0IuWfSamYgMEmfMRs9YpJhEbKUf
J+IwwT0IxKEfIZHYBSM/HnQJ/HAAZV/6vx0x64sH1nS9eJb5KePwFdUBXJv+T3yA106J8E+yy3nN
I3S/cEEKhNgL5AoynWgnnkeyzto5BClCJyzGlXzwTPuKOWBwZq9Xd/YoNiEN6oZSZZGgdQbMzl0m
hldYjhvCSYRhVkS7aYoXffSekaM9d+lXhq7ArjvX9SREeVpAu+CraMjEBNVJviGisXQr3tNXn9PB
74cs8YAdciIhDGryA+ZvZeadigNqHlm6cx8rVodaMfZS1rvYvaxLnlF3KZuYiAcpbtJJaTo7OJ++
7gtX6mgu17oyNK6b07EwcYkbRQyBTKLy5ULQi5TalKcYgaI2/Iq03Ub0C6H5S8cGXuxtvT53965B
jM8pHf9rg1MkmA+OVMS4ZGhDtZaTwciBKG2Xpm8uZR2xaAzydtxvggIoo8KDgOUXZ2iYWZ6YGPjr
vZAnuqwXEQkiTJwSG3b88zsiS36nuxmnRIepFc16SxvurIH29WiDmd6VUOD+0XkmjFUUoDhXlYyV
lCwDVKG07bszZLNJpuggjcXQUzGC8OuL9aKKcoGDqKxbyEAZJ/QF+LMqjjqNwyr79j/UEJ/F/kDJ
4PnDKwDXtKGLY4fgs0LsMlPLzjnX0Zyg6zo2i/jP2m5gf67SgBjNSWcJ4BNWn95/qXYHtnk1+UtX
GtQcg6KYVC3hIa3ZNEZUs/7kQ1My7QY1s4JlBve+KM3/OF4zXCvYQRjY5Ghm7pbuXneC7nTWupFk
8gLareFAz5X1yKfzzWZ+TFDd5a6voGVkvzt/KE0Bbqr+0uGtrLGf9Z8HqN+c6wPhbi1YIOY3Iu0k
dADvlQJ7ESB2n/GxyqxoJtTvKe5peuqHtz8N2vrukuKFAcIX/Ahl5/dnBtaZ96flx8kZTfEr/6QX
FDCHQ6Udq+3OVe4/pvxHDL3Som9ORR2hKA73/1kKaYzMj+oqlwXDpCc41BHIvdD86C4+DM7P+7u3
x7Si4xHYlfekuYFXngCPBeMKi4h0AeNENXfBdxqMXki5LkKRBgaG4SzHJnDTSlsbYCLGHCZpE3d1
XYpdqCjUbUX35khxsFRbdiJKaaovo72DNLh5B1N17z+Z55uvu+EHu5yjv6AzZlR2sIwlw+JzN1DC
tYhE3NysgqrQEPIBAGqUf/0ZywYVhwy7ysrbUmsnVEnR/FCxxsnYoD3QoJ9EhOIhAm9uHJn9HRXP
H6ftZsYtnQZcuOEFRtwXIipMRVn+SaAIWoVVAOlLqfEKblgi8l5ZvPW7uycZ2mwAXih6Zg0Z+4oB
blGWC/asqj+Zo+vkti4WWgRS5Pimg3awikYFGS6GSJKTWl2XvVImm9Nlrz0cXZDYjYL9P8jeVMSj
Kthgyk8uMaglISYZ1lvWghhFQuLqhF8eWM6ZGVOOTdRtaseGTEzFeah9X7mINL+KiXf6TWPzAfvq
3kyZeaPhTw4A3kwuRMgqchJGd4GR1r8oS9VaZWHq431WV0NXzHCrevBO/EW0XBqkT0vzghDdFNid
UW/kgBa9r5hmHx3A/3Qkdm/bv5Od6PK2n5vao3GjpGVL37B7CSoJf0jmN8hF8Gv27a9XriesPpSg
QPxaUOO1T2ukyMKyBPO53S/BveRfJYwccnuo9+m23mcFi7ato6gTwcIU1hxhG4vdYWuVvLXNTNZ9
DRJFbDr+fduvcI9Me0H7fWwcisMXfh8hMqicfXHcn8XmO3WBB4DA1jv59eIuqZhdGhMR9iG7Kx5x
noVMWJTLWDFBYvUY9TOL4TFapWzu4Q6lg0pNxJzvF8+0b0DnNA44w6kWdq3VQ1BzV5046nvJwx6S
BYPiiZ13zfeKUONGXyfFUWrFT+Z/TbH0rL8Aa+HeY11RZNTWdRwGDw61yfm1h3f7uL722od+cBaz
lJY1bWdqX60ANISluPAuyO/Nj/zjhvj2IuhW4v7N6mYcIhgTEuTploSXDNanuB0DZ3mXK9phmcRr
2JAGSbmVUSQKyyfiMOk+id3g4ZFZ4P9GLoyBWtXZjeaPxHR/0W9asdiJCeYFoBAxvS171txECMHn
yDYYUajCYDafDw5Mvrn7ca5rsDhrGoUrG94r2HAgnHGIYw6rsFDFSzJb7b9KKBsJTZEoLbjdsZZx
3EV4KMmJuD7VLn41Zd/wYZ5ys5vQ0df3TUTFjTJPqI4bFPXIZn1xHfa2Q6NX4Ge1/LVNrJ3ofo5P
WXme9Y3l1KUsLWKktIsRwUV87EK5fkUv3kYMAHApXZz3EceokeBH0zxfwXT9Lj+YGimWcRp++060
1sZ+jlxNc4EWxIN5pZk5GNbxmkylGdBt/Mq2LcmXezy65ubRDURc2u1F7HCFgIMcm+VNG+JpRHvZ
G2wzgu7kcmtaun9d7jYNwRk1vsvDhUsdOWR17/yIRC74Wk3kTMffd+e1ShYLKgNDaYP386pJFCd/
dwbrSajkXXZW1AuBmLx5FD/at4MOiFLGvLPWKNJiMi+0wf5j66nborF1WOOAh5S4XnqBTlzeQSLT
ph4C6bakTqci2ij471QSqe0jvm8s6ONs9qxjnOD//WeX/HWdpHEl674WECOVvZGSPbuRwvfhm9WQ
6knABZpnu4bk6yHR8M3382O8yC65b44Jw5CfEuSu9FDq/jGwA4+k9ZSYeJVFY3xtUsOZmiRdtTYX
5XLPVcdi0dcB+dmsKfrJqRg5rV4M2jvqAohMwvZ49YO9uTMSHH//MN4rIeUNT7zVTwDA/loT9Oax
KzSvKlFLHbA7MRRJnlpeMUt5xeoZVGPCt2odNQNykiYEs11XElj1MTLrGf9t/tZ7jzfiD5ethHup
h6yqxywO7XPlLlJ1CQDHXyoni3ccj1fL2neFZQeECLmJrfRyw2C5PKAa1YdS0IdKTvOk6AYpY6+E
ICQIUbi4apM8qnhsFEzhxExwkr4lUBDmYiVZSnzvwPWH8gsevVAM1uWjMj3/69YXB0kHnbqDeGY7
pCEVvbMpu27uxo6JjhA0mNpohnd06Lj+BL7AKF0JlhltgGGbvQC54ixk4wGgR2Rxeav7EMc/YwWq
P0utQ2CgG9iFlF2F6CBZxVR9IMHA54eCGtZqKaUowqxparo9iZ2aAGC9j1P6kea9enRQBG9f5lte
ZV4xM/fdGZdwi0mdShVtOP6TSm9KuiIDcJ4pYir0VywMYSdnXJl3CwhfgZ4CVa+jcr4WxabR9AvY
yXWeTXvmm2XIE8SyGechr3dfbBsm+dINdbG/hsoo9sHY62ZMPgD/a5EcCR4h3G5vkGCsC7jXgWnU
Tl/LXzgZqHMkyETZrq5V4Es3Z5ZZB+riqG1PJo6b1MKZ9M5fmgQsBFqL35k3Xt2yzJiazShMqvdE
jpd5odSvNjpYgJX8NOqtYI3wRKVYQuAUmDm+amOmEh2SLjtVMXZaawbsZmpNUUjmaQR9jgqtqKDb
N44OwSh/53nb90fRT3Vt5DTwAAXNg2wQ6rVipB0WeutWELEu5kXyHQeh2BXprbuU5kITNA5S+4Fk
DP2/9cb4bw7zRkXdYOhzMC3MNGn/NGQ49GFaPTGGYSTsvksufrDAL/3QtI1ViPclfEymmnS0BkAE
FMjVZFLFe23oPnSeW93fr3zw6yjJHF7lyFfKGUjGFrGVV/1d3ULMSOQGDRiDTFVn1uT7CtocDnzC
YHlRGLBush8ZT+LUGaNK2dHbZEkKFMVKWb9vd7g5zXE0FuL68HiGe/BymxSTPv19SAyui/+uhwhC
Nf7LmAB53dd7Shnr8xiaK3fjK3LsN54aE2XFkoBpQPOwF2f3DKVgTHXR7A6oIftZPYgfhEJcYW/5
ZRDi5DGycROK7IppXPWRCE/PuGodJFOA4z/9yDunZk5fuy2U5HSAjBha91N3Zf8SgLpgHRkOPFnp
d6VHtlaCQu/lAwf1lmyUlROTf3W9+owNOgof2WRLugYjnM4DnJl1DkCFdn6zyraSxV06qKPGcrL1
GswVYAu1+Kg3kqH1isg8r5n6OuZfG7y2SEUGEPBY2LCAijNAMbSZ4k/HJgSpYIN9d6H5VZ/yWPT+
w0/Ix7nY0lfbKxCI8NA97ERqOnHR342hN/N8V8VamGIRbHMUEmVJPY+f40eTaA8tmEO2v37DITEk
M7HnzdURhyoxpQEm2Fz1p/C4qx8rZIveT+Teh0bwv1RsPTn0FKDjxwuY0NIv/u7Lh0J4f9o1GJnT
9twceIEUtNeMVGlKFwldiANDw/ZCZPV1bc/15NzVQzwnEnfTji/8IMBK2Sp8zeIKpZ+EYllLP2VE
tl7dnumyEojaLatq7Lq1NZI/r7x3cY38KjnmFSuXttrOHcB9/XNdezarJNmRI4iOCKDvk4xMfRhI
Xlyifkr0PdpjrCgq10y+tToZHlwdKVqJ69dEDckEw/KjjNr2hTUvITSz7VoGMDHx9GOo/BYcLNZ7
tHtvgzcBqIgFWUTvijFaejYeIr82ZOUpCi5E2Uf0ABzG4nPF9cdPisa2K+Y0u3xINnXaC+Zy2tTr
4xHq+PjU+DnEzIpKZAGQQWYWsd06qBVn9ACP9LWyJmfEuSUgUcPTuCPUE6gUnq+Q6hLkTPkSAQmG
LpIO7xgCahE/XW+m6k378hu5pk9DmIxBKiHfUawaYfeUgXWXWziWUaK5gh9pA1MaASBvXyU1Xybs
OgJBo+FGNnwvuZ8RufOzwSOxa58klGn0SKSrOzCBas199KGYJJC8icPCBcggi5WjlbwGFnqt1Wdg
O5BdMCqkt0b3vG7y2zd38ytW5TPUJlcXdp82+S7II6uEF2rhgGBmEAh3Pz5rOXhrm0A91g6auedA
xaclALAhlcN6SVVqffdpYEVNarRkx1Kay+mWON64jZGGMv0gWgsUbe8njNA2F4hZceAaLU8n7f5g
woqG0k8U14wYmKKBbdiA5qsx6CciffD4logmSoO0Yfx3wcyU6rLONZ8Hu36DF4k+4Y5PG0SCwLWR
Y6ygZl9CoY+v3Zo7uPROl8TWbfGNreTIn4yhcA8XXBWS9ZqOAWdX5adrZ7cg4Mo/3MadXXuTKZOy
re8C3GHNKEEZ1NOn4oGkvQA0vrJs42IbcmbFzPweIPqHs/RaC+b2aqWnmEPeHwcG5hN0vqHQvDIb
ji5QyhFf7EWTMhsEeAkNUVdvwtSDICpYWciY77bMUHcbOH88tlO2mHsEWrQqnyW5T2xQudm9JMoI
blGmb6CTrFIs5Q9IqLA7IbnxlmH3u+gsrwCi2FQEtp7k22iraAimeNamX+/XJCgXXSM83E6/w8Jc
M2+rOkYDdwMF9BA8QbFrhBYZkXYvLG9ukyV1jp5wCM7rPbN8Whw7y3zBIEKli3pcVcEHLRcxZrpM
9DojIsmxOTlaqjl7bcKmQ6MQJQFtIJYHovvYRSpNZPHFs6vp13l/NPX0rcRds4flXgy3hL5SZJoo
b+c90aN9yTwHmwuQKb6texDxhSncxww15eytWzSf99MsgRiyn1VvnRl68YxW91axY736BC2nF9O5
9PfjgUNWuLmHQjJc2NzF8t2Q9WYTL0L2gAOHiCwFFy9/0kVU/lM5iPSNeNAaa0qbjwUzTfAavG3i
MiFHs5yoTK0XVGfFoXGiHFBPSTuczFF7jehsBY1cEtxFEvCCYb9QX49IksYCVw/qvSN6Jbu6+aAy
vn4sS1xlCzcyj0vaeJ5uBJG82fwUQ4phWQrhCuMBUl7slVo/T79V5n0TZeSQgAflQjztaXQN72tr
OF4L27a7Rx/k/OucQtZjkK93kb3Go+QOqcnMaQ8f8iMcZZbQksde207ImIJPszbIpJfzXJzg0a72
dlaekysavJVVuyD4Ld6R85njlRovAZsAkAmbhdTKTJklwsWX8f9sKn9p2md/6HXBH0kCPj6wyyTF
7kbzEZFsDqYtZQgu+YH819B3aga4FwHgPzHAbVCnnwiaNpXac40O42NvJSyuxy105lTNJ81Q5rfz
EhpgAme4KIin8RXbVvUbGbtHfRZQ5imlBASjNvTIoy3lbvhW7b8azZG9CA8A/WeDH2nPBpoFVv58
EOKpWShgWCOJTVsmvYwI97QujbkHAc+ylUEgIhG0q8Dv+vqqs5tx8dQlEUVIklQ/GUdAIJX7/YVm
NvGIbCESFoi22iPI0o0gshX3OiK93fSfH0mn9ZJBe1l5xI/exe+sUPEhw+JCWJGzCY5fGkE6fgni
NWIo76pnkRO8vL/hnFkMSfvV5NTEDX/OOUB2nIfpj4fPKdlBIJDag+juNsGg3bOatGWqhtYRxHDn
l7iaACwOmQH0I7a5n9zhx/aHnnS6DFur2YErWXosyQF0O4dywxhF6BCOOQvSyga0PRzaP+c4eIT2
FnpNuIPZeO8cJUO+4jZZRMbSx+ou4LyKiFLVwKRNKCM7fm9WYnLYm0mgydBVcW23ZoIxY1NqLeYt
dtuAJve0ePXN/1zRU/FPfivWljfA+1fCCYaBlxzaVN7UHXfUAc/kMHKvRf8xuTc61HBzdfuHsVW4
siVufS6MyoGzGy549dozu5UWdpMaqis73lqhlZHYgEgC1NIxNAz9YSP8F6UvfKCer4GOGZRkIhNq
ADTv6LGTJTZMixvk92e4b59/41nOymJDpAOYFXZX4ZFVClo1mAf1ZujArlAXxBEIEQAcRspq3P9V
dxphzGefa0NY/yIYB95IeR8JI8IMK/po8TC9dENYpXFu4lkAkh0jr5BiK7xQkAYk3i/8VOu6OgQ2
42BrWiCY3ST0KEVifXtbJOOi8r7LTC+5OwSE9ZLMVK0MCuFZsXrNWPoPPPdcimsaAuyzLrhskxjz
yLxaa2eGjki48dvV1mcIT48hCmpMHolAj3tDto4thXEXDL7bxKtPyDHUm+A+IrL1CSQMCI1tWzMy
eWX8iXBJaRYsws8io56nWPl/FYHZtuhY51P9tRBRa+emAzmIyVcRVwVyxSScl2jStvBncDBz2evv
j+I8nUNeYx/V8hE/LKBd1mYfvlKjgV/t05vV4I0CQNOi5N0HgMPeyOzA+f5GgVgLnUyMxzS2rZoO
wYE5B9oYYbI7fJ+2BoHvAwPiklCiI2x8ZLXCOXgYsmDjXHjD0tLB+xaWGRfEGw/gK7d5IJoKe48P
hn/FpauDScXJo4EGW70X6Zezjk5rJemsEzI1The+kNFtS8VP+STdgvHR/lvo8Nur0gAs5L5Ad+i5
rEo6vRUDbthteekg3n9i1sLeNwxybTVh355cHQ/oLFiUt92nhOZdNbzd9+T5q5SdpgGqUGij+NvJ
Me0hy3wkvlF+0qQZ4nA1in2Foi7EPNhDx6l/uVFjspYniCyvkKU0i3JyINW9fbk/g7xUomrbcS+K
r8oxKtC1bGE7e8AVRR6gwo6l+zdCOH6hLeS+QPYgedzHo1wXKb51nowTXyazLTu849djZb2tPPyV
ZWuPtlJS5v6JTWEtIx9R5YqDWSeuXj4pCu1Djqzm/weD+g1OlQB0ncEFwPOLAuWEXqv1hRlhvIcw
Dy8GctfLGrIxND9VzCEL6H4tQB0wciPYs7OtFB+3odiGmroJaSxAE4l7HU6hUKO6y0DcJ94WGnRT
kVCHdEgZpbGdZKVp3HbJSp4yEDkyr0Lbg3wTj8Bh4iUPJvM9mxjq4fXLHm07r9J8oRyWWFrE0wsf
PSphIIE7adFSPxzsO00Otd3xJunLH+vevejYTt/zklB5F2ZjpuNa3TWD5RxENEjlCATUTV8+rQSr
KQxd8sMkw5xb20jKpaXD6M12MDutnvDmhms+P5h0e4w7f/Ht0ZMdtxj1Yjo7dz1FAgjdy8tE2KXL
wZmWuknaoEnGKyQkbgkHOK1va9/+WK5Tw1sIJwAPVdrCbLwrpYGaBO8X7UlRSAS1HliL/s+tYyfP
LthwRfIwKx3lKGb3w3BT1qVGh5cPXroDoXySSYua7CBCDzyC7+R9hSVSi6Oqe1kX4qGIV6aAhUQj
l/Ndi/2A5uFX8PONoPq6y0qCmQZfBPWb/JHXcd/9jL8CrZbLbNYzPS2q+m8HMyzubCzHGtOv+qRg
mtJXm2JblypI1IGX/nXfWxvcYSkz3QPuqxYIyh2USDU7TcbMXH1cl1xeaQbMVhWQKLhU9I0Ur54p
CT3Sk6ZOppr1d/DDi39C0bmNwiuwANkVmWbFe0gBy9PIHOOYpy5TNqcdtSP2BH9H4kje0rx2z7c6
ZsrbdeT1Rr/8CRyVIYQZGvMYLQ10hjdxNPbCrUdQUpNJBG20I2QQjScb3OTYQfyKm4t7oiPB/hEU
tihBGXkyh9EJLZY+UeKlPFD/pcfZWnfHr2SsYqUXVxcE1WxMBlVl6Sfl/rQFxGVwUa4w5kLQAm2R
DC7xJ7HA79uZa2vQ4TKIc2bA+HYXlN9S91nOStEGV1JYSqjhrstQj488tfkc/ZkLIV2kqTz7SopU
LrtlHamdYCM94GVpkCu8EfuQg8+BFIEhMCejbdBJugBJg6jCTAB5052OFlAVy/8nvEQ0UGgAg1cO
dsRu4ioywFwYuPWxIti4xsfgxsdkuUIAiaYVtb/+qclHzT45V+kYkFY1KABQ+D6pS3HVt3itW4fe
XOqPfyb57g0bsNQVOye/PsQz3B+hwryw9EcX8umBY9VhXdDE/xCxmf8oGwBgEYEMKUnOX4FFsVrq
55REMlHtAcaer+OE6yQgaaqZtFva9N+DPtI1nm8jk1/1DrnvwkBR+b4zN8IEzqaVQSAg0MVttTpN
F1ntAF6nUCRp7DH4oEYGAVUQQq+Rg5EiZmbspIkPwyukSGDsIwLAX/sxqmHzNerED4K7dOHLZ34y
mlyI+QORsfeywIHIUsiX5gBsixlOSa7eyq+sedmi3IUQRV2iTv6vILN4PMX4Nn1/QNlOOAOStOVj
YLWZxQhH1nCuxtRtCmYvHIoS9sAWqnFfeOiAjg3TpdD3LKqkJ5GLxFVyr8PpUZrcsAwc2gpdFdoB
WKVFzFRu1xJvrH7+oLUGoevorH+pr02Jq2O7aQMpcXkqN7wpu5pCb6UQdrI6IB1YU3nl5EoTPGkQ
iRhDEtZ/2dFGX9z6TtPOIMJbbPqGuJe/ScwDSGqzep+IUb6bNnxAXm/PF9eOQVTAElWoUNYjelFt
RV304zhHf7mzo0/t5CZQkbhjtG8kuBDy0GdoAlu7hVgHkF6e4cQLzeJpVGV1VJQdN5doyHYC/HWy
IkBu7utTp319NrKj77fYfXpr8CIND5Rwn7k9SGHYGLN5w1IlTLYbG5OdO+uc95tDPAhh13fkKOe3
5UJwjIIuKKmHTPXf5wlfpDYHFglW02O63616SYorht3hymfemyBGpi2a5SoSfTCmC1RATRD1VWkx
qkJfeyssfJGbXh7JAA80yWD+ZllWikNaOnoz5+dysaURO2ukzP/AbqurpRedyT6ZvKMEmFtD2eqR
qr8NCZVUJ1ZoHHuleAduE5iPB47skqY/iujb1ohI1nYYvnY2HOUJCGgs1m432WSYah+tvEO3PsNA
LxyJsDLPdSYQpKH4i2T9GOe6BUc0K5TtvM9J9OFQwe6Fm7jWWpUfkYEGOXbgsb95rLX9Ag4rL7Po
VIbLxhT0tdCtIfQaBWtm8oOdaCKpEPsnylUI9mkIHzH4jutH6UXdvucAbO5Dgp4N/xCjHRtlQx5E
mbkjItOhDrE3x//OI0YxU5igYG8iLSuh1vToE7SKbqDIeSa/YrY/HuCM5SWwT6LiZ4mDxmy/oU04
Pq6eMu1eO7bwPgV6uym4iZVKnm+fN6oHvXEFs+nFxIQ+oemKyVfAmYjzhxoXnh9qV2HoBn9nGmd8
nR+QqfHX1dE1LbRLgiXIN/HEfiIsTxjg+CK2UHHmiOjoFXk1g8J/2U16HzmXnVmEqwA8A0qSxHtK
Yt3ciXxW7AhyqPO4WgSOasbbjJAol1ynn8q6PnMtWvR97amuVV1vyOWMYZZ3KzKbVXrD/moaGEua
/JfAoa4JCgpRR/960a8Zd9AiHUqSQUenfq2jlCFwBgAQYj2YscQ+I1qwK6ufa85IfG54VGhx7Zbq
zrIOHu+OHeIxdXWI0F7BO0NpIpw4lp9zSl0X6IyJy/rVTfI+GHCQPMH5B9dRQ7GlkHUpxpzTrOKm
ZQptWV5Suu6RsxveSQPHZBrQcf9hvMXkjfeC0cNUBm+98s+fubFeAEnvpXz/1e1qcayA21lKi125
7gPvEADEhE3SIeaMN0igK74tLvtKlbPvz7cZBohq/TEPgI6qysdQMpdxH6mMk1hTmrb917Z+iZb8
ifBbv03cMWEK3z6o+6+tSVCcluydw7tzC9sSKBu/MdjXidupALzEsQd5LET1xY05CGOQNy3GMEGD
aytt5USjAQtZ7T05TMayDqul7nutYjl8o3w/oEExPKPgqpdoTGvSY1IEGg4BF2JmqtReKnK/tI8j
RdSgUUni1IkeWhteVsQQBxW/HXLJgnDNFs7j/0PxGKx6zsnE4pptdx1MQUbp8CWGJq9IjSqOJyvT
VMuP9uRDo3/lJU2/3QCIuKeJvl+3kK1NY+vaqZh6gSVl/XRJgf38v5ZHf+J2ca/E3hLXUh8mDN/5
TTs7Kqe5Ye/wJ62B59B9eeWrE0DAl7ATnwsVKZaJnwUWefifhbyviDu4raTiR55udRoo46aLz2gg
/XZq5gGLEdRGaX0xfsH/mePcE9cwVKf+wlYQJZtkvH4Km6FWtYajlVtkvwtN0VpuPQwwrZQ9/wXB
VibQxAHMUN4GCfaxIR186K60vohKzu8Pg/qXSv3FoAANe9Pbveed3cx4IAlcBRlEwngk93n6qEtY
YC7Pt6CD+cEW6mYdxjySH4ucGRWYH4B1VvFiqT+PDFVYEfmCwiWQRq/KoxjNxrLcYAgdzzfBnQ2W
WLbis3RKMsz8v1XHb3c6k33pE9wDr2Jh4/hensiVEuN0gnIr522CDOGEK3aWKF3Nazz3JCvKfRKN
hETwgmk78Dt7rE/XStlHczFidRgdPQr7qjTciAc7OHLK14OdjFsIHvhWU9w4TCTn8KrR2N0Pvh3e
NpUxPSSjkz0ARvkgXkl66nN9FqwgNZuCyf3vulVq9SYG3P509mEZOZLag2oeEZyYuWJ6p+Cknatg
OpI++lLFMvNSanac3FSrikJKQD8CSnZf16klGjK8ivrEN+pnFJHCPre8Cd9W20VwjEzjLvD9nBjS
N226aV2mxqeXG2NMGtu/yVuDa32mAZ2M4/6l2cZUZcSzr1Umx0QaGW21/Hya8NeSmaBIzX3R5wWA
TgBOLJ83xYpwm5TiZBj2e6uOWNc2nl+7TVqetxVstx/5ZrbWNuvDZnmy81nkVcY811/FQ4yf+4p6
NHuNgSNXK8EGA2SmuzbHyWk2j/JWX/7lRuoOuqpJ8qHj5lHOEku9cDyRiTXCZhUBLWKG63XgHSxm
rFhX3TA5QMRlfq2opa/RWIZNqrpncRVz0Vv/ZDkm78L0C8L47k1uXHI4Qx1UXEsFmmtHPFgDJsn8
MzadlR62FLbEtxADbafDuDPB1O7ZlqHU11uuekAvg2ssXgYpPQguD6EiHQdWyYHMlDXM6zJ+//+W
v4sWd+AiROIW5afa+Ben7ldG+fE1NKTs7pGgZdwIOaNnIxo5VWmC2HBmFPL2Bxh3gS624zkZI7Yw
WWO3DhofOH7FnVte9AFBgw5d72cRZFDgoHCRwMTPzsszgXgVk+tBEBYwjgk7Vw0yrjmaz6BA5kUV
L4Sy5i1tTWg6UmdeWwLlCfccBeuPJKrzVTMa3rLJsvXg87t2sDdXLhKEAuE/qMPKOMGiGJmXHS0+
837ZAhSmEqhQpDJjy1l5yAIzLm9rpcZCQdPm6MdOi0Ve3Tv8PGAtOwBKX7UNsobQvXExKlldVF3B
BRizqFgktPh2Z5ErrZOGo89a8Gz5oIj6Eqnq9ie6TvP0169glioUgus08poHNiZSRBsL2IEf1ejV
nd9KHSCJkEjl6Qnw4Z+L2u0NLgRK9fGq3kpRHdzvXy5LFW89CmaToVG32ZrWYQzT6WJ70pyjpvfg
/jMGd9HWk4sa3z2XIokypri4z3ZdDkfbInJ/dT+OI1yHnNyQbrZeQFvE+UzAXGJz5RLMH694OUEP
5PY16dn+rhfpJ8g1X+iycVabHf9rUg1Vcdz0mnCL6hIAxuIUijoNi4FepmrY7MhjdlFid/9oZZM9
QjeyPF+7wMjnVC2mWMO7Ks8cWnaOKJfEX/hjltyaoXG62LK5yYK0Sxgr5IKYeSROhyo6ayEh0zSe
6cERb95BHuK2dFdRLrW13YoqU/cSRFI6RKC2Jx0EuQ84111djuplLNb2aOFLUXo/gIK4orIhWssb
RIk62kum8sHSZe6E1mhm4tkTz+SvBtT8K/b2JrYKchXJHUvx3rHWu0DqFdJCMSlLto36cS/CcG+5
BGznZO3o+3VDX6vf+W8LCM5FwI8qGbYXm3Iur1nPaYNmcfKPkSPzY3DmbLVVASg58GsM9R7RZkS+
+ZMpJnRwpVA0iRICZ7AW8rK/WHeCAYqXN2vS4g8mnGgfO77JBIiRRoupG8dzY9GbNrrusEJCawvp
gMjZxAXldT+pqftAn0VHGtqn+4vfO9bbjjZMjkQEVoUzK+mUOHGHrDvoeRI/jw+6DvEibpxmcdDj
IPlRLCnNgjYvmA+xcQwBsGR1p6upQOxtq7VR0aLOw+IiLRhdZXE+lhw1ataYNjO1JUL1H2+Abvo8
qiC0A/PWaeBOZT4SNNTEYRyqNZXCjNp4NNqyyue3tMeNDqlXd84HQjrdRL9QNuT9KIiS887e7Ieo
s+/EJULFi75eifrbVlIeDicrN1bDXL3xxtZSIwD57zeq7CalPWi1MSpvmy+EcOrc4HV460vMEa+T
KULJf6905+Cq79rX9qyN3+ADhaqe2fcwcIu8AtWguhPCizOmZo+dVRFxDn/umIkQEIub0qB3XMr8
WqVQ+UTHGLtC/iphNn5e7DX5y/j386cTuZ/+NyUmaWg8OrsGJ5gVkadKnpK86TxI3FJjHIWaC2ih
DhtMjIVm822A8XbuZJBxNR362Z6q3BsMZCLRnKtukalDrpyG1VoDHuuaiDEn2VVHjak6TTJ9O6mX
sZcRjNU3Y0k9Roe/qMFjdsZzB+bxcf4xNePxxIydUMuhCYUhCgcLS2lUeTJmAgWblV8EAhKN9xRK
78s80jAwqLg9LI9xycLXBpQf880wn64Z/7hBnxsi0OG4hIoGYeHEBB1g8+YPTgpxnKjXd7dJL+t1
Ir5dHmjm2c2y4U5e5cE9+tImdYPRJBTiQx4Hk33cEJWOi69HBMJOugPyc7enRKDrmSfED0Wd5kAJ
h9qY/IZ2bthBzs5mdf44MXH4D7jyaghynMRxkhPgHauGeDaFhjruA5vaX64hGI63e/2kqkGPKq63
tZ1IwUjoxfXg4W8/KvGhJcYKrcgqcueFnE26Ph4hyrGXlhb/TpKMPJJQdcRfi48cisM5DyZM1OII
lAV7KfuD8dVXKuothwoPdm+Y/DztBSNJIVggW2TtGTBlJn9AzqxoZwbI4D74RtrezUVqNIGStEOx
Brc7ebhQJWjjTQffE0l4r82MirJeIOHL8usRkXSa/b8TZfg30r5KrhJ15x7ou9gap51BA1r5LUt5
zjMOfG7iJN2Fkw60rAhOZ3zB/KlP5Mv6Mv+wSHWqp5e3M/abobebxAeWewuKESrg9iabnzUcfmJZ
QwYu3AHl74co7AmYpZPJeXgcKombFkvf6IV/eLcAIp9p8x2gSDOhcEvb9pXYcr0V2YjgwNtT0Yzm
/4/Srno1i6GzHeocq9xvJVHzc6DR46wPxVjuEOaUetWzOReVITtxG0fOW0BwdfHFgpuNMfw=
`protect end_protected

