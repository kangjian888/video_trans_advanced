

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GWT/RJdN/UcIKTAhVxs3scTnM63xEPkso8NeqXOmx+sudHjUMJ/qSt5GFjdXAqexLlRND8lEfssX
Q8fYY8TuyA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J+phMqmkYiPgvjvEjlpcdWdxzP+34SmYIPyc3dLXEqt+h9EhMcqfQg7r/svpEBV24DU6CyKyCXke
3gZaY85pXANGRT/lW2K8drptf9l9vYajWMSy/HjvETFYNanQN5XDicKd40/UNr4NV+8K3+zJSD2+
6HJJVC0iWa6RgWieT3M=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZrkwjC6jJHChQhf/EDIYzNRopX0ckXH4NL9s7GZmKhZ5Xuu3xV3LqvLjlAq2T+/3AXtko4HEVfJk
jD8rEKHAwLnqMbikHpL2pup+LY4/a45y7duxNC07dpJvYX19IW6mqYLKEJTs330XVwBLE1KOyaGV
xhWwwqThGo1V39JpBwMcpzmL4YnxHaTlERiq7vaoQpYAMkwdoBVpG9MMAn3CbeZJI8pLk/zNkztm
rMeS9pshqNVtzdUse3pl3EDxWMB2hg/4/G9fk9okekAXBV0rv5NMqf0xPrBsTvRJGO21aW42nO++
dC8am+sI7nAhoG4w6z/WxE1BGkRuZGX4CGhIDg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iexpjlh7M7dlTcv5seskQPlqyHreGwsr94b5YKwilWQsfXW7U1V2aK3O1/+pXS09S+pTH0rKoHNi
ofASVdK1RB4/i9AYD0Ihai7zYaqt6eRX7azypmOnO0M/ZZIrM+63BHWcDodlNlh86PWfwaKQSqJW
hLVuOmY14GXZev020lRZWg+2UhI/Cl3c8nww44erkAvCrpxmrhaZg0s2YPKI/KBqZbZHwn0ufJSY
5EPF28uCCS1urKeejeaSBUmimEDyf29zU/xFd0fvevSdWXaFhwjT2mOL7DranIxEzj0yQrN0jiKy
Towa0uazE4xB+gMrElDuwpcw6ZUMyEBsaW08mA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DVPBxTgKjw13z3lZMl+QMKXV/uHfXNCgMoWbgQb15TKXtTCmkLiaCYkk+UNjnupib1FZuwkbZs4q
pFuDW3Z3x3poQoD+4+Z7IIYAmkcV2VNFgSXWGO5qpHWhRfkulPfZcRStTLiN9EUcwXJUsLi1Rwk0
oFaVSUr3p4Mr6zjC18beDCFomH1w+aZiTDmIDtnqdWVtxtresAhXiT6k51hdPESOpe/yPCGrgQj7
cckAkNk0Y7ums+FtMhs5xsfKLV6GQGr8vql+qoCmnMNbYofWKIq3pY2FrW6f7ZGbFhW+vgaVatOo
wR1vGhSucCD4x9efRbKZpd3HOhDW/vOAo1pd2Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uIb1xi/b1sGS9N5+ge4ctTMaXcuHePw5wBb1FVa9aecf3hzk8F8+/rWvK4DX9IjVKEx0PLXI6xjb
IH/rGtJXdtbDJdBaXxCtQZnZ3bb8a74BAJHYm3BEextG398AX1ZCOiiun/unyz5EkREGrSg9f1qp
tvP1wCaUgYbP8iAi+ak=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qK9lK7oKxV9h/658uwPcMAAwYeLmnKNpsdduH0hJUA8HIiT0JfF3YHf9Z/+4sugCSI1ARr9LlbO/
o+J2NPNqOXlyDgJW0FGjeX+G4wdX5LlxdfSIcRGs2vzyXQiAWVbMq15jqJGV+qheK6QIsLI/qwOR
naZ46kfkwSE8kQXhF7WZE2kD7kLSTF5QPnmYFPP1wrSHpjD9hfcjmg2768Oxg74FqPuAHl6cX4Bj
Enf4+hzQMQ+IcGssYzesFwyeHIqJFbufwMH9hDnmz2bOveVtLUI33QRmIvvIjsEuvmQwCu/AC3gG
UyfxcM7HSiPQe9MbxhcS0KjoubQbTx7z04URRQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 504864)
`protect data_block
ucYHgKzDjK2O5O9Ac/5eyYmnV2yUMHShDyJODcs7KirDfNyvbXRFlkQs3vPmd/QSuolCmzWJNgli
d62oEJ7JpxRmewvGMNahunUdAkmNNY1riHQpmHpSeVDEHz3yg+GSPQj/TTwdXYuita7XME/GCXB+
w9tAbX4nAsxXaNV3K2vgY8yRmHExdeQZOECmgDtqDor6nxBdPa/MY8C3206YkiCV4ithzrtnO6XB
+Qf9e3AKQtiOtzrmtIJRE8Awo1kowmlc2AgdzA9dW1DhMYZL4rQpHez9kNatoX04qVqmRNK4idrT
awSLKDtx7TLFYgPBzcBu4MiobcKT58OWkXdvbBrAZPS2YOdevi/2vzOFFopQOi+laECufcyD4Pu9
qg9GwK+ocInk/5GnRLREzjcHJPG6Q8f1944HP0GtzmW0Mwt5cAVjc9qBW0/vOYnr3J+R7YLpUALZ
yCf6MBlGs6WtdbFE2FnH50UidSXX4gC3LRhD5K2+DLjdvGiut8hhRmug6Qgm8LShHK2X1gYddHNN
wtTySBqnjlpN5efkB/Rf14HesuK0Xm4N+vaLawXctKl9b27UJLzetrzYZK4SK/NhpEv9Dzo0tsjW
RadlK0t9Tmen3C8biyeKUqgxpTVYCmNsGCjAa7e0xWqIDxQTAFQVnQzZ4L4rZoX03owQ6n/C9XQR
phvuQ5uKOv35+Xci/dC4dIXktFFuLv+WDFDrq1SE+GDPprQP8TeRt49nf8dS3i6PUl4htITwjWoE
gHHffBtRP46IsGunOXM9xPl289Cer7MOdyVCdjp8JNyZni7EZWJCwe2N1wLgQuyM1o/EsdAL1lXP
0jB7Ltb/Vut6UiDOIsle1q0XGp/i0UIXpwC1u/TFQQ4kTudDXKVeZmpi2j7lTMPqklQP0XIT0OvB
ofN6AT/WIbwGHbBG61SrFEJhKg/wCUvj1fxLqQtlfnOEpfrhjo3VSnuwjYulGLygT16QQoxUA42D
WKKdwyp5v0I+tZ2xvdb8tq7YF9r7j3bjIfgt3qvwdwlD/ZSmtSep71MI+IKBbEIz1tdvsOPq027Y
7rV0YWBs85tLVGphkLridftHmjz9szhg44/o7ZCCB2Z3GK29Ea375wxB/6tU9FhWRg9XeIFRnWSd
ck+PA4qASfC8IpDQwcmunN4eZCR46YWdeSuUQ033CK/F67IaXJOb0MOCtaZb0jBJa47VM8m60ryv
E6TeR/bKjs6lXgMyMpm293FgNzAPTkKI/4cMJhq9fNtobdZ2W1OOOQ0v/oq03SVNnY9zu+bp4GjK
wjp2ht84HlzBdj2hRVJdeVCOTvvVdbuMydi2+9KW2l8gb6Auyo+gNdc8OhE7hpd7pnhfKxlqaE6M
SnK9B/CR5fkL/cwr0XABRyKv846WP8CFEaz/MG8BeXI6TqCG/+AHwoU4F5ziycavQQN7v+vFeMvL
l0uqQkcGsKnCTPtFu/khDA0JiglKI3ZyMZVoi+p/dMwdyEiu3HtbQbxdLZnnM2YuP8PBV3Ncstmm
FafkKKcIpV+wN0x+ZrXLzOYJL6TWGVvTdOi+CzRFr/T2GsPPNYWrOFkhdsZHIpOoSxXXiwNLdycC
12R8hNAvTPnreQDGx/3jlZMvU/XGAqsUwedP/l45OFQqRxgtse/8RvLjm8kceLhFcwkAHFqpRNm/
K2wX9Nhb9yjucCP7zNPKVCYZG23yoJorWAMs4H1n0exD+272If7Fx7s9kM0Mij4jgDrd+XMTMKCx
a6OxIu63wsQADizBCTDfc7ggbHpnRNvdG87bMPObZhZmAybndavM647FVqfpDOGHvVa3p7xy45IP
E//e6r4rHCcpCBJo+IR7D8wWP2wkwiTrx8q8Ag6W6ZvAPDX0ZWAaexQ+3Yn2DVJU7PiNVX7hlTFT
s0rwzsrWp6vypRvE5LNoUQOvrFNy6wboYenLhfDtmaF60KvdgB2O1zrS9E3N1+gmEvVhDiYGHjkU
rsrCIqDMYlyBmco9UwAuYGBmbfqgFopt0bpBNMRRSI3Z/5ctJanQO6JfZnSUbRTdhIja2HaqloxN
fKOQOiX9VS0CXNaQ107ZMx5EW6UOx8ClyvHe1hd1ElTInILuf3EKniK5XdmOwU4dzR1h1ahb4zyV
47ysI3pAOwq2sCrkpPdvpA0q9GNTziCl5jVP/wUn2x+oUbk2sgRhAi2OFo19pMDL08mggObwHWds
Pj1WW1lOWBKqNJKnNllb+DCi1uwIxVjROJ1yk0YDmnPq/IABabv/V3z9ja0g9mbH3t7ZMKJJO1z/
dC0M0qOViYyvGOd1y7aaqKSX3ZAptYwCoYTT9+ymSzCDR/txXqxoF/dY6v94Vj4oaOFinoliGWIk
bSeimEzidaIIsEooVEU5C4p6nsOA7NTh9HVu/POZS5v+qEUWtQGEFJmaWFVBhuKEpYFcMavTS+Aq
+AwYZjOW/y9VUIl1G/ZFW8a5a2AhNDO2zpImsY5cy3zN1yTy/WZhfBZA+Y7NW9BOU9j4O/BZZlxL
bTVSEG2+OOiQnIAwqAV8JulNXB+WYv+WEQfVx2lV+h0OWvhP1+UXJrmCIneb8cjjz1dgMDgmfGrK
0UNzWlxSmx7i4OfFwn7RAuMCV3fBQh49EENhod4aLfRnpOaLakl6RV+VLilaRagpmVCA25ut7OyS
XRIOnxs9oNXZDsoOGFnSRbkKJ3e96becX/njQyfFXtLRuVqMJb4L/I8DNwZvXFpM80mtuqan4CiO
Pg8Dq5Ya6HpLPtmTrOymJgFA+HDcdmJX0HJyib2FCbrlmq0enCNv+hRies1FWr9eSN60AbGUVclc
CWmVOBdfNPDOVpArGogdn0o+1HqnxTFbn1jNOWszcG+PaIrr4DTbKAChtf70H6vwEgD9GK3mHbWQ
QObOxI/AUKvdyqdVnJWFucNHIHP3Q7Ujwl8WMm5EB98suUt64Qbkx2E0ZEHO5XWUtBaBm6e8eg0B
Ss6lmiiLJuYxe2oYudZ1mKAdtKhs8B6ZwO0O6WnEpSmhrPDrGrX8LiQSjamb6ILOgVEiSXF/XYsH
/sJr61A33x63IdN4dpZlqg/VDMhcsbVzDaWQae4UrFiYaGiix0VhdP5GDyBiDVQq7gJiLww7kRO3
+5IscFKKLGCNHOY8GjmnlyVwgJ8IBzErUQjtBkd69FdwYaySLEyUEEe+PKjM7RtuWx+PC6ZWnJML
ifKnGl8mwiUbJ/mpD3W5Qkp0R6qnap3aY9LLh+IDwqqavpyBV155O2P9o625vCb9BCCPk/a8ya+Y
s5MenmZVl8w4oDqSZo+6VUl8wCXHpMFPrzvNRqm8DXrwmszng5HVrutwXfC63RcuEOy1hF9SLkPc
9eKgAbevO1cxWo5y20edzqBznpLwlK72VI+H++sblirkmMeM/X06SoaqoKagb4jllhBS7cCn1tdP
hINrKJb/cDjoNawPrAFXCJxErM3jQavEF7+ilJ2RSDXlxSx2yeuB/yH/ALkR+7gnE/dLcCiCizyf
A7T3S/T/xhVHs3ELXNlkvOm9EZG8rob0+iazARI1OL6FHDzy0b2DX/NWTQ593OASx9cW5IdKwn/K
LqfFvP7G2JkyhLuDggjj6JAYE/wLB/W2V49QqtXGxVpriJ7C/dUkGCnZvanLpzLiwVp9X0kf87BZ
QJk1JbiJwEEYLy+ye4LF4AJvTPABgpEmVRg1w/7YPShOxS7v2YZgxDEjKzWiQbyj91TqV8BZvFfs
UoAEQuulKw71Fu7O9pMAzlnp+QnQeuTvz5p6r4mxlwJciA4bLQAsrecdhzLc0R/yhaY7kodOsoOE
YeKjvUFaeNP23wCLw74X0yINy0Rk2tovb9UdxSzr/5iZfJCc3EKqQSU9vbQj1ukONgd0YrNIiJ7L
UwBgL+RLfpbmxL/a5w8pc++RqItJVfg4i3ky5M8NJ/npXvIr44F/+gcI98BUzfuvK8/W+cLRCox8
SBpsJA1Sr07k87DVuaasV+VXmlQEm+NJzAxUw7vC8hQtoeYpuxcNJZFKVnzaghsiusxSq9F7eWP+
rCgIS+T6LO6LNBnsdht1Cv96eLXv/jJ96KiQyKHz1BkbJ4AK65Gp/GKnIa0OVncZd26LSsOfx1sB
BaPG4I+ZcyHBmTJpp1MJY617aBZEoVtPBu5iw0ur/oUu/3PsoSdI3o49HY0FcqEN/6w4ZaZvW+lc
32SwcK4spyeC2ie98TaOJ8KGkZmvgKPYuczvoF6vFUgXClniLZugPHiDaZcpV2hiuqykPNy+uio/
/3raQURlRubHzBqjTu4N/rPdP1raq6HZ6pftGbFhSsmh3NElXnr+Ew51faP54GEwaOFJ6R5R/rRq
1CF5UJ+G9AUHaFkWfPgCeO8xZ2YH0UTawyOhG/F50cfZc6Y4G9y3zGHfZySSjmbQiRuXAAq60VT5
u6odA6y1AxkQ/rri3YvnsH7qdfCUkzu3FDZNgjuBOJZpEN/uQ5oIFhwiJSZk3znl1wfJg+VndDLf
Afo9ykJzCj3DTgwRTaBwSS3sWZEJwbNRjDkFfPYwlzC1+mJHGKO4L3SNUKsxOyc9MrFQTtxgdmQ7
PMyfddR0BfJkVU3cxi3RowC53lrSqAe/pP3D/YcoqCe30rKaajwrMk5IiPmPLXCKCWg6HjVt/fg5
dHXBj1tBCemRoQ/MqXsMPKQ7GxldTbiyuAmKDR4cekXwN3tCV2ohI4YkYs1GKOHcwHVauO3wpOtv
5lVjMMXH6/QpR0W7covj7xpCNxYk18DHvQdZKmFp6xiKGi0nORvF3wq6SRxwGbcLcB/KotTFgBiQ
u1g2Lgpr2+gvpCS1IVKEDlpIYNne4WYisX0pSkQUiGYDqvMlM0vtKA3lnBammTDFEjhz5NUw1N2a
gCBRdiK9EX+2hMlO7jRAAvQB9urvpZ2di7gqTrccnN0MoGhnWU3wSrcj85WsHAnuoTDX+zg6krN6
HhJDAJnrXG/HnWYqUjuZFtZglHgFYXppZIMjzkkinZboH18CHlOhkRfBWurjT5l+i7xHl1vZXn0r
1gM7NePnlT3oaej/rYVvOE3Dr2w2h88da1YSUWdkWvv2c7Ytr+Ooiiuvv/tK3c3/vo7aDjPlNpEd
DZnQgP8yXATeW+NlibBBU9f8b9Wn5ymxSlxVoKbk6Kxj3d0s40Kd8ouXwbBhDriJOkgmyUgY0y3a
fl8QnDYSAu4nFS9fvFCu3fImAZmDjaW4W7Y6uxQGWi9J2ZLLicU/uGD4U0VIvvJ/yK9Brh20MkB9
GcbGVLUMCeWAR6v5sXBDlyTrdwFETwtxOXeZ32SyDltPZMF5XtX6x8BLH5Jgp5WMeDmfnI+mDyD6
QsU4k2AN1NUMTAX/wZF8PuiUocOLaq4UPpU2QGMeXRSkC6qcou0oq8Zil+fHbrwgrcEflR69DnwE
OsRJIIHEk2S8APzjHaC8nuCg/smc3/alx/C1ll/XS9u5Y2UNnciD9B7zWRAq5QZMfzMa1iiNxhCC
fHOljIVxYBIVQVSPSl7C2zEw8dLA9718kFrVA7PWryJDL/6yeAgUnmTmthOw++oxVcgb2k7bfKc+
FwA0cKcOeMtRO/tWz0mxBS1Bfe8B0vGnGGxxEFUKkOnqzIFedML9NNMDss7W4wnaPNLhMaOxIkFO
xTAhLQGxIOQyqhWMDpmUzn6Du6yskJlz8FnuKg7l3/LFk8VDJEecDTUqZ5FOp1/s2OB9NQwRkCjR
9Yv2sd1LCXu1sVf+7zzMYPRh/o0LVSj8Aw/Vn7XLbTkdKdZGDo69g+XjDD/Zl+Ov5lttzLs6knxN
HOWhsrV1Vw5piT8b90SN/0glhcWltuMXwQ5YNymcTclgu6h5jUMmEJfQqaJGlbom30BHnSNaxStJ
tk+OwwrL55d8/q69I2xnAO/H3Tr+qiUFa30YoKx3O60FFkDYzAAVDjUBEcS+VxBuojcqJ0T1XMea
QqzdaBZQ/Nf5f6t2upjmyrFlHf9fvkeRNj6LONQf7YHoSqQFHYANR2/h31AGCPDio7AipC6FSMAN
jCWqob3vZjck5bkvX/ey4nNO/IYflGmVhJ3+3DuaRdw4elFc7HMWkFTBPNXe7hAcVwq4xV3JtLZi
rAob9PhQSUybJHbrWC19Olt39C08BeyT78Sg16kBpGt+lFb41l8OmPf3BkDuwB8lx4O4Px8HrZh6
r36Utc4HxC3+hVllcuTq5KsZnIjNKEFPkhVFVlhqN2dE2ndFNd/Ze9usm3k63tWCE+NQhZn/iYys
zcl65VBGWGkY6pvg9tN1YXRlaCm2eCWXku6htaZCv9DSB9DTncd2sZEqU6cO84w7wB5K/opXs6BP
MN5Wrn6igngQ6vR7HntDsi9aFcvfX+/JpnPZJULLH354DXB2jpxwoiT4t/IU8z0Yp5BV2R4jatQI
tvMNK2mbQ0LlFQ9G5HTmFbJ0KZ+NjlSf0xeyD/RIOsOzfUykFSpx/VqGZQ3SvX90z0drxDzEsXIT
zUwGyR/2k89aYS8G7Erw2N2J2UdXC6eTWW66NigJ7AH80UgEvQ34k/HAEQmFLr0LNgGQaWuJYK0y
oI3Ei4SCisq4TutekaloT113c+my61Q4xD5oB2da5HopUQ8RGOJZDb6F0n3C+yvJjg8yUnFreMTg
3ZM4Dbb9TuBV0KLcox/RAvC66AC8KVBt98LmO4/hd2RWU7d/ZA2SO5NSwEYJ1DY5ek9SN3FCEhL0
AdtJmYCiHsdjWNVNocoGElpW49u7XYhAdkJzWsZs6l+a8FaX6uLOKhmRZE/i1kJRY1JjTCAyFSfo
AyiviSZqk9maUVFWfg5qQV3n0s9chbSkRe5Gzhw8zBE6+9L6Q7jJ38JFYNhbgNtaUnxHkyXwU3Zn
AU8JgUdSnDUzRerRWmmBeIcxGVTjbl9pro2+MR0Z/XbkaVu2bHRI9locXzmbzKeAxQ8YrOn67ltZ
U8AVGJaIj/7dnxNuJISaIJ3gI95AiLRt5/u46x80+N3kvP6xECLcu/sU0D55gw5PXUNJ9uORJofA
krKJpsSPn2grE6Oa0myukZBHC29O9UzOasH4Nk2lSTd4I6WWkA3KH/pWKB6FD/RVD1OqwPGgY5VC
r66oI99CDHO4aEXdsFrw0+XTumMm+VHdAfNUi4JRsdkq+c3cScQsz6xM/bV1d7FM7B0xxEFM33TQ
ccN1KhFxlhZChZMYF8sc5QF2lNyB3/l6M5D6oub0wU/dCGn2ZPblAIytBwn9cA8OL35YXbVFCJq8
Ow/hS62emzENH0Q0GM0vY3NYZzDVwlMtwuALACWpEvWVw+h1eNgJc2wV7krM7uQcRaT+fPJNK9D1
MnKPl+jeDOjVoN4jsrkDa3Arjgv44mIDF2dn9invgRLP47bIiRmU3IutekwUMGPmHsSzeYyR5fTM
DkjHf6zZEiDrez6vqlWvWtXus2TZSlsLR8rolpOHJfOVkJ3nSqxVoR7cbQgiBCpdk/OF3se3OjLV
VUXtTuevLINrg5aSPNV5tKpYMn1aFIOprA9KxOvhwTNYYq6vNd27LZzTbP/Bv1CFyL+/TsEIImVK
G6A9cO2H0ILCBg4E6fOhUOxaylV4TC7PvYpCyWQYfilNDMkFfyXo3TOsQuGwIfsyyu5WtLPsguEA
ebplgU3j4lokkwzqlgzRLuu9yJZmDMnueEV7CRo/UdhmBHAGBrAcIq9jefunpLx9Xiu7Hb7PTsOt
nNkrKUyPLwbWr002gdkGIJaK9M4fXXCvYENTkTCCC+C3d3F/1iqpxA+Xh1twaKb7Gw2K8UMBSnFA
D4muBWjw9pIo5tbK9MM37rdFXH5hJLL12hpC17P3pU0Sx3+g5HL/rlriO/Blhg6TvLfV+XwnzBda
jPB7/liPgcVMNROSZkV0ylLHQgZWAuAaVv1rbCJDPdy4TzU9OZ+9DKdTapH9V5xSR75X07TC29Og
JTz+XxPXxZbiRic1p6Ko7oqBG7bIRYK8KpUx3soClvIscpDKSYCauGWpoDduEJD0EE1/y0+XwqD1
lXxaxu09OdhBxMYtnmIkXAiYWQxsuhVLsG0lPeB0MA6GYAhGaJrNgyUV0WDo33ybbAGhek847Ixh
isgdBONY908Ux6Hldmgt/3AaqmO+Vdyb++ZM9+Ypa1kxvC0pBL7U0yJM1TPaRA/tJ1r3alG3e6tQ
++MHGq2fuMHtgO+umgBekWWeFx8KkVgHQDibFxyiiKS4V+l83LepVyLuwD7/bGdwIdmHAIGt3Ptf
V+QaHXSpYN7lwHq2eV1lStSS7fCVoYU+UtvOatZi9dxHX3B5/bcBVs0rrUAn6utEDXa9XKeDNr7o
rQ1JHHISO+BaE9gxwffssH+I6D8ju7ITkYMnmnII6g/pPjVOnrdvKSgKnxHTCoM+SEisd736ISgz
wDdT9qLzOgtg/VFv/slJ1hLCTThRh8HrNsJRp5g9IBCLQTQBdSkrt3YsDhdr2xGUuI0cdzcDZJmH
1H20qLN+xNWthyYamOGs4W/PxSYN/nyWMMc6O8SEvjcfLpMlnCtBmm7JEa1snWCP6jNa7jYfMoi3
xFr1v49zA0g4xkmUzRq6wFfemft7Yz77/5d5Wxjydc99hOLHmRV5TJ3kBX+c28UeXvBg9aIZdBRk
BeUtCYe/3b2zSemXHPnxgLbBfNHcHLrHwL0g924XDCn9pcBnPhPCcO/zW9y8H5E5NEHJc/p/dwR+
y5soIoasngA86+PdwlE0lTI0ppqh1ta8K5WakTqcRdeSxJKIKOPN3QWeg6/rZAe8ne7/SerohplH
ZfKhFSwRGEqEzGJZZmoiRqSelc4IhU++3lR3N0kx3KMkRbgOkvUbf9vFvOBc/8NfmQS0yHobhI2k
0R4TCiUjHd5mAp9g3Vbz84Xy+CMTphmO33NlOn6lpOZnTHEEKw53y2KIIzTgGYBnV4nIZf5vdRcn
7aNKUpBHfjUbJcR9YGa78h4Z91z59qvgtuim8zHIsJVwI4xJp/d27fY+bvX0wLu+Dm4yAKGxs60o
gHy4Nx6wwTIk4XWSEoalgaiQET8YMgRk5V23lWZu3NrHxWn+eu+ENaQxrfw4THzYSXcffNZVzK+T
9dBS9bCMhu8z4sGinHItkRFxtwfwOy5EqlwN2Q6c79wsfdEy8OXLL7Es8w1i85Ll0m9oo6idQZrL
VKg8Bz46XU75QW0msSSpj0wtZPg5ip2vKhXVLAYbgft11ZTCs1Ox7xZSZggXXPDO5QSS68alB844
AbhQYSJ5H3hNC0bpGOvCM6+p9EWjNfg7xgv9+umUZSujQc0HmaVUoxJuf7fRCrx8y9bAaE25muP9
oxpS9tUo4vgwIUmru+UnPnBNKUDr3rZtK8ohoBZmVvOE28t4AcJW5VbDYNZpjMy3bHTvz7xLXtbV
tZu3ax6B2r8fneMF4WrclvW5e8N3yzlKiSfRPR3fAbsyk5o16UYUVPf+uyPMi4JLlfLk+ZAXv+pq
H69Z2g/rrF5I5h7SzxE/WR6yxl5Fj2De9aXPf8ZJBDr6oTjkFYTq+1IwWnBN8g9YnTtt4IpYpSkC
4RBXcAoSOjD2v1akXH5CXWHy9gQEZTZD3toUiI3HnGM7L0zIWUddLgls7o3SYdRUE/dk0ZWAWhGC
RbXZRmvjIc9AsPthi4mCiBLGNNbGwSYWurNtTv3yAY3f8gh+lwnJxpHjRyAspIhpCAMQyEFePuJo
NkDFWh8IZ59wQ0BaVddwKP8BXscC+1eRQluGnA2OcQvJCkScezg8iTHeA96QCwVq29mNDT2hbiIG
QCbMvJIY2Kkqa6IQQ6xWVMmHwqhDMScvCHDIa2uuhrngNMzP1WStbgiJtib9MhEaO59x+3PkesRI
G5udMeaHGx4wh/zL2XzpMUkiVQd/f/y/XyX5z3imAw6d3Xmtd/bCtI463EUPigL7Ju7Ii594OnWt
vrn6OjVM7Ruc3LzX9Rx8ZjinHn4OEaaXVvHtJHHNqL1DgfQt/nvgFB3EV4mDkK6CXmUdxlSbef/V
+38GXxBNbeezbpNDyDscrmsb/9vLG6LGgU0yIEQJYe4+aC1V8Z0pJ4X0oQ5SPEJHMXEbIaXFFCI6
FUdN1SSuYCdshuYFnEYo/KuTj59treZpPz1dms3f9+w8Oud+WhCpRmMrFMAZ6UxJhdNzoUBwqXKs
jWow6SxPDhP5JBiGF894KJOy0GCgv7bspr4ROOllzMJTmDIx7kvJxsXMqawRMF5S4wSyODnNIir9
WL4waRWE+l9SmqjAf11bN0sDo4BAm12rrZUpXu3vY6NIm4Q/FH6Y7DJBUtcZHww0xvKrY/YIFF73
Tx2V4+zn3cwyItK2xO1FBuUTT74Td0b2ZjzOQqzDfzMkUlzx05+RTs6myQfN4NOIwqRoQH2vECu2
FAqcMQk4CVrII3Uy875o2hNZzTvMQZSJWM6obE86nvoJijq0N/AVqNlG25o8x9Zk70bxRKk5Xcnr
oGoeiSH06WJcFHzHIyTrrStUb+xNxFXAQOio5c61mbiykCQxdfM+BOiUEcs0n99BNx4Grpdicmd4
DEQFKez/PY1TMCrmzYRzNhIc8t5uy0P4w8cwEVNzje2ZAYbB5pUtDAvYr6HE2iiUe6F+NWqs+UYi
04p3DicAQBlxJxBtdpv57EPhBtupWk0VpXBne+u3TWfWXcJCbGa726phJwprr1CIQyMX40L5eAka
MwOdNy+2ehQyXS0uuw746NJbr7EmvyDcxN4APRfPghD3LdqZ1mAUhFyYdnNToyWEJFJLqdUeGuzm
R/VvQq2J5hwy6gK+117qYMN9aa02lqKfzhTU8baC2iME855i6yz8Xl1QOLz5+K1kjuLbwbo85Cim
WvQdXx2bNQzpPiuRa5SAhojxslDwP5o0pn9qDBEr4UVLhU8H17a9ySq9Q0yOjbrU0jaB+/FnmhH8
Gt9T/4ABMBX0lI4huD3T+xn0oMo9y2/7n3se0bPwcBxavGq29KOKGkpDmFITC5R66sE+PK4GYvSq
L8aHUrAEBdKIcu0bciengB11VUMCRrairG28lVoGlr/fmiOVZ9hD0MVgqeg18xIJikRrcOpH/giX
cyiYeNnQsIl95sMJ4Ni//Y+gzTNPCX4Zyu+L62PGd0wYcBl8mCtMyf9EiOsC1dNekbfCtXKRWZRe
n6sgxG/N5WaVo9MF//1sR/PDZ+n/M4KRWyQz76CU1SA0NT5ia59JpNsO5mhGJSxupn4hUcXnl6qY
aUmHlFWhquMis1w9isZhy3KKgOGz9IhnAlCa9h188Rmj82Hg8xvKRpKCDezGbPXEEbZtpi0HEQqG
kdm7WG6DzL2NzzZWwI+yD3iB3dBMEe/0JIRySEVB4Wrsch312dEh+5SSAmsYAI4NxEmFcM2k5OA1
VbffbDhPngjzgfECkxw66TqLpZFxkhUhZklJnsRj+VAaKBrZ9yqCv37d/oxI1bpIexCD93s1Hn0w
S4PWIHeu/qO4Vt7mocTpPizaxGNuy8YeZPPUDmqXbREoej4xppZ8kFQgWEmRgbAkC/+uKq4VDkcu
FZ6aAA5Y8Fcj+962P2Cpv5nwfXTTqpYUg8RDZCtlj7GivMPX735DJaHUKP7ueX7SPjAb17D4At/z
6VAQyRyA1Hab9lX4vt7b3jlhJvt9EOBy8dCKaZ6Ef94JWypR1yJzzQEu0jpVzI4bCrvtu+mNyzSj
2Hag/jCIHJophqmiUuupqlIrQjtxe0S5cO5YFSjOsWHid4SJYJAVXRofmZngd4GV+NByhlOXZq6W
PmSfzXxcgMU1/bsxrqjZUcZs5W/8EpGyc6KZzl5Ii52KH2uFmSGiELz+dmsg/9hjEKT3XaXxEEAh
q7vWsW+bQkPVhDoFShUzX9fzYgCEqYD76GFhn+OK4vCUiUIW6ql6NqM1KSKrHO51UDeO3Y65NmmY
3uS9HrgyN0Mxyt4Ni5PhToCwSGcMvEiYFpmFaWzBkAMSFY6HTvWx7pAxmbJH7Zbl4wgcwbyMYDXB
A+61sNZHlMS4yRMp0yKfRU6eK6FgBEvVDyOxXxn8s0yadS1wjAQKsJFFceUB3GAJQeBEzcGuD8cr
pOn8ef8wHLCCnhKVvbiPhxDoZB/XjjAYntl9xFRNfC9Hdt2oRLzX7Ylntb+zAqvH5ZUL6SNYLtL1
ISpzl/9DPuIptLQXb64O1zYWqgZ9FvRe6IPMzjdWBVG6zNxJ6wmgm7ns3/0nmAbMX/2i7wZbB+Vq
DKcdVv5RIuTIKKUuUlKuGSZLvv1e5Lwv6czzXSiun5OioOAKhNQQb4sn1Xeu+bVJelO+YLrTc+ii
dzHhTQNM6kwS1+0twnPgMGi/aWJGvWswQ/NtFLIbBkiv4Gh5ORe2Z5Y/3s0aT72fZXOzaA/wxj5r
iu4k+TXkK8RDuqJRAPZsuv6O7rM7ulODzOsumfIcvnXuyXmAWDPs2mAvXyXWtVaWIFaIn1d0o3yc
v1zQXlLZ2IguvDxCrdMZVjYPPMvUIml5/cTYc0XhQnDBSeCOI2xSlL+Ci6POxBZ++gmJATyeziy4
m42aMtmD6DKNT6+j8kSGUOR1tFeGTcYjl8LB+AlRKqQ5k8GShmBzQreFOuFseKa+ElWF0nNGfOZv
4GFd8olaYYm93lGhdTvjia+/iMAioT2Rsy3RP/mZfVmUeC6tUPqfFw926l7viKvLDKqVd8Yanwku
AKRCnk7Rnfr/7eiWgpKobBQFbzGwVh7YIRtbBmHJJUQ5E6b1sDPFS7j6rYItMib3WbwApfjcHfHM
tUmGQkSRn5p7/paEynQtghwlxSYvT5XNKRixQ4r2vsUOTh11I/E35qvoTE7dLE21G2SUUQ/cOoJF
3Ulup+ppmZuFl1t/z1KlvP1YB548Ck/RbCrTyUtZD5T5ZkxQo971QJ0LI80g2Plr86nhc0f8UQvp
YPGE3aPEN9sGpcjAMh30HpKFEWQ9PKEPiJKaMgCIuHP6YuriDt+RW7OftUIURcD79l3uFHSlAgfi
WuVrDMb2EyUeUAH9pZv6UwOv+4TQowbV8p/U/0czkKvPnOJ+urozqVkG//wsiHUqpvWGdbRTCV6d
EOupywI3azbUxJz2GiuASHzm4kEUCeU9yUB2aaLBnYCKT9a/Pzs3CQf3VzjsM3Lq/9mfmJqMKjJK
QnjOr/cx9SZui5a4W3PkjTOVhJD52jjk2OyJ/9DmFGgCD7gn+23YWcfkLRfSHy9PgWrQn6q6kIFz
Bmj7CwcUrzUxPyRuOl7NhZz3cUN+9P0C3dGRkr28kAqI6jWy/4A7+6Z4tXjjFZ16keDIekwZtmJf
VswAdK1mEdfX73A/r5AjUWBynJOc/qmAHUM497krDkHfBm6c1b1UdNyc7gf4bO38dPIIwU8OBlqT
oUWdF7VddfLPIDLeEEFafT3wxaf+cX5NkwhT+DG74XY6CqwPxdFRHv3TmWZQ7Vi1vyxrR3nGZ/eu
m5D/dS6ZroAGHyzMeVCZ+0oarWYf/dVsgjgweFMoWVvhRBSuY/ZnZGwC6G/vvF2Xg/AqPDkI6xId
gRWNvUR4vyIqnRumhCahJL07qq+D/Stxm7Z+Kp0WtMNpfYEFPl4sKplnKMx6EfyqeiTl3gkP1NTl
hlRfFuKFwkL9MARo18Yi9QhoZ9ORxoE0oB9Mfgi/vlFViV4FgbSIKNWjFrP7vmZarOGCFwhaIaX2
fJlAfjOLAnSmXMo0rNMN1+2/1Kg+Uyg9XVAdAIN0ixsHNnArKp4cC9kK53imVaLiIr7wqb/aLWTO
vqTBJy06dB/cZ5htTREsT0qga9F8rc00lDLoJXcnmubdgD9YuUWsByQNmn3Lh//ktClpLecWSWWK
ENtRaZTgA6UBdELlz7ML/KWB21/twkoVyf2TfrwAaa+cCVhJIHYDbwKPYa40PM8N+ywRDuJj9gYy
x3ROHqeIkiDboFZwQefHTmVUX1RCZ6iSag2FyQR74eb/+J1Ot3wOCgLru295kUR3Pnt5M0nO5AJw
8tZNiZhZO+2EiwCwTVzhGMcMO8n+Xy/Zw5DkfcqD9m3C4Rb6lRhKOwZhsSwWS21Bw7tEoYFPqi6X
71DUgxGHpBrJYJisYwbW7BssjG+9iLrDgwEcJKw1DAtXfj/LlrdSMYWoWkoX6HdEsXVXlaJb/qh8
GttfE0lMcfo4nEqW7ZnLxI5Y32Ml6NPyJ5EjZT59wbGkg57+YF+2IO8uDUmFn63LND8TZPucVh6L
kLsKsC0rHtqSa/L8qEfQjpXuaRo9gzKWwuvpZlQdFLMVMEC/El7WwE4pBJApHbnTBqbXBK2ONQqh
4rwg8c8iLZyJH9ADyOdiCPKXPtDxBt0l/A3mOC/5f9aQCPU/cwXzKgtw7TU6nD4BJ/rQzMfjeK3j
x4LTZgorkvQDRsI+kxB59F9kOU3SBd8ZbT4mquZ8+L2k+nbMVfPRbNsF0HGCYLmmFbBrVDjtYezo
OPujjT8aSRf6drDP0R3rQobKSYC+bjpWmLvrWHJIqJpeyMSnVU+aOx4jyBbuz+oxleIq6F89l3nF
4gssykLZYYS0K8/0c0J10Zsn0wd5GJokZqTcKVj5gV9JROZeArebl68ztIC1HpB0ZBEKJdhw17Yi
Z7iF4UJ2tRgW/5gISFRJ/72I/GQBN0q5ePMlk9+HTYSKYAUbQF75JBSI5Jb0eq+MY/tuIWbCus8k
nvPWaX7TxpRi4T/l4mbg0bxJZuvz1xraWrGhkw8xBI1jhZ5MP4RzoOJ6mhaI7kqKCPbcFjeNcMGa
ppYemdmQJ+oVyK+qZcuM9kZIuyyqUa3yFKjo5aed9T9ALyI9apkX2R5uLzknFgJ0kRz/Oi1UVBEo
0WKrke9gqRBnWFq67KuL6FOolhbmxRAZ0OUGpWSmRS/+gG3PZlFVNw/0q+71L9CuhXADUHDDPBJT
IztiRbTUpdWh5tOyAuVhIot8keknhI9wbWL3azd6mvNoeT0ohTvJAd/cSM7vfN24Sx0C4nKwt3x4
INFspU4Opd42NE9DogygH9DuPZNX6ogMkStQ7pNuwtpSkgbA4TIURgc2k4NDfdozgQ9sGbq/A+ro
IgeYV03V/tr2v0rw5m34K/gYNcEYSqR/Qvk+IaHxA5epIJVrqDHNgnmpXHvZEutwmzv8XEjmedR0
29SD6nWsg6gE1IY9JEsC3q9QaFc19oL4c9x1Mkenuvc+vdBAh7Wn9rWQoWBQk5Kz9s1ESLrrIJ/Q
rWu4xrt4/lQFoouQgiP545fUSAuLRVYpx9WcdstBTJ0/WpItw0zGOAoDSmyCAgVlv+K+zilQ1R6h
srQxQ0PcIP5ZteTV1znC/lsJAEBdZmtTPL/5mRmo5zqfKSqDIFz2goJqUxypYKvnADfJBCEHK+Q7
D3V7UQSO2FKGrEwulMGUqwiSacsMw2gPMCqyAG+2LtMwdRFrVjrjXNU50nYh3pP1VHSw4ADbgl93
G0TtP2Exq5XWEQFJUoZr4UG/6eN/U0Mz/g11fvn2UFoOqZIrAfhSNMoYjwXKEHD/kNcckHe+eYkE
N+imZFkNnh7IkCsFGaUIhWrcQMTLgoHleBrVlho15p8eNSxWDV0/eeTcmokTBWicrLZ5YUMhV2NN
++sk57KLm8pKA8VbSdQQpzQmaGStWotTDZkU+RG+AipMZjGZCtozZ/9LZDLlJNV21A6t0lU15OJb
jr7pu8TmV6dnav2CAzmJ9S1cRXyNFLjF6k7XJmo4SBQMjTWolQh9m8St56rPvNcSNdi6jB3qdKQX
j58IaWnIHvrVlHlR0RkXd5gPxmOcLXmgT1eLz4BqEbVbV09VkzQm57agGU32of2N3Uc9RlnV7Ao0
WIPeb4Pvve5u9jnQZcEkwklwiqyTH//fPTer+EFx5D7OkKOh4LFiBY7GrkYfYZ5uTCFBpp1fiW9R
ci28b/yZLpPz0+K4UyXqYyPubH5uqkev0cnxZfVZqdq6Kmj9SVKnd8YJydekGyRm7vcCgd8gAPd/
0pn40mph1ke68crhj2HdQDEfsbhrBiLW5J3t0/LzzbA8FzJ/itZXR/MO5O2gDTJeXOTtwmNNxFdd
LO3H7W9iVeEOFm3TAyYCYiK31yq6v0cyYCbtF0Z3R/avCWqSajwquOMOdseYsGFeEIINugnuDDp1
GBsznLPVJO3eayDRM5mtf5jiuGFQl5Y/7VKE24ZyZY1Wa3o7w+LlO+m4HXZ3AsVY3EKV2+JMRi25
XTFq+1gOCq1d6BMBEGhgAPxhHK96GharLDBMID2RG6QIjWbE0V09xMHfGNB11avVT3GoH2ZYRsMA
o3KSYn0oFmExpQCIEPkQ77kUkbSYsuToUrsIeRm6ADZ/wsaEMris2ga0QesJfGGuHVwJCPpcvMK+
J6dfgvMyCZWB7XlSacKZwcRCU8XzjnKmMVQydSkQWM5djno/POyl4Lrun5O8hu/PH+Hzunp5WfE9
LExAFCsAbo12EY+Ms6K0DTNVjy3eX5WOxP+3GWi10Ns1ThDJJs8hE5ulB2tjbG/RT8nv7Eg0+t0B
RLuRWsercAfWJSWCsMvduIrtcvI7Xo6OpyMQG9IDBgcwkPHwclCYf8wlcVqeUEsrTY2Q4tpwVjD3
b4CfIa8BL2NWH+TezTwcNm3XbEydXNXXFDL7j6sQgBdqCMxsQsevkZ6+T28RQm5ciSpMDCIeTSn9
d6nAwlYaiGA+qT7T+NQa4kcN4gcdap13qSCZNVv7Cy3qmd7n8isWUFCKTive1L5qtTAwIWbIBDbo
tHzBJ0Jvq/QKlERZkXbZI7jHXPk7jhF7d3vlYzRBEagqCljtm5GEvgf7upoFWAPYX5KrfExbOwX4
T1J8URe2ytsBmQ41zUKra1ZnFbmxPvndmWx5osKE8ip8R6dmuosWDS6W9JsH7etxcAw+CYRVqUUQ
TDPoukn3snaIFbOluoAhzufDtoLhhJSX1aZMsRO5R9gLXDtfNN2/KX28U0OFEQz2yyRQHkQTE6Cr
RoFx1qxM5RNP8qCr5UsZvZ1aqf/o5qmpaDtggV9/pJ2dQQEkjrfU4eEWyhTZhOzjic0+W4L/5Kf1
/d7sZhZxRrE8NFYwSENc8qV9TB5OvhvHgKcpgd2mNClPgkDBk2p+pIh/OXmGkSuyEdeKLYHATBxG
463wXgqZpGDnBYU/HWwDMQ5ZsGe1vyGmMTO0TEYj9PkV2+AtZvlvTblPmP9lY0dESC2hDwZEdWaX
6LjGbGb05xvG/c1KLVghMciNDJgmkN5RMoM/EEzqT8BqV9AKXf9hDe01dTlExnPZiBDTivqKROZy
CMLnvtjBZ6s2jswbkzFx1e2CTopUCdF+HAT5Zjyl/RHzvOSHdbntMtkUdV/BiJVWEk+ZfWCIDg8Q
eKP9XIeXb6U6uffwLDFLCVTSppjNl8204bAUuQH0LMrk9t5G6LaEIf7pgtDorOOR5OTQrJ0vOcFG
1B2Jctx8PMR0TpxUpX5iw0aIoHuBjosnyQ1cOo/ToQTGdFd77pBcepgGYGfwKxX3zyN/dZE4CMkd
doxky9kfcqwqP+O2jyIh/8pheJND67S7/h0fM0cdAf/94Eo5RbQBfN9f/bNrBcrMw58U4xTCtMKC
OIuz/sguqcPKkQ7Qpg3dM42opb3UBsh62Z6+7T5/1vwiupYf7Bkrg/h0t7S/Xjj+KglbMEGWrXBZ
nDJ0YenbxJgiCFOfeTJbZmWDBFvzL4749XwMCMTouV485YmBjQBmtEN8TZ7e6lI6Mm+vT4tLA5ZK
umsCt84B+tHMs64V0jF1K4wUilHqSfpVVwe2TbnO6943mkrcjxBU2nh4kuapEh7k3ZUeckJ2f/v9
L8NY8nkskS5+BWxb39asaSyyDvWKEqyGgDyBWj+Q28wY2ypCfEesMwARMgue9asmKBVNspYYtoqs
pC78hIvaDsMHyLYZAZJC6Gy6nMS7YyrY4VTELkRXhUiuyOsSp9FTiJgE9GxCyy/zb7FiEZJRZ8Ga
f/7VOlCD88xgLudx/NLHnesAwaZARJ04EWT7sfIMOQaYSv/kaTucnDnu2eDQAI6BDFMZS10jTNZe
C7Na5RVxXMttc/p+NCy1sKmgSkwEAL7dQOrVMVMx0Gfj4cBPkChwhVGRNzcHne+mAN1tdahR4hGG
sVBUURu37xc1qJdqpqgEM1gHEs9RsyIZ3N/NlmNEtiSbW2PjpH4D8uHDGRCVsnyHyUqvw6IoAnol
T0R08H3DoC3Ku/MEOvJiAIMwZ4k2xvkWNQrp2DWT02sJ3kNOQvsgeAliqO4bLGOu8+PLxO5HC8En
TYf9/dvRJTzC3TLinFeUM6YNQ3gX0Y7ImhqEiJ111/TBEjU8jHR4kYr8Gviu9tY+G4u2U1sMATYX
oonTBcvXA34T6Ek5SG8s15Kz723WHKWfWZqQyC0gIPPAaM0BEhngnPirZh/7AM17lek3HTvfDEy4
JDKcZz+LR7yKiqTzTsp0ihjrKRRh1XXKgB61MGcW/QJQyR6+DzMGtzA/EpHVRINfcwOVDgEvd9hs
/Ocs3wxDYYJL7RPs3gxTheJ/njdiWbvzFDt5F2gRsreRTU6omcD/MEdk6IEpB8L9UIqOx6eX63AE
abE7HvujMxUt/gqaWvM6IzZcpzY2pljF5IBc5veDebqBsB3+4ys8buZ4JBcy7XD/qJFncRl4m9H9
eBFHZIZeVLHvuxoWoK2/P9JRQ0jlQgVMh9yYr02TGxLD21viVXg3eu2F511ZcKEIyuhqZTujYzmI
i1l7DrxDiy5B0y3joF7mdNLUwmbMWv2h0pZCaVsLWUbZ9BU+vYbMOweqPMSZMloOkcSWDgVEZibQ
w0cCAw/S0qCtZ0Y1YsJumkLxkxnP7+5RF83NHX7CqE51FGpopSPolR6YoOW4uBRipNJZKKDBHYbK
RrGJe5oDsiav0OP6CSRugPPvFl+8BBbC52WU1YmiBTkhDRN0sJTWk+cwTOtqDTtHNERhqP4nvok9
+fYPzx56eQYu6yE/s3jIOcsLhBbYL9ctz0520TRs7CHBkSZTHSTVz7zhVhXce4oMrCL/Rjn/oZkB
hKzNvk3ExfP5vHeqP1XEGym8DLwq1VERG6UBj2YXYkTUaiGvzoT/qfYVh1iMYG+KDzUlekYg6OXV
/wpHUnPj1lKQJi04Q73Q8cWcI+6evny5Z5NM4diPx1cudAeBqtjW8yPsQHy8iuBpiPsnH2A3RnGo
7WTOVVXMLMePon1SaLabC28aoCbiVkuxKpwRQHK4eDfhAid3tKmhfwhtDImt8BEeSinrYGqWBX4D
S671wBqSxzfqQ8HHnIrCQZv4Ec4XnrRTtOVqJp8KRvkgp4LczE/IwWIEV9GnCJBu+ts1Q/7H9Jhh
u8Vmx+APL03jlTb4GvPS9S1lyVO66j+VAMPWpLbIETIwK2mdmSElyFOEz5w9Ai6jSzQOAQZFbv+R
wIDOcESjofpx8W0verFkiiHaW+e2CD9JAHKIkg+ctZGQ3Jv64t48eYkZSjS5AkzwdNvJty9DZYua
KochPfPbprX45W+h8P7jQXjM2+SJSrExILNJwGGWJZ+rH0NXM7CM3C4yqgRqrqIoUqP5jlL3P/Gv
K2p16voejtbuN97nNQyz2NZ8PMpM9Z7fXplPVxOyhAGokrWaibpiSQ1k05g4vkl7NgZKD4S0P3dg
SgmW0Gh12zwkKf0SSyIh00kjsyNAcYz6xdjsD/25c2E/VMrtMq1YTW/it9sitaoXLEbur4YoR6TB
JIqy3968QYPmFBHmaVwIqzXNTUQ9JWMgsl0uScJx4zX+VsgGQLI11pGJgX0Hi7cZkCDPfu+Nt7BS
UOPyapmKs4HjVVnOvuKUHD5whVkWNVfOWnsaCVgBrHIjdGWqNBZIHDAfEXJwjaLGAeyaigp2t1df
Gw00novvAR4v74BYW/2rbnMtH4INHqxbjyrL81fM1CJOfVQ0fotTsoRGMBvTNTXxDg0+Q5Cdblcs
JPtjM+5EnxDfGCweqlJtfTUCEFHkU/ePWlpFnvMiYxce7qUxgZxREmltTfdc+AnLMjVcmFyoaIjy
z/CsyZczE7Nlxi2HqooApe3qPN/B56M/jqn/ZWlzJvMTXFPt60bGC1DGoPOQe9Bf4SYEDPiIFZu9
hvmOHjiFjVEkm79XdS+Tsy+oXuqu1AAAOUvXH6w8ik2wHVGu0lZ6ZRwnxJb08/Ut+0ZnOcsBzR8d
S63EfK/0aJONVfSkpPdmY9zaACMDNj+Pxvu2FXMsp4bMmKxb7QG/CfkW0noi/7EtO7wFrtV/3vV0
olKUlTsLXCSq17GE3K7tsiltu+PH+Qk3lvX0mWBgQwr93GxeKJWceOhSJ0SrDOGOBHgGiglUwEg6
2kenXtFaaor+qa8ZpEAP2XaBITD0P6I6BxISW2k1UP3CHlB+54oA4tqIeiUA/raW5mqq7N//pdtg
fS58f9DBO8Ftww34kjcVLzGQ4cGfPwL6sTLQJ8OLDsi2BCU4BPh2U/RLc/v4Ln9NzrjSQoWpEp+B
LfA81NxxB6GT0/aUVZMdv1b11PpE9FBAYDEDtT/e+Cv1agkaggqSSy9ZVIXvaJVj4boy4+gpswYc
1VCghrBG+PIUOHHk3U6bsf/vst3+Onitqn8DTCzmp53vwW0MqndSCHjNlvb830zGCPXjYOK4UDu8
0zQzLvVICYyRh+IImZVWYe+RHHsIUPgBRJ/P2C6MnxGSwIzYr5AXfiWDi1AVeidPUf70QdIH8vlh
+Vi6p4IW0ndBtpFNNjsMpURFTMnhu76rmzbnEvyyAFgb3ns3H5Y7LRDOFOXldz4XEHlkJxUZjNfB
gPZZT9VnlvyT1OHNsep94anUVLAWu0915ataI/3uLc0PKExibDA/Na4/wsCxsZj5u7k102V0FvvS
kBb8d+Bwu0tr0Jwf4kTQSm13sU94XxEn7kXu7519JkTS50aNW14tBEh7H45D8hIdyWGZL60JE1bc
qZ0JE7hjkNRJNF+nlJ2ORRqppAYGHuUhGMXDQc5fYDRY4qA+dI0LfOGH2TzU1VUPp+dVZ4Me984f
NcFeTnI6gA+dotjf9e7YNX/ASYKIVziRjBxny8ebQ8ZETFfQrkVWW7loaxDHyAZKS3UFMO2zdY7t
N73ESSpglKaLSiWdi5GjHBhcb8bOZyneMDJW11ZNIoXGElGXUKOFMj/h8eY1ngzuJbnnoGAuJVWV
bK0ZN+xOCSocWYkFSr6L7G6iu8bZX/lH+TROAREzGAJq0ajQt+B0iBkFTjJkDfQLVno21ovUeJsJ
XSD84w01C95y5PuIiNbVCG4sZPYEB+wXrAiQOSks4l3HP5KzqOMWKX6AU/JIeykrHNBGvjuAmD8Y
dUnWUGAr8H4zozvsjJ0yBjjhErAS27eFkELeOBubXlnM2m0zh8KVSvNPXL2FYMR5f5kfd+UoWusQ
QMgGtdm5T+C+Pm3r+eA2kcXsCD2Eh6PxlAMcR03pfEDxz3BDPjKMcRk1DWcTlxjYjLTvupUiTeWV
PLJI+nfJgQhjRcvXEGGCkpYOjRwJCWMSD/jGYupVO5gesL5Z3NqgUm4XgDdEsha6PksI80s4G725
cOKNmzkC5hBKl48iNKJuzHFS8DYUOs1/Km/8YZd+caNqxmma0RxeBA9vuZxXBB/kqiQjorAWaZqw
MKH04deFNJD+jdb8c7+XY2N86yiAzRZX2Y+t3cbMucZMl/UxecaJecbqsRh+FVJRi8UIqj4xIOwP
+s2lbJxzPkSowGGeUmjMZADB6BLujWhfqdd1fILpc+1fQf1Mdaku3Q7fUA4U/ylbtsHv9dP/Gimh
ZodWSjHwyzQ29Yeb/wsbqfDZJJVNb276VbgHI9nln/e4hC57m8bo4We8AHyX+sbY2jkeNPXlhMAi
hACC/BOipYNGAckmKTJ48UOC5hIDV45CF9D10loUluLQeeHiTVPiVTaKUO9O5bzG4W2+T1RVPgC2
BRjXmPkXBpMfF3x/KS2EKOFl5LKCyJCEFjgaaBFddexpCRXd9+S/GLz/d/nUv/h3Oy2mt17xUVhw
EQRPq1RWlxBiGmSxp/BfPS5/p2WANoPfzErzFDuGkaLKcIh5H3A5CtVs57YjhGCIUS6BDNaVerrg
kc7GRzLKjQ+ySiH8viXQvZOp2Ewq28nVdfu57P2GsG3yK0+bIzukUfi/WbiGr9LsgKhPyyib8v6T
0i46JBD9SnGYMcQrdvpRj1Gbe8zjnw/vM8W6nPMa5wtrJ2YuNV7jxwa78kEjiF1qzZIiC6cAY928
TkqNg93mgMtEoqZL07eay0YIthnWXBEYWIPddWcl8gyv9cWVa1K89BRuDbTlZ0GNsjZZW0bsK5NH
U3N//lmLSzDVYwLqNsPRuQfV6OMHbPSzJ9/FD2WyG1LWkx+/5q0FJ2MsLyMXs39yJwTaGTnlxudh
4zHV6QLMaYdz/IRc8/YmP8NYABlZ6LAb6sn57422YUou8TZsP3SuZs3Mmv/uP61xUaA4F0wcR4+x
2Kq//rrtUrU/3yUstjgUe6HsSNDt8RhpAa7DHlDnImSpy42tn9jwGPr7SFkeOJ6k1b8IAaibKnZ7
xplnSpoIC83AwCoeeyTPmfCwjHXhE1ahd7SJyYVfEnxU9qEGomN4pnTtMVYdvBV33qVbMV/zIUWY
dcCvC2hYcdJSdL0L2qOTEgBEg/DNLT7JaDPt7NhrE1kCCBStsCjknfl5XpKvh8HuFXmyo26WMJ1K
Rvp1ix0R98MMsH5hvJfq802p+RtOh/EMpo9HxsR0vV/XELIODZVSj3U/FhLx66XHA/iNEkLqXcoi
Gd3OQWxrRHaaDLQ5VKk9OVnFVeFyr9bmTZjEODggReXh+84im/1fdYktKqgzn6KjgAf/ZSe65Zid
l64O+cQvL95IAZyQbusPZXRghjBFxpIjtwvjApyT0fOgGYFUNxeLrM8Shb3mJsAVy6y1yQuovJka
dCQgAx4dFivCex8roJNXbf+A/+o+mrVje0+yK0P4RXjTkuFfynKuvfT6YXXzkn7kMJAMSl9WUPIu
+/7TJzkQzwxg55sGdeG7dpANEcAigoegqPunPKEzIuMPTb5HeA//RmugfndFj+LNl4xO5cw9Tr1R
Lm9G+3Y5JSsn0XJhrtMihStUxyDLBA4lUDXuoGrf2Uxc0HqnDkrwUxlqgjBc2Cry86IbWeo941SW
PIM0Cuwsqg/MTaiK1Xl7R0xkCCmbtlR+ZoqDEGAtZp0QbMmF165OBGY8L9IU/SThON1HpdK7cs/R
5ETF2Zbadl7R3WwNLdNvmgBf4wu6UY7b+XRqQoAZpMggKY8xeMw/YfVKg7hE4iJAY737PmDWfE0M
tHyWgUlTnYfgCg4bx/inld9cY4OUx4uJfCVPXmB8lkNQucbQ6Yy5D8hT/v9PIXSUx1aK5Fjde8Vj
p/BCh2K7lWmEzklnuzS71EiDW/2Q6X/GesOnS1xFxKNWK/GmiQmZTt/HXZ46ECQ9dtAGDaFxu3W/
9zHJzbGSlKWARYp/6e1E9AHuISkF8OFHeXbvOnQYR+iOoN6NjXn0abZAH1TXLFGn2iXqqsF84ZJ8
/JZ1aloV1E5gKGgGtAiganJKQhzwLrRslcNYuyzdfA9VE8UoheTzGhEniGV2nABbVi9Aso/UE6Kt
3mr3OkcnsmmQ8wrx0e1Ty/DXAvc5kOn48S7HYDZgyw8fkfotv6qoZT5ZcFEjRg8avbzdUUzGSxui
73wv9gqCafLA1/zj9j8UzdhX07XMxDAmK6K4WAPqZcrKJjn5ASpXxON+Ln9W+LwzPUBDvyYGqP/G
m2FjEoOhYPRJggaEyBrS+IX44WR05D6oA0cVxv839sFMNRT7H2ARw8wFszvbkQiKv9XTY+Otfp+D
2vdiKj8a6yXGtLmSaloE851Xhobx+cbhxu1uNpT0+DiWu5kVKCaCqyOinSLvivkS4lKdqBL0mFiy
OkobuVI7UaumIBcxltSNX2ql+wpI769ATc7TTsPKCHOdqprLM5t0nf4yJUvkWaSnAyKbqFJM2TyJ
N7wHAjfhywApABRqcG4yvKuwRKO1/DADsJz63A7ghjxFGSgp429pf1JJV5ZemUx+SCORJJj08ELP
5jbuS41nuhKKjFK17mbkKMowQTsrEhuDf/iRtuOtGj8t64nwRTXp2johcDzdxpDdydch5tVqq2AN
TJIBF4ZkRvKTfpNJav6RORLN1kOqCH4ugUEZX/hpUWnt7ChcxWSOdsski1HShGLwTGNpWGL8ojRP
NHsV/hExisgwXs9tNww9iV1Xt1ZEd701H5+f5HSPz6YTGkh/H1kIH5z4DzWlVKHUGEbNexMfq9IK
16GFxuVexAIypzw97E1HnoQUqThqENIEg1QOA4aKHWGbr84mm6bE9OkdjBh6jpynBa0nuhjijGby
o5WjKnrEOuG57/8XTbky0vCWNT4EDVlzMy2rBp5r18qjvzP/idmG0ufIxZ7EVPmFSlNRCmwctoOQ
Ll0a5rdwELvMqsRJ+E8G6eXbl4+31/e1HXu7kXf02KeUqGW4Z26G8z3vrUb9uejlohTVr/M7Y82+
S1PP0HDAQGmcJ2aeb4lTTGrKccPmiDB5J45ZJuDkBVdAeeh5q5CZnPnvyiHWtveUsmlS4jLwqpVB
bL80eGhVRJ0q1FAsPJLjPPgfgQM4rnMdCwtXtQ+Dw1IZ4F6II+xTR4SZJMfQ7Fs2Kli3CJTjqKmg
RbrzMxAsrNGr1zH6g7yUH9ME4uLeWsigu+xhfE/YFPnHwTtVIy/ID8vRf1P9MUQErJJ+Jb3Uagwi
tnYz28gMW49v5syssURXfdiZczKuzSlf7f92V2pmEJyuz8/dvHi9fhLV0SLQcJbYF9jaqkP+hUiP
eSGMvZLjqjVpuQ5aS/cAIWIFibGIyQLA59eYloT+QBjAAEeEWj7OBx8xelox3vOYRs7lCoLbb6ny
T0THEpq2JOIvXgA+JZ9QYf9+gV5qtvuW1HPMbiGmYtJDgS/8BNs6xTQynvhYjwo3o1ntwZ26WCEI
OFLNdFb+moYXcHjHJxf/9HnbxPDEz7IuGlhoZ9WlMDTfOX50TRTCtcgVGXrMcpbFpcIA43ieqPdG
CAxeTpROhIzYCCIFeZG9leflmiigDdlj9NWN2LPBrwxF43x8NKWhxi1B+XQdc5A54pesH9pMJQm0
YSTr1qyZCvq5/bPKvDuFrKDvuMiPT61FIHh/OrPwm/GtkjfBIPjat/ndws9F4UqMB4fiWK3wgsLD
fATXEGeVybKZfLw29fYcnByi9Uf1YjjDUvPn9g0Iw8E4EP3z2UFgFnsUYCZmZtcg2PA6SjTa0l2z
W4lOLschvDZPwbUH5oR8eQTNCa7HF8hBA/VX7vto8VMlcwghhUDdi3OkYp/Cx67mk5xGncm38vIS
lQMcDQQJQvPIBbE1Ha1byPUHemA17u0d9wdOXyX82GRXnPFdqns8nldr3MBGJM5QPZR2SIS3xP9I
iW2nsr54/o/KWsiGv+ynEp1EjHUd/IKRNqEZNf2vr4CDdMb2vsqo0ptXtxFW8j+rkeXJhEMVUZ4f
wmD2wmpFs/0EPbXM2cIQzVhTdpYvu2sSgHT5LvWoKXFpGz6WWoeQv4tth+UK8kbv3LJYXKMye3vs
8Winh4xJVU7IvXFytnU3y5K11EbJT6Qvjp8v2b5HDaLlCdTUiJi3hJq+Nbp5AG6S85IJavl5sx76
sUV8aPxga30TpbdcfL8MAMKteWA34/QM9IKtGiaGapuw4za8o3HXPveJtrFzvCcPuRU7/D2BUtAU
bgQGavpvqQtZboq01NzoCSHPgAwRAC3YURgjUVJI4kjS1D5fizUIvXUHczbmY3YRSDF7+hAyoRwX
Wqd+HS3q3m5Fxz94KfHWprvVYYOxgy9hgixoYuGhO7T46WMBVAoomXTYowJ/FOGIz/hYBX89+Kk0
7sAMdNeS9S8fxDI7n7koKG3slTZSUPS89LRxwArlCDv3Uq3qtGD1+iufiQdGjojJIarqMlruuVNt
xEUGF7y8pPwJUXlSpfLksG07ZxZk/B7MjtIvbINnMxdKoeO465VmAnFcq0BU9BhncWyEaIHjrNhe
8vfOE0UKUSquz5FNiT4uf8J623wCWFN+UiBUvgvAJW0kP7m3MwvW7f15lYwm5pe17i7kXD7DhDFJ
IorM1gpg7gpqICXFlI9ZrimOt00OovIDQ6+1IRRsWxBA+gTFo2f7tEF6gVfD+PHFZbRMXCiQxqq2
9gY2a4A0NBPfJrGxbIMnBFtJKZLXtcazUfuqFOFsP4pvgkiz7vJnb9vJZQq2yTLHeRcBvoyuzI7w
YXROAyFwzvxf9+LWgqLn42SznZlEVAE9depxlNzIGKEy3DFi9B/o5Yjtw4D1ayAqIM3yYlR+N0sI
Mvzm5fYeHuExq5XgDB9+4FN1dMe+8jkX/CXGSGxXWWaxM9NKPgfHlUhe/fMdxLbR+mXop94a+jIV
2H8DwWt7CAgJpi4y47Ft+qZDXbWXMMk7+gES5KWG0wF97GUs6FXEBrOwdA/1d5eIlixmbshgZLqv
gJ9Z+j34Muiwe6g+eWsAB7sqTokHVW+a1nUjdMdNlQDjT4uVAbqBjCPxN2B1yJ4uUtLQ/PkuZigM
aPq0pOaPE5hxtRtAOi7s+5DUmfY1O4k8hwheT3gq/uE3QDxBN2rQ61icsQ//qvXuCKBYH3xsigS9
T98lnX/mDnhoRtbu5F0RwD0LEP5P8Dsv19HTAJJS7INa1bcsiIyi1akWhR/gTgdPYdWqHZQLgmkG
h+qKvLwg7FMx39+pnCxqdubIvPsPlky5v1h5MbSZWcK0jL3ByvY+0+K8K7zPonDiRFumaWmko/gE
l0Zmjknpy0O/nhYX16G4AIxCVgIMGvhCRV4pK0dqsqeIqIz++S3KpZ4ir+huxpgI2tu31qiUawPq
zBmNFv8XNcp98n/RQNJMQaHTXq+tmL97AV7/2ai3zxqR7bt/D2p9mguluN46+WLIBLVzdFjv6Xul
/7U7gqI+eLMfhB/P+Wf0PnRgNFwXid/9gOWNB1iYjT6zXaJuqgPr8BIb4owNNDqqxOqT/xvC4B1j
r8lPGt03D1o8pE1+oF5n8bT3EhGD95L32sHapZ+LqP4rJQ6SSL/cQdJm8hyiUvsHI4VX+7fFnMBP
uYYa1/GRteIiShwWC0oQCe/4wH8UCqOuD6lFSNlCESz+MCNACbQX7V5JLUGVzUDNYs917MG7Y3Cn
yOWEYq1YhJZ4UNL8pnEasiI3lNTTSLp5ngBNry1cYQB/coL5Yr2NCccKk7X2ldMLLw7SK8MC6e+7
f65c4bnF2bWPENmYAtaGnKJnv9Nv7znhD765SiSaJDHGwCCmuUmmQyKe8CRlvzwSHC73izmZY+k5
p1aGyNxXqR0y+L2/mhckYXeK7YLG3vAQMl46pBhcSJ0QEkFW697J8OzRNmmfQzk1BvHoiO7WnqPB
oQa0n9mPBjGhDQYUUlTQ554BMegtjYP0nCCbO1HT7xSsyG1g7k70R7Xw1DN0K66Lz60sFfQi70Gh
6CJzBUWOAynuYuSs0At+WE3QNAoU2nkRyBg/Yd3BHsdIh7WjAslItIdRu0jW2QFeCEdd/28vM6yM
R8ym4g19W6aGonSyy5pMNgWgQ4eJ2mBz3On1/hU7vJXez+Iy3gvWRsu4yiFXNx6cTL55UPVOrawR
4ultR7UcRFla72Wxj2zHbf4yeBl0hHVA/l5kIxFjuL9tId3KaXOdLvhCtNJjT9EPRrzWFq4MIvMP
szfpzDdCMiWeyzN4Uq0cjqEcLKqrJvdOTK201KoAyteYIqMLeZfhvUFobeAtx92C35Mr9eZMM/4f
94O1sVw605GBheWDABWrwAih41vDpYbScWSF1rvxfdp+OQjZxEBrUxrMgFq+G6vuOWgHiq8Bo5vC
whlFQkOQXOgtCm2nXuHcgzMPPSaa9qI7UD/p5GFDew8HLNvLxR59xi8n5e3rHbmqcdt12cbBzQqz
BZlB4Pzba+Zg1xVyT6zlDS9a8URipXszKgDdZy52Xfb4bOD/+eoRfGBWzKVZEFeduSpNVEcnMQfo
tUdy6YvQRtONeazgUgWFbutKE2znlV/89EYSSKOToQKk7rSKV2lwoqNbN83bIi7//hPbE/VAiW4B
5EeQrXsjJlP3x2Qod+5gs4ykdKuJLTGbASxw2KTFwX+pq78o7tgeDuyTusSkH/24DSwtUuP26NqK
fSlUYTXodJ4TLmo9V3cpXlkdx6EBpCHTAphvKB3wbFbYalCeKaKWH5L6Iq9g1Rd6hWzj5CLDJQI3
byhChQIQq0bG+CSKZGDUvRURqVIw7LLh17Ero+vkuAazhFM4gIwslfDGhTyPANSVfzE7XCma+7ca
6cozlSvydZy4NmWA3V0nECeQMaky5fr+tNDbnbaxRVyvCI1fKmd03/4eRxjoDtsmFAzNYBbwx1wa
DxtaZePna5QWfP0Sry3us63SRVCmIsMRofpQJhCA9+6+93OFDrqbbW3hMg09HpjXI2CMc2QBiTOT
L6cDzuZw6n0P8ohTxMxiTqX/JbrKZ/AHo1u+iQdDeLVcCUeBREvuOyPFVBrIzhkP0BgSmJuwfamj
IiZ+7R5UNTgzfxA+w6C/a+NHM9sHpRAMo/hGAWIFoe2WQh1U9ii0iDMVozpxL/0ro4eictLVW9yr
FsMWZbOL6AQk2Z8N7iVcuF+JB+bLe4NH1afawWnZcicC9bIb8SS3Kt0goAa/3lE/aBRdGUCVpm1F
M+xWtLCr3/lr0jEQ8le4krQzKDKsFjMBBjadMlnq7wEIIZXJM611FP8n94pOHC9jSOcipuGOKrtd
1UkaYTm86D2E5n0O/Dn0ORk8WmB2l33k89YtX+0o9ObyxkS3m8wc3Dcq1vpklGOEF9ynn3oG8piw
GJz4sjl1/JQHA0NAgMkBTGFgWX9JQfMBu0Uka/JhoAYLC5e1UTE0MORvW/HvTGMouRoPB+NSy7Ck
vMPwgQEbXpn3+eoJ01eoE9A+SUh66DxVVYHjyim2gLziESPc1sMsCMUkAnYQvOAr3/27Opkrfj3W
w8h3gSUiTAATBPMrj5DEwg4AFHTpa1uW839ksMj5GSNl1pysSscwcMeh/hs9WGZmf7qcUJLofYNW
xJgzomcAxej5WEkdGBNl/oS5/PC6QWfFyLY9v5JFlyKeBI3q47Q/FhAc6Opsvaj/2bNVoJzEc29z
A0affM8RTWI0EyOZRypXS1xXeaBA3LopzXgJd27rGr3ZRbrAAG2yAU49DZs3HmkxdNcGMrTEYjS6
D5v6x4npsM/cwyijauRBkp2/gXBuJpHvJD2bAeLfy7enKBYX/5VsEa2DomRhJAvS4QJ8nTJDQCRa
YnYVEqlyX+7MkOz4k7qZNuvv4iqzQXwKDicK1Qe01KAQLhGfXP8NV+UP6+SF9D0nCNmKeQzxtwnU
/kwErGvXzib0vB6SFRzRRDAHDZJWv6KQDeeoHR8b3CTRvs67pGacfJXoMf8V5QE4QzuQvTDhWtJj
HgBr19BAMC4lWhehwGOeMmfoq/VraCluM3jOe27OPtaMuS5pN342YqJHGc1vD3ka/qRaCkQVZF6i
KqPzZ98T15VFdfHT7mSbpxygXwGVww3ZaOafvyiqGuEOev91x1Pk7oAC1kM7NFqrPgLWpGLyhS7Y
+gOHhp6ATZGbukROMgovu+0MvSSuI2FMyRcWzYNyAaIFkz3e26NU0pzQgf7hWVbc4uXan1bVAtSD
nfs5W46rNlptqBqGK+XfnMLn9Mjm9uuu9IQ3iFOVa6uvsnVUtZrIOpcIc1W49/Pe4KHhXr2fC9Rw
O09hsaHzoevKQdXgdWDP0re+qHxr08l6SMR7vO37UqCllKMvhJgl+KP6IyakO4EjMsUfxasK5x6M
WAHHrRZsFqlnhC00cMv4RwMpUWb9CnlFLVRXV5VJ1194GPLN0ZZzjstWYMDtWZAaGj7c1zuRYpzF
AvXVq5nxUqzqXjJCv7cjSaFBTKtTdlaQ2msfZoAPdELtHL92VXzv7JZEM+XHK86xP+nXVHjGIq0O
8MmNm/y0gt9nzQ7WWmhiUkN1X3uSrTr6Wz9BhE+md/70GouT98x6bWywaZunTjzHH3LQnU8g0kwP
KUhSvD7Jl2MlHE2LkEUFzx5YxL1NmA5kUPbaZ4/63U/bVEQePpgqZbjW1gVAVPJ29kDVMljkgq16
GbfxQg5y17VnfpOQDHCLJPwwRuwJraowVxKDGBZJ0yE/DfvtmHNwIMd26orw3GNbYmz7soiVtYfl
ggjhkHS4Z0E2pM1Uga1MrPCx3UYB+b3or4PaskWT2J97KwJKR9YRqSSqpN0x80ufB9CmWgMNXAmy
NVx3+ZRFRRnstXxATqNVjQOZA1RVAILB9beyz6d4l+GbhVKRQLE8XeKwUroTjaoFaGXgYbizB/qr
DjUZtoz5PTfnTpPGvSSXqeTDzSkazTbspwYycbkOzKpkntdhrdPm3Vt0Fn0Iu1JyyWOXFToSTsso
nI/CjldBFT+Atn5pEL2ZiWe/RmgmczzhBuLNDgr98WsmSPm6aG547IqBZtqoU1Xdy/6GenothSim
S4Ad3e6/iNoIT3iRwKw4dJNKkuPRsAYVQTt/JSgzKXjpacN00dX+HBdpU5PSSogxJ+bc+Uj+wEp9
rSJ6M942ndP5MoUfMeWYAFPUYRW8PdCEAEysGj4o92QneqT72Y1TY0tP+Vkp6Jln0KhBD23qHDL+
9G4BgcPgk6snhrev+cVJX3l4VUkvp3XEhNDCLy6bUyo1qTECTZ8gUOTqH4dsd5fZdl94XNcGaJsf
YTpDf4ktZFHc3SQeeBfQyhr+PPI4U4KS7gGPPlSwpBKDgb5BF06AtwDdEmPtsI4xv2XlTVezfnCY
+mqT8FO1y/ASJZTS0Xiel1Nt7VyLIbW4pzeuXiXhMuAAsTmm7m3H32nQF53ihZdYyYg4Fqp6xUT+
24SF/fD0CmLI0syjs2XE10ZvD0DLup/rfQBGTGDXSv/Ihp4LbDYjaHG9ejY6iOqUXyqlzEG43EAd
DiQ6tD5CshOwaGSgfcUQi1Lswqt29QyoBSp0TaRwiaYfipSD8h3BGmYSSX3djc5r4LRcOtBYek57
plqyonQTeNsKahDHp6VoG+DBLEqwx1RcsIL1R+bb+Ob7pwOEjrxHJh2u1claFWnNKs1spumXV3+f
J08P+fgbx0miSXBrA4c6yH2JHZvJ3cejy0hzht7VuglkbUGjPCtkOS/kkmShU+sgi4BcCyFAP8I9
8J0RCsl/XEYATjV7dui4HYSQLlNfSaq/4fmigeaMZv4U44e2x8U7lnd4JAc0rPdu0VZI0ineBsb+
bldwW2T/OBAoEJBfyZQV3mLeJJr4ujvRjlcTOHsXGHKEFnOYVUClSWoVPkDmqF+K10CBB74Tx6PF
/cD2AA1q/TnME/z/My1a0xvgdlVQr2aAytDrXaod9jELR9tuNeWS19hIifGqAHHioiobpzQ2i74C
YoAY4+ZEVki6KSgyYFv5ePPEF49YSGnXDMgJ+sdg+uG69VUCH6J4GhVjPke8fK+sGSv1v0yuS/TX
9la4Fg7VacIaiTpAUcG1oOY5FRi60XsfsK2hJK9tMRKCZSE+yKjJNqDtvD3QFXWPtMFe2qQyhLXM
B2ZwD/I8Ua2d3+kb7pgbxg3oo+0NdQQHG4wwBudWksTK9yItndP9qemRD76IKECRyEitzqc3KB/N
2+kGt/5ovO511Dzbv7HwEfCWSfaiCUVOVZjlTMSHHFiTgrNxH6G7hIyqZf6moOMHmq0F9zJhvfSj
F+KB19+JTdDgpRok1W6Pxd+yveS0kaHYaerRHk0CIL3P62eyY0l8aptpVcO27e72IxtbxUOjFQTn
gGSPNiaxoZ5+lH8hiJMJ6+jVF88HXqBXpr430gPjcK520cD6G84sA4tLePROKFU0iO3awK3Td+CA
coyqAGYUS8tyl8vTIKeuQpwDblhPjlCzNi8lXiNkkiz3jZU1Jb9rcAuA1yEFUHKZAmo4ijigikkQ
h94Mr6fBvXJMUdUqprYv0XU8/gwlvYKwjGGHdbzym5h9rb7XKcq8pp7Oy8XlcLqDc8rY5fA+0uaU
RQqexZBPBOxmcC5p+90PldVqH7PoJWORTBoXFaI98g+gStDcxtqJXkcQv+HzQQ/iG0UBv/gZjbd8
t/LU7JWmhzsBYzpJwfTZxSEzVw+Ti2Ps3otfWyAmDd1t4RP2jG17tvjXyDFAr47DeDh0bbCZ/+3d
AeSUnXZxT4LaK5MU1D4ZJOCUFkEknC/kzJ6i8bcwT8RaBztVXHoasG9of3azHpTukNjm1D1trv7g
ycseSPoL9xQ0FANmP9tysokrh4JyJCz5WxKeXSdSqeKcnqOqOCUA4daLB5Ef4Cg8q+miCPHUpqEO
wQtgrurtegwFg2AFMFJAxf6VSpqpnGCfb+bRDuknuqUm1s9uHcJ9IZmFIYR9VD5CegOkdP5LTU23
nIne5aaJ5HFijCXQaJJnd1LdKsyvm/x5JE7zd2o0PNtyfOmkwvnmK2j+JQdGK6Xcp74SemKqnZiI
66wn19bw4GO+fiOzNVfL+5TK0t8THuO1Im8z2Yi8j9EoIP9zUcRZOXF9xYXLI6S+Hq+mhPXB8OpC
HR+GjR6colBQ7Tlc2Yk0qhub+tLgoVUm2zE12/VylO0hkLjKEn8lsiOmBA0R2flJDJYq9qhe8nf3
FwNd5JmuQcmUN9xpoAqZ8K/rfgt1LjF2zj09i7vdka+Lgi5F0E8lxcl+zRkOsO+kT346ufYt07+9
dMJEZfS27vE32I0Dv1PIO0EAvz0pD1iErfc15YQaTahxRLGNH5w7R+ZomXKBiZdau7pbystQu/Sf
o+KaLDmWSz0OaEjV04GP8ty/0Dciu71mn1Lsvs7W+SgzJMBa3UbsFrYHqlohBcQaEarWKuS6jB6E
uGOimXH2QLhjiX7A4fkZWYnMQApW85gdGA9qy5ZpJY0jg1GevxxaJ3GbjOBpXHbYBFjB4IHT9fS5
lTqg5dCu+iO3Hg0CAUMIZ7Nj4/mVbtVPZetjThPeG7JIEm7bOGfXNtdHV7fJRKFI5hKKtvmKwWLA
ZJGFZANk2bn4/CDVesBgWM4k0PWjeKv4yMQvxHmT5dbsX3TlO1Jw7Ydu9jI4zhyoCy+OVYDNx7eY
Dzzes/pgevvvig8OW3OmqhEai15MqPyqKzNIeL2Eyqz67+Bx7cFsjBlxFFx5I7FnVjGkMHCr6k8r
yG9uZFWsTFIRkUhPtpmz2OddeiKML+/+srwDvemHp8+yKxGWEFhPhPMjS/nBq41P3vJ1Nkve5dDO
isIDUzPNOuwkqSFDkX6cg+k5jHhsL421D0lb8UxAxWnkjPw6UdYJ8nxtKHfjyuws6bLu+pGWX17x
5ysRTXvCovQ+ASYcN+E6skMbKrJqB+Yu/etcDopbgFKcPtJVYOQ4OfdsWw8BRcqE6F/KU0e2Q306
uaRE8hHFQefaor8ECRQ9Km4//IA1UOr7qksSAbpWRB3kNomdG4gOm+/ph6efA7bJkE9lgsE0CgZN
wQxgK+3ismkwO+lMv+o2co7VMMS2dSuA1O3HFItVPll3lgsT8vboKCDhDIKjtDWccq2b+lnqlu6a
rT1EUzfjloIgLv2hxKLBcungMIXihkTUhVQUnWn2/DvKmKmg8msmaIyBF7pR+ZJOYsd8UDtNXVYr
VbV0rqL4o421W06uXlQkP5ppC7NnwebCV5K6Vfv6V23KxtgDERICE/iQiy/R3ewv0gV3QsWyUuJY
Npo3uLvhEiiwHsotQrewOrc7Na2TE1QeBUH/FUzZRJNQ6g6v4OL/SFVqWmdT5TxtK7faAgwtBpK5
4wvjlIKmtpIDJMQUnycpBbBs01i3MYP2w3wREw+auQqvwMmBYmkrozrjlnCFm6y5bBEBicua2gq5
pDsDwusSnLE5FI6o66E094RkXWjMRMdsqUZ9ugRZYmD2kNev4G01gJ7hFKt5BRpBLwZCbmdgMwsZ
p4/kl0KDVhmdEp9VWUQnXHJDfTp7daKRHLyPkYEOp0zVCd0HPhyll6ZwxcwxY9veGItBZZ9YFjax
tKmF7J1HHkAfrADutOnYbDW5D0iMmXXEE6yYss7PZ9dLqabENmmyBYhf9HUMZp9+NmuE4WGKyuxU
hbkYduhG+/7gccZ5XkqvoAF6LaaactGDDHkPt91js0d20IS+4uJsyILBb8Ooie8BRbMhsK0jvkhS
mRgO63Gyf63VAaPHdJIaaux4e+ub/czH8xJ2BWsHiWrmIdYi0755Mfd98Cz6zs8f0c7hW28vgvDZ
5Wrfm05EqtRcHnPIg90fTtI6a1vgGRqy558yWUjhKLL5GbtbVjSheuhIi7YNCp4KiLL9XmiDOSzN
9sqiNP0Dyqwdy9idBj4cIY+R8131pnOiHpowUnlHod4L7dFIi9Xj+UZDAi9dwn4KmAFJHuVLjv0r
UPyX+CcQZSXWrUQwR4HIXxOgLCiNMTYWEr8F3IOl2UfaZoHQj+JaeGeUGRsUj2UMZJ/AYaniWEtK
HWkldj57NCg8c47ewGECvUzD9P0IOMqnZFQ0KqdQYBetPY8c8yNaLl66cU8sY6fPBnWTVa+fBa/7
K3SeFHgaTo5S8WQT4dx2c++F2sci7THVxG0Fo5GLGqwHlFnTvto0dtTT6hvqax598ibOlKYf2dzW
q7KPbcrBnzkwYteB/I6aAgrL5IpvH8ecWREo0v/Gt9N5PybNmP0qBhvBx4xLwMfPHdhTn+qzkIUK
NBdLNldpts6EbOWC/mSCPz4zJW+QDWz7BNIlxpj0bEHxc9C+/foIuBhaaZEhkwFIOoTSrqqVBnGc
NUsuPcjnRiozZ07TmoJdWr0wX1K6wQti+DbWz3mbSdeV99sqjoiJ8xl+RHtFWuevRQ7HNfi9DNk8
Rn0v0HX4KDrrEqwqsMSx7dodLQs+BZgRqWXT8n2pufvMiccOWQNdaAsxuT7eCq2HFrP17PcV3voS
N3FlGc211tFsKDhQgOMtok6r6yuZNO0gUiI7eZgkBWAdPkQR9mTVzoMdBaqLNZQYQZTCupyTO5Ip
vQauFJmTVsTQu0gKqgij0kLXof/6a196zObuTmxo8Ds5BuAr4FHYGNF0HCipwgvaoesE2lXtPe0p
zbFpnvY7vFF7garJ8cbuE0l0uK6zOaZHsdTtczllZxc2frFuniVrg95Ay1lwDaC4Zh6B3fZz/JCq
7yLrn7+gRCKpbf+ySWokDKyOXSgNFIClHZ3CPx35gvdC8Co5nemOO/4VvmcBPrUx3dx155Y1ba2a
0ZElDyyTeV4WemRY5Wtl1Q4mJrDaFYPPLkWVyZeiYX0RTPBOCbnTa1dAMsMpNcdXrIvWMHK3M6na
dmn6pdh1DAjC9cP6cEsHe3Sd33vEewEBps1amiQLdP+uQ2lOK7tf9NYohI2wQ8RNiB7IOOtE/oAq
j1rWbFryZgC6Pk4uJp0CeBGEdFtOiiF0i13ZUkjqzaxl1M1pbxMC2oFn41njnwu4NlE+MliYj/jx
Hzg7/55ZeyxwCSxmM5FGksiD4yHIV/OfODwSDR6h5gA3t3LgeZXgbsLmcPGReRn4uLSUw7kVSaRd
uIbaQoeukEOqKKs778H2ZwLjPO3sjjYQgWw1o389dbF0Q6E5sO9Z8wFJj57Y6nAk/lKVeLs7f5QL
7+vNVdGwLeWe9lHeGndEohCP5PK4atws5zdGduivY7pKQIJBQfkkMa9qRUWuXy+u9wC3U0CW4iKC
bb26KrCDPAsmz8mxzCo3IC1uXduZw3QdPB6H5K+WbnvnOs99DmSWD6gz6Joc7e+bQNxWvNppXwZt
A966jP8zDWCXFhqMgrQSpgwxPYIW/5+GD7woGTCTlamAakhdBOA8STK04IK0wKXSmMplupqwX3VK
lDJPEBpn/NvRJaGchsNJi1gdCzF9YUdQ0LzOLDP3DeusWaMogmDOfWj+fOSgP8nbyI9o45BpidWL
k0uJaCpZlgPlbQsLOnmNSbzMQVM7/NH1ZeO1lLpxzSlLQxxlHjitELXg3oIUEE28gC6ukpnZgEVw
8D3yZD3Jotu/Gpw5WKNuiMZEGIuE6XlraQqynjMQ3LmsZGpxYkgTXheo2NZlWz67bAEBKsrZuYpx
Nz/ZO5MwiRmELPoC5F9Iwp+H6vA1alSyg+6IAQM787VT4OqWuzTkdRls+7pApyAbtIr5BP8AGX/B
MLUul7VOpvJzPpLjH3WjJjBKZceH2clZdYfOo33lawyH7VgBFy+oNGlDe5W0suLBXCd0yTn6LSBu
0b4blBQ/Yz1VY+AucrtgCCocv93MDEx88O+pDOCvDOSgqLTQ+bt53NzP8SejL2gmqEZdNerlNGSU
m3fPIUVjvMCHpG600a0ZsunNKa4spjTNLP6fmN977x2hSFt+EcLWkcJrMSpL9wDUvGQjgshqg39E
rjaT1DdEzGs9G1z0JVqF+ZPG697Wc1+guFnr7V7/USHsCQHAzyGZj1WFja/XQS5UP8hKDtPLaUsl
Q+EFnhAfiZEfO1EBnc3zOJEon35/ek6UsrJzOXtA5Z8DNHNYsp/Rpdp+0I/1/tgBSo42krCsvTO1
WGqajexGs3rjWqZrGbTglx3hYWB2aAcxxullONl/Gzoom95F1+nt8dpAT2katbAQWoapXIamzoto
L5od7socbQHCSeb0CBrFmYB29l2bnktBCmGQvvmDRdBUuSrHmNZcTD+oID3iCrO3/gUAtTY+Z4rp
nEStrDTFctnNVfQjcVBGwPR4mWxx+oJUzbzN+O99M7G0vdwM6ulOlUAqDgBWDYZeA745m7LUdbwf
GL8G6jABGsiKKU3oOyumXf2NsUScEiBTtdoupi8GArm1fZ/emn4eg1uo1dgWePosvssVDKiPNpfv
5CNkBvspHN7Igwv+G0EvF+KPYeYU/SboOGV97eSb0IHI6K39QyodS8Kn4qe0pJK1uENFSw9YroN4
kT8BsxusTXetkSAmJQKz3XTLWZGTFByJiLc/3aOO+ZDXWaw8gfIWHVisFyD6jOgoZuEoe/EoASLG
Cs10mjee1Obc1IglUVGq/gpSlcsm2yKZG1JZRxZmzblSsnhE6xj5aONY+b6g28VrSf2X+jCVEcIX
S4Nwf1cnOjJBZjsW12foyubTgWsqNNSXkjbAfryAWWZy3pIwzDHFmIsIvdnf6kGBzc0kYQAN7ymH
ecQkCRsVfr/rhCIOiNlaSynKRyjR/+fVWTCkozTrIt9xq/q/BVWyG6EDMEBI5/95aYvp2heVNRtz
ZKhDGpgOc0Fx/837MbFcs7VaLJRKs+7coZJojYCEyZgFv96LTFRuQGGARf3XaiJPA0IBmrR1qNst
KoSvCTFC3ZXdbKI9fZ7EidO+rIbXeZBJeSjDadKzKoKFyJNqRDlqpOefvQpb2y5dSokb0EMvk2ez
eDeTQfAPtqXWRqbTHvIjaO/mGAcd2HV661Hs/Xq4ChzQskDAOfT+Ghy3Kxn1rxXBVPTcR7ganOnv
xhimy2zuiZgYjEiaukja2l5DZc1D78Rk0aGia9kW2gAEe728ZfQMXTHG8iepHb7/hCwnbZFAl4lf
h629dayqqzeFAxWL4VsQ8YwnlnF0bJKAW5BpofwSKtzwoCM67ow4/hWKQZbFEaXuTi/LMz78iFkO
otKL1q1UizRKCS9sLLcVooRNQfx64ZYvc7JqbHn7aruuc+diNZyAHcHsNkPPL7ydKd236FKRLCtt
X2DaN/bPvSZGAimU6AbjQx+yUbljqRIowy5j5b3bpmvlPzLbjFht9A0a04WfF9HpYPKWI6uL1vjm
yuALrAY+6F8vfD7kQwhrNsVx0BXsel3Jp139nnoqdpzkFJMSAQHvbo73DBhzA4FBSSvHUWzJxOTL
IsHGttnW+3zA4SD47gAJvvR+4un8AaZ+ibnnNsxzZlpQ4f2iZjdGDSgjDpvGS3NvQDucX717wQGq
WWpxQdRgjCvvneaPobRrHq2+X55y7m7LqfMK0bNe49/BvF1eH9kwwaI5Ux3wl6wXa0pn6UAjNkhD
mgEt6sEvRAGRxeCxFgpjwBO4ETVyki+HfVFavIk3yX+vroXlc8fXi5d6orxLjyiOJ59sSkLAvoJN
OgmLStpZLmLhXEbBUNt7vA8erhYxg69aqy1R+6vUtEq6NWeg7iP5dkPU7Hw5hUAS9uiNqazVh0/X
5+BjcHiWynPqmbiNZXL16H7FSRTU5rCVW3ZnDXSGPyCUseT1gwFL5msqR+xPNfH/tFVAGghIjtid
T3/b3pUZHBP/3ftINlswAF7yEGsYCxF5Ul/CFEmNBiHF6O8otKI36X2ekSKFfLvqXz/WGJt5O0ca
5eflOp1WPkHSdjsUdmriDrGsjnw1xIOAw6ObStPPxyxyHXCepv523xOfGRRY4lf28Q0qEcMUqPfY
7QUECjfXwkfpeWKl1Abp75g1HGikztKvaVqzt/B8G1MzJk3Ci7uuna4z/koYH/UdUZm9dXzJ1ZZ+
xFug7MfC2qJo89QUMI+jLFVFHceccRnhA1fxxQNCSVwL25bS6gDmZkCfCkc4EtAHWv6HqxLO16cN
3P4qmPs0j3l8iKJj6hyK3bib31TGVMrZiautPw5Z+Q6FYppcbKQMKA7ddl+mfAPytarXgcbAu5fw
ndlhn3CrAGsKa4Jar1vk54IbDVSvga4fx8my0KnlyyJwWDiT6UtRYQK97v/ym9GTMOeMddtqn+/f
rSLVKMYRADqWRwNxzUrFM3rubeHU49dA1nFCQWb+sJnmDy2LYdR6mBqB4t7yRH42HuKACFRaP8l+
mdf7jnBCINo8b/mxZO00izIYTaRbGbUDENdA4isaRLiaxsvfuvgvgmVja0aUDo9XvyRSJpl+J2ri
j+k1Y3a992hKZ1sHfgf1YkOwAB3h9Tn49l6zYpKpXnSp7tEM4oLt9mR8A6J4z9F7mp5GHSuvhCSE
s4cyZ64lqrZJouPY3iFQS8saY91QHpGeGsv6M9Mq/C1wA1IW4HoZ+L2wdSiCbuaBT2y/SwpuE9cq
L5dqE2K/C4vnocB+luNun0OvsSvvXZWjdvhchK+/QXqzZRHNfZQjtlBUQ/40Oq7itxzv9xh4eFrF
sAh36tEpOVOplLlpXB9BtpbbIqbLXQQ4Z3YiXY3UHAzn+k8KRTf8wo14IUR1XgbxGPqMVED1AjAA
zAaQB5U7eE3RAZMh3BE+Zb6rPIIxHIoELt3sAHK8iyW6uL3H6UnepO9E8Rf+coLupOTGEN9obkhg
C8rZ6p4ULdoWtRGYFIy/y8vo3ncXnc5Xev7Qj8PS7edmU02GID/MjF7wbQ5nNcAKtyLvxBu9IRiC
8AES4o3IFBz0LNjs9FtOK4zUIrjJmXfNruZBrnYK+Z2LNpgVxLZvJV8duN4IWDjMIYoIBNlqaGr3
F5WM/3WBkhKhjeehhRcO8Pq9Whdz5ZIF3ybleZt32U3UQbyysz4V4I9zBMYibc81VlA7iXcohyol
m/jwOzCsWyOv7FbE0aPXE1Y47wj7+dPL+EC5ANQfYcORo5LO/9zH3cHoWlUQ53IzMLWT62FciiKm
6zRi3PKLmHWbyHKfjt93VcGPsYKQPQ1O+y83FryDYvjofZEcxFz6AnQbkHGcc5moeZ6nn1dg2UqV
r27sutyA5p9Jlx2YbTmpEWHWHo2AGK8lRn9z7POxroNAVXI96t0AipWs2m6KEoHPknkyOxCEGWd+
qvKfDki9gU+950Oznc3jYntrl1o0LOg3Go9As8gJmn1UDYS+mtos9GvxUrnfwCip+HbR2bRCPDZW
LqJolynfoGact8yS06/NsGWq0HwtD4h1WLnm+IaDrkIlqVAtSHrpfddjgdcIhy5GENtV+sJLVpRg
wduO51oYvl3voFPbAeTS994S67a2LfT+WfiG8GfIFCFX8PYBF7Juz0/NRC3rbmLmi5z0QPgoRRe0
B/WTbIQ9oXpR3UE2gcArVTP022p3lgpgoK8Wv185vhGlI4K8cyojLYVc4MZjWiVArtrvUfriZrPR
8bTWjyMi84dBSIzSExL0peUY4ThAAXfejkwdHuOTghkqf9s5NWUtMCdjIJ3ijSi8w+8G1UwThylq
AKPwHPiv6ysSYr7PS45/fEEkQvzKi7z7PKnxTIXQ/6tnAbjNKOsF1E2lC9Y/jdPp0v+BVjnnrSJC
TGKJc4BCR0lrfkYPuC0xLvGk+GqC7XeuKgzWhjIOnWhrBzvk6C3QJQUS3dT8oAw+/Yb/KX8RbsgW
OjBlezOdIkbwdqe0rFddlm8rbiX9MvxpDi9t/5gr/TFFQ30WzacCa8hH+f/AgjcWSc04VmyZf+Ma
3A9+LJ9Hp7X9rqAcktPR9AGnjBiiJNGbXLtcBt6BXtlsxkC1rcwmt5t4ywRN9sDr5xCebb5NaaHa
tqyzn3VK2DBoTh2IWEotOx8QQTL7Ix9Rye+kmTdhLyA7RjQK40hZJU+IqEPiYrOYrkkphnv2bGXP
isftvO4vDoJt6fDDttwAIm5TKOTFlSMKcqbTF4gTSTyw62Kz+dPZpCRctRooaVN4PWJ4yWTSJVeo
mkwfQezB8nyHXKFwSit1TgE7bwg5i6+kf+gyhJoHPmjbNpf+pjrW3Y11VsW7rfWkB+7/OClat4tk
KXytJCdhw2ZtaMRaZ7N62NHExS2JJhQGG3rgCSMpLse82pXYCXrOr0jrhj9AuBzWy8RnXxcHfFhD
hDvLgpZkMvyvvn/fD4lbyVze64KB+iN1+Uy/WIOu6F6uUGy/2NMnc5Yvc2A2Ne02smEqfCyVmhAi
aLGwhzaVK1gxpQDMV5SLlDq0yOhb2tTDBX0+mwSxTsUbP6FV3GVsQ5kTNpCp0rQPJ04pC9qE4Aoi
hb38g2DBkXXiQ0qIK1cbsVR2wkiVm3InJ6kTlV8Kvhd2z3fcRCgz0gFWk3IJrxczoU7HREk/XK8z
IohxSdnWZ6SBGW+0UkzU+4s8bXetMBQ262Cv2lciw9cnttVdpfIaTtTsh77TDmKa1/U/brOIQlJE
yarieHtUswCkt8PWQD1elQN5QMrXJSKo3xCKpC6VJ0KpkQh7lQycg2vdZehaDZtsyFYw+H3Udbc2
Cr/JS0xxMRGlUl58XurJZ0zFcYeHEZzXJ5eCIa2MZfg0jWCCCUBW+uCPjUNJLkYSowBPEuM6YD0k
X2dZekNgrt0h4AcEAc7iUTCi2zquRMpMNv78NgP6XO/CXJ1l0qCDPG7ThY5bGp/O45jFZvs9TECu
fmJi5w3z7jJUV+Edy1amTLKrWl/9odkmK96c7c0c2n7GnMU6oYfEEhEXAcqREv10o+O3OadmKuvo
rX6R3Zdlwx2CoH/2lYWXAmzBh46uq5hD5HzIX3oR/moHRNgNnfTQVYFsEzgZuB+2eHYCd23UAhGZ
9asW3U2XZdOLHeoSwFDO9yVtVn14W049DGXU9tduu4sgLm3M6mHtDOR7gWXR0ASe9RZHB51oSpCq
VLysEDH9hLSbOJLSdNqrdXwp+IYfVvD8n38xemkOVGTwFMhuCD30ceOZV5NjmTqJ6/aSX6t8vYY5
JY9ILC7ciDJnFVf+RLbEYoc5J52i/oeqEtU62hl4D9sWPzzpQiNmM/YyFGwdsHBL+GhkwyF55sBC
1sb8B316EHd3/g4ttE6D5F6hEKMq4vOn0wEieg/1eGXJmDzWI1hcYyGLkiynbz0UoM+XTUUiwuwP
6I18GcQOXOdB+SGvmjh7IMJyQtqZ+UuOGV2N4SBAJbNX06LsnzaZ0WTh77KGSUe2siwfbViX94J/
YKGGJCoyInmzu3dc8MbzRqhVNT4lVLtF+BdE4j1Iv4ww9EoW6uozOmJgjgEsCrwAdQX2IC+R2mwm
jbBreGTj5mp7dEH4vQeXtaDpmDSPToap4mXdC/o7j4u47UVN/S+p1YnldCWQdyD55pAD//Yivei/
vI3yAzGYGeHdI1npWXTnA/I1szWde5pWCGS6UVk4wdydUuBEL+9izZUgwB3zurzhq74jrC0vLY54
tRp2rv/80E5FN/5ptN3zuDYKRvfPoU/k8Du7lY5YhmQTwQ4H4KKoxAxqXYZWUSr8cTfcbIUtRDSP
3sNVR333qGv1x6zAKZDniiEZcSkGOxzCoo1K0q3enOxFiM0PJhUKtHzt4ZpNwCBbcLojzABfxxQB
8wAlzojXlJafHKQqIq+Vkz1bIwIKOxfgINpAg9MaaTnQJIMTqHOBBtUE64Qxg1jcj/Aun0pksc8O
rvRaR5Zab0XO4LIMivlPq2VxqBTnrdXqIOdJmkXTf2CTovPB8obB/fBnzIUAdrQJtnHPmy/PWA6S
BrU+1bYUyEFjcQnE7wdAF8cuuooaBZ44VkTLTcaJNMU/wqgGW5+Tctsruss87ll6/H17eGfpX3OC
vNdQiGboy71dID/J6SR99flDPK3N44yz83EZb9dgZwK8luTFbDMaBHKLg0l383pD03ctoXmn12Pu
Bz5BUHlHvS069+v4N2ksvQOv0g94cpSnG8y5iOjXgqtn9nWkFLClsNYFTqFquV/YkSydxK/EIu0g
qRr4dhXkZMjTn0WTx1dFBcPyhewTpg7wt2UT2r2XN47sMKCf0YjtuIqCfhBe1Ci7vKUpQEcwDtfS
/BW2hX96kHQFZGmWWrP435hq/aZ3X5ugApPPWIzT2pe9XuynVRTwyjhrlRjbvDH1ta3ECd3pYvGL
EU7ZykKpbaZuR4L1a7DJQ73X6F24SqiDRZ+n2AnADx9tAhcX8NwEy669ETKrkQGYZ91PuO4rOOPG
lfCehdwl+m0qqys+ExS8hzdiGsgqO/Z1REtFUpco+NhHWZm0aAu0+q1pRC4XTajcGDKYdKmCJL5Z
SlTvlcdaYGPzWh29RTEXejRSnCeSRDCAYH7tqyHW5zsap2cKsOKgjEuHZbFt+VPWhcdJ9OLgfZdo
N5pZ/NlYS4vwQWoPmga2Y91dvSYBRog5pOnwEcPDrT4GhpiUWKgnjop1oBrGNmG6R75xrqw7eaF0
f16/dSyM7NFhf4zWs/HVE89QjX/6V98N9SPMwqhaT3wt7jMV/GDbCgxQ6OXmwmqnHIZYpm0Wd9FA
Brl1BZCnHOKgtbBLJ5lFJeO7NMUML73lRMLFOF54T/zPDlkV81MdujqSLPRjRj5FGDmQK/o/+qwm
sdq8CkTCX3cenqF48rsOvNKtkvejNmHae4XCUGjSrr+Z45qJyTRXBgjBL5vZNjr4mg5AYoMW1fmh
iuuRN9qApVXs/aN/qaFlRBjycgZ1wi9H6Hvcy4a7XH3Hlcb702zYOd5xjUvt5E6h3Vk72wJKxQoo
fOYdX9eGDyiaK2BgvXgbnAg3aCjJegAeTnwgkrB38e2rFNY1i4xaazpsIsDednBXDm5Kuj63Xa7j
99t8AhT2fXJ4CPOs2aNPKm0iI1u4JP8jyJza+m3JdyjmdnUAYwaEd91KJEJqQ15kUgmgOCD8TrVD
j2PYTn+vanlDDAjjRaCSvbohY79+IkWta4Pf+LeIrt/ce9MYdm9gquP/FNflfvy8RvKCcCxwRkxD
NFe33wWkg1BeB5T6GYx5Z/qskxfXpk7AHqFeAlFCEFVA3Wpl7T/yWObGw9V8RUDTpyGUIZU0rpT+
Qx68SoQM9JCgTiIU2TaehdSsqXXvv7NMm1cJLIuDRHV6TbLiMx6y3J8223b8DJmGKkj8MIXL8hmV
ofK437fPh6rgypV93fwi6FojodogR8x/TJioS8SJN7VkymSWZLK084IjoUxSaV2BMYSmzyZ9vcey
3mVOBx9/8b2RzytcZFori2uE4pmYML1yh+KFLroFfpBznvvTX0RfAGorMXrZ3OsSdDgQmutXLH/g
oM9FhT6vxhWvYVxsDy9dMXpBh8/0CPYwaltNbKO5UiHvFQnjErka3pfbqRIkDbiyw23QI6mFSU8W
y2fR7B6jBWdvROx4ay0mfZ417ydSwFonkzo7Bytk4Tgy70rbE9TopePr224JojU8HpfZUvvB2FLh
UnCWHIl6/0gAGxWUZzE86YkZ2CG6ptxbjxsAlcFla95IbnvnnFnyoike/dfrf4CAxCsp9gXrE4Zm
QMX85+Bw7dTx5SLs+tWo1neGNpgILS+T3tVUtyDjB6WAewOWG72oCT+/MMVySu2fsEGWOKKeBcJm
F2yAO8JjpTDglv21/XAlVaJUfoEKY1zv9unHaXQIRNx98vMyo+LHe8WYG/dCWo0HZcaz8eCwsiSN
mneuYExSHb0cKKjMYty1W0EWTzchTiMu7+aArA+4xOPIUgvB9KLechrTGYQsawl95fUYOgrRCjgX
8TLi+/W61k2uHNoZdCfZE3oWVrbdec0lXMlfCPyfXT+IiqRI3glIy/fhaH7fxOqSaDwHIh0vCS0M
MIDW2505F6SUh3P1v3Bad5fL3I+RaCRa/6IaYawtSgEgjQ4I1whpGE+reZR5RpmJhTdPlV5cyA70
7y2QwiHfxSvx/jrXAbNhQslRvxtUqXrwICL1Ryvky8/CBBj9IzMXLG2X2jOAld9PYM5eHlbUW0dF
zC4RKX2L5pTmzCbEmqE0W9KdZfbxmpcriFcYUadPqKZxFP0NNokKEgSGzflzUd/EAwdsHT6mRTvc
G0o2tmE1YLbDUPNFyjnILLQOc+b+x3vc+AO4qZwnK2Amy2xIXtcvLd8xTBQqgqZ/q9rIbOo0K2l1
RAmfPOpSCe0qj5c+TQi44YTNatr5kDwXRwlpVtOQkvV/YOkUGqIcg0DsYd5AjzSCMtB3gHmYMoBp
c3x/Sy5q/ajJQi25zQzUTjuObdbA7zraDzmjaZk52B7xxGcrNVl/Gti9JytpKGzgnovMQn3mnwKK
2wHU9lAF4F1ur15H/CEoNbhysxgVRuVumvzTwytRyTjbLkRcS2PpzRcObBfX1twPVauuu5pO6SYM
/wUet1T2wJtGHxsBZ9fURjsGw3sAQ4OhOD2V2whruLQi3GbauDIEpAk+KSmBcmmIRwAoXXmpwDY/
sZAtkZ4Lgd+xKLUBmqkxOZrXQ9kjPhEx7oPyyAOxaKxyqKGD5WzFCtvvu2qPADn2LIFd//xZFzK4
vnSBzwbRlJ/YGCIEz+Z8qgf+3x0KkuabL0Z3mY/z0PAn7eLo4qmbBPkPqJ9ANKViT76p01cqqZgN
vH7mNN90hSvVMb4+a7DJ7D22OrF4yDbSqvXRG8m7vMBsm8MQZXLVKfO3bLCiatyXiWdriV6ykif4
WhYBSwKJiagmz/zHi96kJEyrMSYIdv+G9ziwVzfXOLJo/cJlA8E32tL9afNj1B53B3TYLwXMUAYB
HXCiHUMGh+hiBZl/ccIhsQx3fz9/AazIE/Bpif4hbL43E4j0bUcostO0cgpsHM/Hx0bHE4slAgQY
2Q7DQ2fsvXl0wIeSxvnmTC8ApyLa3CPNhogvSH6oLyHiUUngicazk33OJ6V/hjsZY8PsVZID9lXd
/rpEBm5hHaEscCconPObsTlqqd0gW5juGXpjZHpxyJpqnF6qDQ8zMVNP3c32+oP0rJH/pzqhwhJy
Q67mixcWbVrILirug4pnD4bgrMbAMWw6Rw5BHgMUsXHEbjE8LSKG7G+XVTN5fVVdEHUlU+4u0UFF
zOe/npSI5pHv9B/zBCe7X+JudKfI3/of4HVaA8haVL9KZx/Wvxhc4piEKddvONSyYnSf8O5V5moN
SxHS9e6CXHu+dKGZfXO4JaizBfaS14FAsjUviJhvnRtsxlmeKxYo9XmWTU9bXVsazL0X/U3jjOH4
E1xkIidBvDyFlo4d2lgtlUcbYOk22bzyWzyNhYtPzrJ3ti2ghwNpYGyN68RaZ1EocgOL75rnZAWH
pucr8vFM3vFVSb9DBCzn0IP2b4nuIY1obRC8mjfAaQ97tPahfsqJZ8naCXSVHrCAKsjDU58UmXim
la36sZjG1YtOBigysvPHzTg4DlhqMMJAytyN46SGAOLupuIS9D8lSoZD3G6YfC2fDEjIRWVy3AiF
uRG14hvYm2hVPr6805OX0NSgWDn6l5D0IA00tx/ZaiXEsT5LrddUiZEqfxYKN/UknhRnGmZT9Thj
w6/3UNIjj14+sZr79NtOMXbikaM2OelfEr6jm9UdreFaLzeTCfvS6qk0e/Lm10qS94zmaY92rbL3
j3MqqJQOWT4a57wOslBICTRHjGCC31OmCSNIYLqtUBRe5H4eco3TgLlImcKvoTfJMoBAvlXxGp2b
C88wTy9+rlHqmCY9YFQFaEdDbQPkBkmZHdcRlCThc0tx7yorayDcpzjUzSLLJ3HSJtw0dFoMWSFt
kV4erTj7nOxSQ+XBePfFXzn4Xjsg7PSV7e639t+ELRfX9JQRfpl2ahsW0st7Ww4I7EnPQQ4iqOkw
+64PqyFZDkd89pZt1WdzdkQBMesEoKFuNifQmuDHQxZFT8wnerNGc6SpF9gKQpDQbUPiiGRIMHxA
EDoJDAjkiyJmwWGrzx78iwOiw2FJwWOGUOSgR6iGWpF+cvtzvzxQbV2B2MlWSk8ZGtYbwdmHvHbp
txJgDgUVibvVb5nhZid5/V7oCT03dgX5sPM3cdnXnydcw0KUwIBUcj3+hGyObdpfsHPKI9+9hTmg
povlrdNau5eTPqB/MeSjinBeqN2Rr7JB2HquUOppO1Y8JY8HOg/ukXyxVaA0mkPi5HmaOFex9MmG
LVYLggpxGHKt5KBkIdFtz383/GQvqRjuvcsrJ/e9oGp9jj/rQoagbXr3R8/budYDol6KXwPuWohZ
eG5RdZuzhsv2rQ9PE+/28FWNMUlhOCcpOc5wT5pWhDjeWvnjHwZW8uXV54908YQnBIqWX5NWJrCW
rDk9TepXBWey4CW5LLkaQV6mZiCWZvdc7xPHCAdeQIuuoWfH3+2fNMrF+qJhXg+pJxrKmLJZP2a7
UMWjuSrTVV8RDfm/1BOEefArkYluB1nH7gWzhUvEp4vwU6V/Xg+hhqQO+qwDxUCrPL2RODDyvzsP
oSExCyWIyUe1/SAgkd53ItZYVZJlQjRtb25tD4eb5Wdc2I/Q8ROjSexzUuQZnuoAFzszBsdZBRev
a6rntP3K4rPyy7QqlMYKCiVrfX+5lhzCopXE4hNZ1srC41Cb254qeeFqkm8qtDQWdmAyc8fLggC+
JFEgS/7RBuK1USQNIZox2ih57Kecdkm4We2Zj04Ho42huqemYqThVJFJa9HJH4uJAVu9s3pJMwe1
0w6vbnYduLDrZsTpsf0rI0EYand78KbUEb+nbn7n4rZm0pmwHKvltHOFP+c4DqIT+L5FsFnJnvw5
vGBrgqAcHjFbSZb7f5LCuOfS3owuLRy4QkX/ESe+j3HIO21CPF4PW8VGDdkcjY3WdKh/PUgR1VM6
Iau48umBQB4YFMUrCxNNAAqNfD6M6wg5a5PEDlXNQJG9eKbkLKIdupAqknt1WaN9XyCEQSZj2YVe
zm9A23wCBZaWoME5ixlLlbUou1SdXBK3NfcCTuvKe6wRCAZnbAMklhBmAo1xGcDcKU9YWGFp1dIq
Y8ljl9i4fVmkOjxARSSiPzkP8KMu7rA77hgAYC8Br6ahL6XpYZbuh1Wv2gquvoQ6bHNyv3yClhNq
QQRDd22BuWVwnZI/XLbYsQK9dFQoqeQ/gQAHrNKhD4U0cQai/T9c8U42FmOOUtx8UHDzXPZ1NOCt
wAB5My9ExUwKFby1tdmZ7fQ0kGZFWa8Q8aThBBKFWgb6VG7pEyuAxNz9eNSlQ1np+Phrgr37yMzO
rreF+OScd0LfRvJC7rEexxhl0S+qlx+byYNYQAtn8E5H/2DN3nHglZTWTQPay1Y/IRaSj7RouY8x
dPg+r3XNuQAaUq3IEBEmVbvWcSdVxGbMH+KH82m4JAyTiCHRhsHatcMxXl1moYK8u88SbeM8Dwqq
WdL1btHJfXXeDrO9FKjMHPxm1WAT8+LkMGurm1BO7sSmNillik99BBJ5IUhs4s1OOMKodY3OU0aY
K0zH0MZAsXSf2bvsmvFdjA/lhanuNpHscC1vmearp5mRhsFD9/uUfM4uMrGNqbRNA5Kjbz7Tw90N
ogjbmvzxssnwW2FCTBTwsqMn7KMDQ5vwWfKmeUzDt5t4+OjfIoqo33ry4pILPDrhfgk2JPEmOTca
ePYbrmLCXDal6ISxPeYF+gBTeJfWljgO3M0uokPGqrhGrLWsR6iSbeh7kE/MrHWwBEdDZDk5hENW
iMpQfQsDL3boY0XDXL3Mc6nxFzdtvW9r7iycSq/DIPLh4BYb3FBI6bXrKtl9ZAXJzm6O4g3HyUEC
qy9nJXyBtycIV6SoU0WhE93X3gxZ/tjMBlxI3/Jz6ls+9+dRNZIymcPmvr/tdwf85HY34APqsmdU
5iyF5b1ivtjeNj2NNHPrKnluLIijpL4HICAs9guGoYflWPRZBusyFS8UrAj390z5ro4RNoB4sE+Q
/6shWSGY6oVRC/Sw+fsrV14YcLeeJDe506o/R+pt0hzfvqZFcDC1gRhXfXBAS3F3ZBl5/58nK+mh
YaZz/kLbi+PSoz9CQgSEcgqcC5eLX2rwRRIL/Thwt9oXJ9C/vXPQyH9ReKRFFAXaq3ZG1m8V4L8B
cat6YPyL9R2fI52qtraCSYltQC56KXYfaNZGKJqvW+hDG1CoLi+8blKh2p/ZXO6orLxQAJbZeFTh
laLKzea2JmvFEdNBLRvxSepOaq8547JrlA2UXED2+v2G4QI3PpY4P+R98hAAnd9rlgmCxkfAyL0j
3HMYlITywJbSlX4BSfWv64eQCcJVNN/R1PL0CSnyzVi71emhC0RWVXNKeg8Niz0YyofE2iKr0ymb
uf11vfujady8Y9G7DQfR7prWatHjdsaapJwFMwZ8OrwQw7Bm3OJsOm2tTKyLn09TdP7iF4UAlqoI
MoDVdmuX4ueQ1+yiS8kwxjHjzrqu1EifrPs0aCMMrKyLzLo5R+34jr+n6dJ3p+FB5s6kiwgjjZCs
rAYzJt/O/r+8UaRl3zVvO2uUV7zF0T97QAiiAR8LuhFKREw7WTvosw6fJ0NhN4QNjcpL81Z560x5
iOJfro73UkPvNiEE/awpJ74KZXbfH0B1M+U9bRRx9MtoKPZR2E6cWJONDoG0ngg7JAqN/HsZ4qJ4
++97t0C8Unylz6mfAWwSmByrTt6ZeTgg6z9ZQ+qLkNXmjZSpJsAmcBA2GsfsRu/1zJ/+bTIFRBoA
YYmDBfgZ7N2sajULVLw2QkpeabWvbhwUmbyd6TlBaLtKSLGQ7po1DatL0/taP+T5bUa5Efts1FiT
gjHKbeU/ub56l4MGH8SkuXCm5p+7uGA7gcDdFSeYFnpRZy5mxW+kShCYX3W/t7VbHNBaGMR/y2PE
qO1lo4CLcX1YZVNXNlISl+k1kl9VLmQpSdvsRpE12+JUaFm8FdV2Ic4BpV/W5X0Zc5sSZOrC1AfL
jCn3iH9ZkfcNKCTYgzG7DkASvewkkikXwUbUygqRQQYCrf6j+JvQnAIFBs7NmKyB95WxvdSkHD6V
5WO2NfGjFivOYhrPcqZ0opEB1Q0lkfgZ8DxSNvLHvH27TXfJNvtIH5DEbiJ/zVxR1mA8bGTXm3T3
IOy2/brHfu8Bgf2c3+FZieZuj9ikxWCezNtpGkbmAZOgyKdZHKw2BvNFmPeMmn8wd2P5tWvl9byd
XCxiq4taekL38g0LX0oqcfzmVIOll4s4BBY4o6S5xNEvj8nVCHr66jUXcAb3XMGi6S0a5pFL1DL7
N3ow1NzpFKoWLnN7KK87yMQXnB7HkrPEugXJ0b9O9DyuW0SVKMZeeZs2t77Afmj79iQ7PPmGjjwH
zcQVcSdnYeseCZNhiS6tB6bM4SPuETYoIa+lmnfRlv0QbqOTewNWq+TRC8EXe4ZYFLgTq6Fx5+XQ
foLPb9b0fxOnkCLFz67RyR0rudI+n6vW0c85qnLmG9YMJxme60AqH5nerq7IJ9BMmcJkTtEd/2Ug
ikomYxe5mdiQm4amNtOlyBdAKN28VlHKS7grcrG+D27vY/B3qtMRNNhnmMlZurToEeGfUF2oaPFQ
D23PNVq+hCTUW3sdl+ibrgfSLvQGDexwds83+ORLAIIWEDdQe94nkwqAFJ3Y0m7TgI17dVE0DV/D
EiigGEmUk/U16YOg/mujr31MiGQhyx0a6WMgUfTfAk5ksrryEI/U6sI98wVEnLt3XSlQIV5wnTHW
bgiOxq0hxMOoR9vPsMEz2h9KVOiLf7oxEgd9Q1EROV3rs5q76T0IHRtY4lvFDL11jWvYvuwFJC3A
t/drON95vu+lIahTAVVyrnZeBSDw5mCW3QHqnElreGmtoWwuBgh3Dtidnf2nXuTeMg4s1An91qMQ
8QMDzCceNUoxntjPByk91sEFpoN+Qt27dAuSJcaY9eihZs5xH+x5amR2GvM4b5LY57i5bfDAjmG6
TQXXZ8Hrr515D7mcbdG/L69iCtvvuVU6k7HQUbOrKPHjCTneVXtCSyXmdXP3pNlpZnSWC2+9CT7N
lgt5lwI4MNLr27vtNKGDYt+oyDqq5Bp/SAOvOtBrmGvagRmxcnjrG/oNMKPQfniqOE6fxF6ZNG9H
ckCZpHwCox44ppQINh/ZyUxWWKWv01JnGZeAkb3PTfxr01S+bJ6An1secOF7Bl5FNhBSkDn1ptM7
6atpdc0fZNoWetAKxzj3WE+tWlU3mPc71mcaIC4Hp8cUMKNPx9WMfZGIX1YoO6Jw5CmCeP+0tOCo
pYOmpOcyZN1S22gHAdYivdlPvF9iPRS4fm7lAMaCb1RRrfJqqDjxyD2yAkByPKjk7xnjaE1N2wvX
Ry1NKJ+AuGi/Cm4N1+KmxB495BDHOhRe+HQsvSmi9VozIf2cWLZ+3JryioO27KwqBxSIi0OmIrHe
KuIAqOWem4joPatc98K49hAMCosGOA985YxKlb4hvYLlpX3YHGfkIdU2z/cHDUTspi9QFokYvB2W
r6xjV5w/jj6OA/Th5WhLMbM3rfMWOMymKxoMWsLli/nef+hpJ2CB07B5PW1c2DsSXkdtWibdAw3F
eTY+fF7Jqai7qw5lUHzeOsKrCF6JSFQ956v/KsbUxe4JvHnqGk7pSUTvDy9dwUvDis4d1yZ/cmM0
KZVgj7zA+UF/kmvZeGNKyc22U4o9fHxiP2CFZ2exkaChArBFd/U/2fWaWkN1DlRCL/wUw5YA7hkc
ZYhO9crjORMEzRx5yW6r1zLyqbnjKUOLzY5h6j/2Ww0VZu5mcErAXJKjgwtaJx4OgkmxEYxjkTdn
WxYxRUQfT3ylgmOQCYBjcKIHq/RkjJPnxBo8Ynw++bt3chsS7YpY7g7GiQtn4jG7ohAUvbrq4+TF
xUOVY8sH/mPzfJBRNXMd8qt8l2vugARxq2aU0N4LAEeAEN+M5mQlQozLbI+tS7UavZOowvpfCVSP
QJxajqEn95mAYz20Q6B6LX36GLEQIT/FJhv/ex3iO0xhnizERvkjukZa9om1lYtFUSfySJ4sdPRb
Van4t0ARNJtGnMOmcnPeODG7sJrk9OGzmBKWquh1T5pKXrGHUjICl7pQkm3c2xZmIYIQxbwQc9Ud
xFmiNPryJHoEgcfutRSwvdmVM9DF1TNTaw9ZUSHO0EpIP2IWlfI1a0qpy+TLvzShk06L1je+S2b0
TISx/yF3xxa46O6f9WgWagIcp3XJH+85D5OqDbOZftsR59U3xju/1qk/ij+JtK4GOKNEx2OrKh9C
yfcXFq16o9dG2WYBZ4oTgF242IKtkbxRRqwIJ+o+w55uup2bDJtxekYPZCAIKKxIK7pWZV1kX54V
LQNmRl6qi4WHVWFKk1HdZZsB9q9l6+Ha8xAD/f75/U1zAqF+o+CoQxfwe88vZyCFPLCNTzP7JZme
UrmSe3nPkqLzH3Kk9sO8r8siGGVq42d7y5EzK80/3RwgFjrOTEmjr+t10LzkAWC2seV3PNvPZNm+
N9CJBg6sfmG6ATlG2nbDQieA9PeMgVlpV3yeRz90RK1q6zazyAun9y8czmvGIGskjKSEAsdbOS6X
HZ+smJ2vwNjf2m4ehEqwIx7LtOH9Nn5VE5O4ERsrc6IyijhE4pJ9lPXK5CR+FiqC7rguDfE/MLoM
wVDj59l+oE5ROB1FXbn5O+rjYm046g/Ze/YHfFcdhy14EGZtk9gxsfAkd3B+WM0R5Rw80UMWHSmU
BY5j8jahyeLtCpc157n6xvz08uYz3F+hbowJEkT5GwW6NPiODyP+CJPeyFyFoXnAyZUYXqDeNosz
19ZuBxaLBqZAozdoG8rWUawpGEYiVwfcQpUzr4WzCvjgd0Y1E4sWT7R6ysuKuoQ/8tYuuTumBcmq
782oQWLCVyQ7RFfoqvUJgz8ryt1G2ec85OM2IBBGDEbuSDYaFfD17NYn9FrZv7BOgC1Z18ZOiOuj
CEEWPh5Z2H3isHoRVmxEClaaRmRZagTXnWvhY0dzrN3yN3m/E6Q98ruAUdMbsg6aT0In0D25uDH4
wEr/srxwVpuEeIsvIr5chFBlQmuilQSRDG6g2Y1DMqUqjSXmW6wTRUDnEtX0tBFhgXMs3zUQWNeU
DaHAisBx668sTSDlcED29Cfrmnq87HHI9UUUPdZPhCPeVMW7EwH4tCyaSjsXRLM9ZZ+cYY9DoUJP
vEfNPTqWwUW38WApoCfiQm/v8/B+A9kNGERlnN7g4/XLeAsCuE2aruCUbIfujvX9ClQfVm4RAY/V
32qrjp9CYCvkPV2XaaYlbwWMVNmOEwdZSnBZdUN3xkSbe3RUVjRA29EKEaxtInFVx1bEFs9zEdVM
EFBGBOC1R+0ZNHQDLlkoE3bJbK1IGYBvvvEl8zuCoEeOKD4R58aKsBVCNQ7LIhhH/v9B5D29pqGT
qn4fqILxDPqRVYYKtF2prdsK1TtizVsxUG8Gqu8MGBGwA3OHNhZ/3hFf8sO+ix03FfsPLXpm8PB/
2xP+sL7prxwYpa5zNGS6pO51AdOBuHxp1DU0LZ/Rh/Wfk7rb4gAYW4dwkSEoe0ykHw+7YsPPudC2
eueb5HYfn1KSzJ3apSQMHq/2YAega4d3ZyDMlS98stN6vsZgCa8DkIvRUhxU6PQniTubrJpt+5jT
lNxzmjHyzDnYMq/OecrhvzOA/CUfo66ju9cAi1Zgj2EjQ+QpJndpWhmXPJaZPylwsghBRUk0oQeq
OWvt88xCQ8TpInzazjT1CnlWK+aU5u7fWhptkFXkSp7hFI3hKIM/tMVzQTckhAmq3eCswrmW+Rxd
ZVzgwDx4Z1pLbYDxQtZYfahNi+cHhfhbFnNX8DffUc5oBEggO+cU/h99SN6ts1wiPOfWR1eD8FXd
IpjBtUvFTQ20hq7FUl15vGSMjeqhyjIeQccGO9e7+62Cib+DE2F2CW11yQpHRCdvolMFMtvcD1G+
l1cM9Y7/mK6y8Il9dYjCThAIOwmJtIGquaQgA0uR8XDRhvOE+1NeYB+tsL9Kx2uLEqEYuFUDBBW3
xATMkeXVrZxn4+LcCVe5Ztj9/GqgwEoRZbEIW1WdJ6eoif71i4m9/elWOq4I257zHT+DutI6wIGB
namTuLhyaDm6oEHfvMXaZkQpbxumuOhZMIb9mXShpHfWl7RAI6J2DRdtXWsdYuAP8Bo3t+G91+s8
DnzquVSqNmJd0CYSdSdMPVVnjCy6P4uiqUoAZqVGcMrMu5CtgtideQuULqRrtRoP99MwgbNvzH8s
jepbL5n2MtvebvqQ+dnRj3o9EkiaW1kene0FAa5nsTT9Dj5fzMXLuUnPGa4pzzaW/qFGnVrXuB1G
zAyMe/9tpJ+3kPdZv8X+ljKWZR41ex6C5OIgx7p7+beBxmrFZHXUfY++7OdeMe3I2RtcaIr9dAEy
PLjKdISgDDIdcdYVIL30/iIMTM9xG2cwI+RAWNpIFGw/LpfMvyuVb97jW0I5oyvavZ49PvfrP+CF
gpbn/chOwz8aSaIJbZis4L5QsgknboE2J80D/c6fmVdYJ9PNvrhdWiZ/g4YM41Ep8xCNOn17K7HK
KmqzHFI4K2MUUdcXOUrbKOAiSVV5eLIvhVVtYlW9QT3oBtl+K+sLVutZpfkjioFvNy3KcxffAgEd
2voedq/AjLcQdEqUSF/mk42yguldY04jlwUk5M+fA04Db8Tr0nALLQqskE4+4SSJwFkMsmPNPOJh
gXssRbc3CnSsE225xxfr22RWwgRMk3c7lmkIdsf/Wwj8F4D8Y89rlIfNbpK9cHCichy8y7RcVDbD
Y7uu3mf8X1pNKQ9RkMggOGf3KUP0GtoL3HWN4gf21MEEMSkz62n09b1JO9wEwlBWzDPwYSgWtSPr
F6lm74zLEDy41xzzBlLiG0ExDJMx4mUa90EZBOZsmC+PeFtmvc6PS2oqsusDgLzcvrhQndRTjQ/4
2h2NCZs1JBiO8YtdbuwV2XQiCI1t06A84GTqRQdOMs1ZC8GJj/QHadxXIX8rRT4sRkA1xdpaQQWa
LBh9aK8+NW5Kp5JFGPbG7lbz0IpKI0Tj35IBXA8aw12UoitleuWJKNPb8y8K3mJc/FwWTnA5nLno
Uad0ZV6I0pfGVWvegVyw1LH0gxY8TwEzot1fRb+clHJLtCNm9x9DLAkot0wIwMrI/h5RKTQwbfTf
OYyKL8ZPW0JKIfy8jMMeeKSpJxhFf7Fufw49H1myO83LD8qNlhYujdCOTJdVSkpfPNsVyn+cgdR8
q72EPwTTJfwvhB3zmMsKn8MLsISiUbLWS2gjgozjkNkYGA6Vn5wKOnl3ZRD02U1XKb+PFyo6viAj
FaJlKdT8s0DQpnr773o2vnXy6x7TNb9qU6jqIuMdrXz0+TsuIycEMxDf0uxU95VAdoRaZE1KXrVb
EKjwpf6pOmWAiUh86VgG0zksPL1eo/S8J4mzZr5SUld3J5Bl4oKzEwYlgfnYLGq9aTZrSI7ETDMJ
s1Lo5TRto5W4tBXkVDBl3q3hrAeT9yMGEbrx3DIzEuvh2Z1286J/87stzt/x2pSqwyJ6aOpLfGEs
w8IDER25D0DXndHcABKYWkAtJJkM1Yu23AYAFUBVQ3R/eGJ6NMTeWn3IKx5cAMmOW5MRvGWLKhm7
uTIBu0P1VSwr2qe+w8Q0f8tnRI/JjC/pPdyrcTJcqly4d8K3WV51P/yM/JA8RWrmz8lyTBUmaw2G
tXyXGzsj0QLUlmPzsa7v3Uoig+lS2ezS3Sb3HgyquNIqdTJvIWd1RMKMW+HHfQuf1eZja4stskYb
+ffGXQPZsy2kgIdoKBXW4QvCORUKsaGMOwU0Pk0sB2F89cujZZXLRtB5TsSM41zHjlWM9AEtXYRD
Zy+tKli4F7tZjF9wzGzNoFdwNhFiPBp0BK1oFSlwhkV1MGIe35A/DIUqbw52ZoZZlXGg9+7VhMkO
uMYW3vd8oMHxmRDA1M4KTYhOakrMA+nBTcDFulgq8A8yCuOUWJmyJ96tt/D5g+xnejptO1fmsSgW
85SsSwXJSmaf6QAe8gAYc6Z4EwAWdy1WPyVCALFaCGANNb6RmGfqEx1xlj2+0wXHgCu5rkOSXSLr
MjKVQrAVmjJDoYTkU2aY4CHZVp0jqSZ0LXhnFX/PuHvx5RVj4bwYi6l2YYvFU0A9yGolN2/SkspX
pFyC0GPZJMa6/UAIrhrhTugpaQLdc636LaLbzFgQ2KKhXIWgJeYc9jNf8tCdLldzopmf3u7HGENu
/1nJeXfUAdnA3h1/eoolKPduPxF4Pq5nEN7PYSzrzB+ntdg11KwZhEj4IILxeeLUwulQV50qNBrh
zzH2YiEt5DMTya7HZ+gocpcyhDuLsKwknIUY2nYEnxZo4RoEWtRZp+TQ09wZ5b6Hgw1QPZXnpTDy
2c9SxvjPjzxfXY1szOZxfTwwqm2pWfUcb5K7X8zxvVPw+Pi4BF0wnsRMa6DRMs9NKgnYZkFkO28h
hD36V3idn+sm4FE/P4UBhrzdLHL7Rs+tnB334vOEtXHPyUot5gNunbg29hLIRY+q5M8mnCP1S9lG
opqX1dye9sOtyhj3v8cUp8cHzbArEHgyM5TSIkACNwUCk3HTle+d4zD6PsasHydtRxrkJ91XuTK2
5/9+UHNw9Hpy4udzInyPNUC8vIbLEqdtmL5GzJpwgaYmCbqBQmJfRgtS1O9RbcRAG5DmxrmmoVX8
/fAr/O0s25jy92erIv92yQXnoHowvwiOz9z0yGBbW3ftk7BxUYq9lqDZZLksfLAzy9vdp+fxQdBX
nBbyCZmd5ceBybN5wKXwoSVTNKiHRO5IfkL1w2kzv4QaTgkfMl4DvYbO+AHOXieThapBhkzMxcEi
nbWzd/Y9k4KwS5AUbapg8U79UDCQoLXF73aZxGaVKpnqU1kG9QAbfjSMbF/2CbkooJxUck1gE7L5
Xs+dpTkRYc1Kh1+ZrhYUNokWF1U/BQChIzGn7sTo1OAoUx7FSa9Y1DW6tEsTi93UO/2LaX/w8APP
pjr6WYVD/nI93pJcncxbtAYBmZe5vvE3acF62QwVYV0jDtcZ8qaBlHeV09G3ov4OdIhFz+MGq2Jg
wDqhigpjupEYXwc4GCfgKpDiyvkvqUDtJuTHCwYMZLc49/fz0o851B+tajlNptRGjXbud1O7VdUe
EaJTXTxO2Ly97aVZ36jZdOG8A6AEAgChGAsyU4iaMJtmfMXZGSL3sDZI7rzA1bAkUGSm+96KqeCy
hVHvfTtWNL/5USW34HqrMGssKzow/L8eL5D0SScBbDhpXeXf/j38hhz9m4M/GMfsOKloUFls3KY2
/L+0wTsQJIqMGU4zWlih97qjukanpNd7MZHOM0QCKyeWjAGvD9OxVuQbksbbkH1aViL0ruWql4nI
dPSWeyzxnQNGVKuZuAJuEEG9g82uYIP5OIhBtLiat3s9s63B0C1PKupXv5T9+Kl5cGgmOoI4WYsY
+csioNjjhpRuJmSaIU9iQb3Xk2SyZpU8yclsg4NPFrtE1W8DQ1Gb5skYMcCbbCdeecwYJYCjK/ec
j98jXF2UGTnNVwGZP56JArBuRmrWFS82CLsW64MBgVe7lzawjKB8sRwigO9zOqicm1Gd2eX/CL3H
5GboikH61DkXFBrAjMmWlhtjelJrGJQ3lW0OnXBYkN+ZI/tU8y4NixAz3WFFmuZQx0v20woywO85
po7r+kCMX6Eus+J4uLIubxnO1ry+yLT+NEEYsxVd4uAPoJWVES40jLg3yXuAanub57t/XzSKUROm
m1GLrqK/O8vnBvoE8kMyq8Q3ZPlKi8uQI46Tn5EfLzMAjL375ONOruqDSPhpLDqIRnEbGVvvKXhC
w3mDv7nQBI1QQTMgE0EiQzxsnUuBXZhLHqZ3evasi+x3QCv9iYUvzAboqyNB5XZkOqc6Pgx/1Ale
WCYIlHkdW0Nr7IgikWG13RF6vUT2AuhetbpsSNnvryQbsHZt0IWJVSmLUPX2ptIYQE4ptK3oWCqX
28/PB7rxHuhDe16RqhxfsLahzYPPH9XMfJfPaQeNpxQFQDK1gyi2LLBwmtCia4+bLfPOc15qVv0I
f72g/5KqCgxdSmlfCSFCSZhX+M/7N3LR3Ed3hykz5NKrf/NLaEt9FUaIlCjUHyHk/5sCTevYZ0yk
Hg1ikjER3dnKlAk6LteakliCjQ3v0rEs9IKKOkR/C9zys/1K7+n9wMnxRgjZuZMDKQu4G1wO2TKq
n/B8IulH8jZKu46/w+PtLRutc4ojfjwAMNauHaVJHdIIDFXCa6YQzyzuy9ZSlEIyelXdL0m/JINm
JAoXWIJIu7rY4rHKOoIKsvbyTDuew1DUxdORB6lP6ocVc3zoJgqvVzvuzWm2hoZiLUeZhrDL9Tki
2v1sLbvQhr/b/cvDGkto6r6UYm7TjRFaUW+BIrnIXU2uLpKqOR5J/2D4zx2/q/T6agVDQzhS+6WY
Hk/XlVWZMRKo3Du0x3KEk0DhLthEm2868Vu9cB6cj8TU9JulvcagPuUS5gSMroXLJ8jzF+Uh9fIf
lwtcqvHjZFzzYlh5rB5YEXjH8E7QbpqesjTSSAy3+cSpt3vNXkgbu6zej0hh9INhkjCS6NJmdu4q
MzqwvDjknE1gkDtyF5VSXQPNAHzhzjoRNPqi9RFPyk8cLvFKiVIYLppceKENWVQA5OC1C0DxyphR
XglnjHIUMbcHUJXnGMEgC2bGEdF9PAFjFw9yFV989PixZvbVSly7lcZd+HpxLzsNJn4hJECToZ1t
d+9holhF8OJia3toN0XDFQkAsBcK3oiRHDHtrOLNIPweGgIjaFhU7b0zaMtLf+8MzlV5JZA0hYcu
T3JR9OIMCxZGFnpkBeZQBwK17YdPAcUrS1xzQRwlZPCc7prd7S/N9z5yoyjbyovUSV5YknafIu7K
f/y4JMHE6xp5dF4HZC9DURnmRjtk5KYmgDPgg9AW0QiHZdStP5GQorpBTLyk9MxrvXVKBLI5DWUn
nf8WFKOpfoSKTnsUQdQ5f8mwzNarqYGnOQVwqtUDF3MGnYJ3bp/YekkjxPgK1PCI91MnvkRz+1DD
r7g2EoTy0HRFNOAwM/8/a8lkYf6S4bzHrZHh8LGGDiJO9WH06SaMt7mI0N36HkQvhV+lPGcX8WxL
QUtf9shaIfTSPevJZwVGqETf4t3KtmWSIexwuQOl52Zfu7cqjONJOw/0RNUEKyXgXTRc9Th1RIyK
N9wKetfZzMm/x/qITWNbmirzDe7hDZ+Ro0x1VPf8Zqjs8p5ebR8d0FsTt8aJK0v87ns/hNd4h1BA
1oFgcZmTrQEbkUAlwQD7sYJl45B1RXbGOhkWAYFJqF8+DsLlxTnvH3ZUmKml1z1ckYuaXXc4QAZV
A+ta9KARJ4Aogj3rc3AEEak8zN30yN3PanNpRS3GilY4/odUKr0hzqOBc4XHtVuX93IFy+8oeS/j
oqvtQz0xI2So+IXIxgVFJDI7UEhIb2u+ZffL8PUrdVuwGDNr1FUcJrrKunFkwBHmFnPEL+1i1ZjY
g9/gvfEP80I1w8P20fUwWKgVWpEdUY/9kbCbtzbt3CWZFitMEp3m/90zBdFiJtBBq2TMYoxDyWPW
3Y/gYQU9l17blwKOgFDC0wuHbVdjY2oy8bba4+Qg7TB9brku0CmkJ1QZMVzUICADUNECXKQ4vbpX
1P1baaAoE+PGzFI8raP6jwJBoxRGaonWlVcsHGzWLqKQtxusoeCImMGD4+aFoeAdSv6zVcPJDxiy
F22EIGzJtNdMDsZchjwHz7NzRMcn6taxvfcM7y/PAXCosIffrlSQ8AMF3HcIHdw8m/+Yfzf3BtLI
8q4qIMqT0PS/r19TLNneROvAsPPBWkc88wlW0rTBzlnVG13n7kLq/zMjdPeXIco7gAstdBMlusef
DTmg9YHUB2+6Fp+3Sl2Fb8gGyKPbLf+jjFvdsH8fPO7/p514BaL17xgMSIkUQy2ot2DtJ5zYJgrU
PLYhd89ZRKS0GYR86DE7ulei0pktIpr9jHBrCNZEgEb8DZRDpxHde7y1/9Nz7PoIwgXKjZapOp6I
NL2qHwEY41LVsjTZJ2fT6S0OCm1fFHUoG3vlbOprlf82Tjhc7fsDYPzyPGbI2wltuoPC0p4JIcVw
iPOcKOc97hDVAj940FIFuJdIzXz1nXNKzDZn4K1QVu3f4MWJd+EWLpfbvlKVUaMAVgD81J/1ZO47
DoKdAdmXrRc/518eyaSNF8h/NuNX9pNZrT7KCSMurSRdH+2B8xC2K6h6AnlF8r3vDUc2+k9UbI0R
OwhDby5vRNOlRSkNAUHxWgB0L3W72aSLKdNJWVwK+3hav56yPkpKYTfj/Atbm2E4xe6CRoIMcHmX
F7S3K7TheLivJjvoFkYEosuOHG8F+tx4p/W73sFV4Ua3HGDZpuTJBtx/pONN/mRDGy2wYkNQFXBo
thYWGzjTgCOLGlQSL+2Z1aZkcgEmetxmAffeDvMXDcRZzPSWELqgI9eAXzzWMLzI0OattwGQbP13
sj2YWGgprwKvfaouWmqqWbmgELiBMru2FHZPxkJ6Ixlnyson5bFK2rT/MurHAgCfo5dmRyNCxC3z
cJmvP4vov9P1eAg3AIB3p4mPF9X/ENXsFurYpdCQ20UsUu/CnDy5WKkS0hdl+MnM6aeBxZXmOFUp
h0eGYOuf9FJRfR7DBVLTXnOTjC+/+89eQjoKp572QQV5BLosz+Kvc/XNgfLbkKkA0OIz4JQzyOMd
PW0x3aylGWLQ+sCSS+sabcIWzoSqxrZDWXADRujJVjJKqE6ymr6U4BGeqnszSC4+uoYm+Re0qQHd
zRobUPR1ZKt5HU9tjAk4aPJNJFKGGQKaBmuN0mKGqwVit3XGKvUh2Yrouii/qY+jqpcTcQUWKKwk
17rq9qfPkciXHwanRlu2v09ImVKhXDn9TaNaV8J5lViMng91H3ROCX+/37rurdlYyTy4oEHxKiK1
rk5gysGHbUwbOvnhZpl+Wv6qdwaEWkXa0KJ4DYFaOJsoY5dQlSzjENAFz5ME/cF01tszk4fpuuYB
o+RgiNMDancfVK2c5pruTr+isXsAEP7gVP9JZw9fNEz6tKNg4arPMiLD7pJQZmC2xvfUv8hR8Txn
v/du8mRhglXWQANhVyNOnheJWbSl/LjMOi01/Ihujwov8VGbvcH5RvCYhICSRXIrKFwjOsOkvfpd
KVD6hYwR0VVBYRlXMxRueb43cTslTnKq2syjbX8Qz9EtNP3MhNro3bGBQHxcLTx6Dw1LjqhMjZwg
FoB6SXByZvBNIfQcqwNyQkiltLoaLVmvgFDM/TPEcAGndWcIRqv3tjxL5/jZERWehb2jPtpw/2nv
s3z4CVxpQekZVX/Q0M1FAaExl5Pw2tvRmNB+ypiESiS/h+o2pFnkIRgcCwDYz01dNjbIjoD7S06L
bxmsqPilhZBU4sNKSTF7iZnxQBz6F4J2lXy1o9sDq0o/+6K12Y4b+Ny7Us+FpSPHVH5uM1IC1UGt
Eu2zC/W3tcBegCwzhBCWso2JvA4IF1uURq3O93IyMqi/btrkSjqFMsVEtgA7m5mhNDt15JwhmvLx
lQcdYBt3w7c4FqZt7ubJRkOhqZbnVxrIEKLLoW0rIu8xbYNaWoxnZ8+jHnyUqhNGP2BU9KCYjHZ/
+GUAHvdCnIuojiqrxMmVHOyGu7jOzzdCfPG7YYcjrS2jbqrhi6KoLoR8z+1Bi0yXuXdEG1P/wLQs
jgv+gQH8c3KBeYDhASFSgZTT3NY0DMn4B2k6u67LpUNP8X7sjWTwX1/g0Ol8EQ6Rb1S7CT9QiO9j
5FHsMJHx/ZHi2QO+uuLadaUqsrPED759KmNo1bj856D7NRXHntHHLWwkk8FC1rvan4PE2zWW0ajm
1kwiYdrYZzd21/wRFh7SFhxgClpFhvTc9PDuPAR+PdFi4a8pbsKzZoTxQEC0Bu6vbaQX/SCM1kl+
oriyL4APW/AM2Gd889tb68IUpdpOSsrVB9VksRX/jZlp//h+5t92qIvf9QNavBclQcd+q+uZmV/U
pr/BQD0IbIzWTACD9waY5TxxKXqbb8zuYcjtmtdOsootY1LvTxl/b+tfNzNaeBmGAqlUOJ7TpJO1
awOwvrEdF2whJAyoq2aSgRx7GgljgQTN++bk53NdOHuj6nvQf3pBdO4TLnN25nzNiEwFRNW2srsx
CUugLggvgM4AX/6LJeXFUcyU6fyignOcnh1xWEu0IF9z7Sz3qAdJpS8puVJmu0YcaM9nxqPQJh0y
TRwT23xRv5vcyx9811AAvqiQridAH/PWaz1yjzNBfHHsA7GfPW17V/K7YQjvjlcDk5+7l9IKG0xc
FZOqFd4SoqMBedkV2BdxZzmncwFQpT/AP1+fTmcEEM5Bn4Z5SYXMLV565291OHyvm0LonQDO/KAp
5GAtDtSSMY8n0mqqpk5UXkhMQ/biDDBLZ14WGcDXwebVVqhJQ/e2ohTgb1LtNPo8/SwQvlBPxgq8
inCGaEoL4ItQLrYO75fvO8AQ3SGpnSrVkyMZ8ZH0cdlLxcr2hyFGEWSQSk16T56BkNpK2/VFNCZ7
oZHUceeAe8wFFi+igELs25eAefjPy1sOaMatTd8ZZldYl9ek+NkLvZ5exY00SbHWSesQ2N2FVR2g
XbpQZH5pWz3ecwIxmohTkrn//HdDflzuhzFppBO3TMsB1kxB4HRSn9LKEWMQbHSLTi/IiZhE8nwM
eEEPCmXRW+nIv/nnfEnJl+9b9TdIm6MXIYJierZkGqVYWVeXV3Vbt0nvATa/UEzgRlk7MGTuCqyy
+EdHbaXMPn70/rFRfukuf0BSjCjVixQa8tB1E/gaKxqTrA6ZDcGdBPRD6qaWYz44txebItqGL06n
G/7nWaTQGsRwt49HHZ0dnBNcQhTF8vA960V1U0wMlIaMsiNQampEI3D8NbemfM6dQYmCuH1f9Cbn
cl2PQjPFINrFCMPKN6HtMMuwiSoWjJDShzJLW100Jq7OQzHIguiW8R9MV36N5beG3tZinHGvXwAi
7kFlzM2ekTfHUJsfNKpv1cWVH/OJxP42UjLlqhOxO6A9DW1yru2UCLZAHEo/jSpJ4bb5LqGr3Zc6
ti6pXKbhICnS9n05TONcMaIBndAiS1oKAE6Q8LwfTqgqyq9K9uLVDsX+krYOXWRyOE4y+L1d3LCm
HiWvkW1KZu/l1+q93CPyaeGoFhxgWTc1oH/w68zESLFyDq2xPEaVav+bfrM+jyu0p6yyLw2x/90O
vOj+iAZ7VQJabvoptfVDjiDaKjK0+OR2+xqj1uFqIUtV9PJDKXXTGU1D2S2I0MfzpTLWhUnW5XaN
hEXWURbxyDXURqY9NRLNmXa+eny7Y3Yw5xKn5hNetgA+SVSP439fkZhhePF6hHAaFMEpaB81bwc/
+BZexVpSXH9gNo0Yq1Ae7zK3we92PptVtkrmVyuwYePb4mxwcPCA1844IyYpJphYxpxOq5uGRuep
x5Wq1s9sGdDo1C7ANPKTNIEAYatQd9g+BpPoKXzNkDATjN0DIylAbVl7socZBm48WY3lNg3vkPfm
nxacRa25Btjti8ic9HilX8///UAU6gBRRyZMAlAdHXAlXQPC6/DGD2yqgIKTzJ5IyjQCMnwju5zW
PFfKCK8GgQXsLH50SGTUNvioPzDvOSp3GhEONe1cjzgvKNMcJ6mEGaFy+HnjQ4e85rLsu8uPVv8M
23NewkAXNp/vSjyOKXmtC/pwXmv38/fTXFZD6OgGgD6XTfN8xtp984Uwx1LAUyO1e/Vb9kzCRBw+
5msn3AfMLkO25UjkcBt6mCS+30Ro2Lw1wthSCy2bryHfk35JW65jfDQWLOfe7FT9fYQgyOZWgjBI
jD3YflIjqDtOdV9MeLyTvjsj0RdjfhFiavP6+L0VdCYts25HPMe3YYSL0PAMhBK3MVDc1/i1NFJZ
gnLcZ+xVB4wisjD//ka4MGNQAYr1I8J1yry2L3/B/5eNDYyXi0I/1btAQKqhKdCfmp9hjJNFGeB6
HQuulN//7BeVM11zAdOcUMA5+ZsTZi4hAMogULehfJjzpuWQDlkl+lgF70hXBADEw0WESZGbGGGR
P6gml9eMfelwfXOI6/I8ELpI/ejHSjbyUjmkTDObmAmojR+w613Y7WVsJOHzKhaZAaX/j/gLsXhC
SflvyxNJjStvmEchQvJ2dRfzQu2BmiKYYSBiWZwRfGy4oB5umSY+Kdi7Jej1RPnLzhGpaRkHGsk4
gfOjllOsukf8qSQSeMB4X8KldYwogA80OFeN47PfZjOCBxu0f2oFfo8cyWcaLMJleSSK2rfCWX4N
hGSSUjhuo31HVyFsL2BUm9K9PmPhJJ2m2cwLMEku0v/Hj9VdSfO2UvW81OHnOD04TIHEfaLWBxqR
RKahLTT8Vkha4MHWlvHs1eppcVVQhuZgPdNxmLvYT5U7+vjPCj2it6474l1GUd5L5dk8CeWt2Is8
6lAKpFGBDafSnLsF5TB3WBCm5h7JJzJiEjAdrNMIsnvCxiBA1XyjG9HmC8qRffRzuIOhloKMv0FG
Zmhdjh2B33I/m4tg02H13UY8cXD627z4gqPJ3v5AB9C8zV3pbMjTcnQkr6VAFai/GDw9vfhzkBSE
fdq1oq/sv/l0lJt92nepXXzHZ6by3tz+tmHAtdXtcXCBUBSMd6imygphVszlosCkohwkl9jZhrS7
m0YOTPkZoSq/IwOaN5rAEktN6+3Ky21oo2JPJP+kAciL+ahKDm6eguN1JIdrD+rIPphueptpdvnP
72il1r8U6b1rsyLmE7Zo6tvGa0DuJ0ndpszFmFqv0BS1u0WNWTWDtIsDnZ9X8JeE8elxMEz85n43
tlMGLm16eJUUP1Br2bK2IBZtGaI3olFyvywpFn3LijIuVIncOoJEvtsiw4nYSb/aDo0iOw7sZxfA
mM45HI8sFLAvPYsaBPD0k0xuU6z/zns0LKZaufSAYr4j7J18wzajcdqffhWNSMAzFZz2Z8/SmQi8
RSTTRDV6C+cJQHTakXDwZA5mc9KfVc+RPceb0od3guvByuPcX0UOpOPfjmTrALorJ1V3OaFkbyvS
LDybxXi2APkyYN45g826fe5N4ifu0V+rXomdf8zyPcKHJjtNHfSTFSRT7XM78KfWJGxtDSQTJoJR
4UrW+gitrxGyTGC00604Vr/Od1ecom6BC6VBvQ3U1iuwSmdN8aoWODW89ILNktUazzj7ZKgmre8q
Bh0vySpb+Oj3d/s865L9yAab5rNZ7n6Lo+ckX0e3RKVV96xVoNnCi24+sZ85QG8IJXpATmWz9VEd
8vMbu4jL5YPCvwwMyTt5TjsEwT2BEsEBfglPEoSOOp0AwTJWbuvkbDweB6PewSJ5IjV4X7sUD4Ji
ZDLek6RYuAgHYNdnFfQYHzqLkcWls+gJ+hCXG8cm7O5z77xL9KVcLKDavt6OWQJpwxtt0eot/RSw
8cPRiP3DHh3Vd67aLCvQ3JNbYObTiIYo3ZFl5Se42OS4UprKeoku1JZQZVFjwSpyjoe5FldGvYnV
9X+zMoM3v21HGiUfJfMdPINB5oaPxEysBFMjoHVpIPIKCINKmGbmeWvcK/5oL+ZDPoRZUJEAe9la
/zXUFGaS7DrTqfY56gyx0zaFoRrdbg2+F2E6rN3vSmZXMAj6b57ZfAWzamhbBiwLN4yHjxlOO33e
xwt8S2skuglMP9phkkBk3Y0rCc7PIPprjomiYrlMxgYP+4nU91dFgUluLU3y5+JqklS1+PIYvti6
+JgIwGxUU4KyDyUms5ySpAl/ug3o3gTs5lZ18qKPYlzspQBx6Bs6gKwuYVJzGWv5yMlv8d2ZViqv
j7Hfe1A5S64tRLNuJA0KBvGctWqU8sD3wENSWIg2v0U7jbowMd97zGoInCYoV9arBM7roPXb7he+
nALnmbLfn3wRJlj8TsmfTqGAxT5y605AqVnvqwUkBXFqIX9i8dc219+04SCqnXgc7NdW41bQGuCN
yPeh88RN+nsIjwB9JMOOZnEjXrcisxc1IEoohT9dxSSbH/BqEPFo+EA6QT+4vhAEXE1qizPgy9/Z
PwK5G2mQnY92vUmMKpJ+pmVdUuckfeRLG8tpAR7wi1JA8+peqMwhHXDko38Wn7F5ZIKCZbihtBZH
PugY2XVxzyV3x+2umwhCLo1QTbWTctVaQ1FdU6y3g56uoc9rSjBnUoGu1K5ukZXEXEczvZtT4OJP
qiUK+Zmmh5oj1qZ8/4YnsVmXkeJuOuQi7gUHH+BubBkXhrTYhJhiCJJKwPZBgWTRIhvkC7k6r/Lb
fYqB3/TWWihgsNCgatA7F+7xZUWelL7nCKjpG5xPuiwaV9SNSwzCuVcqFTcBJDfOPfQBc5zCsk0E
gH/j0YL2V3k67T9cBwuByUooXI6z84zUA3A+1TUTsgZ0glRJAuVwQzZWXfOTI3TSTMjc+ykeOcal
ges60hQAX6QoSW7yvBmqAGrouw7o0U+AFzdZYSmTcDO8wDkBq5bqUT2NPnl+Jr1GRVax+WuTnAfn
1fQLuoYFAtoltsgxeUFynHFLqUtWPYriacsZns7knBc/chLx4LBoPNOcV3ggwLRsruXRhdJsl4pY
thBN5axPlRO9dbB1SfA73Ua+5yo2ARpMXbWgAHO3vEOASH03gdyD6ug2apGAjZQvlXeqhDaVl+pB
huFQQC8iCbFluCald3rxK5Oo+RWTHfghdbJorgrbC63nCExLSRs4TIwqh/bS9kRsdyY5T4idzWna
yrLM+PubzZmjj1a8tETqtoY3/95egeTAWd8L5AnU8G9kmpy+dKDgJBUcu75/3b3TV2ACP7kb21G9
ttGl/KEv2ffSYGjRsiUIDcX39I7PJ4TGxi3HYQ3PAZqtUF5fmcPWCDbL5jiCWNJpiXXeeobx8wvx
Zs4GA/USSK4O7sfds5y2SpG32Rc/fAzLKyY1D2w70F2L096ED7XNzAsjen5DMiFif/nZMgusRml3
ZcFV41Uz/912m1xJto6l/yeP+PuZSxj0qF8A9sJLMk2V+5/Czc1U/+y4WNvFw8ZhUN+TiTeiovQ0
Blax4QvDMXqz9FMqHn5X7zljnb+oz1inSqMx6mWu+qMs/wv9Esv1ZnIfr6YYbZLprP1CUDe9UnYR
pMkFb26dekxCDgLYQIlbv6BFfO9hpNkSDGgZOxQMQ68a5bPtgjyG9F9E/PCbzyAxIyA4AB5O7/sF
sgEtYvQrYTVlngObFrOLmWUKXNKqYSPdh6x7g9z8ZL6aqdIXwGWyaZItBOXIIlHzCMJoVLX7EHuM
/GWV+5F14jVai9WCuPxChKr/LMLxaVyIhy3jKej/zp2AfnoR1k2gnbzFgJH4cXLIjY2veLHVtqe6
xW1aFKuQENzdlchiIuf8SN9LNNWet1f7q8fE/l5HTM0PgR4VwWDdEKbM5d8D5/5uBbBzekotpwte
4NA6wcUmccw8LT3iR2NJB+/aoGzIA679FQZDg7PtrcmRouWBytmPwhf8fblqZ7MJbEgXrNB2Hx8a
ugQqt1r0+Uqknk3zcSThjC9gGfMsXM0tsFC1PNEa+VhR0acpmtRaMoUemPRGWyL666ZhNTzE7z01
BCtq51CG/ieK+D4uOzMHnQ60Sks+/6zDvb7VJkEJmXnYlngTKWPm5Qb1OC9yVNRpn6cPk/GDa7e+
ofWhMYGkv1v/d0pcImjpc9kQFKX/ay0A7HSyLKVuQWykK/eKGOrxNoYLjqyDQe3cWLQz+Z7UeuQq
WiyjHN8mqePBwuQ8dFxBtUIg8z0hItAjyeDrGFrBSSaDtyo8oO3o32AnzdI7F5qZbGMsKZpcm5Jx
BLyQBSW3K31JflVwHzMJJIV1jM2H3KDnzFdWRb9YZEYhsvWqdseSwUO7lzi2ZzWlWQXdDEzwWMJu
Fiq6OdTMpNaTCFE+gvcGq3gCKTyOmNYvC00ulpKrsdecrP4JeyEiNhuEkTkff3fn2Cw6yZ4pg5M6
o9OCoU4LPdIkIsE+D/m9ITaJdpbKp1eV+G3K2UVaJyphV5udUJAcB/Pf6/kiu26AhibH43OCfEBK
vMeLcK1/kYt34jKqD4Kjn5T2Hf1rVZvrbam1jgFUIKgc4RbcX4JVm60Kk5xNTogSe4KmwtVsyB1T
/Gc9NBhZzGIJQRFBexVe1J74eU2O7Jh+SUVMrXSrYO/3TxQwMrq4enAfM9u9T3BD1u9R5G4nja4R
xeStKY1BnswqhcBQKwwk3uSQznUiFJuQqyUO6vkqTFzK+YUblcdX5BkwU8AFKKDV5EMvehuugtc6
xlfG63uak9UZQh6rg7JyS3Z/QzggxWZOI75SIeSVcX7rd+f4frQIly8/Xwr6KxGY0EMgb0ukRJqR
Z1NZFSh5e7U9KKeveEgVF3u6pcOgx5HxIqdBpUobWoAv8OkMI+z7HGrd/MGvhzSml5vhmW70zgRw
0ahCqiMj/MJ7v2v4uZ9xQcqJXWNTbnwGz2ZFdTjEPfWcVcTjf3Q1KbzfMrQn/X9WJbyTJXwkSucQ
UHu1psH1EgPKOrYekG62QF/Sw2b10nL8cDwYcHKwfnfmDHfGLkDLtgQENyxoL2NtiugdTSU0tolb
iLzXHhOX1+aM4LHqGyIBcqJaWbIJxfTpV3EcoeBRJbsV5JZh7rDLX8b3pEjxKRKfSXanbOz/jaU+
7LHm1qb+ad7UtxchdCsEKMirE5OQ9MJoLX+RKDxFL9WLce7KYSpyI1Kt2TWvtKtqPtCNKxKOslt7
CpT1Q5XhKAsSeFmt3GKMtmkV5yjtHO87O5zwWWqKgtwn+N4Iubc9n99oPQaVKBEAZqNbUKaenPHn
Pyzmq5SJ0nZG18oGKvl1NTysSWLkkBhEorUc9pkLLkhCf/pVfCYfjeKCES99K4Ijg4Z649TiXWeW
KFksJpYyzIbvtgP9fDcR7gTapkZsMc3Q69ITCHa7WHYnUN6AXGila8ZhOM68bWeRr4LRNQIV2Dnl
zfS/hR3OxjrfOcC5aBHzaOHGVniBbSuYYEfEmXncRMEhrRCjOR1rmbC7FxxFagKfUy0Pvv8NbyWk
7/hoE4il4xlCa57JCO2zXrS7jSgi2ygD5wQfu/fvqxoWJl9MWRxoNt+k4K2MwDhqFRx2t9hw59WG
G9aK3deq2LMIWDlj3hrGq1eIdTng3/p1vrjC5tFjM3YNf/bOVFmvwQ5jwyzIzUhrjcG7ioK+Q9N1
p6ueezpdLHLcPI9HPh4vIudit3d4qDmf9k5WoK24WEUaBorRvktPeWcNRFi8VCqFz/1Lk6c+AKiI
XUnUbPiIU0LuglIjuQa4veEf8yxemncFnHcLdOihVO18ELpmUePY++UU63/QYy5sLYjoaMwb3IY+
YZSla4OHlJZTwPkeCnBKSALzHzvr0f1pp2IRXdkVietCahvX5BGseNViab9f9EJi7YxIMwuhfHqD
9tU8EK0uUnKeauYSCdvE5Kgf35/EsU5/eB6Kh2Pp4eTLVY7q70qnHF3xdpligyJONASNm0FU4DG9
WYEahk6iyWK9S6Vhtdl+v9x75LppRZrA20uU4m/MyasARQRJ+O/qMZqUE5z+PW/gSShEjC//d9ZP
J/cUCVYsawG+tLwOupy5hy4VAyqIyqaNza+zrxJ8G0x/egA6+kJ8VtduNiXPQnkDrIN2Z8OVyz9Z
0jYQ4qywZyc0G3gyRJhl/7We81SnNv+0tY5hrjN1TnEdn7U4TszDu7B8VXhwj31gY4kCByeruuRQ
ctSyEiHyYyWH0ZU1EVS8vHKcZ3eFcKmrkuS59Qol6E0mlymnBs2ioopy+Djowc3NH8GtTJ0Kwx0T
YGh7KobZdxz6XA9WwOhVR0XIJb4QTdJpc1cCnZXUPZx7Z64o7ogCBenuVdL0lAKU7gHuS3ErdjMH
/vEdawFBPVc0fblhtFQ6NgNmWC4pmSk9CLsyUbIQ/pSrabTJLZxKRjJNlnVl/6kbwyayB3HizNaM
mShCQQs/NUOx1Yi0/3d6l7vC7I9VmW7BolIuIxGSai3C36u74KuNiSbvkrWkYk2kr3YIDDhlVLN7
ElR6gIXpX3GixHtjrhUtCc64pxTAqKIAnsYurFCqoVT2MekWHTAVUHoHxKN76sFevh83ioHQP3cc
0xhCZgbtHYlBvb4ZTW7BaaoGHv2r/doeNcTWMS2FrxG58GWdnOsXvC/tM9JhviPyk7/4M8BzfB1S
6VmZMzqRqWIOI4AITo0YW9/lCzF3ucO7h9vRTUcaHlmLXuW/9hFFl0PVqVh4KJqUix80YXF7KiYN
+XHbvENeXTlijNfmDNX24pC8z1CEk1aIl/VeaOypQwujZEsLlVYKayvURc6J67SYh+bnAewvfHvG
OUwUDVM+P3JdOkCy/63XPNdxBS1ZuuYNGa4V340CtovzN61JYHkm0FhKHiOkvAkFY8s/frlMvMpy
Tjt5kJ4TIL+6DeaW7SJANYs/uSrD9sD8bmZpftc87Ujh7d6/LvINPOAQY3UDEE68W7F5Eob8BG8U
YHy/HFl/VtjbTGkxhsel3/Y5rRYm7dy20A4M6nAIjKv+JbIh7a93k0ZTecM7Ndog5VCXO2E/PGsm
3C489CgChpLf8lprpkbnvrPPuHguT3iKtNqDVeva7SsM/ti0nykkF3gBxxtEwJf93JNX95okjkbI
0PRhh6ugNKntm/6VZes+lzKiQMMUPe77J3XJsipcHEIT6BwwIYsrCg5EQhpwMYR7sYwYltwCNeaN
Jt0FME09NGEg4458hsI+Cu7fAyNUI1nzlnJ3cJ2p36s08uifZ3mo9oHe4yiVboxjfGlLltJEs5gG
vOeaZgZtoGn1aBueVUApQmilVbSOqEVb3nu4ccve7glTk5K6yHpoeJ503+6pCzNxuliEm2meqb83
eQFDv7UkkwW5wWhlwuD8SHpI0vn1YVWsqRWLYbJLosm3PRk+VsrrO+9XLhrPD79W9CEi37CFyWTH
yPUEsya3yCpAlrU16jEmPJ+2lfx38faJDbUx1XPFTETHpz8VJ8QedSdg2s8P6/YeFexRlJ0hOgeZ
t9V+Bx9aKs7nWcox41QuymlKtvdNHjy5Zrg73gf6USvQs1p7mtollyAFmVQzMmEEEXcsNgtYKRW+
WOe1vsWxGijp2VnmphVvABBeAZCpIxIkNhCT6vAHfAbP5VpShJhJYUt5MoFiyRgKQ48wTLKHGoQi
HHtaI+YTH2F+9culyxsPJ8AW61/Sf9llDtNyWulLyVy/whENQnNeXtwzHNI4N7x7zImi53IJkYJ0
rw+9kKkkaXKMd7b5YrfNPDaBPmxjH25cEs8QjkmdeeU0iFV66DpiOdjAcBb5QXA/sl8dVz3pQ6WG
Dhb1TfTER3WymmCpt4M+f1iP0SESfIwHfbcZfWBzXNH7cGAs6MZYrPkyqAjdv4J55XlzadIMIe4C
XL1Fv2cbts/g8awwcoiqWwnbYpe3I5+TVUcLmdeTqTh89wTJFLjuN26utBcGv/lcS3R/QdUHOG/s
+MoTXazEZdwOopA9yBJHZ76lppeFPnMW2eWsO2dYK+2eMoyAXQu+7xYTIJtzRjPubYPo10iqwxP6
yh3mawVUvQf5uQ3wV1+75mf9pa7VvvHxO3QMz3ozHiPcj8dxG94F/jDGnMo0P5g55H+NaXmNqEx+
vqqCeSAgCy4TBRqP0B1YNzbUfTfuOWzf86Gg2kbj3viv8rW3zzOdo4Tc6NN5dO4D2baG4cNOAqYL
tQEU6U5KFP36cPqlav+WM7AUB/UsGhbpY0ybq4FJCNgBz96205UvVODp2gJougvZxojmpmQvQdzD
JxVXKaKqAqY/7+oDtxRQ7MYUGI5WnzwEsKCKJJ7As7gxNxtWzTvU0Tue3ClTDG80vZGwCzmQjlrO
M46iKV90nG3tux9B9On+Rw79tLUjxaq9GMupYdzkzsMTQO/OMhZuIrU5eNoZ8t/xeDwVcoDMr7sq
uAqWH/wOw4WrjW8OAIII5Ri0Ab0EfnDPFKwuI2ZErbX6GyhzogHmq6dfV4MSn8XThxN3rwMTrH2E
JRmjVj0/+qNGKVqcLYSK2OxsATr+M4xxyoIPjL0tJ4I2Ab6vcF/pQVPd7rwZfeZQAjxndOgwP22B
UaSPFfLiH1l3hPHZQuZy1HhzzEPPcfdXf+SjGzIBfVOokO39iCe5G2YxvOzQEzu0s3HnF6Eoca+K
bu55VTqtehSbutpO1kaVdkIegZMwbvxQMR6Pfx9lId6YaPelTLXJn018ZxNTkpqi0m9KavBJJuj0
4qjLOjZRCY22ENjsihrxxoTOLWt/I9n+T5/3eFhoarnYZPQ1shzSwsvIvJhdj4l+n0I3BaPGvdZP
56k+FdsL4+m/tJzvbjnhCdcpnrBSzcPE9431U81OP+GjjiPpEkCl1llJQEW6lQn1U6QvAWyUzHJm
H74c/Kbs5G1+SvVk8twvJVvo5ikRpMLLKMPaRrzXeMbI32OmWeaJLSKfPHD3OPaQGdjojo7we0vR
YiIFSjeETgD4BhlMZLb6H0tEMDuXjJ28oPp71UHuLG9vAI+Cx21JDXeWsx6IEpFayXlEPvJjNfqG
GbWdsZLmRxLmtpKLY6f7WsZ+qcNqLI/0FECvhX5I1aTtEkW3AiuMYWQhZ5zDahr5CZNJI5MjjAnV
Y2E+EuUoSk1aU8dAVRA9o5hp+ZyjLLOnILMs76vbf+bN1RO77z5/FU76KcYefbn80RmRMjzybZ+h
jzHuqKG/dD5cARyG78XfKWCxWX0zEdsy9ZDvLjjTooTcM/5XNPUz+mKwviyJLcz7VclQPHuLqE6E
EnoPtBpFf8NS94tJeN95eD1GcSt2/scDfTHCn9J77snTykZYZdDjlKfxLPl0O4dCvuAA74PaZ0zZ
OW4KXtbyCTkW0ELPnSr8LOXEjP+n690rFXhPgD/aVQll7RmV/iz6cRcfTKDcZCz91ETuKZ7/voxL
0A77XSIUI9TMgkpS9iCYPpquWQXGqte9xRE62IQRDQMr+QryR+2OtBb/7YOaP8tN/eGaaUNxEIs7
oMyyr0k8FEzDcwn+2wWMW2WopGrfKkMpiQgHBxFQvF6PPQV15yNMN46cMcsyXFVrDFlnPbGiQmbm
TopncaJfJKUzo/taAR7H5X0u7bsnX2eflI6U4nUc116AQq/v6Vk4n49prYur6RcCKyWcWIf3KOHJ
F+nujg5Vak3J+YNw9NfvGt07y5ap0i/WAw1KUK179E1Ip+/HiOIq39CZjpWdXgYr+qAiIEFyNlOv
nucphHU8DRI9l3EdbryW5To5MzZGYlj9dGHbtDsQEKh5bSRVhE8IiaUW+JvpFY/vvA3HB+deK1Ou
VeUBcNbG74VzlaSp0JtHkRqLXulEHiokCJEyEKJCemF8YTKDGk6UJ2biyGGtjFZF8Aa0PoBHzO1J
8C1PynVngs51nGbPu1DA6pLWJ37qDmB/67FvgizF8MForsdIFTvVBHDZEM05uNclEQWOX0wEyIgi
K6LW/r9kWCaF66nGU/NdQ0xVU589mjHNbcc7pZFezRqU+9GhvCw3RN6hjSLZHM3+PAwvfRCU+xeq
bBF6jrQpa1SXO5yT5OXJroXMYxINBJQKZMQekgCdh0Z4wrpr6CRZFd2iUxLbXjVia4aypjJ+789j
jtmTDxsqv/Zk4iiziTkuAIYKqJMBCqUmAuBsOlJsGT3WwtCOYfhlho4fEkMWt5nOV4xsCRhsVC5s
SVZkNKTW1oZsuLqwy1L1AIR9Xg/j+oh3Nr3yp2zZ9AhLhZuGzCHJmOzi2BhFKqmOP3j+3eh0DOA6
rGZMMLSMNdB7w+a4x10a72ES52/tcUE2TdlePu/hWxxpUpip4i0ym5emW5+NJSd/QMmIycoAYddj
WJ4M1TAAjaEmrzTRJXPDF1S+D2YoaIlO46mhxipsAZQzi1ya1onsOImqibrYLhm0X97O9AXtvHQJ
JApt8KnMGldwugPRLA8zAhAcdI6kzUF+WMcKXQliBU9k6WM3XzUpLMPtc8SVs+YnueiLMAPeXAWE
xLdeBS2SNm8qdKOkc5ldCX6Xo2nGQvpvNC8MLlZATaoE/vh6nE1pJuGTMNitwoQotZ35EDFam+H5
b8QOgH6+A+XlYUJ2WnG+9tWeSBaIW0JXF9CEW/1ttL6ApuKcJAmt+GOJWlenZdq4htUXh1rZPa6D
nqdYh/kphT0mT9L88xz9Jh3kWRlq4pbGgxvOol6C9ePkrmafxjzQGam6uoSN6+3HP/Nw5EwJ97u7
F07xcqst0QlOGkgLtLVOuye+k6bVS+URp16Lkg0aSvLQkqyH2rFgrb6NmbT38un7edIM3+EnCAsA
4l52DYd64bTLCAvQ1YY3KK3aJ9g34DQLx/Chuh6U9hPc/MwpdW51CBixmCdxOn7we/4y1drYjAO0
D2+VC3quJIT7gITc/DU6fe/zC2F10iiwndCpSUMd0//AcBVKb4E6WL9a6pRKyiJCGnODA3ou9kos
fl2mLMsmJMnJdb3hkkfRLBJP4mvXrVka7/HCCkcs2h9RT3qvXnvcyZC86LzHdoxzjObQhlVG0D7O
016OGUxeiH66cIG+og3agx2aq5io7391uBKUeJkE5R9jmVidF1NAGv1cG7VtS/MKVM+AfnWe4HbY
OSDi67wxjtV/cPWzYQztTHvxZwUCJvQT38UCLkzxf5DQzI6bG3u9yg5vRnBP3ePLBxxTyR3VrMyL
MXHmAiZqqKQVClRAn0Q108ll1W6lRJXexTG5sfDrCS17kcBcQHVIHFSsv49cNsoZk6TzIGWXTXLM
ayiGee03I6c4Jc+CYIZICYRmDcm2UqXCW+Q1NxFoHWGFK5YNmZwbSmbfhtmgaY4mgMxv+iO17OG0
e5WTbzsmOIFfcvIjAZF0EX1sVeJp8skUxdK4Ar8Ft4uAxRJHk9mBz/DBtw9trQukuFhA/5FtQH65
wLHKFbqkAfLjrZeC/fH4rGFDXYNAMSx7QguTxYxnXkPmrOnfoZKrsKN7idtK6m2bUd2nRoTDlSHC
HYh5h3QkUUmm14kqOWzMBxWvq3Auop7ZARp4xo+CzyQTSrAuF4prYu3qWwA/gsa8p7V4TnA1TXPE
RKG01cxg08r96ZV6XQmSJKWohmAuh6cdo0HFc/IAdGDINLrJjy5doCp+GOWiV69B7RCHxJVA7xyy
zaEq3nGh0xJfYuSwIN28f5RRZUVxVdT/3LbUJ1pA8z+luvsBAKkUFgCXPNY3SPBvazJdL78Zys0Z
X7RZgIEM+nfiuqQPS9C/yZoFruTl2ByO8EEdBi4uxBbYDx0Efaz1svU4cNj75IfoRc1dKkO7FPyc
mwI3Lkv3g6HzCO2xpfgmMS4V+84seNPxNwwL878lNMuQ/yP5wa/4GDhzHnsbWUhj31ZDJk6ky06t
dwLIiOws+KFd9QQM3y2rJ4ZWZ7sOpBntY2fK81+EyYMDo9ImGwYBus+qjKbFzr493pItwaNbjk39
LlEs9QgoOMsC9H5avDTH3YwU62aA0aY9N6qwQEAySHtJgBZXbrGsyelmHrHz60CKQ2MW54LD3AqJ
3VkC/RV1L1u2QvgJc4JQJcRVaELOca+W6e3SGVsbTHJHIuzXSpD8WIIsmI8BUH9/2pMv8XfLKpw8
gS+07hAgS9WBuqatKyEcEmMLg/hVAjS4Cii2SjlrcCZMOQDPWuCOcx9OMivdee6gl4Gm0LS3v3XE
B/Gfq7fTt77whYf9Q+HEZZ3p1rhyE8wh7SRWiWdVAVqSt7UDgp2j53Ll+GASrVf5/W65U6MY9svW
H1CmNRfTfcyEADsqAuhl5xRebV18Hoq/hScNnk4zLJF0nKshXv7RMZGQlvpXiBp84uhajIHv/z7d
EfW96YB6+k1JA3FwKuEuQ+v2jXQVhzidiy1vNGar2FHtIEYFUcgvd/UxpSPcI0KTz2M87shPWEiB
7R6/rWH+ui1wkr0vV+atL/xvtoVwJ1SO5C1OBZpw65rLroxFhcVCdr3KMOabc5VQwUxvvIEXEvPF
woKqsgiUHEnmO1NmE4cMbfRVSUnKf53V5z2B5FJmgWoEFUhfaS+x36lCftdt0wF+dLDJHXc8+mIv
KjCHAGEELFZ9B4GB59kojxvKRtqdAbGgZ5wE34IhmMzZZo1JNHpzcF2bR1/IX+mMMDjFSOsB1nUt
BBV7CgJCb7CAfqAtfWw5MNawp+b8puIXI7XLHFQxRZniMwnAFCNKzJkQs8BiRKReGrRSiu30TgUZ
Ka5BkgFNA2i/+5C9B74C3FwwLFzcmgUPJzZ/SWfg/hYpDiAyZV3X5VkuE57O6L5/wd9dwMvG26Oh
8pHp2S6BECC5kQkeSGmx0YETDK7C2Ye9WuSgujj0JxTdaZqpgWnVoXeQ6oWNpy7WTH1dko2FAth8
6PLzkYMo2JW6zrQaXtFlLjWn04lpHfzOYRIJVzMzbHsrR8JaY38BbM9HHMhZnrbwFt8mnNiphxwv
VPPI5rL8jOTz0jOQVHxKMFlrytDCfA1R7iEeM6qM9bk93emKOf62NRtistnTOuognTQO0BKfLDvV
vMwNbLwO6XALVqyLnumCDRqVgT87JsnzIML+W6VKNYp5LatA2qwcOVsxNFlh2naE0DMd0ZMtEt4H
8LRY2NGcc0x7XPcnNK3AiJwqMQZvq7LYeqleBvdMlAcsylrFGoiwUBPDY8Naqd7XUf1q1gJuK3X0
PjKI5qcT4ycIM4xMuVe6tv4S0gq3ao0Wn8VV+4f4DPa5G/Z02fv6xiJhg6jAiUgTTm0bRbv1cY0J
8cOh9h13xeNjAO+yLfuSs8UJzFOoNf7ovJXFUGOA+8R7lw6wYFx2n158fA763+vj85Wjawxrd9Mw
BF8K7UUMXA7SoHpmRSvZK0PF5boENoykfm+Vost8QNIAP/UEYSY1hAZbVBeDTHGo1d83QaPfnoU/
KLkKGh9Oh50VNRhq1ogE9ZeEMuI9rN6H8QOi2ODNHaVWq4lB6/e4Ml/5RfzafyGjZbyJwLf8LQx+
Y+JJ0XE0WD6qViyOL4FUF7C+6pYVWc8xIXKuhvpJDqT2ew6/vHZUExxsWp3ZTQqEucJLAPXCW3Yt
j1N6bDW2ILpQbTHu/QF50GhgvtcDiUGTgQIZm6rDD9cd9dSMT22tPwuovP3cEFp8xoYBhOCSWzIg
yVZPqscHqLlduCHWIOauI2D5oQTQ6824EKmhtM15acQUrBQwgd5xnIsRMnQdL6lvtDJpMwKXyLa6
6pTPLvej5Y3H1/QMdekzFWrScNcYqqZKTzqFCvPJ3sUwJP5qVZwX7XMqQ0LHfvGLtzNeQeOpWi1Z
I+GuzbhJsy69LlNpSA+tTxyk3UFazX469uTHacAaU1HvXaLRSpA3L6FidBWK9L63e59UhQHk0FhK
91+mgdkAphmGPcD4Wy4FIa7CjGiaHEZATAGK/Lt7XmlC6nPWcAiPpvw5XENstBmMSba5HsYhs2CL
GWWGMivPodVv+f4CwPd9P9AJivxQbu1ulvw0VzFpQjEcMK0j5GMeBkmcLPf5a1hLc3SRJPsfflzW
JEK9EjQyPonujt6+vBx+GLhvoicHZjyexJc2HDMtpw/UMO38keifG4qDHJFJy6+gNvKFSZiG/q0V
NSsKjbiYgNEKGqm0IZzvuWXP+WcLLQKAbhazOkUjji4MMoG6hUIDhj0wkN8L4fXCBR4O0/WjRRgk
ffRn8IrCa6Wq0048SOUND9Rbbt27+5wxWnZap7y6lAgutx5PBheFWVMJ7BfY3BNYujPbDSKuRSlR
CIwZpu5kEKXRL0J2WecqlEtT4GQJWstGBAvXxk1bZp2qrCcph4Uv+b+8uFLwlvmNuPr9cv6lCT9J
nlpz+jF5BRMiBPpakKqrUNY060cKN114zYO2LnHyF732mbI5U7jBibukHFgLpguOqM+87Qi4hQPS
h90tmziZ/FXFJoN4/47CPhZZ2ZeuFhgTr3pYH0HhbuiyPIKF7XjDYr0SeCqhFpnePolRzABAa5OQ
avZ8CwvT4TzGGcxjgqFIS9q5bmmJNfdOm3n1QwlA170htyzOp6xUSquz1n3Pn4xcSGVHRjPHUls+
KC1P7zxiJ0TIXmsHag6+J28B5EZQ+1/quJIq9lp+B2msaiHlFtP5STV3zHMKAAkYT1tzYIN9pK6D
m2Dh2TBEKq6YQQ5shQfn2tmBeXqri+Q2jo2+GqSyT3MhoS6+f/GDxzv1uqbddV/dDaEti0DhK640
eXwGZnEmUE+mub5rrp+5lKMrxBCMc8rU5g36qwbzfbQodRtdCK7GkFtbuaNvdhvZwVv/VdgnELmG
lyFp5OkJEj7MgSlXFe5zCpTEv1kLfkD5HF8ySKTfbIfHgTCbRAdtWnCy80r8czKnYyurUAn+NTgb
KXVXIeS0OG6YIqQKcCpqfvNEHqbZwG+HiIh+YVgTubetLWF3E/g+Mtsop1E+vWmZTkxhiP/Enxr/
l3usbnKW1Jy66ruaTVOT5AxD9V1S1fWtclT5gKfODof3Rq0B+CYlLfrSXEC0iAbdmfFvYSf+iQoj
teK41//0R9yGg9C8by6ystxlXI3jZ/KklNtrni8uN8sw0Ud/PjL7VHVpcAthmY1q8bNwk9Tc+9b4
5N0j/4P+Ut/Dhcp5fBSopomgzCJpcvqlOJMvIAYzbqd+ddtsPXWMH8VKfj++w1j8cU5vas2p8G/d
lA4T7mnWuottLo/JewD26fANou3YaQp5HCq4AY9zJPen5Y1y0FrazL9bUxE8jGzPi3lu7UnYmZzi
kXLdTnbRu7Q35UEr+2zaJHALMuTMV+Vk09KgdS+gZx67PIQWiDnRoc7lSE/pCeUluKiKL2aVKpTe
g7lnh3Os8dvPUoA3KNYQ3EGBLVvcCgvctA3PfKUgHR3hxCbwIo/TX7/M42qJNfRI7PIx7kgvGtfh
mC6S4CGn5djsaJddDypjeKfIap53548CyV/TBIzB78KKKqzC+iWDz72VDRS8JduQr2fPfT4BB3gL
dapUgqnyITvpsr24A4PhQvb3nN8cEfCsNnFj6R6o1q8SeNpOxBhAhECw7lw+EajuyeeBsxqji3k4
QJfwp/3QyiCHauLTHoBjy3vUlCrBpCpv08OdcwXhAAbOPRyYz3V3LBWwD2MCxTQhCAuDAuEE1yJd
g5UZq4dBOHO4o4ObWGkdsT2eJlF6sSejoc/1VGZRDPw4/5jBHAqvm8aqkcmqndt7YVIRIbtBmuwZ
mTmGYnZQrBC48lZG6TmWgJ2cAi99zMylS6/eui9ZIX8I1yXs1Z3255mLb2bn2wfVym9wwzuV/fOW
Tf560NS8ZBZHQFyIR2HykNhD5tlmjDBjIUGqp7tlSlGrTcN+CmbUPcqxQAMPJABtCkBynMxGqStO
KSuUx0oGKRiYjBylrhss32R/K2g1rKMvRDsVx7GKzvSXa3U/FUR25uhUmz9mrKjyzG39o7qaytLr
1MrhOb6IbJPFX6MF+YAwzvKks7GKmXpwqATB6Qkqr1OocEfNlYAliaofsn2hoihLXIF2CFH90Vbz
PeMzzuBxdwrfjTEGuVkn7GTZxvugAE7SN/opaA7yIUfLiwxvLTg5Ih/W+xflK69HsggL3MkR4ryF
awqtZNV8F6Hl9SyoEhNsuKYteqQmuHzaX2E0rQbFqGURQp3lUMVSQ9e54I1N7K+CAlPocLaBCG+4
79n/L9gGyjHsyXJJsddOD8HkDLKxK7wG5RBJHHHxS1wNEcQUln7a8U5BvyI7Pq0p0kpmXItEKTrp
49EhkXAxKkki1huMAZmH3LjtZa/moqHJA+VWYvxecVBphuiuiRq6Q2MJdaW8RYPmmwLFp5UK1okj
EaMXfQrXljAb62eq3M3rbEI/SVxSmy+lRfiWJhsfFfW1DouU0fsUUHuq4/Oto/uNS5amL8X3MhgM
WramU9MvpxWfXR7tk2BNIdOkuVuZ5jO0HhqkgDW88SkB/HCzCYhvP9hZxn7iybPqrsqnZNlP9EWb
Hf6KaZGnMbo7H1yvdqnNek5JMZ0DAcYiGn1zyZsY/hVBlxhdHB67Qfd2M4kh0fTCueketU0r3xo7
s3eyJnYp8P0XtM0veuqJNMogJ60+/EbY29rsTsTdzvGHlxhtNEer+mHDhNrHZTv16Fv++uK0PwXI
wLSph+YmbrSccJ1JkwI7uCtpDb+sE4ilxqWn8vWosePVPR8ZaDUzvVsu+O//iZ2UPgB86qQ8t401
r68rg0nKOKqt8VZJTX1LVAn2l3N6+BZAUFin9h2UYynbHkj7n/iMm22zHfvs8Ibmn6DyzZQVmTs8
FSiQfloE/o/4bNT9gs6SdECXiASbqcQ+JhRf6KKFy/b9jv58O81O5rr0DzFf8JFXJTVsO6Rj15P/
jnF9VWDgzIki8rM1etB6uDYU2GUDVujqfjzZ3bVVkvEwIxD6ZJNr1ur61UkiRd7ZJimGZYM3xH3W
0FnDqdFUMb4pRPCCa9DSjcez3GXnMAj3vU9gXChTWwS8fN9RUHGsDTW5Xim29dhFTqE8vLb7RvNu
MLvpnBb2akIUttgwlTT+54x69jutynn2teKI4w4RtXLyRr+6uSE1VCPVBbT76IVUH+niR2CoWkgd
6bLpY2AguW/a3kGF99IHHZ99NG55KbIWpdPEEHKb+d4nU7o1/s0FaR3L9vagTK+LYJLldql6ZxjG
Kft5erwB+aXDAf1RnVzJNtmTIWivD8lEYAT/n4r/I9BkbEjvaDPHzEKcqJgJkQlhwTeOU7UuBC2h
5Rq3DLKUJaVJHTbDOc1PIT0t9nrtWElv6MLZ5PqlVoJwxvCbfANi9W4J69iSCYItluDDdXzOYlVM
dGjzpKaPutY+ZOpBKYG8aF9ohFAC34QmjO91PFtO83lIzmo4QThbOZqNCbfCfRog2TPFNJxwB22g
R5IjuTqrU8x/Vs4mvxVBBL37Bkirs127ei+OwKjkgHRJoQzHigYIxbv2YnyWggflbdffJTArBfFp
o0giTopFzCv/srr2JktYW+Zk0kGKTU4+AK6Oy84tTE52Cb1jQEKvbrF6O3kfh1cgAu66l0ARJ2df
eDIZTAGhz1hK1Wii3jhOkmAWX28cLBcWSlGzo26maWUnEgSl8ztFJZArTMz4GX/o3c2xxML8I1qp
KRbrigczhyWn2uAReBMVraS7xdafcccnvb5ENdKDEk6IPPZZMCROOIuNLx68u6JquKyiy0sivyob
SSyOEinx3bLVtp2Atjt9aAs3pYgrNlX4qwWt+LwU6y2Rh7O4BCNMtmD5tgJLExE7qPDjpsg4DUo3
ZwOjP55i4y+yVpAQwSaAoChY6ANeCCliyk1GdU5TL+yLRt7C4TuuqQH7d+MhJbMB4FEzIndpSgia
sfhoyG2GCpMCQvPtMJjlgnblwmh7PFIjo1AGnng9slUBuyEVWfAehZy75catiIr+7r0L3wmsotfn
8xBE7kRgTD2Wa8R7gdaPqlxQ4bkGM0yYEn4zviufsP8fXHMrHBBuODCZzkXajYHc9JBihvIdZH7i
ngiElmblYS0xICbaeF4SnDvo3w2asgb1TVbP5nvPcGKtT3y7JdJ0777HAoE94JXGj5wQa7MzcZ/c
7hMJChdPEOoc3tAzJB4E7hrtV1re0+ZU1VvYZbvJGKFRxzmaV53mvkXIlQWWlmQfIOZY/efSbVNo
wQcxpc9sw7DbezUbUAUtC3FeRN1k/WoYqP7sbmmTjZal1K0IcUFUcLDSqjnJIrqMUcFF4lQ090QO
4uLWzMOgYZy1Xavics9PtfzLM2hbR5on/WOSx2CGRtXJgwB2HiJDCHNA5X9C2727f2IY5p5CUDf2
XBh6wXDlZ7Fu6fupiZkE4p8cE6/6mFUY5Z900cbLhGiOZmnfYmzbn1pXFaneW8iUZ18KDnAhmzQX
qOSCTn0Za161o3cB3Pc8CkodX9cUfOwGHVSE6uAPp2A1hcI6h5LNzxsEJ25QUq+QAtxBjnCDMnsr
n1x9nOq6Qe2AP24Kpg8jFLNtO0bO+mo6qdzCReVoOJJo23gxxeODeGKDgxxIi++IkLKqQ0Rn0dBI
73mlhpsmLNoxi1jxoShe2QOG7Oj6r5AfQMA+IIeEAaVrl2i1lZd95Offe/PQ0tLMfumeZoDOMuX4
MBAwd7SgU6/paDdw6PYtIqQmmlYNexTkPrAGX/spnzJlyqZ3o6LcrYZ+fwDJnJvnV71+LP5fhyfn
qRSeec2k2SPnnV5bfD9UuEdCmHAi4ZNeQcR6TvJA5sBB9L5KT8u1y92tp01EgAeNGDuKW0+aouD4
YtLSHQuzQTDgZZ4yj4tM334pCWVQz8Ioxc1/hYydZEhHy1C2nArGtiKCxBNOgaM1AKzTSpMka6w0
sX7PEgRpvv/haROT9HsZdbehrK66TnXTutYmtSQ7tdNoQbsoRrz2AZs7LMiYFMARSA9CAftuPF0B
LY/I+HYjiOYW4ILIhrWrJV3izXwyTpf5agfG9vN/AQO2laNkeAQOGpnVm2QJhfA/qsp353bSUaso
268kDi2O/JFvuadeadaK5HhRdt242gG1ebQ0RDBvdk3I/bea6v9Y0hRVvdHABteQMp/SfQgEyW5Z
jJm5b8M8USjmAOl4OI+g3C4VFjIwih211wx7s1GkEPxTk/QioKz2Rk9qF3dtq8Jfv99JjvSqLQXZ
Dh3ojzkZ5C41VKjYCbVPGAaT8rVMiLRYPbDCBMBLNRm7OUSxh5L1UdrrXagt/i1U/9isdXWfqaUF
ZFvUA0K2MFIIHB+97NTI3oqRVKOFk7kLxmD8UvAJErRwBgfQ5IN0M49NOLSaQTxWU8kPEkP39aI0
PX42swgfArAIP4490bNWNbPgFk1Q40u9r4gvngjk9rJ6CfIYMNH3OFSI5hkybrAY3EKSteTyvNZI
YPWKo7we5d+asPl3cZm56nUnZTqDN94x0G0ArzoIGu0+6A7ZRfNaFNPYxy9LpicfNY/7eeg8VAFT
8eRB4exDTTSAuJkwtbWy3BeIbHOLwpfTlVIyHRbN2Eq82yinydAmrx2KuO12GmeVgbtZOvnicpNh
L0Z6ikgTrrVDEBDuLsMl9nTgIGCqSd2TnsuULTs7O6ivv6kjZ2usfWelH6uaMMQp0ligqgLetAcr
H/gVKM5KY4AuY7ERle3aRvYmNPuRwFuNaDRmAvKne9vxQQwVs1AjSniPBwSYGBTWVCq63b5SQ3wl
Dth8JskAwEnGjkv5rZj+xBhwV5cZGdORDvW6bg+MHeULvlUqDWi8GUzEJGtvQ/bIKRZDNh3Z7arq
pB1T2bM8RII2aCUi3XrQeor0nbPJlQqbnTd3pOM0ABm9W3T2S8eq6rdHSz4s0Tnao5nmJf3TlL8Y
l6SH1iuXaRTmRyiZcFBgxA2l5IGyLvupP8o9ZQsWC9p3YCThL/lQXvK6l1Vm+/zMyzCHtrcjAaJ9
s8HRHjBfz6e8CHrWuwn2m0PqU4Yzt4Ho5eSr33B25iUFXVnFcq2gWjmy8kjMj4uVRaQwW2j+v3FO
hpv1wkKpMjALpPS5OQGdoSq9MduzGwOiFm36Hz1zYx7fPNqeceRbJ2UxvVRYNU5+XwU+ce7OloEZ
Wtbu/o+rdJsSou28rgaMYS/2VfD67Pl+sIVdsYmehz7H5995UmszCfhqyUi8hJohx3bd7DrMxdgV
5nVVrw7Dkh6cjusbRka60JSC674jOawp6LY/IUgu3xXOiO4HT+DHIuCvFAVxVVvGanjalTeCG35H
+zhPGt+JN1WatOWJwgGVXJjiqn/LAFS/qL3lgSB1m91ODx+VV9+YOIISovyPig4aCyRi3n/PvNMj
5draGK+ei+nWFeZuu8FfasEcogoSiHDs0vu9ivU4eGxyvbImxLgydRVaTE5AY9ybvkikg/S87BPs
N9dJsJ79wtESFoh60zw/yA0+fmQEZNaWdnTiQQHOyZI4KgDofmqcWI+KaEWKRAKrqumtEYcctW13
aEsve65FlF5j43JDclThl2IzURNFbsPGHcDH9u4k9+39N9UXBgV/Wgma7fD1HQR++roXhf6rfJK1
hrF79ZmD+qA/zi+b1nYwgc+y+AmbO4zq8DDjdz8lKk2FovR4lackHV/QeVLGDc6uRKeIF4lhKAY7
Ls5oocLsCgmQ1bCx1LTrtO7Y/lH3XF7CflR1Ap7x1CIQ3S+LN9m0dVv7PvKlIVwBBrVN2tEumIL1
5zGqMiK97HUu+tCWjOXH6diFgQ7OdO/UBdbb8Y6yij2ZNHH2z/9yg3PhxavxKaHdFu+i0Bk+76X5
BJQvq2OxbJsI60Mf7iQin3JpOAQKnXBiEhPG7j/tBt99MpHcHAxvOWZcBWUTu2W9yJaCYzWIcPSv
9v8fxpd0bd0/GJTani2Gr4ZbEYyHY9uxLWF9+PFuE/Dz3D7nreR1Bz2XjrbMUkNzpsykg/pb1Geb
LB7pfWEEKyiD5r37GgFIDm0ptMk6oInfg2GR6J7CwavcDgllvuz/4/g+C4sYMGs1e3dMe8YFCkvr
2y13Z/kTe7eHgldsh6bTG6eUUs+cqfX+XjpII0BFrMblNek8xk5+TPSWbcONuu4H3mVaR0d8zwO0
xqmouFq1A/cChaCn3rTcA680a9AGkO5L/o2eWUusml7LoRnHvf279Jp/7YdSyA0R+FxEuCgnOBS9
L2pIzZQqtMv5PfNRTy8PLsHnaGmfIAy+c2k7kydgGZ+A0DxWA6/Y9tJRNLvXQ4ZJQQjHInGtwk12
q+cjvyySICFzbLZn2XhyxS7/JpjF+aHoGP7rXdegAbY8BGto87Au3IT07S1PKMN+B41Y0GYF1IgW
2cT/Pm0b23qX6wBTfA9J/sHhT5F+fr/d3Rjk/faScfDUvmFUzeUY8TddieWwtG+vvfLTMolRaJoQ
RgEnVcylyoYSiheI0aFnva2oM1T9YFWEf5VoBmjaaoIT7SoPVbFXm/EbnbIiQoZC9bLQeBaMdjUU
UkacGIy4JnNgdb6kwEATyQWWrUxbcVr4/oKpkxEjh6Y7WOlkuudbEdvD5xf5/y9L03OmUqU22gFb
eJuKrVxZkZxoa6lQEsvsFuiT1TJ5Ds9SdogZbun6BTse5vuOqkjTlzK8OikXHyY1UfMxgoZOjB30
Qqh0jWEuHATUbQZI4UZ1WJSR939Da/m30JjwmR+KmYKG1vPNFv4OHl+X/2RJkZfcsDRpBpPoaNl3
BsjMestCRw+5upH1FbJRlJyFHOrPf176i5knIuQJ3sFid2yf69CrPfH1as44SZSP/d+TDIMQXTEc
UK/aC8ZGNECYG+nugW/5c3tK96stqenTXTBzgZ0+0LtUbJEMQmL4AwoSdZyCD/rbLz5En1kbrn1J
RIZ/kicaXnNXOcNp+eFYmg7vd8pp+W9jEE0fPC33EdkzPvwWJhTQkDb99NxYNJN7UCdglWCvLU5B
HStTrgYpqye1BF5S9PaLF4qY2FsB2UrNeZV7oKG0oR0VMFZiJdBApW7dJ5LOHKJ5EumDsjIctgYp
6qhYb4Mh2kLMMqDOxdvhzqmASok8aLs8JseXY2w/bACFcz59aFrFIDFHOLRJKvPLb1SoO2u+5sEs
DclZM+Y/E2VW8E3rtZJNyVNMPrEOUoGigCcK0NWcAQQtgEzhBQuhzpwKt4XmzvHBKJMo8beq5GU/
MAdV76NOvJZtFv3woWVaOswCTWfrn9Ky0WKFJwaSjQh3KNT0h9K3lkL9qJM9/Uiozp8tUamhrH6u
QewfVC+SBrot3LaENymIXaW+pgjppJKK4EdI+C3jtoWcARBfrOH3Mn82+4+LTIZxmni+3gxwkasj
wjImLahtPqqFFhWcG+yWZYeAx2H0EkQHMX4WzR+txPtyT7xn+ueyVWeREJHTlSPd99V/20w7iG1Y
SIKxIJO1MPxtNwXHp6INqiVlMxcJwL0V5qX/T3MHaFcwzgIQxdVIU1r0iumDdTnu6yFiKJzle6Si
w8ScnXfCm7Iy5yqxwjf+gs9qALU+C3IOJPSawD6JcDTxZfyKEIPNCcQS2Bv7t47pIeOr2r6Htjwt
SlKXEAkiBwXpN5o6FPg3FZGQ3BSOgRrqrx5DzknxiWhplauFJfFZrTP2Sr2hYTICiucJumCqD/cI
05PsBTxNMGNrBtgPXVqYP+INA9BtYTzfJjDUXYkLjArCTDQSoqMkSqKLnunG1mF9LjQQZIWqON/N
Y5Y2p9GN2amX4uZ2qg3NHBtKnXnQwKpRWS3JPyCmyNuftbdPZcRZcy/JPvFLg0aWsptI8DvIRKq/
1pjW7bu3aSaOxfyMH1JELs/znEjJyGiD09O5LszyNRq09hCJ3A0MgdCwp5mA6zmgbF336Cc/TiDj
taitphvQHA94me7kAMaGj2DQBLQkKqn5PDHpm/PDyj2LBLjsjIm41lNsvTSToZUJdF1JhIZoGah0
fp1JrWw+vxhHIdp2u4qHsNLghGm0UqvP/bXxX3D68/hgfv38RjcrYQBUxoIi8CJUFgYWfBrzBaN3
EpbiHVOYE7nYN4M3Te2EOgAxCNQV7ZcEiTTR/6i20DuoMmgoH2OSlu1UEbjxxAKQKCUp/f6HdE+f
61ifu91YWCZMS7tqX+PLG1IfrsduOUQgZQ2fNCQLRg3QYUa3OiQPr2jYiS58AhNKKenFNee9/NEG
N186Qt9AkrO1mMhAQ0PWZkFP4DUSNELSk80gejaDbc7DqPpdheZH7OfArA2hbrpZqoEJjH0tmsb0
XRbNK9ufPqc0khiDi3O2dOTqIolvw4T5U0Wx6wNu67jha2fYrHvFaXNxYrFXpfYcJXXsMQKKeekG
3+/GUmwmJOIFPs7M9bY9/GvwkH25ZGmLT8o2M32pjOXrFfC/1LJsR6KdtkDtcLPuoA3v/eUAFGXa
h2rrGma+3Ed+S5idmxV+6PIDjrZfa+sBn3tpag9ZmKDbxf0A+PCLUlHYgqycu7HftbMx+RxLmAgE
ztzDkVcxJgV1piCW4V4oGuMDPePjNK/f9XxkTAlXTn2Z/zGm3Cv5mVZBmNFLI2xO6tLwFwPkAhDI
qCDKd8n/+qDTSM3Vgg+1Dy/fL91Wa8S9nJ+V4HEO0v2CeBYQ6GYmwqiO6vfsvGIAWASSxJsQKuL4
3FvWqW5ByLQm/YMysbRrV6g7HYixDG1S9zx6aztdKe4Y0DRTb94jYI6lf/STwWka1GQpQUcItHKV
dV5wy+48csmi2XWAWh66BooHqhbb0ZNHnFHQc/TeHQo73DZMrJOj1syj4yp3Pebtawmac/5gAg42
O9JZPUxHX05fUqCaUy8q6xOZcfh4cLOS2tNgpkEXM7pkh1Njagp4/384lvMh5Bfw/Vct6doCoiXC
xtfLOgDaCf2AWp7IAOAoHgAVJ47gUZrJIx+momQE9oDilhsMFscSERdUSxv4/ZYi4KgVPNSI6oDZ
O1GB7kUrD3e+aRiyPJZX+d8texAGFjkisIwMONYmQE+jVCsUQiIOvLLJq9jJrJLas7niI/fVtze0
9jtkykQlWT0PC5oHdu9xIgH4LzaFl/EggoCqHYGyIX6QcMZGcrBPRwBDZu0qQv3J9UeiRRrPLJaA
jwCRE8OQJNJ81mHMvf2vB8tzGpJHAH+dm9t1rbng6p3HSqGCbq5TkJYiTVL0zospp0DSvoLgCDpc
nrAJEbvIAWuK40+BbHu3XRHxc/i40Ul2RxT2IVgbhebVqQq4z6JsZE/bMt20+8d5iZI2eDC/PY92
r//JF4TakiBv4exMytXGKgEGQHUk+8v1U5Wnje+T0UPGFJZrhf3A444gHb8cX24udObLy2wZ504p
PfTP+3ECalc7nWKQS78lex8WfsBwWBA0kmSqMBcNq/3HeHAlZ5ZXhmoljEq3DKgQ/eP5gPRRX0QD
RJdG0apegCPYS0CtqyECUTthkjE0XqQeTQZNuPqn7mAppGlYQd2cOwGsKKUyit8Jf2Q2kBNQ2IzG
EuRHws4MOnYzysv27Lxdy62L9/f6i80y4ARILlNNBjQG+pEypwXMZkO/X+HQ2rrMmjTtRZAWNbNA
udCek4sQDLMz2B69djdO2lDL+bTkCHdNLNqmuq7tkhnopwIg63jzZHUXwyciq6aMRaLsmc4HRB2e
eCcMfdsAb/BWblyJrkzHCOMnGqA3xjRLt6LqgmePMpD5jMYt/1vz6LLh/tOdTuOW2pkZElV78yHF
hRKUldgSinVNViow4jHW6UYy8XLYz1rgd9za3AQ9etx5B/QKcdlz+tgP3JdhKjSWaCpJzE11fwZ6
h3nCr3lPc6h3sC6KjRXglvmZf1tmdAeCOZ6j3V1/1usygqhqS65w3GlEfGv4iNn0oxiACKg5Vc5H
UyBPELFQwzKFntVD+p+nEbeGv0RrKhztTWffxX2T4P08zegt/jw50sfIgFyKASVJCN6l1OdMy+D8
daKtGWzLXZbuBXsuhPHJ9YlJHOJZaqmOBilupTIY9TwJhhFEP7InwZEkweunNXKVrTgq52TaOkq7
iM9QxDD+IGrHR2vdgcppVZSrHIs0uWbu0AneLPbLdivR4XzvNjXFiGdTyLJkcljhe5aKNLDi/oAC
vr3k9PgBvf3PDpGfSLQGaHDXAGJdibx0RnjrSM8WeusCuHd/aJggSTakvzzrvIhS1xaqLP7FGP+d
jyElEC9E2zImLJFUSBO2iUd1Mf2en68SNUjAg4nAklQDO6J1tQG70kNYE6VK9dHRLMYW/Ypnf1rt
YD/XmsSyK4H3i5A3zdAAPNvHVVpCpD2C03k3qHRpFIDB81sEbjlHSukzhclW9DSP9E/kAJCIuVEg
hUnzqL02hXX3F4W53blYXsXz58406sbty6NYWfnDhrCBhytyJh7GNmPveUf5J8TsI9gAh8BEmZd9
dU+ewLOS6gR+fKwyFwVnRAu8/87vOc7lUaMl8elqw9nbiAKaOeH1OCVtffxH7MbTNRZS/5COkqrF
7yneO8bXrp0fmV//Ir8sxt5pXWcJGHBGnwUNeJ3ewB63eAgDBmADkBz8TqLwkk6Qt8LsaJP1D80R
elAVczXDT9zGhxNVinxw9L8qOQKoQo/PQvp1tKDxuFSndkTBJ9t6fkEBI9efw9RPO7qmRizuCPGD
ElUpfxWR9ciGbbaDP4KIz88FiMC6w82TltSBVZTpEH9LYeT1iAuLdpQLFRXz/FbAn6M7D5AD0d/E
yuKIQOWBURtMWWjxLZRO1HLJ8lzJF+bALp6ur6IgaSgR58bIuxMN72o+/q8euuREZlMJwkGS2IIU
dCyUC7mObKTswsUxaCwA+rtGqmPV/i9OlA2ymvOkXc+62c04YgiT77XFlmMOx0XqTJHfa48xs+ua
7LN+XFawy+7+qhFEvI1t6lfjNJovjPbLSR0U1RX3EFyx7ryHvPouOzJNOF754U5QCG+lJw8q+l9V
sA+vEcvJjiJcd97ODaWQSVjFNxAKWUj0FML2fo5r3kWhZW23vGgO/MrJrZUlv0NbfEem7i4q40/W
VwzjjAeEREJn7Z93xyAhkfKBHHrU48hIxpgDKwsrNywKohuurmmVSW5UBbFLvgAZCLIVeswdLJJP
JhCvfOHbtwU/qJ3c91cSNP+CoGEinmvtmPMVSgLKVKRv1v77NIPuoXyJRfrKmBCwSeB7ekYkkEyK
BtQnsWLcVsa/5qhm0G7j3q+yf8lfeQfUtM3msMSXtpP1Wt1ycfOXqMjrLIwJBVU8ILTT9re0ylTH
5NAw4SS3mQ5hcUbezrd1p0ANgVHKkpCh/QQf/VI/jm915Nv+i5JtuiDYaf8n3O1ABaPKQiq+ykLj
6v5Q/gEya0cjx3BxAQD0DwP3jvIxq0cnBoENf8y+Qbh5KI3Iun2z3m/b4iIIwZ3ITKkOuxMGVl9g
uKgxxpOwHdId15WY307mfAhYgCP8rzoo5Tpnld+Q1M0dux789IoMvhFiEkvif8EU78QBPPo56HQL
vS1Kpa4Rt/fhIp5+Y6xCtGHlLtJFsL//t1tgWu5SiATVx335gwGMjwzx1+egRZ4JrT8THrPeAAZK
wk6pQc/Wz8fAyNBuq3SXbDOLl2VUmRtTrbf6vhjligZgog6JCosC5CKZRbdEWMmRFCGL3EcOwsPY
pktXf1ErYGyczQXojGNw/Yn6oZ3PpSWknpq/GJNs/VwO68o/Q7H0oHWEHKGdHlzlWMuvCK19ES7a
Zk74kSl0XmMg0XI5ueyodvNjmuvpoGJ6m9M4BUEYEAn+paC8WxAuWe6tzGuy4NI022Xv4iEK2VYW
9dqhsh4X+N5uS8hSLndexrbbynVId2AWdO5RMYpjNH0RoAaxNAWQ5GlBkncJEapTNF/XJkJrpfDh
zSHkJowmBQdQhYbktzMkKwv8LAYIaUEuJR3K3Rx5JxF3l6+oQ0vXoeBUnqS3PieZ90MIHsMfR7y8
zpirWQMD3zmfKnAPM9DTV7ZGLaE00pH80QQzec22PC2BDEnXGH5/hl2eCWKQfs+MwiiPx1MNiOS7
kvVmcIl33L5NQaf07VoLlZIhPdwjmE5xCxww5y1xSPvNJQA1qgcVv99WanD1p7j9MeQ4G1nPKVKv
V0TevpqrweN2VVE3fp82JJu0ivoK2uW9PpUeog4p7/5M+d9u3/T4+gYcdurjN2rBJqj+8Gsl1995
6nYX7rj4U7Rjv5pf4iKZsOYuzHBJsE4zmcvFnYeeg9eJFmcwX3ohV8ahL4jXpnR1uV6rDOJ0QfeD
Gxi9If2jDUkLhGT8twXkBFcFLeeRAMFDnZUE9frYr+AW0CrcGdSkWjPoi1tZ/hnDXoNYhO7rSbY2
L+FGnhYYlZ2yOWUwW8t6QpCfYnEEwkKhfos1/2FN2+MDKzD6KCNytTunYUOzsyKPiFiQ0Jr14fn1
7yxX5JUWPi8CCX9QcyacyiADjEgZG4mcXVySJmJ86t6uIog2CICEfhdigiixWMnEmifs/DDSGd8T
3rkcxxYZFxa/1pfDKZdlGv6gOA2Va2GqFeWBKVg9dmV/wgJpQUFwJxxztpkepXdC0YgOEj64f71k
QmjIYVtJM9lGmzIn6BNaeQnumWd0pdIx9PqnfOQQRGkePIkECNVoHaxRpAKCVndbYQvjnzM/yhy3
7J00THkD7UwjKQGF0b9Kj9RCfVrKTnXaNKDiuaTz7gGXZHxsFHNKOtGHNgt+h3DFZPrUZAC7h2v1
ksH7D9ZdHtZ92vjsA3g+uTpIhlYCvkzypLmddJJEkiW/9Pmf/uhgog+gIdE6tpKpuCdsq8FxdNBb
ASTZWADdHtpaINmwf9UiWrv/qQmyKUZne8z55b5X+NChEx+hYlogLXshJQWAoYZOvkL258oK59fJ
yVF6GUGMWMcpJSddQxNhSl9ScWBVM+qligbGffQBZWGHctsAIiGN37H9XrcaoyWiUls1BdijEYe1
/5UIqApLtx1E4rkEf5XZrk//f8fHTyrY8cHOXxosSrUFVoyQykJfTOCvW0v0BNMb67mB27+sqVhC
KwblGZAIU6xDU1NaxKEa2OZ43Yqe7noVWXhKZfPEiVtCBozPI7IvKflTRK7xBY944rO9ssBBPXUf
fTRzSOh4/sGk235YApmyM6dUJG18ZBPLheEzn2pYMT+3RnFpQ+NGBdWkFf0o91CFi6nNKcPqVrfF
/L+pinZ60T86Jh+gd77AOsbcZk/x9ug8380+l0r41U7IvXJXRf/l29BtOu0B1TlnwEIjj8D0rqgc
H572jGRUB23cM/cN9Dvy99L/fCQ1ggkM6a5dQ5TYl1FJbsItgGy3az5+dxii3Pup6gIY/TpdSzHd
j2qpk1AEX20s0csTRUysjVv9fLLwGDaca/FYvjYkMC3Y6exVsF+YxSEi9H8TM2leyjZrOfYojK0j
cz/oAcfIke28zJ1YbTNkk1qzgIRuTFvxoKniEPKswTAMxzjxvE/yTVIyqy+DFhUIxi8xjz8fK5Ay
CGdcKMNk4zkvVatfAcWHTc8FyGw9DhDUxb/JqD4/mihayUIDm+bgucPprZ2q9ine6otG/WnFPw3w
9+IytIaY31pKWFKtcWnw0lZBVOG4Paj93hIe7QyHBdhOSiR1Hth/YSmL+c1yzOL/tWsdM6mzLV6M
ervUg8HWxa/vh9zUjWUdZF5FrsM7b8xJwnLwcmAG5KGBch26/nvnaz88tdW9Ssjw2n0TrVljfiKf
OuXrpIjKPPD9vbMsmF9aNN7twnjLI/cMX6/Nx5vnqFoy++Rnsdv0QKYAsnEQIVAbp47b3rLFim7i
dbgXZVH8g+e+JWUYi1sZDAltn0QqEkbezXtgew8doy0c0Kxz+vCRZq1330D2PYGgGn08QNckrbrq
Bqui12AAKqV1gsrTnj3JtWWggNV0qmTpxoJhuHwMV8KaitZa/BMClZDS/mA85WwUSLmHMdmumS1D
+EvBgcVlMsA46SXvxM+8PCYT3MgUta0DxwS3xY+JLpWONjTUF9CY6uHztPtNR1YeBN+TMunY2Sh7
pd2xyB/QwrmyIeyb4/0fZ6WTL5UkalEzIysLYDWVBLMqnz/BS/ZDZx6XKi1Jga4JUQHuQ4iixEQt
uShrdqvnmxnTSnZXkdCw3TfbmbPrV5zJVFgHNSvxp9GGu/pgU7efJ0Eo9ECd60c0WvJwgjhThE9g
L5Bx83Rc7d8fD57TFwt4ez7TKIj9cCtEz4BlqWHWrmvtWAXrCmjnU7FLQje2RHxPuGWEwD0Ytz5y
Iy2J3WmFdF59rXKvDqdmevb7WFm6/zjJnUPEkZTZy0elTZi4KuU+zAe9TNvF3jE1iHTcsoe5RosV
m0ortmJes9AKQ6249TQ9PVRT6oBygbFZLA+EeeAQhkXjsgFpsPoPkwS08xEKMWvSLSlMNLtppRiM
Esi2nZgP9AMNE6Fh9z4jZxAdo0gKhg6cuH7hgAnYf/+aP1FB5h1AW/LBT1VnUz11v0fMeWUtvRNV
Z2lxzi3+WztmdwjbZmpCKUknLiGoCUbxS8v1OtqEgZh/1a+Nks2GNmFiDZMjLeXu3l8JOSQ+V/uQ
Ibp90S8HrnkYqIeN2i1QQLokJxFKreh2mxAXQTllYvex+e0PTWVamKBUCKVwbJMMiDp+xkapFJ6h
eUTTgVb4FpXjibx2DTH0xT699/026tJR9awKUXEbU/seiSuGK3QUe0u7UXGCqUSeieFZlPQRAMLS
es5yK6nQZTuZsUKzxL4++R+IY/bgBN8gTaIwcvFXnBducgD82+2l5vOGsqATb6pTZDSb2DFpGP8r
qxfhDJUtH2NfKkUywKRQSydTJXQb6X9yfuOFPl0b611JQly/vovXRGOTnLf68zANcnM0RtK1uxqY
EcmA8FJ4lkgOXU9QX4HciTs9VjwB9gYvCjIUz4scPVHTKGD6vZdiVDVVz4MKSdEKPtdcO4JKfaVh
NlCJhdUwmj5wpa0j7aGWVRU0Yd8FVYzoN26KBExmtC9MNxCPaKQ7LaZGXFIrtCnKg53VepX4NmmU
iDUdIFkgyDxdY/GrEb6t6FhYW6OEM0IQ6G58yw27O3PuVTIYJ7fYm4o6B73J3Oyn8rn86HDlrfwp
JnxSaBWJ1h+jsy4l333c7q9YHoMky/PHGJyQGUascYWxPBQ98vv/cn7Bd5sJTbhsk1pb/fUS4Ef8
5GXD0EjazbR4KCsjAjrcuXHh3KEKUTEDtAOk2E1HkNXvWUpctsSYNgNY2LtEc+z33WRnY0Kf01xr
E/vlPwXMNvqJg8GZqoJIwPJZXC9YC8BEbbloijyHTLZUQvneaNFcr+W4ZeHuzJ6YTaG5QHy1oZIQ
uNHeo5XfhfbseOWt7Urn4hkG1vRyn3BQFfva+Q7PxnHfK14KUFUHs7m/QZTP8Bi6ErhQWiha739/
KryTBJS9EkaXBtrMTBqcAihKA6Q2pjz2vvcCJih9Oj2yVkrC6Usofy1DgDG2uD2MLHd422KqVOFS
Cg61sgBnZrmTQM+lgtQo9MW/TXtpV3qvMQ6TVBbxEsGBlYeO5F8oG+uA9TDdMMnsZGYIg44JfkQ5
H26o3mLvVvIhv7YHfXR5zXys0W5T1QYJEyt/DuVNHadscKLODd8ErjVAGBQDg3QjVrm6e6N3gA1q
XTXX53A29/UWgJ6kTrv1TaY1p2IglGEs/X3YPFTdMcW+oPig0MTNeCkc63/rq/29tNDXc4ATHAAE
i5zw8Is4g/qTsWuH7sUKHi50lenxXhAYYSIxxlABOchDQ4KoMhVclaMwDt7nysatRbqf5+uWmIac
/J/CulOD7WC2p6RPnS7SORXlaT47K2+2ehNhN1d7tuXEW9C7ylIQbpMA3uzEbe5hD28GhqzF7zJ5
LpvOuY6sgqCm8uBQtHVaP7bBW19R48xKZfETjt6IOkXL47WUvU6qPlhHKKSHtZNWYsCOw59ARcM9
n8mdUPOZQsOMx/gL3zhnjhla8GTps9LZnByAPKpF4yfRS67xHVr7Iigkw76JzOVfrrCWlVci5GIm
MeeAG9yTiOnAilZGEnjsM+X2AR7UnZk+aGkpwJbCs4407G0KxS+rF9oox9ge9dGWlOSrr9UVDffv
FtxMHaXYEDgc2S4s9kOSI3VN36f+I7bjZUd23FYuVcaLU6aPHd3wFFCm0mZ8Rrl178x8vbCI+QkM
dFCiXOfF4tOOFits7VoGD1Bs1tfIg02CcpT1X3bAtjNkRPiVNfah/OA25fjIvEPfB5IyDpk5iNi5
VyIx+7OhxtFj9nyibcuDwYwlxlK4yM6aN3zslgiIQiQcktAertYBXhccjFqCiqhO5uWpZsODxIOR
yN/fnNUPNyWRO8H8v6plo84B8URql8VcZR90L/74OxAAh7pbTRs2dBx7d3643bpcrZm2zEPJW0KJ
HKMxfFDRP7KnVzjvZ94Zbt+m/U0Mcb53cXa3RnUmTNmgEUzDZ1PfSDXx9YKPhRN7ut6ArzkSl3Lk
RzUPwmtwWL8ZQo7JrOGYlyPiBH8LWcRfNI3B/mNwbBSWgDteXbRbheoZJLM2BFSI8UsoDnSQLUnl
pPLZbWXtmwvKME6fz3r6qZWwjYZth9z9vo8aryrDfxs8HigLhizk2kHGSzHcu/C5ptT2UTcN3ti3
CU/0+/z5wPMtlZyRTMjTVLToydg9JgYlvOYA3YyTjeiIQvZjddJ2t5A8PtZ2lf7ow7WQSiLcYUfl
9A/nWgn3Jm5ISEcLqgvYWvIH4YkEHlYlrJpLYv/Qf2ZkfbZDbse6Lg+pbRvTN+neK0u1Mqb/OioD
4C/6xAB9yd75Wud0aoyLOGxjFXV8UpwiIDE96b7nn4nExQTZH/dZPW/UZI2zAMzrP5iH9cJyBUAO
I0tob8be3BAhzPGcdzsYNvl+6u/C08u7Fgw5tS0lJaOniAbSUy7ha/XcD4I4UbzS5EtV2O8JxmLx
KADhmO/mSQGLBm/9cbNjmp+GFH1Yvv4okvmwqkX+kGxMd1AsyRXZ4Yhv4l4R77qa2zQLu2ElMVtO
Bb4KVGLG22qhXBx1uNcInSmYH1qhDcmO93YSi00XoliahS3/SZgbQOklk97EWYvTUHHdRTVUrpJw
Aj2o8qU+v19i9qlcqs8zhOsvlIQlzauiXrlnxBvqNbzs8RJEUHRpXxf9nXfu5e+gLlmAvEO/JBQz
mfZD0RxGIOvtwOnzTRzyaNIPDom6aK63FGlbKZ1NG4itEbM/DgCGOJ1hxv0hNxNGiuagj5x7Mhep
mZ0iCUBhX7Yd/1XaIzDCa9oHK7jvO8WOIc62+5fraL+X1tSvLeD7cvZcc75NFr3DqAMdUoSYiz01
08NiZVkhSTTg8N9SxkqfCaDzKEJqz/jWFgwaggtJXHWB2nIbvWmyELPlnm8yicTEguYDcNLlcDB3
pbPqJ2vKw9sQCXeGczzDeLwuA6n+5qOsZrrPO0fXdEPaBtRyr3DBVFpgOEowZIMQHjKoMhXXYQzh
v7WgW5TxRLYjSTBZPFRyOFhlRHgTgudAb8QZw2AesahNuRf85uOK5jL9VZmE1ie/cXDczzYRhC2C
Y8ox5XbPMkSVgithSs8yHLuRwb9IWhcOQYyZ34nkTmXxZV4oz2YXy6HC1Ex2QaJhoPWyPP3Td8gF
FSzTDsKDejkKN9l1KgshBGVnk5jx0Ioh8KePx786QagCzX8u2vEjSrpSKEcwfvm90tvRzQcMqsKb
v84fG6ZY9xL3z+Je3upI9Lc47o1tl8k/Ps8S4LmO2U+EDJK5ba/t570r2xJaj2XkRjDUK3y0uZIC
1m2MwZbbzZyEK12sEfcW1vClftSgaijjchxH2HR25oaZfHUhpf/BYWDkjBBB2Sisq0TyqJnDtcMj
MCi3AxMNZ8PyysLepqohpF45wN9Xk6tzDaBDB+URWX24+AkZ2Iy1oru2KE6YxS6TS6QTRTxKtfjT
B4KGAcZLX681jUZ0AjG28XbJ4I3FSwRWPWn8jln0mDOs8B56MhpjXuuzyKwlgn4UmoJL9vZC11oy
9CqSSJ0AOi9AZc+AffdqL0jkqYZf4aJVPOAZmfLIoPwJxaCVLo1y5kz2PLslvJgSWSszrQebFxFo
ahUqFRIIuJSPNLrdvfIk5sBwnHc78TRc+VCAsarhHbn/Nvwc2yX3RU/V1o5k4RQhYxRf4y3fJ73F
WU1JwN92KSyoMoNYx54Rj7F4oRItW8sHrpDMVa//1Gwud2KYzCtja3GwvCc5bF7LX1h5B42HJSNz
IgncD3ugBTnNHDLOw4Dl78StHpJBEWGjgziYo4w1J53Ib50+Pb3UsBQvvYBHlS4cSHqjF5PlKzPH
BEByOwKZjjhVJP2+Wuj7ET+y+4hx7PSQtm11d2ghp+0KlGtH2Yv492AWC2QXKOebN6PB+SYV8lZO
YDmpefhi0HkfLn2zZAmzu5PlTCGoFRym5bG2+J2c3BSE+VFvqIlCu5lbKONz3dT2Clt6Ps4UTzoB
BlXvWAPhrj16HCoyfvYfuI0Nx/DnZU8PxPXubGyvz/x5cLQVKiAT1ICKZrO/evv5pQ+el2Dh88xH
azBGwwphHH6HmETsGNxN5TC1X5aNO0AihXp3jAHziuvx5lwjFtG31Upzb/kjRPCEZ1b1zQuPkrkB
z38+JZHsxbTKLWIfnPoVms7s60p1kYJesHBG4aZTQeBZaCx4r7Av6FJKbToZQ6aWG1Ue4eYBTT+s
zLD+uwRNzp/FyFwPeWqwzrY+/FWt9wlMnROh2fzgLdZgV4rt4TY8KtKECICfnqRUhyFmwpks9jpq
X8MvU8vW1ywOQ3soa8FsKzpFsFSgiWe2bK/3plcmgMC05PbRvuTOljTHhEpG1NSr0+YmJjRfTeDI
5y4dwMFkQ+JvUFCN6AGFlpDFiHRfcAPKv7SjLBLPF/VI0EDBtH/OtogajG62BSBFi5wtZWLZtQRj
JVppTSJBGOmfxnC8FyUlfG/JhJbAAdF7mW5cGdDBqPWH7+EW9/ZTWaMQ4RNuMCtQ1nk+FVTUEPxS
qocjM6OxeMhWYxi4b9lCJBhSEnstMPHYti5EMPv0L8bgXp6Q7imaJomEDZFzZl5A4QcD8TdU3TeZ
kv45SaJHrMf7kyLIt6oFpKLu3qTCc/z4W79CkX74+66OcWSOxm/iVDqnOPsTe6B9/ubcot7a4PZp
3h4mHsfhPLwtUAeqqm5KssALv2A4gf/5ZZQW5qpqt6UgWKvNjg5Rn6xOdB00q29sUYZR5Fs6WsFS
oHkznxwIsAkBuxXPyh44hOrUvg3eU9WM2GOtepNUIknIMpWALP/rbnB8QYKojYTFG4NM/6b7pWuM
7o/F0uMx616M0tOZHrKtL+brRQ8Eow3g5LFOFOGiszIJq6c/9tBqQC6flC6fWo1yVMgXWXIKpATG
DoWydxdV0PI11azHVl1cWT5g6OvMrt1lFQGzubZ8HDqEDjOIe//QI735j6qciBr6N354DWJb762n
iaujl7N5By7xmSraBwxeRVkjhe7XHpQLw52tE31Z97dN6e3aARWtKHNBQoJ95rTKJVf3ZWtnfNFk
TW3LH1GXvmvbBvq0P975T0P4ZnMZkh7I7MPXFKRN/DWCFWpNCKCEvJWpnvlzg3QuHwEYZDiE5FyK
/nc5pLK9BYa5d4sknon4u0dwF1E2Unxj/iQ2oVUMDvyfnui3qL0ThiEwnldoKTrMzoP2kv248vPa
51y7EynP948MllDu5HselnVyEAhwKb8QcZVc6z09RWIdaA7BOtJGX4oa2g7MziU8b79V0h/J/c4F
G0Ge4HVGeIZuM6tkUyUPqIak4AXZSW+EUoOQcJKnzfsaa8BYkQ4ASOrBE6gSQOK/QbM9ZQmmfz+e
fGAaIDf8+jqRLP7kvJ9uSS5B08cebmd3gz3ZeYfJQ9l0J3i9Updg4PDifx4Dd9iYFhUSEyQ615DZ
cbUMFWKy6VrsumidhpKltVK4JdMEOrAGT+2o26ngNy4UWKCxUv8OSteb424sl7y1wjUGKo96A7KD
EofaE41W5i8+6sUBJZYmEmEbJ8rLUsBYNFUbrSCKdNP8g/CKTs6ZwnN/CVe6AZnU3++AJvb1dT/W
ULzLcIBV2q8U7AEvHLuya1Mk+7+PrsVTIjlIt7bwIrFHAhB4x0fHOXYbCamWfvpkn8Cny1SeLZRP
ddGEj5oPNR9Ljofwf9EtBOivPME2qCUqI3/tAfK/t/qf6BJbdsHCOOKM7v59BF6DBloepyfxplIk
0IwOKPiwh+PkU4mKrsIxDfcTMXIJ4J5n/FUyvXk0kLdMBwBc7M2uw5w2s0h1aCN3LMjkpWhdK16N
vIhbnxKag7/DE1r6sbU7Nlt1PzrKy9zBaEgjQDujfwb5zcvnfwx6orS2C+fasC3tBKdJVmRSk1xr
5Zb33wibJNNkoMvFT3H3KK2gDZ5oAWkn8xQIg/9t55fVP7zWWlcW4iZjuCJil1TiD4yaZg/SnRxE
aGlNBezO1+MLGu6fjXrtAbn62zDh4sVsj7M/PumK5DwCfoEcsRhz/VQuKfNzIQOUmEmRgmQFd2zo
KhsGEA7L57jH5tRc477Zwk9YJvbXkVwgce06QfpTQrmyDXArDqm2s+mS8uNfk7RXd177u7QJTkUF
lYYJL1Y9fTYMcfzdbbEO5pY5m3V0fYthm+k95PBHFuhz9GbYhQbvurCwNU5vNAJnr7DkaFRA7CCZ
ElWqmceaq2MF95JwqPXfuZy8UKn6fNsy1vRJ7ELL2OIWIeMm9ea6U1ZupbKyTZz8qWGpgc2po0oS
AOc+hC1lYBqkeY8XCn7CYqeYzMKd21NIRfKYqO2V0Z/HeCHYaqxqS+pYGg5JRO/O295OBI515Pds
wZuMQ7ci9WJQUVOij8ndJHkbtdrmTTV2hUQr5w2TCGiZL7kuPGAGeYwOVik3FmV9j5UWiSUzcA/x
Rz0pKhEBPiO+Ralqu+SPE24tNkbCXB9KUc0sQ9qeN87uwju3FJU9J51cmc9n8Dn8mzlcpC7RB9xu
TIMsNwg8w4I8KCJ9QlJlyk4VykkhjUA2f+VbzMtd8OBg6y2PHL5FwsB1XiaVOIDuUQa78/4RB8QG
2QlGyoclFlA+U28jQz3L5ir06RTrdcKZf2Wqs53+KvOTRjPgK4ceLtJet5IYuwb10IBxKg1UzIIa
Yr/Jv0SG6iNCjNmLoJ2PqWyzDy8V5x2/LXnlqg+Rq2ArDai0cMiBcSAV8FhL9RAFQLF9YB22iRGW
7kD+fg2eYJF/Jk+0ZHAJrsHf7BaCVl/FbkGXI/cTDKFtcmZ7eatiplvQVmrfHuIseu6n835y1DBn
7dXJyOdwD6+1aaIIaGc8xGcFc/eNH5XN034weuyikUyxLb/9czhhVC5d03BTy/j2i9mhF+Yvcjdd
yEyGxoujnE/vzsfPHZFTF8vSitLsE284AlnWdC2zDBe2swiwHyIRyodBWDIH74emdI/QGlOHrZun
6L41sYAI9irkILcLcpMQ4XBuFIVGwP3Qo5mUWpII23yr2/vE07PgeBnh2oTQtzrjvHuV5FnMRo42
+kRRUC3hsczEQRmJ7gMo9+p6dkREZ0qVQuNy+owycMrtBUqBTinzqSGitw4NW+cTb1u4DghlzLww
eWTzeYrNpE9LPvYMM5+eh3ah04mJkZ1HuYm4LsyTFi+gw/VQURBRibx5CuH0AQ9cioxydneoFvDo
RrRmNla83niJxlExuWjlVXobINd08+oXqBPgJ8pT1DyDZHk8lfotK6j3RRmWR/RNYic2ItOm4u+8
V70Z87vPaHerFokpPjinOkguN9FD4nMYgKe5QKQwzQkXE3VDRNVumRWaAeNsbmi3s6d6/arOP5K4
x6sKK304Ke8q5YgPlH284EdojrXINbRpWZwdl4YMBSAVNZrBSz58avUmCaumphDVC1mUl+cEIswT
v/4ERFDaWpy6KiReafqiBLKwbC3g79S0X344Wjg7FWR9cydRn6ygU30ylNIDxjWbzFKc429IuTjW
9fkFWXCR/o0coqL+NYT4tJmcewXIfZE1x3qZCOTXX0Cl0tZ7q7MZnAOv1X/6zuYRoTQ+NEfEBGUL
Vz9SOOgikJ81x3zZdspYrGsN07lSx34RS1Rhsnif5HsMxV2bGqFvk2mejywwCKuxbydTsj5fnEwu
NLpFPHbq1YSXG2gQtSMgVnNW2qCxb4/hX7NL/ChuBuafYjHZf63cVQPPoWfK/FvlAGDY9n2uu/ss
Bvp0W+rfgXwn/XefmNlg9S6bhNOAbDLWUnz0E5P68kVRAVRjYbM5raEszceFeNjtFQTOZfTrupcN
6Cu5RkxzdA7N85cBqd2n8nARvCJYRtre4QHjf/AyvkfyBvqZalJCWx5T8y7JjlbHPmU/6mOzjLGk
t5jMOs8AEea3ArUSDd5Mg3Fbt7y4BBStuyx9tMDlGlZdsa6PnuKY2p9aT9nalj9TPqOBkyrAB8af
RPJK+5M7GZaacqe+zQ5bEhw6bBJbkx8SHqF9D+rBEyERLxPIsQddbArjDfWJezBrh8944gBZN9dX
osr3ambtwe87U9tN0l6GjX0LfaZ+ouFC3/KxOZnahWP6JBdGPemJjnfi1LHj3TaObReypjgaJ3o/
KF324o0Y9t/6ogKlGEb6/uxwo+2zhGI2HcR/ePJyNJuW8aNoxr7hIHr8EVABmAvWrhi3JoHWuKyj
MsgBxuizlZRM4z2wCkGwcGaHatxXfO4sJefVWeLspD+RfyfhVjxbscgkERdhBVz9NpKL9yFPu8h+
KmMsyMdjiFsZTaRyi7t1A2eGpeXxDV1T5bYCzE/W6yxLuHmG0Y4TyCg/1PyVqeJb17Fc4HmlNgUC
VzJa7iSbPEwS4M8ALSIcjiQuVeM/vOuxEQscDhDaBhj8YUGDsU/Hj/OzH+giVF97IBiI4fYPhSg8
5tR7z8wnLNQj6wXb+PlDYffLr/RkWOlUdMBnKLjQJ4azQTGJGOoTXlLymQwk3eJzSvuW8dWKdZmZ
YisH8LV9Hgcfr/esJG1Ox4ByoriTDl09vd+CeYMm1kJef1EqCuzglKxPVVFx3yjHYm94GgRb17cU
eMohE6ihJGfLdbcJwmteSa9SZbdXAzEd5dij5Y3odXYqLiRl004UWdRK9os7roraOdX7l+zbtTAx
5FXL9Hx61IIvuhG1FTJ5kdbJyNr5DBThlwQUo6VSRLHW2ij1jy1KCEIvoUA8HuHJN3pTrAaiDe17
HLdCe1a5XeQvitMZM/xL6I86XmXoItSv6XkSyhGIruqQ/cQXULBStnmz1497JdItJlg/ke7tcPkr
h/RB5FX6KJJ9+llkM6zT0GAkGda2ZhIaQzTPudCrmwFGs5W5NZcVT40zGo+C+bhaQF/jvIP1Tk2I
+oi2SVkqQzYwiMF5INkIVHuO3KOUYBdcRn+b1lGTJZXxOe7C2BdyY19fo1u/ro1UYLwk/KRCJn1a
yO5E1fDgim9hQ7AH4ILoTqzbuMARlk0ZlYYu2rnUrk8qppW/wKycT/tPaPqKkaSfRN5PMk4JK5tT
chKKT/szLPcR9tmF2KwWAY/suJGQrQfFrKE63/QbBQas8eAnVLU1xPREUkq3nW06yqgmBrYhF9mp
RTVZI5OwmADv2J17PXTO20ZZmLNV96GW8MK9HEwoFVAr2fUJAly9CbwkBzKkcss0qo5YTvf4/PeL
9QvE0a4IWFsQdAZk0iB/w4TN+FxgaMVN9UutK1joHvMc6iMmduoMaKZDZqv+g9B1CCRYdyEDaoN6
aG2K8Fb1nK8bcr65SPU75Mu4zz71Mj8jDQRcM0i0QRWQCO+vxz9+EW1olOYXYAHXyHUF4PRQKXhF
Y0pfzTt+JtYrMtVtnZucbGC7OXQyhH9YAEr8/j6hUQKi8GMdpNgx9qudbhU/tm4Wo6kR4GW91kQZ
wMXVP1gXHEq42necngOC6JckLxqX9Mh8y8Zs+bncu1lMijbkiAE3fg2yn4vi9qayDB7ZH7oy3Z3q
lBN3ofgwvcqRG/v08Fq17Eakd3jYJEsbjwxdjfVEnIFq1vM9f1t9dSy75uQ8lVV85++TbnLOaa4o
g1g8dvxX8VxXIjfm2o+ok+yjNE6Mh9iFxplIp4l08C0sFLAx98QzLHs5lKyt7r5DtWt/+dvJrRpk
H2paYG90RUJ7WMBMWp3iodSCKKnsuvTPEQmGGVB8L0qL5LcGje4uDrorIX6nXDOSxVBY0nX7r6gy
/gAYo42N73lGx6wh48/Cqmg5BeE5G8YlOz6P2X2Q3YurDHbMsbakysFSC5sQGhgxBUiBu7iRaw8S
QqjZEQ4zx0wO5T0VU1WTXt3vksnQS97TtRb5tCSw95L2A/ulfWmE4Zg8rNiUXRzbmuiKQFmJTtp2
4cCwqZOPT7jdvw6lWFnaWnH149EwVuEwUPhQ/r7MTgdUNCYCvFAJJGjnb3iQ8ptKe2Orai+4Wtqb
HkmDu6s+epGG6+HwWGybFwCexXhBtGN21+xrBk/phSXj/sd5p4LR2GpK3EaRiELRWhz6gHXDNPBr
EVPdoWbio+bn4KJFfYnUVoUiGdQyjgmib4Dp0Oqc8mKPhfa+VjMUDrwakQxvpMR34y7GFQ8h0Zt2
JaYQVPxAu+mywKB4WOJVEWyvjDaRuCZaumMTr2rxPz/HqL+/QaxGFX3l1fQVNgh5opd/MvF5gM+c
zmjHv/Exp51bvY16VAVwjoW+7C9bv1fwrFCWTfcYTLhBRLSsDsPEKi+n0mupvQhfY53mGMiJcqFX
v8+fs2JXfSGNHJ9VfCUxm0azdOp172YMY11s2jzNDC7b+OONLd+hJdSeq1eFbnhDlm+LMch8OKHH
cRrDYQEfDWlNBjZb4pzVW8sYLINjl3UwQ2Y3xgnRd/ymHMbKzaFZozqQWCH1LPFrDCQacJ9eiF3q
fFyvoFpGMrXpPkRStOfAsqz2Y7YJJoQdeo8R97n9NrKJqmMuslw/rlaZ2CXnU4l5V1RrHoPkA790
uUuH/B4QlV6J+1tLa421z0jmSoKqB1mQZmRGbAnen85uI3XcEasOf16xe9Z4vp4xB+LObd1VvmGH
3pe45Hg14df6rJj8RVIDvKgqJo+KWzZ1t1eulITO4pSYMR6TqeuUROgNY0GC7yo3kOhfSRSlz5q4
YE6a0Ml6mLIbivowqbjXmVXmsSgbBTQkKSUYBN0RZ56GbrisyzX5RZROWhat2EA+A2NgzPAbhB43
SUSJGwgdkLMroFfyguY06hC66XfWiD8Z7T8bk5xj9Oyr54g8TbRoFIvsIADN2jA+rggVnS1jhss0
SLu5eT1iOPdI2yH4qs1q5iYJZDGtAGL+QSDOg1VzgbZz4LjPvIuwr9NG5/PNFyHXBiim9rIQoure
Hx+MPSq2jt/tJ8jX9gpihNhbSQID6956grSBjgviT1bDiUjdsW0jx/l2c1y8KP226GmwdQOPRRP2
o52uxqzTfyC7+FQEwyM+l9aoMq1plodIv/uQ5NJSyu4osKzKQsyzFzVraTXWLyMr4UbQkVi2PNJI
MQlU33Xw8fkER3Lt0IFL3aNBirqIUiGHpwBfoxywe4pJm7Gl1AaPyeRAvw/zaP10GW9v3AwwOXzt
I4PGMgxxF6ZkAwwI1k30os+GQHy/uAVuKDW6yS4DUaPJrBZ5UQrcFsgWi3TXsKtfYWGqeDaTmzHq
huZq6FKjJ6OACyRz4nUNwcZG4oT/D2WZM/FXCxPI0Ddf2xC0rYLjrDF0euW0DIS/h1dKfzukLJgO
ohcrJQMHnctCM2h8UM5TEYg3yOyEavIF/6ckdoTySQpRGFz/IXD+zDndciI5O/I9p68OGcrykHsh
blcAz+4i1jbwTRKH6M8QF96uBKB6wXV5+FlXV/Ix8nqyx6Z2TZOyAGReGmRZ/lI3YawkTMcVfKbF
xeSQyZ9ol863g/h93okXGzVsWgdbE9xujxL/gThn/kqHAePo+bsjSYvgDTZrf3J6lLKzZacYhD6d
rtfCNQyClaBD7RPh46KCqNCTsCUnqIpOuJAloBYNNMS0ZV/p05Y/dFajNLHluiuwa1/D+bVkxafp
Ky71YmSZn13dcFbV9loDXGumfu3Unb+M9bMwKs+rX04dYRA/0RwLCC7vg2BsOL4YQu+mT7w7M90c
ScTCLi6c9QFH3BIRKxgoIyXlhF73VNyIgDGQ11stOAN8svVevC4QqlEl7CEXa8T9JfWP66O9DzJp
a9peeJlrUi3++Vq/AfUavAB5dazETjil50cqA8Dk1Oh1kDTEIObz8Qi/xvFa+FCvt8Yw4oxiNX5w
pqTv7oJAY70pcn6e79XFD/8kg41hzhz6+7+8A3eP87K33+u77rsANGHQ9clJOgUYuFkONQYvm/tk
C5v1g76i89x9Zdn8f3VmD5Z2tdRKYzDKWqhRW9Y+UoXxIwOza3Q+1MyTUvTpOO+H6EFYRnuPjoN5
HIykX5a1C+Ba32swDSts8OQWUSk3xg+IMVeaYg4CTwdlpIsUhfqdPffK8qTvMXCu0dROjO+LmMWx
j9LMTNYy1dNttBXc0Xmtp3eNUZat75TSxBySqfAL7dUgIcE4KASZ4gEzkbzpCx0S5WU27AEdk1oS
JP2Xn/4WMZLd/J1oOfy7S/AxN92zAEN5IZ6TD/iqFVbUXBeoOGwI3cXFXdcWk8lzYDNUwntLQafL
jZW/vjVaXKF/P8midVTVDk44CIJYYN6bQDzKhGlcDuJJrf4Z4X9oQxi3gGK4dYhqHVH81SAgMdOU
UxsRvnyyXbV3xFHJ13ctvxB7FVMyYyQ2PVr1rmEYhd6dqHV7mgXryi6nt9cmJL9RajoEmujqnmRs
susFEJw2on/+9QkID7FidWaPJ0pENNDNE2kiEyxY72HhQR4RVoduv6nC53DT3bB6fIqcVkYONFlz
67Won5iEfBWNOXXpYJTtjOHAMBrCwO9CJGCMvLH1oBd4CMMtayBC6K2/n9nxOUEGcmIrHyPYtZRQ
z2HFz1eJ9yU3i+D3JwYIaDoEkO79ge4KESc7E5lWFAbJuIvQoqw0K1dNqcjhgP5npnBGpkCP+Yst
5SLXS4LXQzGDIXCAa2rMQHJ8pzbnMbcsOvHnGK56Mh7yOxvBFo55LUecoBZ2yt0nX8UhkiDW20XG
xDsn2pcoPnqQJtSAxIhRScLrO5sWwbGuJEGyaYAmCd1GbnHs6Cop9tTpf6IEhTwmV9WMbEg9NbiY
77Scl1ToaBY3whThZStOa+OzKyVHecYlWcjlCpnY2RoURuHdRH4g8EwgtrVLjv5iOWKivCaY4m+R
ogFZnoGSmBlFXx0+IgLrV69m3c9nGzchYR9MI101Qbep9MnUFRFYSBXbeXpjSRvDGDSI2o9jHp34
YIHjMwytFSz0Yn+dmPlpQa+9DxpKhPLWplmqVYX8zAaO1GdnFjijeo6NuF9+zHS+MUcO4tPcGohK
o7D8srzl0LUmGLy/FqqEBCKEpkgG2voAuw80BQuo+SYMo+MGQoA45zkCFrh3jgarR6rTCqUlnvT6
7fqF2xWUqvQa1Hz1rzaOzpK8bZ8bmbRhdAAwAMmTavQvEtUr1W0Vv807pdpuNAhipLkek2CdhyCN
hMYYvmYnKEyTIGynBXSFcnfs4umf24+MtCI7dbY+44najRk58u1Ntdw+0lEhxFBQfVIr3RgW8f7M
9e8skbUZ7Hfwoz0IFe7G4YEW8YTLWrU+LBVBTZRKRXoJtBVjULcUGNjbaf9XxWdhq9xuIA3ytAPQ
ZT6fv0VbnNvndqJE81VLiUa9lrNhvE0nOsxOCZP9k9H6zctCdLHgTLpF+gXYZM/mekHnmTRfakUc
iv1Jy/lrXo8QCGywZ9dwE7b3h8TON8y3okZrA+uFh1/AdlcauJ6PzxyPYJMJ/L/9ziYVmA/jjP8D
nlV0sgzkwaVgC5I5l2bwJLf/T3Oi3yWCBc0CTVfaazk8OhNW1AbZIFohQi3oWp5E0o/RVvGv/i5g
I96P6n1+fjd9lwHFCBlZn2Oix7xj2h1MQ9tR3nmpKzK4y2ItwDnikUTa0h86aWjr0PiKwkPU20sm
HEKuOYQVNAMZEmrMztDDckPSzyblZ2tH6xxsNuONBC1lX3p82cu7W1D3EyIGsd8kFHsjICqQUjIW
u8W5Rp70B3FlhAeImHEl5IBmFq8L/mk/kN++3OSUih1Gg0D1yQdbYh50g5b7ceDQSnOFgGGa2Y1u
Q3eTo1ugPygMt2cv6a8DlykcxUOZIvuafEbQjHByDCaUH9wtb9+izbZDwFjvQEuJu84jztlX/HA0
2O50eEtgFEJZa/CjRbAx8+QtxKKYkRv9gZzZz/74CWWD9wUorkBNzsLHRx7HoDBgQqmRQGS6QNO4
9VONza5O5xS8HbICpOG0ZIvRXOV6TNtFe1YGHdW3YADwqhO+OrxYZDufSaASYNHvHVYhGF43W1Pl
sNmdB2uGSE+Y1zJgQW+dRLy7cJD8WitBtAA5sAHnQl6sp286kGN/89RmhpfM2lXWI7g4sGLpSYWq
AIDo/o3kkTwsd1VO+V6RfyjYjOpRs5XEF8V0PikfsswxgSRmVv3dStnjKFqZ/SMPkJiACkpnjojk
MC+8sts/ZtmStnVwPL/E91WfKuQR14Qm1ucDHpBBb6hRjt+MLe0tPPI+mb/nq1vVNYtMkPW+YwzZ
cdrGs0W3f9qXb4rcee0EwkVOqnyL8AzU6QIN6l2J2XuT5zK2w3KCTNfS3u7BTBud9HOS5a6TjJjY
7fZ0gERxCyFo8XzRnZO9CeUgApYuwJk3P0L6EHBVoiOXBGnx44FVwgQ6bFY3EXVuETUOyqSDZI/7
9FSIXDvVxjZu8onByrA88SjNsPCN2TN4WnzABB36z+wfwnTRLajou7wjtGKyYriYIDG80YgPJHry
ouhcMAgEb21PhbReArOON2hNV6mzfZnjvhZvKjynn1ECr/IJNwjE8a5z9xndTlDWfBjOjBwCHFHN
ezPCxWfxR7YzoSXP2EYpQvvJTgn/uG9QdB0g4HZjSe8xAklO8mT/J41KPLHx27ikNG59H7/w3IXe
/K83pPnb5yGYdjSqG70KxDWC5cv0fGuEAl+ykteI5k70myG/ElsKxAUkpCKBV78lrXdqSSlOyBas
JNFlK6ozInbjAs7EOk5XZmU7vulDWQIICpJtcMU4LI/DKT6rnF9PnkOIDRJOZj7ZAAhquHDNvEsF
phvjsHEIF8pg7bEtsu7MhM77JWfBgNTD2hlaOqweqx9x8o67KhoZPxowGKi31Zylh9EZD8jYt2wn
LMa/5rM3bQoEcLOw5nIpXD01L3b/n69dkFchH3drZ4j+UhAWFg0toxuPpkmWhpjAEpDBTsL4Y75g
sCtJutemDh9XBEu4XuNYN2CdtFcrRekvpX5fe3EBhGQW9foxML6OVWroK/dG1GlqhoVSEK9+vbH4
4xmezNWdGnJLabedMC9A8DHTnPcXCGPGYWUNLUEQXXy+PUnC5omkG9esLuUcpJ574N1GmLiRXnIT
+N3OM71PkDt9cA6RBIZmkdsADvFPHPSs/Jhep98Q4AZ3agPu2vaxoQdxnMUY26T+Aet8CDQj39sb
4HKVULAEJ5jLCfA0vKeTgF4pvnVQkcTjXLSicZGFHkm4gk5gKD8kvTkxRP8LaQS2R29JOJroXdI+
6UjMd6aUkIJ98F58KGr+wCueN8CHYzeFzb0/xa1mMIhUfUA2BbDEoBYsMHuioIHJj+V49xO44BG6
KSmSbqt7GOCIMAF0Cz040H1iWf5wMf4hfDPA2YRb6AJyO37mT5LVz0ytwi9SBpPuFbcjFZefCj0A
rEBt8b2jMqDzbBbyD4wmiehc2bo3PY0i0DPkVQqnlk8b3Y6ZnZwG/UgE6sqVAtgBwSyz5N4e6hps
1TlQUwoUcaqkwClwwm1+wIeQMBp9mSmryvrLuUVxeAyuQs4T8dK2sNvPbE1TwpRn0fxIHotCPv+G
rFj8c3UqRrlJlaQJidFnXMOCV95ysr3SvjxUrTgE/NUFoScO/Mwq2J6AZvmrx1hMl83KMVgEoxjl
nHGXLtmNKvaKmRPRfEQtwJjlXmtvshNUakGrfEUpWPeRApOCbdLCmSvXQno3jj0T2i/neF+8ONsU
NZmj1+ip/H5GZK0yVMivZoFhttlVyxydvrVwHq+qHqeIL3INqcRCxIH1TWC+I1b2aFf6Ykn17ey3
HIisqPl8H4McmG5wXEl0iRoR6aGGVAYjyzVrveuQ9LuRE8nhCrKcT5cDNHqw1ZyfPkmW0PMnJFqy
adE8PEegheU/KIjlrqW5x59+JkWpFhi/2/kN9JR5r9G+bxostXsP6nFz3Wi3MBwOBLt8o4BIenpa
IKm4omi7n3DtU7ZXX5Bnv2sPnobLumFVMQs5k+955qBQeNhoZ2a+3rnlqN7Z2EhP27c0NSfa/+56
clc1zoycSaqS9lIfW7duh0VBSIQAA8XOBaOCYeabyG5NeWBfxBJC0MgEX/NBEyCxAB75odW3dbXe
L9fihd568uFv148oaxNho0Dc6xkJT7okkAvS1czkVfw3wZlIuxshuRX1OYn/eAkJPmmfa80FjW4z
weyChdhrsBp5vqlkBCcrvzcDQt4Pn9cjVsnChfsuyxq8D/ZHlgHkVsBptyISdo7WfE30G/Xb0Lw7
GFxB5ephlRD++GmJl/JK6mzxHllnISzWKmsK+5VRn4eyPLDhKJ0oQgpUSzt76wG5ga6eXZz+eZQS
kekRLlJYoVSS7rgAm5SoiPRFG5Olv1YlwWbzqPCOMY0kYQEhvT64wgj3G+/SIzSy1IDedgcInXNs
cZbf5keuUUoZ4Wzpu00+vCbMtRUC9N6s2COOnSbo3SIaPJpR+RLeGoU4Mbt2F/vCWno9imEFEk3M
96U3nF2HoY9k63IhdhUWKbsLdm7Kgd3mukx0YifBooDxkekviEc7aJS4ksnWhUm6hHxiYspBV5fB
PgBMkYnjeFUUA4KxgfmWYSeJz7l08rrrPzFO5Q395I4cLSs5lpIp9oCFBQL1p17qmLj96A6g2ZUe
saEavawPbP+7FrZqChlUCNpqJ+Fdx/edmwM1BMGhsWkBf4ORAVkr1FNiZrpBpA/W/DbQ1YjrOXYN
I6rgleUvbxnen5ajMxUq3kcwbXJAMMovabwmTyqIzyuzZqehwwYGEahQRA/Zg++6mNUQHW/+yi+m
OmRGWu/tn9ir4ZMag595i6ejIZjhmbpaJs+mjdaZiKizGtBnWRtFQ6I2IU8QKQ2tCGPFbZL//gEv
ETV97ovrllc3WJn6xF0agDEQ/HnPnYpHNSsfGBuugg5wWG3uyiEfbyaR3B3XesHlBXplyMID7oQC
vJ/2ShqJNIpgRGDKvs62RZfqpezELkmn+YmaZJS4rAwmFuyStwBZjg1bX2p+jB0Anj252wdxYRZE
nFqONYg/nAcYwoEzECUMY5TSdUef/nEGyOYkX6fWatR6t+lKf4LRThOdenU+ynWSHaOXurpQrKN3
5vie9Eu9MycvGtdxFr8hgw3Iizpver7FG8yrRNwRZa9FbbgmZPRAtm4ynahc204kWEBveq4CmO36
qSO2gIZ51bQABuPmvg3D3p8X+6wF6m0FUpm9W1Xh5KbVOlymxytA1JMD9AGZtNBOmDZL6ti2VudY
zsATSEN3iHPIPEsRxjo0B9IEOWxvC/HSjIB5GETaph+0i2N8oYTrRfrZUHC5sQu3eipdTdP3pxTy
vBYmzjAZMv09QeDB6Q5lWnV+GdiJUdVAZUHLpAouH8zrARJBiQfb5ax54RIvGYN/Ct1Hmw8KNu4e
qUes4sk7puwOo3Ht3nvh66H9pWFVYs8Yo0WN4u9JtBr+prwLlQiqFPi+YJE4J7auX9Qp8QBpF2VB
hSI/G1J+we8+3l3Mw/j0tNQAztgTUtBFG3hqeGIUVJ/116qxcL9KFeR6IdIwSGlEvyE6DgIT1Hgp
4XbY3QtGCarCj9+AvDtuRs+hPO1uRLzsrY4j8+2+a3PH5zXGEEnaiH8EYNBDeGKhzrLhglvSO4mQ
BySjiMZsC/w6yTQ3eKINGyGGTNnM6d86QUDTs75KIIKBMVw01bDET9nZPOXf3weOrfhnpsFvFkIU
U/gehaebJNms4fcrybtoNJAc6MVxTShhrvAI3bj/HxhMid7shzz7f08imN67J1eRittzxP/nMghZ
52/E1H7Byvqhq8qYAlYfRrphdvRDovVc23azEWK9RhWDw5hUtrCwwQlT2mRrTbT42Tfd8YC41OJB
BtDyjoiKxiI4ezsWv52tIEX/h6VlpV1i10JyTLZcx6i9pORZNSLXs2uLmBMPRuUllpAW1vIGgm7Q
wzKT5F2lSbAA7MkCZ+1zphQtI+gomObLfpO7703v6vsy+/gX8cjx6HvKld+4RjlfqDi2kCm5Q4F7
dzFFe5ygoa1O/Ad7PmFGSyxqxnTwNRH0v71Z5Pf27SehKYpXrJGVBfNEreyZIMgsc+sguQLQND5T
4jY/po5BvNX9auaSnjz5jurfrSZ9Xy5h01ETEUghSjlA4q568MxnVtftpiLghB7pBUvN3jrW6/1t
EtYPm29tddpNsFPF/XDYajpVLKV1vvDPQ+SmRwI10brH00E3J1qo4ddKsUMmv8Z1nF4TzOzebOaK
tLkaMwMfjh/1EGW5FetBmpzwD4cRoJR+Ty7Ge5R+STrVVAgv8xyGpl70J0P3TrPtZjZyeI1lY0WV
aO9DRNw7Y2LS2zWKGrHiMPw3JmRYqvDLCb98ZmvkWoLt3I9EVsDKc08P/Afcqkb3HQxVdj+LozxV
uSwwjxnoDmXDkAFXb0loO6GyzACuLucs6+UyzGjbD/SKDvNT6r3eNyLhh8tspDzjpGdIkejrpxZL
+anrtUylR5Qtf9qKkvtuPHhUjSIAug+/W0+DkDU/HJDutFli8/xRwWthFSr0NS4lkfEKuZFwp/wR
DAjlMl569losABNnrxcSF/ksxM7QkOaHTi6W+QZ5MuIjWQT+sMiKtKAHPpcGYt1DexjAvgTTnzbu
0y/B9T6NcmEsVXDCAaboYXW9X2kh2+qgXB7D4QViaO6rrnBhzfdelmdcRWQj49tJqebRR3r0DFRt
7fnxeqURBmFymp331x2HRWAWts/+KfUJ07B8u+yQLO0oetXYpGrv21dpzbH2Ne82w/a2jtAZJRbl
tuteB2OdJVFANbfJ4H/hjxf+WpFKXUufRuVLkMzYewXT7kz6+hpOQV7uO/v1Ck2tbEX0hkNY6l4Q
6DN6313qnmAYRoNV4m7oL5I7Bg9zn3BNHChHUQaRccInKVpw8D/FuS+N7zF+045YGpSjIwc9BsE/
aHMC050QWHEKaqVgho7uQENkxZvTCsyA58JrqZZ3tY23RJdIbkq0A+Tm840NZuskk/yWMO/av5x+
yEBluUk40wjUR0bhzwuYPEqLMfsDKMbZuLUF6WnWVSe4RSuNnG75Ob2G9wbgZM4EdLW8ocmy+GqG
UKSJM8BhhgBPBKwm0pWNb3FVlT6RBbiYzh4M/BOSN8F7r04V1K66gKBVV6tMkXrbC4dt5JteLLGV
k3zBnDSe64MC1Eeah1RgVUH7hzdYhujuKxfG7tAYOB9/bAOzEJfkXvlC25ss2LdJAHHExyau2eGf
2UoC612FMMJH66b1/ab26ohla9WLZVqkK2935fpCZI8cLP50SAJjGskyttD9XYNlRZ9j4SE6zXDn
x8XvF8k4bLIQXDXNLEl0LL3L+MU7JcJlbQnAMekCCvzU6fHE8YQ1ySTa8kMNKUiu8r+tc+xQZ63O
HaGqfAbEdBgw5XXgd3mDAgnhKz1duf2JCZwnB7QC7HGC/yKj0AMcg7Cj55z3gdPlmO/om2LnciaV
JT1FqBd3ODfAuYf2GM+/r0J8Hz5/MoaK/iTP7g32xuanAZ5sV+95REB3QrDwN7KFoF2AqxrdNIuA
CaD7Ec8s1mA/beomzY6DSkw9hSIjrBo7oktGBUN+Dxg3SmwjLvGcYgLVLzSu/gmjW0RGSWeVAO+y
+IdhsY5kwWjACv3SuOgqMUpklZewpuqayszAQzO4+l/seCljuh5w1C+ZnuXUf79pyfByaDCT6cHv
fTvUHBZB5bIDTr7ypkMqQXAEzRiwc4RBEzWvzXMA+JCw/NOdUCWZ1XGE4Exky6p2gLfBijztZNsP
6r6yfmJWM98AcAx0uYyAoxH4pZO28P+6aQEdLq3GsRgorhPIE+M1hw626hzEmMj7Us+Dns5OhOAV
D9UCtbnLeZwQvrsCVFVyDaGjv7+3ObvqxRQTHsWU8JEsjVYclSZ5UQIGZqBrniKoK0jj2u1hFyt+
/I1vZvpHlCWAe7OL8syo/wAyelQvJI1GGfQMPUqAWmgoBBqPsZq6YcDcIAUC2p40YqGhDq7r974z
IhsgkO1NZY0q7C95NQkulWwbQZapxwwwN8DRdu+iRMNT2g961dnK6+EQqZ5hG24qOT/ARRu3KVx8
OQ0PGknKcgVf3eUSYSevnuy6l2nrvP1qW2doiL9kMZbCSjgTsYAYHc2l442jOhwY+vpt8QzqazYe
+iUZ83c+gcTSrY/BJXNlduvZw6gRv4gVd5UmiNvEZ16p/+CgZ3gKKz7UtCAMKEoYUMfTa1zIlH4S
pY3ybJvTS2tDufjz7mTRTg5+RzaHfD92IKieCh/KalZm/4EmSMN8hFt/aw6D2QPz5BglpLk5b+nz
Kl3gEyM5KWISrH4ZVIU3Iwnq7hkwUHRJ0rOp8JHhqqm8gshrN5FfeRlu3bgGcc2/0Ta4kfVLKm+E
5gfgLWepe+5K53LFLhp4u+0W3ZI4dISU/Ux3/1v3eOXodOjfLu9K3tepJ1PRd155+UkJARAGl4vf
lucmnCubE0N5vP4kHzqRj9TNjY0VzYuM5oQcbie4pZdKYaOihcZc9AIFnsZbt1zKurDcgBtmJhtg
V9zWSLzYxnajn/IHntgPnpNGBzIFLWEdIzzsTB6fZ6UPE7h+/GVH4a76Nxq5SiXV8VBm1moLHIyE
1qrdnYmIwLdyJe3M055smdH4HzaleyLnH7AQe0auho483ydcp1NumQmc0W5xxOH/s0FWNPEWxKHA
rplqytqCoXZ0uYwWQO7g8I9cmHUnYtawZSF1ri62y7UpwhfDuc0g9XXXcnp/TiHEV7iRfx2AHTM9
kq04kaBecasG3KNII3P5XPTVObjIs4DAQ8HD9txgXmxiKkBh77fmz7m4ND16AiM3VgZGvm7Y5FSO
gY8HC3POz119HkQ6tV0Vcgg+oqVRrRAm1NhBWvjPtmhvA8N5t9EPEA3PWEA2M/x1YyLMsGVIgoZu
Itey8PmdjFeXmHh1kskRPgR5TgXRdC+JjWx+kNwWU5xGM7UvvVXkV7YB1Ns6kKdGAV36qAlGQFgh
hvnmR53jLlkkSr4e/C2CCCM/HykLGrP48o9U45T1SIhlEaPDs/PO/iS4esyfP0siYYPRsV+jjz1D
O6jVceo/ghluEpIH5d7LYd12/alIy+IRr+eRjr/W5o0DylrIE/jJ9cRAvBwGABMIUsZmSFt3iWaz
lU2bq6R2M/CoXxRWE6RwEn1ilPaLH8JWXOFLcq4Y3rHC5vZa/2k3zoBLbgNZ2VevOK0rBkFvyOZ4
utwM3hDqad/oNxmzrnJc7Q23M184tE897gQe0rabnCKihgaSKwVVU3Al7yOiaop/WyAZgwIiIzUc
kFZflDzDnbvIolbm7cOYPY1bhnniIAOGkvpBgD/mph0hZi+5uyyKL2IXA0HZTYU7pQrrzdwKCu0d
FjlUyhg6pz6prLRzIvu8ljwR5lw5oZi3pBsu+q0+a6WAudkoxDku5KKNyml6L3VxC7uSFtYlkAR8
rfqCQQ3a4BL5/VD5M6vdNv95fjRuKZYl/JW55xoL1Kol1buxqyJoEFtxxCDfzPc5DPVx99hHk2eS
u8enbT6eHXz26vKSK2cYlAhOvXFtpRVHTQHsdQkbc41OVjLkOqlL/kMn8R6nZ7Eo4Diq1slTb3gv
o03giufzZjBiU9it2u9qs1QV4TyXqW9+SzXjWJXFMnQZyzJ0OX4n0Fq/nN2LtCj0pY1InH9aZPPJ
sqkL18JebqtC56I89H/BCIgteHkokeJXgw2ovQrE65w6fNdxslePmkan8pcrqSskrqqjm6mkIyIl
QhXcOAYXByReDtepqgT9Cpcmum3Nvx+rh1bQ/GaDGs8Uz1ov6iGGBVX1ZshAIdw2APnINOjQFKFH
70x4wxev76Kb+qKjCbSEUBHoLy82WTM835cKNNLOxVJARwAdxdwM8fXd20olRDppSzGGyEM/1+1H
hdzQePANHxxEt+7JmswR0RPCxMbBOoj5DznBCFTVk5N5nNWsB/ucxqD5ionHYom7o/GMgwq4OH07
BHeDMnJB55OH3MHj6AgelrgFifq9gnObAKc2JICgCbA5uLSmk5j4LS2/tM+kDDa8ovwKQLzhzgi0
DFNvc5fCaOyL5/X8cLf0qREQ7XlUHEHX6FpLjYWsrydYuhCP/w3cNkygOpPQ9kjbreFd1KgfOjQK
0q7pg8pqIeT09M9GZub1KPxh3vq+NBuzWLRjSHZOOURJPdYAkjJYwhbTLKswFTv5qhrYxl5UFwIW
nvX11ew20Jtj01yswz5uc3zT0YIsnCOV4psHciRSAmcb5FhAGVsdzCYsnXY9mEzGfBw8ChJMfsWA
rP6gL4YR7QcwRBbiAlE3CO1GZqHQoFAxX8MEvBOkAtA674vllLMzYD4+hRrqiLwshDTk/Hhlj3k/
J87v34OvWibxcAc8ebY4gpMh3Qh34R64g73GmTWRrLRhkrIxKlSVFPYZFO8mDKK2fh3bnS/ut3Jv
LTh+nLif5sZKthX1W4MKOiXIkrr3N1IpEwJU+Pu1rN8/EyVctsRvjpoi4hDYiqD0MF+IfQ6E/SaU
Uw1ciJBRKshRo1nzdDeNGvS+cHiNoKowX8Py0mi/rFWoWnkWGWiG3PdPUEsAAsaHVOxJoV0P9JiD
maIGgjr8NY5gkI8iVIsbr9XaAxFd7WSWHI72Ran6xg5KHYnp1IyTpDzIjmQYB3WtF65OxD4m0Yvn
Tx4YOlX5Jb2++nQFTytUaCq+h04V//b52ETEPvoKxIDdRmkwt+Zgx2HRpafPXAAe8U+OGk+HZUO+
KjfVs/8IY2IlqA02c8qAsNbG/KGSF8RG0fiycosbOcnIOU4e+k48YsycWav+KBpw1g5mzLemFU+N
vRg5FGLmb09pFgIfBaKjHYJauHFU5OFGKit9TjTOYxw17XE/6yjHNiIhY0rcFqTBoqBedkL5yhxx
+aBBgnYfEqXn9L7ALoR7YiKx/hKAcTqnXsPDcGf7FpPcVZQBfRBa5rKdew2Xamax64jwrFw/Q/5A
w2P00/7GLfTykbhXd49UcbAd3+Ev+F2NYPn3eLCPl0u2NfLWCoxMt/qoFuZ2dkkBkkuekf96Ta4+
i1/4h/OLXcYM2SHI1SDe87v+O5DMUDPd3ApMjnK5rJ4delNyoofA/scsSScj1jwfLuOW8kHh1BF8
g+UtyX98YgechaFmNZIdt8++qJjmBkM2ztdi+47rFrvXS1Tc/0C+0A96z7I4+4uzgLQ9dWJXQxR/
zFEpzdA/3sOoP+CpTC8p3pfVo1qnb7wuI4+X+nnv0KLkpoeuDU0FecLhcikJGD+TFUrTwduedusN
cmLF+avxoHb04Xe3A17Wgj7pYkKXz9DKQDEIcjyM+MyaUrUJJt7igLFcgB03l2T13lkAAD4P7a5U
Vjeab7s1lYLRZP1cx3rYVUywdJt8B8CFiEtV0Jy+/YWCq1T8ZihD6KQl9hTl4XajRfECOigSO+aU
N1rvLGXJozU3Bhnn0xT0NNY7zxZzSRRgL5Ca1Sp5jdtCgnTq9GI24Dcu7DBdSgrg3b0TM1aOQre6
rmEWVPRIreHPC2ZfKuVRPhtXOBhl+9c87b423vkxO3NMS8q01Y3eOX52b4tFuJcrgqa70u+26xjE
rU4iqDVNFyIMb7CNHVywjXNbyQfx35QNTOWGKYmzZNZGY75WNUP6gN8tPoS66pa3VEF1yfYsp7Pd
jn5BIIxlQG+tD6raNEYl29kGtfm7w1drAMyjPmcSbK5PUi8XdEG8oxSXX3FfFE2AWOw+BhrMrfOS
1uljRlBq1rG0AFAqCwhKJWjYfMfCtQ8Kt2lvnPZ8PxxJa58KGJN/qBg+p+YXc9aCgTGdS4JqEtqD
7njjc0nCwqS0GUepxMgVY2Xj2aBxfLmrEP4S/jaZ9C6YcznTEzq+xbwCe3/2lK2aqucdO9SqzccH
Tys0BkNiWx+RdQ9XUHLrCAuOPkvIz72hTQ0Pv4nE+vkn7QwhZ/6V7rgWhH9fInYEHCVjThrHZ6EO
iGz5qeeHiwiAihAvuF2cHrvqwk115jiXHp0R6sNFfZcibPTLg10DOAVEaYHRM1qEJFKxfHXJsE8T
vdWZd0uDhqqKvWS0D3RZ3//LvcJ1S/ZB/592DN+omkwLl3e3X/QGESTMGteIhigsomuMLf/5OuNv
SvSj7qaqo9HMhoxrGCA1Kr1+PDIATsDUrm8XuiDiCrKTPVx8GEKZgYUVNGfi4XqEVgmBrztG5eQT
E7s3eu+yhxzlrlgv1OM+5j8IkC48cB83c5FmlOmYizpmotsX44Mk4dNPpdhB+ugJDpGMKUxIJlwc
FXUYnaAZkRbeUjkLTldW8V58FGja/Aq6zncsnviCeFyOLE6wUB9vrUWPkeFkp+S/sjVB3xbYbOK2
4MKwD5elShY0N4wCxPb7TVJuI5v0fTJtvX3KUVQEU9zWnPMbppVuddPGeH+DoUCe4FtK8XlFMlep
EmeL1XtcXDgLpPoYnTxd7TJxH0VC5nIgmOdh33CIrt5+eH6hFC0g8rgzv33uaSD90vtqlPo6sEDl
hf7bXBEV4L0NbSjffst67+eg/EWL8E8iXb+SIJ6fg654Ov2I+Heqo/8x28b3wKjf2NjnEO4NYS4u
qVmS+9g14tJQlFW4ONxq0JpSak0gZNePH66U+fXZhVPLouF9oxVlDnkngU9quLXti/gmJzO7LbYX
DzrmcgPYhPHgJ3aKso7klKE/xzVYT7joj0CD4xs/GYU2V2adapEfROU1uW1WRS1bOzHBLkG2og8M
UevOGXe7Iz5qOFvnjq7+mXQs9Ir9ZCZvNNQi1biyTzc/p/Ky5oG8bNUadCJJ1hXVaZeGZCl8ehjj
HaUx65sog8qDY8rFSp3357maOFQQdm1UxCRoJRwobyQIPFvfsLD+X9BW+hY6keZVKpsczToPkW1b
2KrZps4MAdu8BWoBD06jTW3UCHZVxMCdXk/1WXRkZt32Xmz3mke38THbXBfaZG+e3+9HQ/8tuDN3
Te5ExF57u2M2vW6rz3Ac2MExe1qjK2hwNkhiOf0H2dkH3zQd4de7E+/+aaS1d3k3krg+EVBgKElQ
iZ1sbgkfgOOXCscIRNZS2vr5UBpkj/1pVOWwaqaZxWHxTEIajiaottAU437+hq450zdvuRfj20HQ
+vSSwaTdZzSO+/vepKh8VmBXX0Ktjs9xOLkv5WHWnxkoh9onmyKuGK64uAaWcqy0OXm9rmauqDND
uC04Y6+lFoDa3DJcr0g6E3c0p1W81/pWdcmI611rcXhnqlNpXzKqMjX8qSmWnw3dYSmjj+qIjHt2
uXtZm5F51/ZmjNJSNuuBl+L0F6hTpgahHuOcsqW1ieuK7M+6OVgQ2UKgMy4vcW45TZY8WEdUAB4T
7GWn3I5e6blkML6kD6acYG8h2q9a8pkVkDeIGII7ssd2CcBpHUzh7fy4J/3AUJJWH0AOUDR8EHsU
ynihkMWP4ATuajqvIDQyt0+y2LO95JL4IcvDUZwBQBUaL8Vtoi6wjFRJtD7gaIpnUBEhgOIJS1ND
iwFD6nsIDR6vxXpgBeT+Vxr84lSozmRJIDaf70hTelRrhxGwwoIysQCyNmZT3Yx05XeTET6MBBsL
LqVvXB0vQo21gdkrm4WjMh7T4iq7wCiEUSZkT2Dx0KG6cppyTbBhbCbBb0YzoZRN2xMBvQ7IoC4k
+lFkHoCzZDUtUSxmFXqS9sycuEJQUSBsppmWocz2JzSxMVsiD1UCE2YCG26wiRfzixls4hX7XZ55
3L3DGSIcGnAW7k0E9/smBPD9MreQIFlR07xvV8wUE/WjuvNhoRRl+JWdZMeZRb6ue3gBW+rJasen
cVmId1LwGjpFAanMBO+UyHSOR8lrEQgUdQJS1GeIgS39KqXY88FtOH0EitDiyB3rVb0DtHdgBr0t
zKsce2b0mBqZo4BFnLqOmjQAnQC+79dJzCnrlmrlrCg3B5iPsQul1JVSfBM3c9s5rBMY3fGaiJdb
heAqe24OMOEBQwDMNb9lo0w5691pV6HBCC3t6qWAsV48/n2eEgheBOFUDHGEByP+a6/Y4++dwYTe
BEt7Ig2TazxVDf09iD4yxIrBU85GajrUda8UNKaGf0MVdCl2XA0hayXVhlP0WUJDwiX1hu9F+Syz
2HT3oV0rtz3fbwGnjmgIDTXiYqGuYMRo3thlbUoHETUJ3UoiNUzWT4YNDX6l5Ua3HVTlCsxIc69b
/hGRytOrGegeJQ8MBKT17FA/1H/rLnS+jw3nbxWLYYLZmWw9a05IHGY7JW0vW6Yc84nEq5bQqG5q
aYCegD3O2JnMcX1MYkBTXG1769U+Aw9Goh1y/87fNnibuC9l7OBIp8uUOWaSV9eoEG5CJkxw0Jtf
gu1MhP1SFszz35Eyc0TW2s6EEriJZ4zHMcOyXCJKzXwzgwoyAO44YbES0hBdM4W6nXZO7UifEtww
KAa6fOQdgI2lgD347ZD+4LrrVHcp67xLX5cUzv7I/lkodNxo2c6ZaZTO9jRAru+uBLnQe+9+Zmre
C8Pnn28DGIzyNtBNvU5ANC8S7qypS7yhWMoF6BXmfCXELWvNE//ZJSou3aE0cdd6VHzC3ReAj0LV
3Hezec5D0/l9ZuyB/H9VznCoVwXHku23+1LUjQa/UxbQRqps2MIltpu/8sE16hXNtLtCFBVIqzpK
/cGDyizn1vZ9gv1Ndrl07waiFRNAXMxg99g+C/ZLS77ONh8WOnLjx4EHyr0bHjrfNLH786Y7CXeY
avl9avCBP7AZDerofCAU79L4QQl8Lvuy34h5MUvgRMldJ8qfZdH4ySl28LqIUEzl+TQFn/B3evc6
PTNN9L+mQELOexdAwSZg4TpdIN435766fIVHU/3Xy+ayOM+ug/LvDFO1GmZsGsxX4AVL/x4jdRt/
cVdpRk9pCqamKTovkVUreNKNCXGFCpwVK8yiv0jIqUECrQAjrYb7UL30XD+VDnMeoYHJPGGjleuM
2xi/3uo8wAHOBRYSKh443j2g0/jwVpYpNK1ZWuPGBd+TCQX1lukHZ1cgje7UGjjLN7bsxxekncXc
QzWfb+pG/PKIXhYPUfW28a+d168IxHOtOzH7gbK58+9xIqSxf6N/D8mevU+M1QB689crNH96Syv3
t9u9xhkLXH/OxY3gX3I7iGD+rOLoUFC9hTmt2cpZl5aAOiKLXF3YAQrq8Ou+QDCnZM/eUZm5lMzp
BuOdA2JHjskCpa/gGGZYk0W06rU0ESQSHcBNF3OxGvc0XH2WAhp9QCVeU2UxiSGzLIqz5VADDfvq
8J4jM5uK0p5z4UIOMiofwqL1SJu/fa2eLMz/oNPUNce6DLN+y4CNfXdqnD+aOad6R9+wE0VMxl9m
+ScGSdxx+3yYV6ebfxZaIgsBP2SNNO/eG36plEMsbZm0kckO/p5ODQKf4pV8ZwsYf+RE05Rl3192
wjScJY2bfCg8cz4ix+12le5yEEqqF+h7D3tivCVsWxOXuiIn+N8M1j60wtXtIbzIGGLg5FexD0np
704XgxYt8JKXja7RVG7OuB1uej417+xXU6s4iyfWghE4fl4Z/hRIuDzjuH3E4x4/HsAjX3phPAF2
P/wGCV7BO3T3SnsbHxP+11iDFNjo3aHHQ4C6TZaCs58OT4M7JUMnJJmJMPRoN7fyKkq+OmYtHwzk
dVdC5QfIKlrNSmNrRRneQIn8fLA5rlllBTPfYWHg/IJC5SlQ47GHEY2NTIACGQ0wx5Jk4OmPOUO6
7qJd24T5qT2aMX0AXOl/M795wFG7NA4V+nuYZdgaeelkubEmqB5Hsp6PbXS8OrqQEVVbtlE2CCYw
r9NGi3JzGli+lyPUTzNR/eEoD+y4vwCVwzUnYMWy/JC+e5TLcsGx5AO5/JAX+t4Hf+Ol4uV/KaNd
oexV8kW3btMRew5Z8UJHjq0x2mjaBmxARROfSKldArF5hoS5isxzvIxw7hrUTQmerkTIej47pJd2
q7EZUPMiP80fwjARjZBGvAx20UU9ghRm/zQCoOl3tfHwy++sKKVr0IWDbNIOkdn/SmrI77PgBkzQ
6rABz0LUuKih/87raYgzVfho9SM47gfhPQ0M/QtXoz92kIGPKUPpjoOU0LBl9HxZGi50FCOmLoDz
Cx+62vdNGWO5hFqvG4HiIkAj+V+egvmy9jhybleCQihnFE/NUdiDA/iYttzquDS0j/+zA+JhmJzw
gGRU/FiQ6s/7sieRgJZi6llOSFhQ0OdhUBLPEmbpJkaQozp89X7hPUnzVnFNT3mnR87CD5BdcuYa
RKKmiYwymoyNH8PQhjjyTVnefhABSQE/w41ApF3bwoZ6/X/o8cxTXm7OroGk5JwRlLzr8R2znx/e
4cWWw4qL4dwxRI0NuJDnXFMixjwbsJfgzuBAzSoNplA7ZSFCpHeDXqXDqGgsm461P82M060hMZ7R
aMCBygMD7eLOtVTU0fHw5uTkKARyTaxH0PJDauv7DcVm6gp6YeQF4YYjTkB9uqXZnvgmrqCsl0Vi
OZWKZPv7deUjOsi+VRC7rJ7Oa7ZXDVc+QXNYuUcTBmwnPoFgSQOUwAEcdEq3si3LxWJ4z4M+qxlk
mqgO5HOE8bDnpBZetLdguhJDRPbroYyY8rc3swdLa6L+vbyiqtV/A6K4hpgBEoTOjvxARoT8HNZM
At4iXuNR5wjHuwnxeL+OBmEz6Du/dxMEdJP5rFMsSO9d67IiFZbpIVwUY4b8t/iFsUePd6mlwLdN
LK0+IUXxjbetGMMjKqaOA2PrmTqZPjQLINw8jr3405pRhpHrtweIUL4FnrChUsVRXB6QrW4qRnoh
PhuNPynT2U0X9IJkK9puUQEx95fSb792tbzWZxDmtJVi1d09pmoilRi3cyyAwHjAWhxPRI1nX8tX
QZeTFGLVhjxCOoWquYv/Yan0rGFAlJcJMIlf+kCViBP7o0JNX0qlt8m5diR2uXk7TEsbA0ehPLa2
+QU9FN/w/tXBJqJe4CnzlSSIdbwN6MK0uflL+DUlhkuBHOO3uZHQg0G+tQp10fQ7GK4Yjw4/cnfO
DEalxhZd/b9biWiQd2sn5afABwgX5nOjy1jro2oPQneq6EUXXUzgB4vrZgza5CnOvsrKdRAgeGrX
yNcG+Iw0mbInlF99d25xLdrnrxxf6Z1tSRABfOt/XmHgM4d15rNpUFo8MDYYBOkFEj6s2h9RbtkD
T4SjtfMxO6lsnnhM/iMbhspNPwmA1DbPiv6pbL7oErT/yAtiM/9avSlsLA/qmDSwxZkq+3qeTlB1
ILIxLgpIAHug0Rvn7a+hrz/tyFyynzka6pRATK3zs4bp1HrmKTwcxLEgQy5qcOSlasjLNTgM/T11
JaW6sJz1x97p4UhcPbKiPpMmOlh01ZFIGCHAswq1JyRVx9FjETQPjkqQ315hfmr5+M05J5W2a5gZ
EjFQvNDM9xBct/Dk98qTZ4znVBxA3ezWpu+Ew4rZWeh9TLX2qde1NezUn2UzFD5irp5hEX6J53ut
JNgz6qIS1pbS1Lhr1KizKEy0r2qQUHcuVncTxSxPE9uYLXLEqDifIsTHIfKg8hdvXPUpAlakOgmk
RDzKkgdRmSYRVCMzWlD9OhIDjn94rVJHTaU9HFDGRTNtjmAqDy7Mcun46yqAs20eQHCyW1/oMS9N
fDN1Jej8xmXYT1aPV0M+/VfE5dIyximaJ1SYG0Pp4CD3lJS0kjCoiIP8SbN1I7syaMX3iwMJsZdm
pzvGr9220XFl4ObcBzvoYeayW/7n7bv1+4jivJkXVIu7N8h/UADNrKEFhOhK1Q9w+69045X6RuLr
a3ED+uNuNbobSzLF7ETsQgjJ3nn9ttZp5pv88Nm9h2ji5SLqfIJZAnml+v9dwyXSa69y99uyHlS5
W/wHK5wcyIAq/z1w58sXL4oLk0g0wUr6Vs31UJ3Qc/mYdacCpeW3pn9EwlpeUueBgLCqVN7CiMUZ
cMIwWzaTmmCxQIuBFNJ5KaKbt+a/h9jG/QKqMHxLndArQNS5gEKowULDoPK7ODd7YEaSTWVQOV6e
3KXYJkceqbXNR36lawVVgQrultQp3BTHxHnNi9FSplPWM/Iu92lRoayr+pzwgjZ8CpfpN0W4cUSe
r1HOoA0E3iBDntElWcrqSt+4l+M9uMuBuXnio4FcO+GTUR+ZHDnD+wg/uv1zRdEz9JS8+bxnCCtc
EHR37u1ZLjm9FbXU849KJZLjcsLxxoqxwp85FQ9hv+TWTxunnLIiTB+UHG/dfFBwJok6wK/h+zHV
kkI3giUCIlW5nv2N+6JODH4Jmypm1fbTtOZjXelP3tBGMhVaOyzE3ziKWGwcQqtUR8iLSg07Bmu1
3j6gjGvcIC3OwI5d9z77V9bnnpojhGM3D5bNxeTINOeSoy/xvjROFA0Ot8Xqeip8D2ICrmYcr9q7
Nfl+Xzt3RYbsbN6Vbn6WvUyZ2vLqisO4PkJSyvwP6vbcHtFw5kbfKJ7ufHkQAoqU1tz2gFLUfk/k
CSzOerQx/MjlUu5Ze1cglJZ4uvnoLaZxXJ0halMFrLe29vM+qgmpjeOhzb/pXWIC3Lx4yY/yitCw
s+Tmt7i5K2dp4DFtM85FdPp8huMn4xdswDnpoi6KyTvY6Y5GwFcwkyrnPYzKDd3xRnomP09CXYJk
pM+QqSXQmD7FtGSTNpELxXAUTbNQYNy6Kasb+FT3w1106V6f9hrJ9zb2RvKTFzqP4fhP9plp1zj+
4uBIYl5qSdY97sX+nHjHVl7mxQjT3dLeeIdNSmLzhHhpsOHNsrSk90JAgFY45Rhu4Ookkv6PtZ4q
yR8WGNjmcAbT8mLfvFz4PW2knjulfLCfVs/N8Y6ABG3CkA2SVqLHv70eTHrKc3Sfz21pCgaATcBx
H0uguXXUqJCDxm0/r1bHcyZerZuJOXvEmzHRrdG1v4gctUYhUQAQ61oraOGKNiIIK8CBslM2oHAk
sK1i0M0lvyJmdMIlKtzO5cb30GBbTUo7kUroKvVOAp4+blOoZ1qACsD8kp0FNASxaPBFMEYrS+7l
kDD943ZCcJSoh4nmVtA4KKv3ZgVVhVbBVU8g2hO7ztMLEDRkLltGE6iMaNUb+ftEhN8lXLjpDX0z
FfKhcIAoHO1w66DUZqT7wCR0dcB6PI9lqovDQhjHvgHjIDTgVoqH8jZYn6vUszZ3ULlV0B7gmfTS
zxPMWfJOmjNCN7kkRdfpVOJMHrzXvMtR0edEl1x3SOwkelnLzrqpoqJagJpux6GwBokAF1Oia0dP
MU4ZnaFu/Oc0C/Nse12Zq98XDhTbOhQF/92p2SyzOcxr81sxdeauNqfqWawaU7YzMXT404XIR7GS
CvuQNNunDw6ZeblZWI+eJCSEGy4YOllIvM4D9dlnq3x7L6/6b0rOudyJ/egy741NN4mbIP+FU3Xi
ds/ok2is6w1pagH7szhbpir15tB++NmM2u1cnHRHY2+d9UNzft9/SAsFzh9E3AloJIufUjVFZY0x
OXfIMkzuy+UoSHbjv69sxw8sZeCbIZAMcXU7q7QBuosM6aAqdUwGx02eag+LCmJZ3Z++RZclxzso
tseSvSPQVZCiqhSI4A2qVnULfgWuy0The9OvAFgt846orPkHp8iPnLnFTxnF4DYxs5d7Y+4qhiBL
4AvycYaTE1upYPKq/EoeQfn9f6Miw8DUFb1RVvnypuwTN0N5UBB78/TNXTZ5NCyvWLEYNniS5t+7
UBm4+oGGpmkcy7zzXACONDwUrQ2rzFrrGWRA9MSrS7OwhyU33H4xmGpAhZVg1/vM33eO1nH5tccs
SXrAYTLB9RJ9ibTbmRa/ZRuQmFxNhlT7bCMILsOc7PrTl2fPrUD/saPZS+dWdcIShRcIblwLve5E
fszP0DOUbbveMKLfEb6b1wboZfappXk9nNf7ySCdbY5MMpR9yFLyG7cOWwmwrsOr6oS3GrGJhCaZ
NOhzZj9daROo/RdbIqsSPohKPKiMbaaPPUfh4ss12NZMbFp91u6bqCQ6nKEYZEbhTcCZNLIe9Qr5
NZ0NsbG9QEaUJ8HEmfgpgkVXl4iravpBJ+Xl9ZPzaLAobrBHCNbXLPnS6bG8uvxgU42ZiROizqeB
v0I7Wf11JfiEkftEvmmmqnoieQOdZfQ++62+K45cVm1xDqwLNEyNNw1szifzKK1MrVssRwgGU/iM
9s5UY6rSheIZ6oRVCobN2dhSbdkvaz/MC8ynKLr/L9m7oFibAq7Er2h+Izac8nMKuLj0f/JrkfUH
00am4LZhh3jqVLSCuM1lG1pSfq9EIRtSSrtofgc2aRsL+8M2Urcgam2MUZzHnEIboKs28DDTmZvH
k9MehHw6AFQUSMDgGe6PXi+FMA3RQp/B5b2kchnbGUnYjSwuc5joja41MlwkPCiMZAAvxFhXO0U0
vKHrPbF0gKO0YOGAbnT5lWUqpHrqNGVdxelcYBnyCQO4tW7uJAFRJGScrsZvlc5LVeV71il+5FfS
z0rmplubZarLuLjWqpO0W21W1e0A++BpXBq/ELXrLForZYPU8wq28jqkM2xrOk6ljnWNdU/xcZ6A
tQo2XmnRnglRRpXu0uEguZx6+65n/p7qeI9XrLT3qhNcuAjydyKUUv6t/3+FoVWcdVaX/5UTxS8d
uUuRLLnQVjiV+s0mH4Zptx7ti7kZpUbD53TNHI2l/fEsMiWDAaQQLCiJXeTJe1Ykf5EMrfI2HM+s
Za+7yzBzyQt9E4mYjkvv2k/I0IQG6h/ToQMPBiCZ4/pRfPkohh0ZGbuSFDLmSoBJPZALalJGJF+D
r1WLz0Uqxt+JnUlB8seR9P6zKdNXHHeO2izK4Rcd27odl77wFR3bWdQyMjsvXJGzSPnxQ08GDllS
FvtzINtsWHx8pz8A9aZNRzWVTFqN7aLRSKg/aEyTfYks5nk9Lj8zctUu1MtHln9avKefV4zrftEw
i5gS2M+id0ag4ljASYmLu9x6iV98JwhUM/iexdhgYaq5VguQkV3FKbDMD5NMcT03xUVXJV42cfJR
3gV20A0XdleiyNRp0XSXz8xXO5+jgPCDswYZbvYTiOIFIZY0fB1j/QhpZIWj3KpeAQxk4trHa8hJ
AH93DmGLkK6Y9YbBnQPQAw5FKKAESD3gAZZ/FVi0Nfe+/cZUkPYEze61P+uYqwIKIRiqrTYmcbFs
PSABNNH3i1VsAoX5xzcSrmEZzGriC7qO7rrlIkMiZLyhegW1jRuHXRx1nEGZF3dD+P72JczfZF3D
gy5Qc27rabpoCVlfJ7clRnAc9fdCR57Ft1y8ok9zXpUM1zv+ORfcgrZYpQl7iucb5LH7aQzKSU66
45OSxdoKjOhMNbD2USpD34rV8JgNyH5EXM9DnciPk3LnYnAwo26ygmm3jWGLOgaCpm47g0VhGPqy
Q3NVF62HqogyOKGwLHsxCBwaDooY12zRHlQFTq1HDD6np0lySumculfl3Y8EGP6WVXBq8xkjWa5d
/4gZgN/qyD0KGGPsrqbSm21fORwdboSlUi/TrbbIBIFilxhC0f1yzyn2Ec49hC8aEL6JDKm7CDSE
EFTJ/pPNIF0eu6RdnFt39C5pAcgMbaj5q4gD8TWnooXDaE4+tgOt8OHFdCf1EWw66zSVnGXiOvxq
pDBnL5oDi9yk3bWreLC40TtlEr9mwZX97YF0FS1obERYETdpH133SdcPeUbd+thxC3AOJLn9E2P/
ebmu84LWvh0qfI66ObzM+TMf50i1XBtl3GYN8s2T8UPwK5d+L11Z+FA8EJ83lBPhnSOZw26XKfCv
Y44LdTnl/obcdofqZHh5IB8YpC9HeYbsLL31/zpXSz93yzo2Gc/x+Hp2D86Nz4Ikrb0EqWw/oP6J
rR84z1OCJZ0OeYQxwnlE20HL84TPUtSATtHOtUSsTA7jDoXo21bIBTSQTOqaksFtCW8ypT+/rw4I
hlzlMZBa2S2WP+z3thl48kY3Z2XvkB8BgWHrLTQfNDDNeLC/DHeSY2UwniDDIZ/1M/z16GAfENxd
TBUgNbwwTtwlLm3RVRknaSzfRVjq5neDpAQgxNa7dm6japVnF4eTBEbPVqxk9hylBcSdn3EXlNJ8
JrIP8VZF3Oeetl5BRGypQx+h2Fa3o4WgZ8DLlCDyCWEBv9I5eBvx/TU9NXFTMqurhvUQN0QmWgO3
k+gW9vDqcQn/Kkrgiz62KyzulJddmChisSFlZuezvlJYG3R2VLPmZEoK3ZtIasrVGYV/Vu13bm+H
1Qh6mk1+zsJjvglggqiz5IvZPCukOj9D6Q2TkCM5dkS8eEXQu1osLREp9j1GO78Lyns/0HEniu7y
2YlKCTsL/aUHsGoTz2t0YDlzhdx9sg4S5rsOpKvyF/kX/ZIE0vINLkJuGfI2NhSrpL/CoJOvICXp
8a+uvYUvlzjrNgo2mmtUohnSQGsXWvqeM7jC0ekEJ9WygGCW+Qlb4SeSM2zoEdBQeGglI7wsVdv7
OvKMyg6bMW98VfvbaNfproymlSkL2rvxkErIz5UtGD06gokT64wEt3enTRKYfKxF7INLCwwvbIek
XYhsUb5ezW89OgeXFuW4FFNvNFwGK6otumSlQ03wOHFnBYlMFnPEZ8U9b0D7xObn6kRzzFVxllIo
Mc33WnUN6N2yGB6uI2MgItTcUp31GgoeP9SdxxYJ063x8Dit71C095k8y92v5285vkGz8JMGB6d5
KaLGaUX7pbt/ERt/Qlm/uMxx8orC7olekjSXuL1Tca0J/BOJaT5NSkez6sS6Ejg/I7fn3DnK5lVT
RpOPqsbZXqvd7fPnG5cFOzscGHltpePry5nMzPoNYKJz4bX31NEmKA9DouvVzX3KXbnDfSUnLoKk
LvRG0tugSmaCVuirRBXJ0uHFiHzc5J/5KkobFq/EslnsaPY1/LI4eaNM7zfZPZFA2porNaNE19KG
HNzjFTRfsjoh2hAOwvY6Pbu/P2E9t0Rx5NZTReQwt6VbGvbpNK3n63HLKLrZ56mHWoC1o3GFZQwV
cqz37T49KwPgf3jSpnxXwgmEW2VJQ2AVybyMRKHeC+DkNcEQRP69tnnVSMf5HaVEHb647s2OE2Sg
nXmbMinBxJcpdlMXqoCThTGG6UPhAKjao6p1/01z3xz3bMh7bfNI4lg1U9etAy2ZtNfdY1YdTBYy
Wu8j62kc4a+5uO+cv1ZbxmnLdXNG/DIQHbzC4s0ZPRIgExfqJOaosZUcqzwD8EkAnJjJpxmiCdod
MvslTuyg4IPAiBXPqpAUycZx5IUEfzZAnLMZFXzgPZHx3Hk+UabWNIrGZy71aqmcLGD5UmwXFFA8
3/izR9XKPA4uVZYpRDwCRlQbOZLhWMLHU1vWdabqSucZA0SM4kQICqOQ27kGwUwo+4tKbBrThep3
oIWynodYNKIyEVmihSSf9t4ZwCxkcQ5xEKuvXMIka/tSKK0it+DtQtDhjpzvC5mPfi8WN00yDBbS
8fkMlnhVPaMWARIVs9LfAQfvAP5o1UiF4jz9qsBhdSD5MrO4zGnPbjFTL/9ciW/9o0Ql0prPShPP
4qZfM0XNNXvmKO+LMncHSQQLXvRG8xTHghmrKlFibsabVcPAex34mb6gSpOITHi5EUX1uV9adNN/
rJjZg5xVgo7czGDj3cqzyyFvZjNBBpFxieCu9/VAs9Tv/iJBZHiicP1/iGrw0yvBwyeFiEMkJrvk
OHjwiLTWPsJU0hI2lwQ+on9AfI6j2tptx2dNKpsGkHtBwiTWfT1Mpu45pgQoIb0DWMACYawQPRe2
PyH9uoFSIqNgUU3IvxKP+KmosSEhx3qcCcH81weesCPqS1k6cHOuGeD8uRoL7m5LopInpOX40Gtg
23UiQ6S1Qmk5akx1C44sQxkyMIZyMCCvz7pNyEJUk05M1glsT4icXuZRfMJeYIwB1eGmVQgOimZs
pM0r5qzTQmt6nMLfzoyiPSDh3gvosru3DezsavnJ7cuQmsfBaGAxo88CJNAaHb8dGcM2zcwctHyG
Dfe47w1RO8fbh1s8KS6Kbrah/HdLY9qptBQzsFrjy9rl+Gt5pulVbjDOhQbXNfSQs3ail3b1IsOr
kqqxRtzNgZid5lUMIstWYNUu6p429EBkHIXJFL68veG5oNdHk9qY/p3LhgGGl1m27TP2BJFYpbWP
PRKVeeTL+mgpYuypemw01x1LtEqvD11sL3A3knn+PlEKWQnEyTab27Ow+akS1otOhZQFonTcUMno
qy/cRv5KPdO3MdjDIKLXSTlIjrL89afFnDZlZorPCJSIJUXpOZ+waBrL+Cm/XeBLquBZnoA4b9oT
0iWGm+UU5MrpzEp1Ur8EBMXxAUTFWwAXmQhs20OHuLIrd1B+vRfoImCy3+suRC3Aj5++w+2vXPQG
gLSauoXDoIRyfTn56PIOuWfzsH2XecV+KI0R+OKJE+ScalZBb3j73Hh9IyDt5t5GA9Y+pBIiiTlt
s8UIPtMkz1pbDK3BtFCgKo2rWpMnztEYQCpQEAD05RUSYAj8v6TUp2doiURNUd784HT6U+pk32cg
ItnA7M5kOvLNuWgHyhfAo3T3gJOj4ux797CJf/L/z0560oZJaiArocX7cjy+hsvXQm99RE8LUwOS
W6FjebyQKdQaLKO1BRHAbX4OLO2UjXPBqE8pf9zYY2BiQh04POlP+e6VF8JqcXokGUmFJTHWJXDW
1HQU1j1r/G2OAAKTFINw9bRahuh7wDpuDb1hxpls73PZwJtnNWPK7j5CPLckCpKQHR2jE5jIo3G/
yOQY2DfdLf3mxbDl0c/kZU4shk55oUjDdh8DkY296KynuiECEc5SNw7XUg7Lshtzww2cmXjUclKQ
GmbWdMLMzHmBeqaOWr5FyfdWOe/4R3XZE7Jh4iVc+LoLQAdQHGjsLJuOSOfUBlxCZJLDuH+rmZck
3/fDqsa2WvhZgkm/y3Y4GiiHxz5kjxar565ePPaGxyiXqSWJ2BQZ5OMBvxdMVD0/VrhaAfpB0FWA
74MET+f8U7B1nAS+D00TqQavVY8kYmu/V9AZ21Tu+ro+XQAeqiNjkSWMGQoVk6gzv+Nd/t+oNiWh
HSqMGPbQlaUhqhzmZCAaSSY0LGkvM0fNcP6lVoIoBiyoFoMKc5vALCP0Y1aDHiTmy2ADY80I5uCk
EZAVqqgR/dXA/Z0PdM7tm4d7xbph80RSve0nzGmyZG1onAbgA0hU+DzT/56iOgUAu3k6BygWDOiO
W4qo8m7YjJZqPt6aBo7T9rYuJfNdJFXiznOn0JCpjbmN9x9r+TQP8ctTntJ4ZuBvg7mqJ41LYPWi
C8j1YRqZGXblTtA5QcPDzEy0ALoTrzzJWoB+aYqUdrM1Ms9EIdUObYoxu6jkFaojIhKvmCjBzF+E
DzgBE/toYQrIM7ksOtd2QGj8BhSd/2Cn79D2vlxgIQwJks5+kXbuYPRmfwNAP+5N++A3LRu141Kt
hO85nP4HNfk1zfqXlLGiwuuExxv3GG9N/MrYkjYb8OIak9qQy89aD6V6p35d6uYwfdegw2+Sc46W
ibJevKAUn+5dP/BpmTJ6hjcehgDc+JiAhdgnlElsXfNW1FekwDvDAARF+dOi/n4sAIAnc3KUGNxs
A6Vfv02h+ZcZQFw76Oj8vv/zEBMeY8beSeNxqk0ZUptDdHF4RIylqjWv2e8XYmAVrm98qxvDssA9
iz6DKF/KJFtzi/riOWORP0a/p5KzLHHTtBrAZsxddps015rW1rOgMN9QJoNg/Qhn4LQ3q41yzhs8
oPhBmEe1u9pASY4J7zTHvwGHeXgO9Vhl3Ak3UgJwfARn5zdG/ssxkQB60+k4bHT2KaYE6Etz+KiX
Obur1arj16rsqIhCxTTfCQ5navGbebC4e6RHOrTTTl2luqCiRia2RPqIVtHzzaJVWj06xXtGOtWW
GizPG62u3dQkIa9/WWvyD8s/6W3ZxSvmVV3bsUqh0m4k9XY1fbHeRV239CB/jHNNleWe877s1an6
utugQRrHzR+r3a9dCf/Lp24lUCRVh3zONAzuBwv+rLs0wGHizYhKoyYGM1JONSvv7J+Vkx8HhEaC
1tvUxmseFQ0a4B5yKU+3tpPnY15naW5BiFYRuRmfOFVNwJo0AtT0Bcnw5A0ad0Y02km7qSszy9Wk
yWa5U/lqNzGAwHf3Xff6RerKSO4iUKrJsiBrxt/v2FpS7cbtpjp5L1J1oaZk0FM775nUq6XqPAfv
QHLVLbZB25yfJhNv5F+eHcBrkpR/rVlx08rhoMRf+4MNxmUAosoYx0u+lz5itmhBUkSV+xEx9FEQ
3a+7kewzHW7scAswJ6a4ZQePvqbnlCnclzFIWs01dBhM4EXZPXypLZAtNVfQS+zZOjjsl3pwndks
5NYhOASyGmNZiOLdCJVFiMVWNF/BXJug7f0M4hNTea0kltZCgUnMBpid+UCSATTFcNquYeMmgh+s
bJILn/ymigHUToRa3XRbSFWwZjTf1CN5MGjKe4Ou0hwAa52cSnCh1057xXAY5Yvx1x/vzfXMguH0
rwWtaAl0NwMumnOyREyvgWLZ3Vijt/VKbQhbeOkVn8cnkoyMGut62U6rtiIMwaUIIVbuvjL5THa+
GRZmfIYvtr/N2qlIwoELfFda2Sbm6NLZ8ItMPNX3KWN/7QOD64BO/bCDIpxvqdGcibcz26HyxU9R
VmYatG04AtORNKfxWJjQZJW0I6zv90Op0GkLYdQsm1t4PHO7s4+Srx88rgivjAV607IPE0dTV4DQ
trKJBnukg9tAV+hKML9W4Uri4NdqBr/FxXu2b261o8uHadh9k2uGYZ2TDs2MAvErjccIZkokoY5K
LvN/Mhzj6M6yJTpIB8iXHA9CmB+x0YyCoYthG+iYoypxirLZfSYCHl8zngfgCDX1rMH7buRvy0xR
rmzpDnxxLLB83AkxuE8FHj+qn+2XuIm3vx3Sjk6YJnCujaWLgYaExG2XzLBu6gXu/WOlytqH09jF
tgTB15vTiEBnVupaitETCZm1QDM9hoIjj2A05XTFrxGdMzU87CZIvwh3aBcHno/ekjA9OtBsBnlY
IJRaXCwoj0dY9hCK4Vr28WqsUR+3yEWx3Ir7ZfSDsbWk7XpOAxa8U0Qz+LoSxuY/r0YHLwQkzwO8
PQpU5m51DpcxCL5UWxeheRGbhWQHtg2MFnyfxhSVZ3uDXeP6TbVnask4pBTrY1dFwp3ShKTWp92n
Z9sHJBHFWSOOldU/932FSklGyGN42y11lSMsZ6Lk/Qf7t5e556Q6w0ndCn33wVVgCuZdbxInpbp3
HuzP2q5SiPRAHFOHhQm11xsUaLQ5PbSz1p2R01wl+ZiYxH75W9OwT65iM7YgxQXxS7pAiaz0A+e0
BmGb3oMIFSsQyu6zIwH5Bp4390tyJ2d0dc8Qp+RYTJScppmlJiFilFTFc6DcrAXWV0ITfp8tOx38
wLfff5rUKA3IID6ASOwWRf7OQOztbW/Y05twSwgu2dF30/xqoAeHmFHXv5M4e2b9eFDs6ieSK+S8
ZZ2DOdIOvx8TYu0R/AAl+lB4fN0aW4U3tjXyigqTKHCd9NTx0KV3bQjN/DmT5xzrGk4TvcXE/d19
8aZzHnexFnK0SMqMyOFsfc1/xdT9ICYM7Yvtoet88gJkK4mGjFUnb169M069f1RMyAPGZdDWuB+V
KIPK1kdMfyHtojjW8eihuuMbkqaNcCgvmWSZDpQnZwUKn8eM6Oz6JSdSJM9Mn+Ekh8g/noRsVP3X
q3O6ZptsJYTWmUekB82m6/LUIquv3ezpQGiaHneUKOSL95e26NH2WYiWIodUurUvowi3trAK/ij0
paVjkvH56Hd/AgIzx6Tugl3kpYHHlsjchz7uJAlN0VSDrg5ne6gl79OZ170X+rgk7aQXcHBugKa/
StegwFyC4aZnc4RQsu+gNY4WHmgejkL0bOLuwB4TzGCTQrlSoy3T1P/Py0kv3aaWMn5/KF9028bh
DCwG9rfmhA1mmmOaoswV4FknEn3kt4FmQZN/cWOWhfcIrKWDjL0wxbXIDE2cSWl98joePkIXzOSc
ZF92GpGTtsGX2JBRXAOsw3N58nvBL8M0Juv3XK5ISqQEU1ZgJu88UGaBE/6z88REfYa1RBQRQpJC
rXrMXG6HHQvHHwfZLuWo7vELGkZXH7BqEiNJ0ys2ctZfFq/M2NgVVP9KS1DTqyR3JjMS8i9fuCZ4
1BduarjD4AzNoYO3zeVgnUxidIMtjwm5anV7InetiwSmfkmh8TxeGggLTOToKaGXL91FLHgw4KX9
ym7DrBrhldnN/G2Oi1+Cmk/iglQpIC0M6FdQVE0dGsD9ky1M2srKu5FywMJl14e3tWBh+A12VBko
QHofPiSvzuccG5CwEmitau5SiPoY0PHxVWjlXGIH40r8mXDkSzhNg+g9VSiTjfJ/uZQjdLJlynY/
AmMQu97VVS5Nq9hQaZtG1/9ZNf60G0VNdi2xvH8IWX9GuHuSpxRvclQComwGZfiNKAy5lweELZdP
1gTNRN6ZlejHAqKyuildiFG/qIzcaIf8paf0NqzlANfmLzisns010OkGvZK43InoWDPO7YODBgwL
NoVPeQRJbPokqVZETRTd6Rh+m8ra6A1owIHe1HSpdPVjUYwvFG7KlWRgf2LbYo9rkN3YqQx1JP3n
YcplHw38WXt+0u6e0Jg5ghFqdL8NKn/AxsdTgRlxhllSYGsKAMw+MpJRwQMiiI4GH8TSCiCcOhNE
H2Rfx0Ej+OhKKjE8KfVaAUFZi69orfefKvKKTGPFCIKlMOFaEWyaA04s6/9VaJbfzyHUoIvuLj1f
yMIv2uL4SUMHk/bdxRYhhCpqBuyiv79cjRoYmSUDDmqdjzLUxEW6E3yyZ8e7NG3puVfxzfBAehua
qyF4A7uc+MJrEceS34pRceiBakisOb8WzZuH82YnfoSbubvwvr2JNq2dfuPMZZ7CQzmKi+INTvzC
lCymeCkuYi5Ec0ntPox0jO+7DhDirpPXDmc2yKe7PRXCYVBpcr8j2EpO+plZKvXSRaQsYUqdLc1K
7h47LS/dniratRPCYgSCGVOf9SeLq8cWAaxS/A7jffdtBXE7FYjg1aUQ+BNMBMet5h/Mtxk6c1eJ
mQEDIyUFYkgZQbcea+FYBItszL3CThCu2jRsNOaj0HYZr67Tas7UJYjMvGBIV3RQ/nbb1Qqqf8QG
vNTsV3+yWAEzDcuh6MzdCBs2xvzPe/JvtFATkX0X8kAQDTzpxUBmYpKiHGgUbZRETVppWDzTkoCE
pNmhdTGkBJoypP+URX4fios54ENRk4e9KiozDUt0T88LOrdTa+2hUexVMRqZpyW3jbOtF0Gl08pf
f5mAbPKpRNH58WHOLNj6CN8UCPPnnnj/YYNPq0wM/8hQ4fAM+htFfBOB4vpIJmo19HRrmPx0X8Ai
V2LBoEOVpHYkI6VfV6v7jRwGOaPkJIpfGxev/ymKjYZh/L7pBRE4WkQXdRUZJSCpho7tv+hGlg5N
B//YKe8m9i1Z+33Xmk0mZeqN1gSfKi8S1Mv+R68lORzSBGZZoXKEESO6s0jVLlqaG/KPdmsoU+Pp
kFONUILg+zpJaKeOjTIWypO8MX0tsNbyrAg9ZjyQ0gyoqruroVPhZCpxTAL8m62mLGwne5ixKLrK
dPc9XYXnI+anPcfmF10A4MIYznO1iMCLDdvV763wKUm4OqYOM8l4R9e1XxccR9H4MHs2Lo/EikeB
Ci+rSzhktIWeWl7rkOBHT5UyayzjBoth7xfpoglIKIrKJ+j8mYoPwUb9Ta0NlcKmayTPqvVAv8Eo
D0yDxPIl4ueXJO9SkkNaPv2F/xkV9M5SGmcY/CPo0HRuapfrg6BLANJykHLQuJzGcK67bohCbUsv
ePwAwO2E6dvaT1jlFi55CLurQRKzWhlHu/9pUXsYaMUu/uAK7+fEt/8DgrN/BkcZJr6cMj2hGDR0
C82M9fcofFicw3GZNkTaM2YxDll2p77PRJDvsgOlNadAxNUDud1SG9KVCOJWsP1wm91NRm+lW5BV
Tw9h9jBu8glu6ML37qDeJrXWHzpkn1hQQXApWUmpJl8OEmmuPAkFBbyAGxJ8cJd3JVxCTUd9ijJW
pJinspxKikKy2aRtiBp85xShREp8o5xl6GLrd+pNIPtbSpxcAEuKTH/3YMYtJEvfVKSkYHS63aSy
PgDAYDUy+b/WYzwar/wUsGnlW7jIzbpvvK2vlir392OVijkp7KSYlsXbjeY+hXyt+dv+B9qnVuRo
Q6CPqLd03l1j7hf7893bwwijkIyb0pC80KpjgPPw9U4Bw/BCqYahQlL00iIGmW/PQxo89yXY3fCX
ld82ucP0ooIlNb78wYwW1LsSd6xD8VUIyKzigZOEOKf0J7qgDBZywznFmQinhvkElfWTqWs23jCg
x6gZSs7jgmNS72YhHndrSapb7jdLZa8ji8awTm9bHdLEFvYDF7BDCfwzMJT0iWU7dvfqwThSBqWS
v8TsA8zw0TIw61a952PAxX4oaXqPYNiNIP+3tm2RZAaX6j54NhpjBcKJ0z2YLff23Aw4Oqz+hT4y
NxEreW7jPZjRuuKbGNxs2pI600wbyA+4HHfRjWY8ZfokIRmAGag+WeKsLUFv/2M+5j+twYJrcYr9
CKt2gGL6JR0bVmnoJhiRtoMn1cDmaF2bs9Tz80vuZGk+mLOkEqTuQKI/e4gHx4z9nQWspNrY+WJH
QoqsOluW1zzFZ192YwTa8P24ruYpf5bndmPkJG21LbpMV7uJ+zeXvL1fYmAKpDQgwdjkVsbd6tbe
Rvmku86UB4Tb7cCvnwClJ2GIbx1cDLSk5aVDn6+ZjgZu2DMtqVnEZGU2hj4SpL5pFQsRRwtn9Hge
CA/dIIZiScYDs14hVYr28Ej1+sW3MjwqAyvKSBrgBb+5ZZ8AIpka0n0u4PBVidz2U2B7986VHF1P
vd8dX8WH1jJoMpi2VT1us9N0heDvWLNY4dd4zKGlOJy/6/bhUH8279LwFKuzkaWzWMytzIH9NVWr
OiS1Fa23JeTUCWDeWX6WzCw2b9GZHXNuqnrDysl+v9Z5ePFKdGXUrzbMAMoH2UWd9lHBtd5vsFB9
x6M/EYiAyHrhDvckP2FvKybqQmVOS6SStc00tjn2c2hWbIDXJQNLG+GhmIeG3IgxYynEB3/BPNan
7uutCmEHQqK19YWZFmNHDkMw7aTMNOZZZuDK6RGY+DaQFdeW8GJWSUMmk6yiR3gYQrVueiBYBVqI
Z5uEMRolyBt0MpO8kWTLkrDgpTQH7pHNRS5WHk+Szz8EncSTegETHM4QlEa7LfVaMQjqOherc05k
igXEQwnokJLgFRdhUmntR/ZdQnOHXlTp5OKx0AthXt+ikI3FlcQWfTajRIV4rzjZF47/7J1tPAhK
36Gx8IZBGiwGUaUaVWrkYG+UelWOjBq63YY3aD/6dCd2y6+3MDtv/V+aoQS2mPvfvZil7mZzQkol
CXBxdxzuL7OsM0zeGiCn1BSwMGokdIeEi9M6eR7mJL/gBUgOFLKLNZBKqdsmEGssmJTRtAIilZDg
0bUXidiNz25TF3IE8QIBin7F+zZMB/BdWztDVoJLgemQDuRrLYSwFOAnfpxBEqWj+e//J2ifNhZw
JkfXnB/k1rLHsqxo35Naob0WL+pHOh6SK2NyByo7vDYvHwNHPjfWPkAu25hC0Z2AXPzTm2zGldG8
nstmsZpmSAPrIXo00lMlrCnjcElRjRp/wDRaikrw1u2X6EhNQP/hQQ3zX40mnaZ+D3TRU5vi7suZ
saPpuIXL86HhK0Eetz+68xiNMOXE/XhqJxH7sNsvtuhSX49cLyTJa+SOlPsC+sdeSGsWR1K+ojiW
o3hRcsyPwX+h4afbvd4JbX8gtC/WeXcNfyhacOJCg9NJD+H2rkNviIS4x1nqwgk568B8nDaJAoRn
pYf8p3jYJYrisjSoj1en8dcB6i6nD2fEnNQGK4eYXp6ArHtNmfEZO4Wb/9VhSJIFOENGozMZWeDw
+L4gz2UdXsBz9LkRDQ2a6K+IUocEZSEaUXzCKd1EuoVvDNRLL7iTo9YSgEfNxKW+IYDmjVHYHyEz
vMKsU4/eSoaoYQUof81yYpSaVwhqQZqb87Ms4rGQ2LRsRgEoHjwYE9w8W6YyxB6zcmoIkJ+ufO8G
dCk9eIO0emsb7tSZCH1rF5cU7i4FT6eCqrLcCcNdv43UCzDjok1LiBgXrTBw8ZXRUOjFHMNCNHzq
u+rs7otuDcvEfGIX5KSuBkwNf1fSgm4RHiAYdMA51SuYAnrY6L5/trbJWQSgF1LX7BnBmcNCUxIh
MKxJAyp7msRn4Gd3eE6dYQEle98GvwwkBBjJbfT3a5OHCx1FpE6ZaY/X9VYF/YKOemcTgOO7Yz+1
AHa+2uy7xUH6ZXb4/KaWHq8XYb5L8+yjuI/0/8jrPnNaJ1hYr08IoqgdXWIOx90omkXr3gQumaKi
kO4w9lP4/FoFKmM3xsOvkbyv/zBeNf54yS8OPwmijpLn/sWO+v0D5VONoOkTiy9lV/5/B53DEEIn
ppyLe+ubUx6bewF0xOBuXKNaRaTr27iAD8WsvvMACJUrJQ4oE7FysbU3INtPmn3nG102wnnfOa9G
q6fjs8/stunZj4zV9V15Ks0BICBKHmWSWhR4ph6H0lvmbB7EVf/J3cJ/5BpExe5MvRM6/dfDO/yZ
Svjwr5q9ksJxlBl1C5p6IWYQW4Y+DyZiC/Ru6i6XTvtz3wzGvRB63osbEXSQ9SHsk9luW4EwEKZY
iYEyRXN04l4PvwdtnqZ8mXiJSHR40oOOeRWNyNIRE9Xzb8kshJo8ulToWXKD7+kg3AA5BSa6Tj5+
ULl//ocr0mbxUPGn/bC1xrGl/c7y1p/5Z5NtL6H7Ka4/cnVqpcOA9YuS65Y73rAlmww/CWDdAE2W
K41rJToKNcmNL1Gr3YInvMpFYO02nPN36BksmpMMDqYP20ALWmuccXtMVrZonDgx2fmHnb8xxGPu
2YIAttIXSGoYxHOqQiHbuKiJw+aPLRRm5A0K1TDlMqK5gu2vU/Z6Jzwnip2cRBGpA7f+bshbbA5G
t5imUPrfpADkSZpRSyZ0brh6j+2b7fBs5r9SyM+3VNrMPplx82BvWbGb+6+AQv/DCWdPu4y8pdzC
0LoBFpU/nVnRhFvaOdNNl3UePWaZo1oUXgIMN/gAp/YvUsn9+XUVtio9oxyvGoK0H/DxZCAFOrRT
QXInqLjxzPxskH1O/ADg3XMKLoiy/WrKCnQ5SzETKd7oDYy2pqi+WLTuB6crv1zIZRDsYGPGEy6R
Rl5iO8PtbFp535VPh+A/unQuZsGBYHTqkvOf+u0ew3dJ7+Rrfvuu6+oaGZFkoUjvRgIyWja/oOrF
oFCwqV2VwFh1g1Fi5clNeQ1k6qPZ11uD35aMEc1iYDs+8qAaeU6RntBAsXwE5D/9Sm3VcdIoUZ8s
xGov4TfCeRQG/jT0YChGKBY9rDLbmkYuNWi7+8uSqSaAKER9Cpzd4J4qObO399IpUHrFcpvIcyZG
SydoArBfDWCCAUTSyL/VWJpV1xq65GolTYvf/6UgdYUneDhBaQi0lx0lkOT9Lw1cOxS3Txr2/Dcj
f47w9jWt3kY+e+uNSRV2Az/qfVclMUlyJIS+DbU63M7hYk2RUelV5A4BsaIBv/snzGyKpfYxx0Bc
L05FvcINL1i5NhDQyiBrvBQwpbHB8EqUzyOLS9SPyH6mg7YUPa5CFNhSN4r2sXNkqJCvD9WUaJV4
y0/9NhOo3yGSfMlznI8fp7vsiD/YdVAHLaaJS90Xuj7+PIr1gZ1ihecZvusorzGixjaDDx8BUWpI
UilWbu/joEFpOnXM6BUZegMnyTIyzRVrfhRbboE+SPK/WAMUA48KrGGox2Aaw0IVllhgX1BWEEmG
/JiH9tjslScOND9dPAS2F5JbLXYNylxKgRHnC+vlMMD0IMjEOQIVnoS9QKBP1rhA4gMaCvnhgLxY
/1SKM2tM/ijexPM7yvAbxWnJUMnha3PFByRE9ZuI7ftLgfLLln0o1oTuWZP3CB6TvhvqksLVGuYP
k5ANzFs51u8xx2EcaL+nm5eQ2s6HhqsSEChDfqMB+evf/XiZ623bwnST+V/bMfVIhLlay2rS/LTi
hlcRJr0cbmMweP4SmTzYzgYaoUNh0qRoU5wm3dBnoLqfoTYG+XGRAA5lEO8WhA5bd2mHNnxDQtrl
XZxJUfBnBkGVBifn/DxhPX6EoPUBa7BJy4RIXWJP3Z1m41B7FK8MtGqudMj0FHMKEW1Ib4A8o43t
U9nt1CKNKhDJiC4HmSnWj85dy+epKaHUAUblWL5aXuFOQa5URgB0fdcy2SDuexwh59nxsFxn07eh
UuUfIJvLAYOOLODJIJ6KhUaucPTLQvekpAtmvVyQ0fv7ScHwNFxfFhMLUyckfZM0LByZyakmKKHg
+Fh8nddaBaZEo03uSUqYC5zWdksEXGR1OpUYzltY1gOPeAhfeJaZPsHmsYosDk2CvEJGH/T3YhKZ
uxZ8gXkqLAtzeCt/A9vdadZ0f3Ju855W2UkZufD8HpRqutGdSLj5P1N0+CUgSyFSxyRx8CVgRkdp
kQCnxBLzmyFmOwgP1klEoWNhxRH3J6GcjSqENDueyUsYSJoCpIsbwj5YdgXNneObITIHU5wfxpB3
bf3fw+WNmUYmof2N5Y4P1KUgtge+M+p9J7r/OVjt+RdQW93ErpjW/Hu507CIJVH74cg6QZKYDbyI
i/MQQkZsGHx3rN0cITTEw8p+xkY7y5E4DRldY2Kf/gae/M0lJ83lzUytuBRtj7B++bnSLjfbjwV9
pIDWyEWECb477ME2wIGMSel5Y9fNYh/oAItVxGRVjpLTL5DwkM5mTLVzavRnfTUImaujDksEab1a
VcvNmCHrucsOu4t5UJxyG2/71dqa8Rfyo7LhQenO00ol1qEQQxh4COaQ+CoQ8Ff2ujoj4vJCj3HI
hWpfuwAq7Boe7mW46tpAvtSyur7PVmntZnhiECQfWe2PA3n70jSfZ04V0UzlRpP/hkhbcnVOBkbM
P61DkJ3IPzeeIkc1GJcvmWfgdtES4URWcJKz9P6dNqH+J4JeUoIfKVMu9W4IuP6OvMq7xCpGpWrF
qeUUz0BsLYYJrErYJVyX+2BrYBBh6IFh02UyypHJNruPdQy1QlQh8m/XqSfh82OCa8nSy/w5guLg
zBn4yUI4jezZgGsEFFjz01drcDimDYCJjv5zysF9Iz74xA4JJEFI7vKz62SqZzZj39a7ayHrE9LP
KlKZUx05PvZKZbqmI1Zgg7/y8wk/I0GeoOmQyA09HEFA1tAlJzF/ZgIB+RjRAkgLTTeXjZJgRAcU
JymNqEFp/EqBo1lkJ4cyVnrFiCk06oK+Xij7D/iCmroQjQkDw/tsRhJ5Zc03QfY6ECenO8SBBp76
biwsjlXBr8AywFQvXC+/SVy8T/MXkAodBC/A2rXT4akq9NglKaf4hqPkcQJ/C+whUh0ZSwzIXfnu
yicui130uxmJcNWDrNHZv8EXYuM0BQ12z9qT5bM/CPdTkwsAG35zQKcaWEhrTMWO4zUnI6BhpDlf
nY2okfOvMmSOlvJ9XYN6mZxDC3mOEPSclWaCQd14oGT4ZJgAbcy6jsdBiT+kMVMgEQo5yha1wbnW
Evn9w4407P/k2x0RqvdL6gevlotonKoj+SRD9wRyYRsgp6IF0DQFlYdGWmaK+e5BP7jn1lF1lUOE
+fKtesY5GEvJ6FWJtRLH8mWc5M5x0enjrWu0DAtUWtfzhwNgBkx8r4S7pJrTKClmMqUhH4C9B9+b
bdmb21QQp4U5PPxAdO3ziKKx8liKJYhzhmtPacLvu+GCvtzFm2I2CFCU8c5NIY86pybVEKuA5pSc
YzHhq2H/DmVHgcCWz+AVUNcdjkeV+G98qMOqp5JST61lfoaPr05k9/qR4BihQ6KS90T4qgZBxRhd
m7WGDxLxvMtG6vvcfkn8ILHmrWOUH5UOs6hy+SF/4aBq+rsBXHdUw+gqicMcKu9HF6r/EQgBl3tS
kzx8xrT6RAqLJtUo6b1b/8e1wlZzrHqrkwjTdv7NcmXwvy18FRMuMBCBzJxcDX49MD2otrWZXvML
O8i9uBZUo+Eisgks4zXsrcD+VCiprihMVTCz0Gx7MO7QTGWlBN/SeUeurCCU5nRTp2J85rTH6t1c
GVFJchqp485gMO2HaLVL5YgXdohY+8T8Asxn/ck+njmGESywTbXNawS9HvGqRWzuw8ZWy+m9X1dM
lA9WotqN8DAOUFtCQyAK190R+ytEQbZlvkONDODUxTi9wxdCKCmXcqO8mrvp0LUbdJRX+hfJnnnJ
ISKGDP0Zm8K13ienGn0472FuBNDC0WYo0drHQpBXkyQs+4yfj25l7AG5Gc4tIE57d1srHDktSqcd
6Qg4oeV6bsdHDKxyXKyRZrz9hajBvrZ89tIBzimR+gScOYY11IWLm2fD0HRuKvIPo+LPxO+64tJS
vXRLSlMyvFFRHSJ4QvxktLqKjRXcsLNgHnH+GuzWTkwX5rcD/CdGXwJOGn7Z7W+BloKim7kevvOB
XyLFCNZzg10BY5/qU4J5GeLdXHVx+vgGHvSFk1n2S0ZeUX6qS7OAfTWTtIlOS7ZjR1QMlEQv8piK
ElnWc/zSLzZpGNiZT46LxTVpYzHN7TK0jLj0Osu6DYPxXaOXtc5xqch18asDF0SOMuIYtaLJvcs3
FKrJq+XO3YabP5aYN9nS4JuMuudwXzgtjv+D8354fA5CGhre2sjMzmnOTSJvPLJLzbOlAoyPF7xR
ljUDzC1CjOkem7anblVL9GstvH7ZVgOan6CK5BQXaR6rKJyRy5KpF1mmT2lCaD8x7LXSd4Vijoux
RmDThwf7TrgHUXayWWgV9lAmElHHlDYYcEiH1zzMo9RatPpnXLxkpYgXS6nxqK4IinMooJSUdhSU
NGQpdrxAtJ26I3xSRhRFwXdPwgjfX5CmGFTNJbPXFzMyaIj5IijVvTylfOb+bSz17ESPBhuT+BKh
N5PL0RHTWtGJhgZUbeOdJEOVwT2p8SRFgkdDmXoiZ+xEDRYF75VVOq+WkyMzd/go/5NikPlqKYrL
LZzedzQt9qfPG0qaIy1HkHfGd3mWKZpYvIkwsGbGO2nwvXBLnlgunodm4jxKI4fuXyOEgD7ZX2Sg
fK/TmzGGf/825oMWDy0oJ86jxtNOC8BkyYVpVm4a/ROD0VD+Vg+mozJif3L8MGiEBeMAN94DRYfd
APIEzdMuS87HLD11sCG0D5Ht5O4c8RgkgSPhrzvSADO/Q84axCZsvdP5de+IWFT+F+vlxdowgdNk
59UKJ34Lq7Qha9sPZ5ljAoBTFsWiTtMC1nlUG35YmyaTSrShLHn3WSXOhGIBM908O4HnX49/4GfK
A5GN3hfViNj07lZdv8J9UEi8IHFT4EVb2uqF8hcr34bkgNSP8W+/2jHtF1UfFo6Z30qd0axxYGOO
dq4bHgTLoBaz1HUIefH6RCr8iNq8vrC+f8yB2aCDj4Yadv9XsYvR8KA3JfKObPErGpQc//0ytTwV
IHtDMuhnfLu8V3D96s91aP3/IzgoJmzlllY963GzhKPl1LsFdLI4NBd3jbnKhgvtp31bMIPUKK57
M9L1c+j09X1xvi4Ox0TeqpTbaZLdJGDWFq0VY/XLH8fXsJHhA3f4cMv/IqGnRT0t9377h0AtcMz3
w26tbGV6ubFhrQhXHOXFsDXe8tTbTp0Qgrisb2OxKSlWwKQeDwWHFoyASbFDzWRufTspb3Lpjkfq
Ac3RCwB/Dm2N0hTgX+DpZdcwVe5vd77jslrZQMYscTwUo4PkiINc68Kph7pe0uerwDaVFa0zQ90J
wPaA3p18FBBLkn2W8AcVin1/npYefPyPYnxY6OZooFTICVOZiHAXaVAdqxph1jhJ1Y4FRuB4StwT
ZGMMrxQ3Bev/bruU53qBQVyyz3JG8AawwLXNq8MHvXKl3tBRvNXwWkVODFYx/boYYo4iqrc/8lo6
0fFe+oio+XFvj0HK3YpyWrg5RtrotHZo2WlqI6s7Lpe9o1UHG84AMcLsTABvt05wV0geiZ28Qid7
614W2XLUGlulFOScnH1Bn5RIWStHFFfVmtqqqP5vaK3yweUNdn5Z/h3pXxO7L0EXhusKNBrHnaGy
JTS4UAxdxDCIW608njQK0zN6UXM7F4nClI1791ZkaKiwCiu0zzhpBFRe0T9NszYxZGYrUxjjcIFk
DroiC/Sx+kNnNZesaxzEMgJjwfWFOgcAqbdrg2D6mNbSaDVQ2cFNxw9yoN8ljXSbgoEDABvoNVgj
OzZHE5W5uUybSBxgnpTrI+dZ3aHs5SJYXt2JQsji/udNIcoyn9mOwmnoFVfDfJytOnDMplirgssG
sDvLghCKIDnMGHVIpr8BDu6X2VWKVfAMu9rcqkBmbo4YnRIcsvNZ0Ke55BI1EBo1FvT8Cor12dlG
IhhRGj/X5xkuI6ehHrCWPLr4aiKOzfhiFzyZyx6UETKekdn/IvxgQjm/g8bMcsMwEpNQMUfl5PuD
3JrPrUcbJKf3BYo7N2700ZqbB8hcVbe3Ar+4IBpud0y7Hbn5hxT1uEWP5kD/J+Fo+pgcnFpn0js6
1w0BreY3qUNU9GRSe35KYE/uR/gHLpJTD0u4vGi/NEMtcLO+/bVf1KOr24f9Jd7p4MnsnGiA+Lse
al3tSBBmtvJBGzulbeS4TVZHzjP9FN4ngFE2rYxOWKfeAzGL4S47Z//oF/xE+P7x8oD7JhdzWzJe
rthSpoime1RTQpRjHK2eShk00KSIcDDNkuzZNfbPw8LuRcTy2wnza59ti3U1YosUPmGUZhdezNxz
Kobnmpe4aaUIiGqQlBJrHjytjNsKSP+Lry6Z4LIqRestyiWVPb9ajwkDsMyDSUtb2sUnHQUCGXbW
nk9zRF8ewrKEIltU2tFugZWKZUGb88CFLyRYKL5Nw97vLV7k+tg/Ie+JsgFDPRXJ81N0V6KS2s3e
Us/59tOqUDbyr6vi4JPbE7Tvst3wbICCtcg4v5u96CqO6uRX6eAeKtfXjMLc7wq6TtwrK+fbYRDc
SNsDkqdz1tTO1sqGiYlD6yYCVx2UDeDTyAedVVMHwuSxas5YhDjJAfDRCSTi1weHGc2AnWbid+xJ
KgO1fdyqk10iizufKHMkVEniQ3da259HcA6VI7ogh+sA/U5OmYsfzdmJgLiwbDKpAhej83omzE0N
E9McP3ZPfwCL1xq9f+AJwlt8YEe3zJOJ4Vmvls7LSa0Knn81/UE7tdGLNyOeY2bn3DPob6BaOZp7
CHmsyQ/4pbWLMOsXxjOPVIuNWstlQ9lQO5M6pufPr86fjKLBqC6KLM7DEvRPi2MVOWGLYmQw1QC1
VtY94lXQczlqPwjbpFqa7WiXaR+IBtYjy56yscjQNPopNO8ur9qbKTuldLB+c/ewYYDQxyNEzPSe
vOHQv17LHTj9ovP3Nz1Tyyw/YYyyH+eAsi/lPY3jfIH4t6je8dR9ULOZPo7exhdX1cQlFnabrwch
UalPssAlWExgMu2K6FOgGl7iio9aBK2W/srQ7FDYAe9IhR3v03mbH3jnH/SMgUXkk2c4xOC5ASyG
n3esEhpTh/cFjJc1aX2ztFJWVlqlmaKEm0sP3aMrgPhimU53M6BJUYLmEo/We130HBoKr8YTPn6r
9Rz+of/szzB+KtOcWr+8njUp1+BXDrsvsZxogWUgPxUFoZAzHBxCBZ/AKOE6sTBwwI7WG0kjFqZa
szdnhWm92h0ZErSzZ5amfFCE5KvfR9VIv4hpd2A7e46j9XnyFOUOc1DHJsvmU/Vzq1P7c73GdjPt
4KQS+j79Ze2VPHgtlkP4FH+TlL9QwdmG9E0MJMp2IlFRLH8o0uTKwyJILsdSg8tWx59Q22zFM3zs
wKocTDXbJh3RecF+9GcITXeD5ruCJD+3Qk4tmvAtMvfOElV7NzJjA9oUC3r9rATCYHYdcPO1IRFb
HMpgeM/Y/pmoDwag3Ji/o/TVNOMClh3I6XhsdNRDkAu6XS4bZvJhEnkT8+EMGIAyCTJdnfiDMIty
dCooJiMRCyHuCVIyfGrD03zrhNYsKt2LVPv+jAkLLrfLIGO6SEA1FXzSiPHRLbxxPscsMOY87x1/
bgPbZoO/wl+cFfgNOPhDd36oY4/3SCODf9k97T5gkBJ8EdwmMHQV9QpoTp71xxvjMTgA4TIlQJxv
U3M8OM+RK2/SU0rlquiVcVZLjztb0TmD7WlxfaHR2yU88zow+yvBiN4BXxA3PGZ4VSXKjLB6ZcBh
B/RvWh/dTKhjOQ71WfNlJPiXhRTCqLifkBXy33LeQN6tyIas081JoZS39tPxlKntAaVwe1y+XSYT
uwd7DQJcjc/+d3bfLRo3pfg78G/pxra1sfrYQjMwZMHBhmAx6pJTKg5US4B831YR7e5vhB3TBCDP
ltJiAyPISccQSYtrEDbmiOVIhBdfy+s/MH+ne1tZAKT+o/dHTP+gtTxDDt2wi2glSBDrPuaPeNST
8o1qNvtEmKrjfshbsFk6T265McKertgzP8NnFhckS9YS0kEz/1GR+XQudhFyNqIjAT4+gy0nxbBH
VcNgK+33/uKKOXGl0LZJyMVlzrlCkfgZIgylchOk3U+HRzPRIA1acWLDycniFKkYK7uph9l0C/wq
+HbxBAqu+yEDNbsQ00wCDujK2qxYgy4IqQihBT+BrjS421YlpKZKWzlBspC5N4EbYuu3yKeecpWJ
7cgB8OiI0CIwySKFvo6uAKvV3nRXQB6DUy7Jz9SAdR5JYEQ/td22ch3MFOJmi6pLyQ0R6bPlAJ/D
s38SKH/rDApm5Zk9+mFMjmAM/MJwJQGJAanj9wjSm5G3pb6nMVtyFeKsiyOR7u5YBCn4Eb/HbPYV
aYJtmHqSQe1cGBp7qTqf6vrZiaRglMw9SnVVvJPx+dOzqE7pXu/emdQxU2E+VXjxVVXGcumlQBTT
PbwBoab6fayA7pxxaYNesOqo5OXR1biY9bp6pyBWetQS84BvFDiyjJqwYq5RCG5LNxTGF8b1kVbA
sYvpmkq0P6n9JHy/vQ5YUjQzZPyIQaqcY7ByrraYdOwgGch4wx7qWEHC/YRreFgUaJ6cPxwer+Ql
n3SXe6be2zDF58tSubJE84yyuoSnT6f1DHmhApCA08egeLGUMuobwjxl2v9x7lIA1c3rI6nZ6vkw
PI3jITmOMD3/NIkg1Oz15so+57Jz/pAa+6msC3GDfo5fr0FMEAfNP7NUexOLZewYSGDFY720j7cT
KTH55FzyXGc0+rrQJ07nDj+CgBWeZQ7zPy+NeFDy4NuUCcX9OpwS04axK1A8+8FoQyHrCjJ3mxjq
EeBvex6D7QxhH2wtf47qrJxKXaiypSDoWZXovu3zlZfjtI7Sz0z1dWHaL4GUlqlwbePmfZFEp3kR
tVbIXg5dVEj3dRzCQS40SUtiecT+5lN/lqN5fYe0/Ba+Cw/96jbvFvQYezsy98YQS6fPm/2J2uOk
a5X4GzEqtezN9gXdio4/JvkHFnh8dMggUHioyLA3Vef/2BD74zsXZ0bOqV3wd8Zhv2Or/twILXM+
v7RB3vwsMcGFO3X/QDDfIncTAGpqOdI8a2Z8UI1ztgmSCsx0l+uI7pR4dmIS1Jf+WanV5xWUQqwY
cbVPk3/QRjeySwie0WB84wHPpniYjGU8NGZpc2xxRKVjqGGNeGPKYmg/z01hG+TEItecg1i/8Xxg
qZ+qud1wUok6CcqA9kWfNoFVoSFGZgrFsJXKtOCkLkM543vUvSWYKwfNGrUgKBz19aORM3KWkexa
aHYd2PZkGbuXjlPCCYSmEpqfR7ETG1UDsXKi1kfIxqjiacuF/CSrCMzZZ21m+As2pAC3vo3l1HCc
cVpzmuXkgmCeJCto6fekF0zyg0/aoIDSPs2BPqI7kFTjWmT7Z+gkfIT8rg+Tme2/r7zbS0LBSSfT
R3mlxTjkHEvLBiCOGfNxfoqLsQEyV9gPZ7kdzjxZzcUPv+ODAcMfABkSb7b2PhPK8Eg9npJa1cBd
wfIaQ65NBR+on2NmZasyWL0as6JijiszlYTf5MJtZDfaDEeZDmIAkRvcShTEWV+L3M9Uxqq9gUsL
HghoFv/vHXD7C2LFa2yxRlvrX5iztswk9Mm7qFGRemuFQ2ehhEo+NKMYxOpmiLCwnOP8Gn8FEFj0
N71iuHMpRVtvSQ6XZTYOgD2TBAyYsRNphfQtiguwmsu675sE/dvpSSyVHHz+Xn8WanSxXaEQUFh9
FA6hvARisXXQCtxvJkk7zq+DSjoyCOM3ROGR4xLWRfxBbop72PGOUwwb3W+nArqov9ZvI5vZr3zK
vbX3a7fcY9KjNSSW//+CE7oW4BX1gXAUOnq7ZDLG4ldwY11qXlQjxLE3HUXKHr8saB2rsm+iALd0
mVZyFc8TzB3EauCy7Pw+aSaQjY2EYeHANYT1zCUL4+IEb3NHC0ECo05BYH6Uv9GhmKK0RWU4Peqh
+g+P6/W9M1KKy8iJ6pIU+B7xhmQTFY5LjyxyWfrf4ViJ0OeQ9crWiaF/M/YNwsFF5h4mUaIsTO3l
ZGpoAS1FMWvQ72mtjpz50Tr4tubxJD2C8Z3xbacv/S4EJ00sz1llCGRQo8GvnFh+/OVFtb3Da5pZ
Yr+vzs96m5jvoDDFG5bXDK3u2wWdW5qUV3PqKN7N7bKoi2ehXJwJDiYyeNzjbOPdiMko+Y3cOAQK
eOG9IGxIpSopjMXxLh7GbydKwqgj/CZsNgLhVaP7L+NzSSgsF4py6KjbRjkX1sa5O15nirj/Otej
Kw5AlgiF1ddmSQ77AZaB3KhHnKXIxVVmHcElLLZO6XuX1WlnhaKAqvkZfFvLeOibZiI2B4H0GIoL
k0PiOrrl1Whp0E/4iUeDnS9M3zwoNZWVD/wZ8ox50ybjva0ycPHJBws4wvOKKRyLCZj98IMg9BzB
k5SB0b6Ew6BQOZ2QCiqUMYuLwtC6tu7n5smNc7/C6BEMQ5yzqT3jKOtw1jNaJzs1klKOdf48KvjG
cuSPHkN6W7vA3bNphUz3TV1Sg87sJ1LQnoyDM5GLW2sQKAJ3rTalGYZhUcmgT3tTUaTO1VUkNP14
yj0fxjq4bKHI/iUEw3Uj/hxsMAjExDgoLw9UGprkNn31QhBd42Apt4x5QzsV5aKq2hz9BqV/M/4M
M0EAqdcjJptg6agNWMroxf39KM6vi3urHEkl9d4Hiwrv2Ca1s77Y0PMHoepGET5zuc3YFomliRyY
VdLIvvOwCQnK+CXPXfef3GYzIIiXvRz/D40m35naasVqarlv/xWWKU8teQS0Prt6zpnzCXJqnZ5C
BW6z9JiNQ0X9WVlEbcSH6EBQzR/9ldvRFdIRd+RqM3MVIhriVDZDOnbXw2AND2f9aXWwlcxnZz/W
mV0cEt4Onxm6Ijbbzti0mO8onrt/ZtpTXgu7WZORxiDf3MNoKJ1ntwgbL67QBAYo8tIs2ySecWBA
v6P12OzBCD9Aj5G+nFDxWhefau7DpFxhhEiI0RTMwjtH/v1Dsa37XDEm6g/wRMPAPS0zdSo1FN5I
AqL2g5RsnM2Y95AWK81CF1fhx2SHf3T51ttcEgqHzlhDK3S3y0mcTKCNE5zE4kM/jfGLdxMrbDYw
FCXO5yZpLxeuG4D0Dqf454hK54B9lB6+FjxS78tHiD13hQ78ATCfXc/IwHDJ23F+GH+dFkyQGoQ2
g3nHBI+8aWHVJH1mYq6gBqhUD+oI1550Dvc5/N4xI25S/nO9jYV/THt7zGXeYjMIIQyfv/viJeFJ
XFlR1l9ClBC2fhMp6aiS/AYFYUW+Rz5kTg4kxMJs4Yf97C7zwQBRhHPb6yOUBn3Z6YdWX3TX8RNW
tM6w7anej0DNfBo8P8dmd354+ULBcMOWBPDMstdu79Lj5Wjanc9CkrJZjV2KZFLYF+3nox7+WNYj
WxRMiqV66DnF51nJKT2EUJE9lKML8yzf6clLpSZKA20EYHoTNubLZbgnjkLDwleCnU/rMSVAJCyp
Ezwd+NG7f3f9ONwAxDGSu5uw6kH9621vzgcrYzCUlA/vzmOczXyfPe1iiokvzOEZRlcdSG9EnwrQ
W3uuYP7hhUzE0PBXfnQrnZb16wRgaVJPIKzqfklGsdcR6Bw2f9QO+fjaRleyO5PVM2WkgrMELobk
uCI36mFtsZH1zuo0lvcVkmAhi3EhNJPx5WUfNyxJeqS1m/IOT+MfRoAHhFwBHo5shE/QwKNF9Y3b
mXTpNR38cTS2EGekuy4dj4LfKvUdZNicejMCtejk5W0szy+DudUlvpOFku4QflhdRqwJ2VJaWH1D
tFu5XpgpxICJxAhl3hkdDvYGS3S6jcKE7hzdosN07os9Wp4YPq8qfjwwr1vaH/AWKjAePXJbIhCN
wJJeAQA3JtYePMCI5rRVwIXcfvV5ENWc141fHohmCfwy9XcqOUAvoe3+TcWt1EWfnEOx1OYb2uoQ
HWAEk96qck0f56jImhFiunXm3vLV54GMek99CtUBtcuOBhVEFbMyQaXNToMfvUplQREHL4axp5+6
STNWW+vpvvzeXFb2sLA7iE4/1ctclCvahKq6Pls2qPmDv2leEWxLX16ttUFGbZk7QgczzHcG6vIq
KQG09s2Gfrdej+6g/xH5bwCQZotZYcLVHH4AZtSuNI0U8dQWOfKentl6+/mRHgK8jl6zpNAqcWqT
XxrUoITaiPN4z8P5IhePriCeoW6r1xzkq+rhqdJUQ0Vyq7LQ6yVDAwfznrWVwTDLPiCt7QoXulRN
YS2w0IyzpbpAgpMAP8RC4JI5RAxBWvYXy0XLqsFtyYRKRoB9U0+6yrU4GOzdWusXtV0yBKaPNFNl
CtuufMIOHLH0SSVvOCPLQwAqfYQpU2+6X7qbHUe7FcRPSucsEm3rgWaKz0f3GIPb/gJ0y8SgFwIN
uz1K7CFpkyQPlt97+C24qjsCerBw/LjbPMyvXXWuV/iqMdUg4hxpNh6chnRDBVg+V5kEJeuVWN6L
CzRgNtS+Jv73fzKauEtXk2KBDpHCwNNGyvURELWyzlOU1VJzkc/QiDIbpa3qS69tZ82pKu71PT4H
6RFBqGGyedukOTCzYqHutBa9VUseifcvHDlo8Xb6z20sTymJ2L6/8UTUT2hLlS9jfxuOsUZrvMxg
Qzj2qDLosEBjzystHb70Rt5wtSA0gqxnDYnTenlGCL7/zJxi3yXWvrP6LkrKn6mmxi46+OCyVi47
KmN3AzQmfbvsQNYx28+rSYntUYFSipFwK2tnqVbgwqyTHQTynFkb/m1RkH5dpDgEW08XNDRwPDya
Eb+b0VO8RDXTleUZ4c+6I3IqwtAg60sqxNR6kNTA2mODvA6KpWuzdpOuRevFAmH5rzSv7eHn70pd
qfMG/hlNYa8fpHLMDqX5TQR+nVuXutRwtAxYGcV3+P7N6NHnRGM2N56Jme55ulEtpYvN+3FM+jx5
AfUkI33kY80yhwOVOOYDrM42faR1dfEmUrFKnRDw1nprygTk7ZIYZB89LipLtIGyHbNenIAXQv3v
ecTiU0AIB54lKk1QzqhPH9W3HJbuH9b7hktczde9hMkXeOXgHlGX6646HBE8fkds2jDkYTuW18Bx
5QukyuEjcvaP8RTYVJFfP/hOHOAzpZK6HYS6BrFmPgvN0SE39E9jmmwxF1Zjrq2AADQFs25xkTL0
P1+InQIaRdExHhIRB2B3A+Unr6KdlrB2IEYUGkaxXuoAQOrWgNLNn1SiWmw/DFtxwXGbQhlIwY/Z
PP2iZGiA3ucB91jPJwhFZdz598xvWO+L7uYkuzushKlKnyz0+DC0jcFglZc4NsJpcFCtDiDqjSJU
frT3HYXpCNk4SGXt6/wYDENfKr4xuB9jPqa0Hz5o6DpqeQP1n9fqsViyE5JK5k+jVxHJNgzGRh8S
mVerF5tTrZ5XOLsucWJEBAxVtyGIHtwIjs8FSEnWpyTBgglshhbB8ZGhLST1lWycLxewqV3k81el
28FMWfUf8BjPYgzqz1fwsTYxZnVCG8ScXdY2sVT4gm5ShRzBCn7Un0qtv42hvV0qDPYKBn/mH5lN
TlsuDbrEVvvLiTP6sbtnpYbcS7yiw2yYfNXcOaDUP1JBzK1GvPLu/P8g94XC17H1cuTf67/rvj8m
tIVn83pVyx47/RFsspQy4slSjAJ3hpJGsS8PEHSXRldTVpN+c06FHYXvlphZSIm5IcQgYVqMOYK6
9g1RDG6BWttJUdWtynYJ+p6W98EWqvFnUfAqUGMO8d0B3EKKPBCfTmL5a5peJuvSO/8N5Wo5UXO2
V4LVezZSW6RV2nMhH/WvqFdswJ2pSai9v/FFoaFQxEqzzB7g6geJ9oA3H4Me3ElZ7zdQvs5o37xs
oNFdPWPtEEo3+0JricUaksFsK2f15soRZHFrR/WCzgKxOzjzQXfeKEGYdlyU55NuQYC79P4ERD+1
uyKBpseIxz63gxlcseML1KDQvjiGH6h0n/W4mELKP3pWwVKXJ878xkD6GUOseaJt4sL4MdK1vd9t
lEnpfX29EnsFbFCTJ9jYhECqhV2+iJo3ZLs33hWaP/2V9RC5p7d5wQUQTNAAsSNHNi9EvW+xvwJQ
TLfnqmEtSP89iP5+cnu3fADKoS0ZPYFdCIliJQs5kJQ6iQF0IUdI8MBqouH9QfONqrS9xLh3vw2+
/AX7j1kg70yIehWmpnhmo56Ej/i8x1EOpj43TcymsAt0h2km5bn+vHQ7pBx7kRoZt2XgzzldsoFh
Hi//eNl/whGsPlzMW+f5AE4UpYn4Bvp9i+mEVDPpYux4We6Ik1/z+Pkbi1cNH+W35I3yg4E9RRVI
nH4BdVbxCwFscAKCnxkYzFudHEgAYihdQf6xqOUUq4hBBf0pYBAmFq3yL5GJTZvZ+oy9Q7/NL4jm
iPjA/8tPF4GbD6xURI5Sd5QDIVD/8GaSHQmmfyV7JAqHwQUnkT0JaC5w0OTaW1+mBClRw83LCedM
G8fteMmWxt7J/1Zj6daSmlxd9vKC+wMMHlbxaKM+79OB79ZAaxfGQwTtAG72FY66RCnQWms5DtXx
miU6OttF+TU2JJ++LDxilXl/Foh6cpwhW5zTRtkJ37bSMB8Ll/RNTMRnt02CZlmVOhvy/yedcWW3
do2XuCWWWe16yHGpfQ5JZzgqtq04RcResaC0UAfcoZVtfF7Q82iAPevizInwby2HmHi2LZaC3l8y
lOExmvqcUCrulW4SnIwZSY9HMAwtAUz0YClah/YWDWiQY92f4XAzAhG3UwZPVxCf/NkcmKypYjQY
/QYgv7eXcL3ZY2FopemVrxoD+jLh4bbvPF0xzB9+uIbXjz9dhhlX48XhcnQ5/YC2XZI/Sf+Lb+nf
7pjq1e8Pwl07PXI3eCTeLAoMx1J0Oi8W9ilvy+DbnmjAD+dCajzFjsAs/tCWqZVVMJ7o8gTnsCIn
6mmcn3fJXHN6lAwYoWFlwNEEH+UtJ4n2tUWGNLsf9lKzGhYgc40xhPp4O+kRaY9GR5jfIWMRbiMo
gvxxy09ogzn6EArpK1vdQABL7oeaZIYXmAQyqiNHkSG7S/EmltTzczR2ZAqvsAAhOcGpniXbuHsI
ODm7Be0nvI78IGgfglZIJf772R8vJvv3OWVhYe+9qXkv07/uFYEGJdzsRpx/K0xCHKfyiBIZef1K
JAvEd8BSkaDozbp0jtdZfndeQQhaUQq1kFqsGxtWSyAXh3huqMfmI6Owfa794t1ks4Ln8/ij2mta
kuDm8R2SggnSBe1q0MLuxhtD4H6NFaw8GA6B41oLrBrZqlHdSaXbXYrdFEUpUTWYKfXWzNAhYe6+
x0ygCRnmuCncwsRCfycykxCYBM2KVGTPBz4ZdiaLpxjmnLQNGbpY2xY7tmr7VGSg3L56+dZ7EA++
S65UWiyBJ8vZzmCpeJoPLvZg46oUqCqlfJ7SJxLAOhB9goarfW3eoNdx9nyP6a2TQiwZHHOaIrov
Pved8nDT7TiQjSogPhSuSqROB0BwRrBHyi8LK0k7SA5cfGdNDK6C1IbedX93TJFr0xJwJEPNpcL/
KqWbMYnouyd5QAoj58kMdVOV8R3S7Ee0f7A1rju5FS/4EFs457TlFHZLg8oLk6e+YmskF/X1JXPQ
zrBzCSMaFXt65W3tm8GYsX1bW+3PBtouMP9spX4gCfhcWW1U3vjNr4X/dFFHdunEsrPZSs7DkY58
0D15NhHa4uaSFrtFvM/KnxkLx1xfIVJyd42XIR0EQDasizgWCS1kqFaZHtFhS464Ij/FCzxKFHAx
OUlx8OUk9MlEpPwFiev0kfM7ZgnvQeSPQKq3jP+Wcifz0HkLXJawRMmQ72MKPlVlyB8/zUa4NMkK
/yHdmUKdUjN8PKbUTZ49eBAZfrOSYIZTSOQo0kHIqvyLDTDViAlweUv6ddHo5piSsCMuFpqt+J5M
8rGRTx6tFlvJPzIUuC/kZE0qFwzf2BdgUnk/Q+iOxODm7VLXWrnw4aqiiy/aZxHniK8XHpWFJgq1
DCplMhbaA/shvscAFfSlJ8qL7ZKpAnPuD2CjzlaVb+NMxeFSCXvSvP8lO/N0r3evxH8mcxMj48b4
iNaBRKjzBaCymKjI9yR6Obx9IJZLc6X+DAaIxMWTmI3+z+UcdeJpjY3XffPmA5clARapI8z5CEeQ
jGXUMAPJxXqBEhpM1MKTK/t0tFFWj9V0jM0wSK9dxf+rEQfOkXKdtZeS7NqKebKS6KLVwYK28abo
n852izVId0+8kV+7meRe0CClsi4iRlD3cC52WEfSsfc174JfmBkFB2RHGlEifWJ6JkEepsIcCqPT
RAEIQotS/W7itwuC1FTz2mBJiIMNHzzhlIHgzzoDqB/vZok8oDOgkPMmjHfLF93H8Ur3kKtYt/B5
cneXtdoQdU/O24FVzAjs3O0dQWX7PT2zLq8HYMZN8UO0IAbdSyz0W4EFfzQ2zAUZkw2IAinFqN9E
mba2VPRX1fIogpfmUCBn0tt7Fd/8P/9m4AxuOZhtldrTPp2PDi5zMA6vsiUMQFYa/DwA7HxwUVRE
EIa4+7X/Dvl5YJdKl/cB42/nnJamJglwl46lG1sTtUGiZrRpuLb05cberVJpNtmLZvCSFWMSPrsd
ZCvj806IB7083Owa8anLao2w0qoHJxaFsLxAd94mOuxOiCeDq5PRPWsCyKWNrrZHDOE5tDz7/gdk
gkcRutxkbFEfHI2Uiz1EzXm7/40JHPaa5aZCh+pDoru9n7oILzpk+YfApIYgdfBUcmUY1c7ozWUv
WCGUdQFy9Cr10CpR28bGjynfiE783G53O9v/ChXzK7uJwS0ModnV17FEnijFfFtbr7764y8bXKnU
4dQIl2lq8IxcEEmZM/SOCQbMh/v33Y/NBcgfT0+vDTIshlbvw1WH1VuKfE8GHTJwPuF4h3yfU7wD
ccrV9CHysZlzFPK8PGXcaufbwslQoZAtcSucdccPyaFoPi4+L364FbJzOuMxB752wArQYVETITD9
xiQj8zTn8jlbiujsla26PP/jWiKvuPevCGiOjTBX3AyJ9MWOVzDS8+Au79fGchLY+dGOdBFd/18p
ZAfty6NoLfQgrH3tXK+3oXqZdJk4tK+c/BLtENNGWMoE2PQrlQkDENPUEy9KmWQBVYdW7h4ehb7Y
mp0rxi3CoIkog6W+alBd/3l9xmney0n3KfXb7nPfTeFpzBWPJqms53uV7An8vKvAb3MUVTFq4A39
Mw7dgHb1rYvW/oIbsP7XyUbwPmO4jQQ/7jUqTJmsnJFoKl/YdFIgrgg//Hv5/rLmocgxBdzSKXo9
049HhK4oG1CwS/KRoSZz+2fH56E8WyfgFWEJkGecKGyvr4rgRhqaBYQl6x2CnoEhvSS0V37hLTd7
FnDVJETbwC7Rmwkh7FETbCIbuyB2j+suTfuWrmOfsmI5odmeVjAY5Vu/LRYxlZACKEsMmtiKMTWY
IP8p/rADvzvNbbEzQJPDQ3gkhN4XQsb7O53hdGnPJoINHar8LHr/4BRn+drWSQs/xXlycd1haVyb
C+rYv+pv+F2kvVtR8jOJC/SBQb6AWaofH+wLyF9Kx3oh0W0xlVrL1SGFfMBQMyyc+GN/BkOcMuBj
83fqiyABY1Xajst/iCkKRczjdjmnBPJn+mAPQRaKzDLNQJK0UptaoElegWv+Y8el6V/BZ6XyM1Xc
/iw+isSgiyc5wsX4xJ/fsvqV52WlxnRfpW9/fKnM31TFesFRwU8MOpsq6PhqFqs+Z+F1gYQWDFhn
9CxBLVvpMcpKmyIJR59NkrYW/B3/7AtE1iHDTsTz5qGiCp74SfZWCw02LBNoFzbyEDEqQx5Fd9sG
+aoDm6Qk1E375LAi0QAQwX9/2JSKeqcMkTopbfYAkrbJkgfTGD38Ax2uq5TbltVRYbrRys+NYAmj
LkuD6KMFAGxyEWynPobDFlw1WmBNjcmn+mO8Trmh1oc2hVFMRMMdpJFvMoSJvgPNB3orEAguXMK6
URzEjahmwQQftOKhsJ4Y+9iKd5CuCK9knRMLT+uEaYePbxNNKRdo5JI8io8nOKNR6TlnQQ0egtXt
pWwRxoizbZaNv/oVjBewS+EhniMdEQYaD+n1UpTJ6UqZbMNFoao+9wdUV6F4iuzskPc+UrxFN0gw
LXtvOIvt1a1/Z3Itm3vcAbWB0+sUmzcxt8M4MHNdshPraVK7EEIna0TQx52d4laVp6sRtHp01J8P
+AocJkqkf2R8coB2FwRB1eaiSLacZjTbMTDJVMf38aoUV9pKspE+gewSdaZJ5vDtob7Fc9QCBFhS
tG/uZ6E1y2gmq3BCkJ+szaesdvUMbv96bXK5vaKjktTmx4kx+M0fPWRWxwKBJ9fsDtOoiG6uWSXH
nVsTQd9TjC9ZxrWbEuq0kw65JbrPu6ohVuFDD/tK9gs017cAJlAz6rTPIrHvRwK0sltaujHwKbNt
ytL4bOSYPmH9eX0ZAVno1F79DpSriVDN/nomV58iF4y51tQvXIcJth+aHi7lGoTNA9elaBFwc13/
3gBgH5FYH7s+pWun7S7+Dcc7aPfxXmsuLn9rgx3iVGm5Ofy7Wshm3jbpz7B5Z0vXv/kPvx7mYUs4
scJr3lwKnLWCBnZSJsaBzORKMzq4qKDtSwtvBxiaTJzVAWCmHSPpknNZ2BGVJwQdQ+eNOhPG4qRc
3XLEtRfI773s0oHYiOaPvrq4BEKv7M2OOIzlpU/2UaVNsKo0TtDgWDIWeQbXy/TV8xcBW8YYKFJB
884s1KJe8dkn361zrZo8/j8tngCVUtVvMuPnBIWSUfOar43rRgv0XP9+Z9bEX0ypAUITktZh69Xs
U85Cvxgf098vMiV29S2r4ayj1gd+ls0IAyQsD6vKmqTlbSR/zTVehhl+/B/SqeTktTWCPTWVJ9mQ
X7KTCPUYo0lPCTkaOpz3Klj5gYxUhA06jB6C4ZshOd5xqrieuUkOtpt7fkIqEm67qSFgA5vsPQh/
Y/JWtYIa1bjuJx8CC7TkRyVSyBXMXePPidbfV4bJUOr8niST6ZmrR5aa5NqVW6KCXs1JMPhmvVRg
dWlOhPCK2HLTXF6XE5on8Hi7Ci//pFjS+YkJ4gFQ5GNX+ZSvr8Se4vjp92qcONW/2zSb7GK15Thj
GTw6u8sXHWREMGQFjlXuZZeAOWUwbs9bQWzTM+wMNtPPMG1aX6V8o/b2ZfW4LxUx2xvPd+0dcmmC
NPrXDOeHAHWwsYuk6FFY3x6TrPeZhJ2r69gP8OvfQVgCsKcsb6kftbP6B7H7oRJfz02AziLKI33i
0/jAY2VXLEb4g0U0oX2hkBs35sp5eXOQoSTyff3n0ryvJpqVOyzQDBwOULg1tJNR6sd+0gbl1pUs
KIBM23Tk3MVQXxK9z5bIDs/CPfofJ3k/+5cCxdDmfNXIidEO3VByBygYJpr4EpxlwbWhu/8QRiEf
l3mHmqY43KaNvYCE6Nyvi6eOzy7JBNhMfzHXiI2oDUK66kVH7euvNsFHyMHTu4ni7atAKlLuDJRD
GbnJAxKJalA8r4EEnDDuxlhY3fyIQiQY3Hc/XMU5GmscOxi691HnH/uumdPqbBMYw6Xy2mNDrfHP
aZ3RSnPSiXk1d0Zb/Or/lie1XkLo+8yXQetLC+zuaDYxan9GMHMSCmIfxpYvs6z1HT84mucsLZFh
9MBNPmsH6UgTaBoWkVXd3SsFO/bMigSROI3TyZwZKjV4ry2+AcykdKhg1SRqMnk8lM3XxVl6E31G
hlFsUqcgl2KncAiUBWn2DZAI1E1RIKh6Gsy26yeVVQB04wE5uT484nie2eKJJu8Fdf6BUxBFGqKP
rfbBJahdbbNQCFqSRObc3ZM4lasnLawDMNdb8BqQpqtbaxAwo+Mre5tSpKTv8bRs/zqSxZawqkqG
bFW1reBnZPow1a/wHGmqRSi1IxMP07heR90+dkN31iOHHAU0I+A8F+HbArVTMczBpkecKdbgcHnK
0RZRVfuyZskxxPj/2a1q2tBxVLL9PNwzRMGGnwmwyvhLgXQSiXN2sR4K4E2iWF44T1ZlpQdhh0ha
tJlTV184YYXR7mIRP33qQuV/qdB2MDWs/kINDjAoculV3rBvN09Ol2FzcAzQxtI6Ul/wsQkR4BeQ
CgeHyahds5WYkReMZJKerBQJVGu9pJ7ce7+fE9jRKcbMwktf+LiWOVRp6FAqKQufe2HXRGExCpiT
TyzXgw2z0kCOqUUsdF69LC3ZyCPGhaoJbVe+liPAOg0BhzTvcFEv2attfdXFZCQcPMcnNJ/qN6+i
vLxa8rmaipzuN+USTlSXHDBX6AkmbGQust56qg1Y3B3E1YIG27Lacj7g8MEK7Lywt2QHTVskc+AT
u3V8MeXrT8aKokgdo6yjys2yU2q6NXAKiEIYcq4BaVtsJNNu2fHLxpdGU61XChnQAMc29CJqrwrQ
kJXN9gJxNyaSUGv1JErrZ5lhIMn8VinFS80quDiqm5AAhve6pIF0QzsMMBEHnB9ydmw75PC0bXY/
4dBQVFZeH8Z1uCMzAD+15n2nJ0RhhP5LXp/dmBzQed1EE+xtCOh3BrJFIFihcCVDNxrbQwkg4k8P
PLSntlL5Et4ldtxKneq1VY63BrmUAs+9yaP15zHkER41iY7fAK6UFCUZ4aeD9HCEgTJWZiFgK7xb
twtwBMXCb255nHuRIX6/Au7iKX7yeaIRSB+LYSJr+wymHPrj0sIQfZHxIypmgLJomUdMICXoD9/y
k3lQ52oMu0Y7lz2kQw4aAhRZwnZo0nxHyfoQAZCAfYJIk8ouzrAy2uqnq8sO6raGjnglw6573KUS
IK9ELTbB/5ro+GpS5XCFK2zFksYWmE7ZOxIK7Rw15rWdTmiqEXfhCYT3ZtR9uAsTdOZzabTMsyWO
6GtfshTKpwLZl8SHskB1+DldWsQ4A2UJBepy/wHt5Cn3RwyyEiS0aCCPJj32mIXKhJT8SsLQmckT
yvE6KzFl1yhCQn6ohjTgG0zpaYC/txRNlrVsn+DXaD+6Ci3N1M8VWrXXg8WFVY/GXh5vnLMT+fHP
tEH+8dlBVAYz2R1AddG39S1On/LxT4PzRBNm3JkL8zCIfG88lKOo5VFyxyU4Nmpr3oiVtwwbLf9A
DI58OpPhmBYvl8Q5v1E7S2tSwDYhKl04OkdKpUIFtcirRDYiS06as9EBa+KkcBHfVnnyCdumY7YN
D2RKvK22mNyKWYvs0EIjwRw50uWlb8HWN5yHcjFo4Yyf0Avh/I6xLT5ZUi1MSvKv8/Q7tnucOg+k
jgM6RNKvXMcsgoIpFskS8o8tf6J64xHlASjPWlT3kjw63pDRmd6NPu51bobSRuyFEuRDh3L9bguZ
DwPvt6/QXVanNRIpF0GT3NYKm7I/6BzdZzs5UrNAro5OVXR4iPgdJ8aR6q3C3SPMJlfbMTiUUg/e
wba4mms4BuQPz0m82TeFb94JdlNv24rK4XXHEHXND8qQyHMUbNgYPAss499XDoT7QvyoOeK0/+vm
WhW7WxYyMQjq+/r1XM8S8Utqj/edJIYqIpbGoUd6bhxIv23anGHUiG05bEjlHvaUutOkefn2DX2v
cm4uMtltyxE8N2WGwyTJrj9yKh83Ts3JSwEJu19MB+8NExrwkTBb2A0sVUtinFNqBpJOQLkvXVL3
4bNGbn576hx+RH3Gp9wQ5ZapzKQ25gh39Ydr/Rh6zAil2nsY+OQKOaP4tAXkz9sVd6jiMLBVWK8y
BADyciFgZY0Prr2ULpFGCEOPLbxXJ4+H0xyZ5LQ2IEB0FcZTARKlCY3gSoL4yxUaJWxB7whNgfMz
GpWQ9O3fOJ8ALdOtX4NLf0aAbLMHY5GmBhflTXqpKcDuL5KkeJuTAe0OFFVuLoubFQHhYtEqArZl
26XEnlmaUri1l2d5An//fg56Jw0BNhUcP7GgJCXx3GFcKiluBp8aqyXHfkl+Z7u0luvLdKUba9Op
x1KT7DomSuegwFMI+m05IAf9Ix3TRGOvtFPiWymzmRfvqoolGNsBT9ptCFtSoY2Djzas+zxAW2lo
DC1bROt8JSFgnkX/CvSOAQcDZoxlFFU+RMNOktl3P4k5W/tppypHWNWk78xI0aX1GO9r7BzjVdPi
HGIHp6k8aGaG535Tw0ToE+7Zts8FRT/tg4IFGbqtMA9X/xMpYWNrTRC37629PM8k6iHPxJwG6UhS
TpDTyljO7VrcGTwGK4ZvLK5EdFdA+wGLkgHHfBYStWNFpumZ5CTa8pZI8il7QeYd+p2bjtnXwueh
DnjisRLD8LNcE6BATpZl9QTj9Pg9bk9/Ts5+PbqX2c8THd4hAD6tmUyU0Z7sy9rTPwNXMJqPANkR
bpSpayt7KBInj8DWtJ9zmdLbvivOVyW8xbGkrr4oUW+5jQjUoGRMTO0W6BCP9T2oA39c8sP/4GHg
o5ZCdNysKIL2RTLOislHIJpXyxZAr2DS5n44r8V+FekWKsCfVfovmbQQgjuj+vgTwtHzDGC2m2T/
c3KhIt7Z7dDacM26CqxnctPCCSMJRvOmaiOrUZsPf672RizhtR54aLCFOT+N9/ITiF0rHpdU0HVm
/l1McQwLORjg5i2pLjkszjYQpJmSV2yXFOghQWmmNyqh50xO7RLuXKeP2N96tQrPeDEnGB992mWK
2ssonAuZKtohg0+JAS1uKvFfg+ePLv4qOXuTP6s8DWi2tMFRgImqhotdW7acXVZUXo7u6YjDW7RV
+/CasSnUXfBmkBn0OOUNJEypnZxYY8r7luKMTZ86kAlTub1H5vcaJYIinPTK1ihAsbbA8pNdFPe6
F6/Q9QzNvABlCQw+BBjaKA501NSvcRbXjJaaPTve2yz/CPBkxXvQ4o5e4+is+oFqJZcbeJmpNFLv
2Gms/TfkDKtv4hhznNSOry+k8GRapqbEo9PT1xnmlCHMTADHul8jAoknEKMUlROsWJsEYdKqqAbD
hH+BWwEIN4Da314Bxc0kzGh0xuQruZsst7sZ6i0mLhpf7kpsg2mHYZXTNPOQiKbF+Bg1jGZ3LVPO
RY+G1zDiHgJUKZD5l0LRCgrfkmgzZ+eupfAlRc3DDAUGJ7JIAPmTXsdlosl64UNH/x1/C6+21+d1
AVcgWDKkc4jFpuk4A+QlbPZomtOyiLqQ7diwiKyKbpg2jNtdUCDHvg9aFgsV5towqFbttdpFFPNA
jdoNEhSmwat/ozfmY7upXx5XWY0rpcbv2mKzKHEGrmX4Ckfo9tuw/jaXVJpqlIvrh9R1s9XX2KZz
cCvc9K/N2/NimZhOMlx2Qnm19K3rdR9IDQ798c+S8v6k/rFozkBFN9DSYTrDbtBXa2Ly80mPxKpz
OYiV+C3GlGwxYoLMz0kMfm3v6x0mkEqVhjiFRtzW/IAUw49jEbphyXVGLZfK/LLQtoo0qYzoPBym
IzBeQPPwetAsmdhrYmCwA1+QuVhAS9R+jWu1QbBcbonFfSJn9+XsZYeASRDmKlCZ3+06ZByAluWz
3ZKnOe+G3PrDQZvnvO3TvnnOZ0Jjd1KzMuNPD394kT2JFUFn9W1nmIur7EEq4ZJlujKd+bm23znm
2H7EKNqtAsAjyPOUDSvoBG8RBzt7MUp//wMm3tktQO9KoYz6n1NyZ6jSUPOK3AVHpBt2g77Z1gfu
/rUT7V0k0A8l9mySg45a+FI98ygCMBXhvxsByiZD6l2kwYIuIdBxsM5hTag89kAP/yi/bBVJV7NS
bhMhtH7MnyQh/PLED/lCIp9WCAbL4kV73oRgMWB3KrUj8DS3D0A1KPJEp956k6W6m9vf75dIkGcG
srRx36PJoI3FuICzw6fXe7OcgzoX+H5M4Z7s8tpjnunNwgUPx6MpcTGN00M0fGqzvceh5+VPmXZ0
a8GJ/W5f0EDtUzihxy5Pz6qEoY05iwPu3oA24iohBAGkjI7e9Ddf9iKhfs5qHh5x+gNM/GoQSQiZ
iuRKGNA/ZWL4F9cbICPcIG+yXHj9FXyUsyVa8fJlrkgE9RBwC5lngcjkLOX3h6iNHvSCGtbbElVH
betCmHMmgteXlQsXGnU6daQBUkNjTdxtJQIRMi2euAHOMn9kY8YdE46US2oz9NXKrA5y+asBjj4B
h52ZNxmUJEGS17U7zUBVIMYLQl4ACdtD2TTDyP6lD64dXuCbYE58NhVE9IHgujtzTA5g0xmThLcG
4ZMw8k+UwPFOyTme9PEX/bLbL3OfeyOIejQp/QyWo2M0NJ37DpaBEh+ItJL9mg6TnZ7mvCYO0L13
69A3pMJzJ/CsjuOH2mLNtj+YYq5JdRmpIBMeFeYRiVTC4Lgln3zRdbUZcrC2uy6i4TwXFSNW9vPl
v3mgchIbW1lJ3rJils7YlmjdZ3Mf7Sn2Xr3FXoMfc1nBhfe2JcRiMSBNp3MECykSnhIewcrgUy5G
XQkGEJFbgToxAtaw9VFyyrCDV33U38I2KhUbvdOl2H/uEAyDfsZkY7WBR1uDIHJkovroE5G3eDhP
551h4NzVKwKro1X5+iDGnzDzQHNXj6GEH4yVzAfvbqjTPqFakBUhdwlUuh07Kdnro21STdjomTi/
DbbSlq84+7DzWr0V7oECSU5rNYDtULoutaCYmQLnUaKMejM2cG/s1ac3f39/3Sf4B/5UU1tkSAbG
7XUe4ilgjRDxzm0HwHyWH0gElmmBK57WK4TAj9B3Ae9ik5Ljav7Bcddp7J+o3vNTn9bUeNNNRu+f
uLxyGV4H5Y4icoV0XH7t628F8MvWrndIGIYly5E+eFsU53+NH7JOkMyw5vKSnryfisWDksfVH6JB
vNNkeLtTZvVrRdEuT4+pYzieooIgcrfL3eCYUt16s7cDoI5zbLMHxUmP9sWiyznShzayayFMihDV
C/i2sx0RV4lbxaNLDZ4canGZHpIQviYdgBOJBCIfkQXRn/PlJB/bkh32XRW3zhHctTv58Y43hvpz
dtDK8D1daFeczy+RQ32nnQlQWhi9hopl+UTdEIzRayyNsehsp2dnItKLU1F/kxNgyj0plxHQYnwn
gcfu6/XVVLQEI7ppxo1+M82a+2U85B+f7PT6z7tKqU99QGiNO7d3VYaSph0Zxqi/zuxjRiSsu8cF
SSMIammI7fFyJuVnVf0gDIGd8GXoa9ayMAS/DXpQNVR1aAzaTmQzhMQOVENhjHWsBs2vecE8BImQ
UBiT/pIOuLNkpiSMDnOjtc6kMNG4pMTNObRKIzvzsd2mqZcrtk+lecTGQ1TaXU4QWGpzNO8IvjuM
sYvz+wz9uRe+OroWeSBspgqW9OybnFkRHsQ/KF6SfCA4u9hZUF8rUT3PLIpwjEp8Saxz8CIGffQ4
qOZkT7SRKoSqVOTD8OQGQRtUPJOJBZlfaCqlxU8HAiaToLVe9d1O9u9eSzp9qV7p8T/gHYmGuD7n
Vn/mFvhIaRe74MbWeR4d99VnFIOt4kjkUvdLOZHuOBqXUoN/xYeGHt9LszGFbxVI/TJRO2kGTMlp
vv5cAh1aLsq8W0L62tZGIo0TNKRYOwmEfvYJFNF3jpBhIm6u1hTiadCLN2ZP5S56Enrm5LlGRqjq
wZjgfWEUwtXpJR0NlLAYjdOUH70ufWWvF8mb5LvV5TMrBvHYiO6tw5mCV5F0mRP6dlCO7o/IFvPh
nBUpA6/+kPm9ayXBwJ84b841mNdj3rYDOXYEdjtLJp2JR99rwDIY/P9knuhQL1Zz+SV2ntDz/ZPE
StyCL0NYh1u2REHJzhh1Ju1d6xRejFomB6OBadzRidu8350neVkcJCPr72bE8z4oLTwhVrERoLcH
yV4khDr5YlHLg8ZO/t29VA33aSDTNb460Bukrn9DUQVUUoQy5wt6H4hCa+YB8Ab/dvkcFAwu66nb
5BF2MYCu58mSTQ+vBf1v+wrsAL3K/0kM618f6nEbkvJndX8DQPiIOTzlI85WiMwShYVw9SvHsdaN
ICCcAoH5Fkr2Lx3hxp1ylT2Cz4IF89YiZvh5AXAPWAOdU6B3jwV22/VDQg22yZdWrjT88y+26+0K
s4S3O9BqDPLppWBtuMTFXEG1ZbVXH0ktDIr2ARm4em7bqQI13OwYHgHiVKxp89/8r2aDq5gU35R8
qFLzxQnuOjPP3viTI7J+q186NQ2vxHbDw7Zuv0CAgSa5yL2zdD3rQivoToa0WxTh+BuRUEfRlyGO
wClb1f8BCdYlEpvgh8fQD4e4izr3f72P0WN17JhhU/nKEBqP/C48zXCILIRQV1KMkiQYxCq6Rysc
hCqAqIU/mlPOgwVaYaG95etq6tpbCfIDpiqB6pANG4pWEpCmoE89t6tmlE1x6R8NJqEhE0+ZzNFr
Gs6fXlgDWAOpNOvK/ThPiTCY5NoWXFgEOE0OIBWRrJuAe24EsJN96N+K5unjGO1dIb6FaB6ITdT8
oOOtrulN17DckNpjaIfGkglOZphLZ260jHGo3vhhJQNamMpGBxHHZMicdgPywUHx7QoS5q9WCmZW
2RI48tmDY2I4isfxV1G2vdankZHliec0oWsT/u8uviPCF2Scpz20JHpje7Gb3J0geakZCQYDylHc
dFvqJzgDJNQU8paaLU8WHiotauL/ECmp2AbIhY72NdRdIbEt4I5i050ZvKV8kxqMoS4ibKoFBHrL
AMIgTOev10NzvMrPyo2dIkxH/51GjtR5FsW5z7ayH+OsygTmxNkscYjlajWViuLByPt/K++sl9f4
PLIMEk607PtJu856MHU2qXeuZVWdTTd8LZjMNO4dHnJBY56BZNhe3hLizo6NHqf0Dp6I7J54x3k6
UZnus4udlvAAFF7/3+DvOqCkVZfDfWTbaIFg3WnHtm5ZRhWjxMUONerCGBtEwChC7oRZ2Ylqd8h8
rkHRVGxPDHe8gSe+P+9/VeUYzxMhXpxIwBWwKAWRSoEMYV11G57ldqio3MLCtG0wW7KqMtBLcqLv
KdmUWmSHoD615Opi+F5XS0uWVb4jdcP5B64tHOMBphD3jdKtP3QgHdlCuz/+JDPzJb8YRbGgmi/H
xjStIRy+BfLrKMNgoChDDVBB/u7GvPBNtEfBslVfKKdaKTDMhOUT5Wf3KYnsLa7v/Qn0f4aaQzBh
90peqCUIAEm/BNbfBYuVRh0m/ivt2++zcA15jJjNSibSzVbtQyZlZ58Dii55xiptkhlh21k9jDwk
IgXPTtB4kFSowCOno5Rc6bT/Q+WGaP1GNFMITSA5xViwGxOxj9r4TI03CN+N1G5ZKsWppKBCo1eH
WKXEQ4Tqp3//zV10KOIBgCGyf9+vYYj4QwL1BPF69jbp8BqjraV6MwfRUrgrFzV+2NpHE7EWJvh5
nivMh6Xpy8bKPQDflMOeRcpasqA5Svci4weNL4sP3KcsRGPmR/XUHOmq1U8FtUQuJ0ql3GSaH6Du
OxIXLfVvMwAQlRrKJCp4Veuh7vxbawH6pooALRvQjbXHkw+Z58jDsAxPCbRb1d5Ssg7+ZTnGE/fk
Z/wMPVMevQaQXFWIlPKFeYbWQ/XgjxTd3g5S5strb/MsaavDjzA9uhHa1k+vcTrU2uKRg8dMa9MF
9ylCfLQLOuw2u0qspOM28PiywZO7KOOWrJvFE+U3/HBD8jFnVa3ipJYzqxSQN+QaG2fNMWLeh2Tq
zVadqJEJND89tFAEVtU6lVvSkRpcvVSRc4i5I79zYl2utDJ2Rp1+pqaPssoI7nHN1XUgF2KW9DYU
S00z1UgfyVZVIos7DgCi4PcrYDk+O/eSq6/3D9P+wI2WpDSU9s4tgsXQ+RsusPl6Id3YfsoepBuE
YN8aBAEzzJIqJool9rMmzQZVhHeVG2RqKhvGTBBRwT0z985J5AGUv13qiYWef+pP9ejUE5+uQBdU
cZZW7ysLzM6E8jP1dAbcI7+LYruHSa6eifn0EyF8lAeb14DxEYiBbRyCXEh8pC/SGsJE8ZV9rPyD
KxImO6dVGD6Zpze7JmXu4vJI703Z+mIBb5HYRjaxDj9+ZAjEQ02xKO9+TRWmurcr79HUO7V5vV13
eJBBm3foXSKW1tjyuVi83r8xrbkOb+n7hmkM9QBdC020ovQkl6PGr7fGGvjEaJsMJVYuGoogIBBK
lNZK3I7c09oo4RSHRdEbbrsp1NfMRHLrXrYQoqKa/ZpWnbZpbtuZcv59iACE86vKr2KqI5oD2lBL
7nTIJGWJQgXrzhmT+fStd4lIEuPkMpqbv+APxUPl2yE6gLhkSAdxl9rr88hqftgAqlwhDozKyorE
6/L5geWuQzRjt9gUhCCyz1Gf8ypyGn1hb9+r5yC/e226A5KxZ99vv1muUYZY2INhvSpWJi/YNNBf
a6HsDCoCiNBifIjtgWsjGTJttiiBa4WykytflNMMDPz14TYb+gmghFJlBWe9INGIm97vecqwkN2y
9oHPrfnM6L53DALHRUPCXv5IhaEPzkdN7XsgFbWIqonQvqUrbX0sXdz2z5ocfy7uUZHxXQd5z/nH
uDQIz5zYiW2G8rWywb/ItkibUxjUCacT7GCV/L+bGhuWgD/UT7aKXmSZHeTDMRr8DxMTJH6HMnRl
PR/MYG/UbzgIHzr5w5cae8QO+sZ9GXjitiBugQx9ln44E6DdKGlrMShh258ASA9mc5T1w7n2whnI
j+wiTHkk7B7ABZqtGRmZcK8WQWNc/NYgtjtEbtxd57VuPExVaZ8R0xyJXVotAjjTvRpad4buFMYa
MsQB8xCFaVmSrewbDUvTrQZjtfAN5oDeM9fVBF3DgrgtrZPYx7fkfiC4Aat4wLYhw1qnETemOYSh
MpAlTeuVGFLQVBrW4JpgXhrc3nEzG+yD4Vfs3a9IOxKDOs6K1fj7KuxQCo/wuCAS77z3yLPJ3XRh
hk2ckxLTrS68upuf9uyqiXPvPxZbOt8Mha4u48BOOtFUWT+zitvIdrVPyVKNW9ESw7enNoJU4TQE
OJHExZ7rxFpmIVVuRqtvpyqcxY7egOyBqc+3lqV1etrwLqmas6r/BkJfvm/7Sgy+eTRhgURwR/1e
hm3ifXrd6xOujQ0o96YpRCkr086DJMp20SlXANSHBHFUiJWtr9He4Nv1bc2MdVJD+7pEhUdmeSc/
L16FpJpWIqXg7k9F/IMipiBLlAEnJmnzO9I1O0UbRTujbL1QwVy2ItezhkolkDP9XGxdkB74Dcds
CczTr7km2yID0myLuu8Jh3zBJyoKLOKARYzDTpgiQ9bWKArKpT0Qhs6QpIjkfcjTh2YWaH8t0tY5
c1dZsQBrDr7iNmjmJj9KK5lBOF+LrVRlJtUw3Uv7YG+hI1066c18m6N83ZuatAwYImb1z4QzuHqx
doQbkdkO0qT+QEvVOCH097NOnNu3h69CZEQIKzHyQowIPG+QBN31tKRyGyFb8OioQ3Pk/8tS80kX
YnZ4xvs/kH7HaW2rs9WL5MFzpWGiI3XUbGQyvDXoDERjtcPFzCurLoHYhQZ39uezFtv6d4Eqa297
V1OEFQt6faSNOSXMlmNLIvV9fYlqvzAiq7ombplT9JrKIko8Xv7ThdLcbL3bwwiZeE3biEc+YR7m
id/eTZJiQOpTqdu8+010oeKWzdHMUg7SddFke4gh+a9sho3ZhT+X7KWyKkhNNbhEVOATj7unlu6m
yONKw8ANscW3+ipzu9TVdUo7JUoqgRO95B8ISIMvo58ftyKPYF3zG4nyxO9QkA0C0YXq2wWEGY0b
wA6VbC2NY+tcEmq1l7AVAB7cq8yeGlhGzMAl2FFcvVlUK79SS1QQ3NdOi2IpgxcJT3dmRsG2PC4X
L9v30r6k6Q6XP/LQsgcd9T20uBEOkN4ICC9Q0KkAZzjvWswXYDQirlw0WmuAkGO5lcH+NqsqBPyN
0l4PssFi8EsJs8Adc2/ogj6W64WNi3eqn7z6Kdm8pI2jmhanh6jh15JRxbpv7r3/in1DbSMO6U/V
GA+FfKUL2mCbuw/7747/NZc5IXV3V84JJmKfr3MwzajauldS7JhleiYCwtjCxn5Xw0CkPG19rj/M
Dsg7U4u2A4BaBpgZ5BXPCWxcBNzWBA1m01wjoOSZoe/jTu2tgZUfbCo33zWnFYT22ao8MSw+5tRG
EfdkGRc5js0b4lmfdEKA2xRQB9/0uWPWSrmaGFSpmyS3iXcPm7h+Zd9FiO8NtVL9Vsnp/3LtgMr0
XpqDyRVLat0sXE59kYjkgVvLTWZ3mUZ5/wcY6omIk+GZDx2Vsg1IV9QDwsowaMv+1IJCZQyLNBs4
0Qd06M9Q9Zcdy4H0hN/PrektJ7gbP8pNP7FR/t0Rvwc3IJsXC357qwH6oZpvukTqGkdV+gbZ0d7h
ttYfFic+rY3J2bD30m5/1ZgGeBGiaoirPSuJmCk7a3iWqYe7Cwmal3/uMRpQOAYrIu8namv4pNVN
MoIJELa124stSCFtBVBne5XYXjyyk4aCNYGjJ2o10Z1XHxLVee5nUHbI7T8dXLHs2/t2aP7nnlrY
r+QzWXhsdizUWLNNEWOBxwW03uAiA8UkXhJ6fJSJrhzGS4Lr/C+a36Wf/De4fXWGfgWBaiwoJdhQ
2BVjrbWlfuwKHPcgA/6ssej92u+ZMPj4elkgrQIVzwksfmZwEpdnuFau6QaIpzmeyJr3y1dQeZwW
pZn7mPEisltLWI2kJZGEWZa+hV2y2TJ6zLTdKF3etAmcm/L7R2YhrZFyEtKPFaOyu1sGKSMl+h0+
RjVGvbgko3ZWLxHZrNq0IS5Ee1GEO2lZNUAI4L1eoPrk3EPk3ew0artPDzKAq4KRXknNQK4F1BNT
rq01MzVvW9rUa9ptoL6JR/PQAiSYbDBps1+MbDnsmysSQJXkDK+FNWEWp7pE5h9BBimdaO+HifLX
20atyHOj/Sw5oiVfNMyLyrCuAk2ES9tsTQQovCo58zjMTt46x0lFL+SUpxIaXzsEU3TMf9GbnP4n
tGlM3Ahtd6KUDWq6eHhTvwLFBDIA8GaEEq+2L864q3ow/nThB2Ny2ccVVSJYOBe4Z0MWDy7uMRkf
FpeH5OK4FvNDIuAOFPHApr67gxWnYu9ydz4cABZye5JY3Wmv/hlSrie+y/y8+axcmzh9RWTNJmnu
UB2EnnUXmjkm9DXMv6/cO2bGx61706oQMxsCJ6YOWjJ8n/XkosrLGzGhd4YrMZKgYG9SAAvajFVZ
+/Ylta22SYM9ieuQTKAwtekcDyZd/bdPlDHnlx3HQI7ekz8zcnDQsQgP5lXJk9tXeG4H4qTwBXUf
CSYXnyoQGzNw0eMQS966+dIaVWDmJr9fHOxDGqrOZb2pBJmExshc0oQOQbC1yLbhEOLXtfI3MRuS
FPxC30qdtprzy/0qUb7ZWqxevyoATZrFVM75CwTlzAMp+JlXa7Xnwo1jYep6T/dOp/ymD1J/ELjk
fno2dqmvc9Zw3EFl1L8zUvG64iNyIibHt7SLY/C3F1O5+w1yeIFu3RhtTRh8Bq1DmW5bKcYJhMtF
LFzx56vy9hppWpgmVc6jLvxrUTGtMd8A3B/p/R04tZ4WF1pHs3dtERzBBg2jrtz9WtVWhj+8gvnn
UX15rTLp5w5NZVVkYnjq48dCHHp3ddvonSP1vb+oHRxVXanqVXRDVmL1o4hdJrmOIQW2bRRx+8mg
mR+7Gq/bQo4REI/C+LD2VIjI6DZnn4dg1QVjMgJFyGgTNAzxSMDjakl3pSdQmQ4mF/Nin0g0GoDj
3dhIQIdN20zeH5Zpi1zYaTDofW4tgCHNYF0KJUbbKMpM2ubYjIYLbYKWPAJ2UBOpmRPhAMJ/W23P
RSPHgNXO02ashRQDmjDAEqNH2PPzXVSPagGc65McoSR1Xqg8DdwsyBQAz+ci7k01WknOeTCrOmKA
LWv4DdDThBQaXKSprQePtok7ZrZA4ZsozAdyK/19zthQUtWMHgVOjXKjrwakP8lbA+fYpWr7fq9n
7LXt+OPbESI28TxiqJoZLkkFjipQr9ENnvhBFLG+Zg70OsrD0cVt80WuhuBhlhabarn+O8pccVso
/FwN/c19qKWKTVd+Apc7Girr4IIob6ZeAykaka2FSf8ovepiXjNoddHVJZVtSPKpQ3L8qc+XlRoB
VqLG29H79AxFtFSOT3vBae0vypAU9PNe6UTWISHxRPINRUxxqNF8pBkfb+GtmhgaEfhvy7PF3Vjw
Uz247dqU2McWcLkfLtuSsruQgRdaaXu0vW5pOb6IdEHae1MpMTDSv4b7TZse77e3JR9puYINM27L
DrysEHFOSX18RcEpyrgdWpYPvQO2Nc42jMYoanq6ykriIuMyZmp0gI5qEQyE/Ph729rbteeF1R/4
0pL2DGz5iXMvBQV1ZRVD0NWWWpNZYEvLebMpVsMhQbJScU5FTF9GI402oRAgVsM0ZcDkmhkrq9bq
7q7k/HrEm8UGHmv4AVTmJ+OxZy2yMdHh1GO1Fsfu/APTFq2fwG7FKM/ErOHDd+/8AossF75UMGEO
TCAOOaWflN9DSER40LTIjCdBvjhZ6aq8EH15km9K+wMz27neFuUFS5vkp1jyROx62weaoDeD+abc
dGUcpclqOiWg3IfBCmhdRuRKe8xcW+1mKVCLtRkxW+25e6qMCEdDrmxyHxSqolKY+jK3gGMfUwtK
X1Uked53ZoXpTQy0G6zvDgHKrizEZqIUHclRGIiUM/m01tPgKCWbw7e+l55Su75Lnz0AP6x9LHhe
iAcysl3QpXG+1QyT5KDC1BrJbIKfHXVGhmLCcp/kitaqK++kADQ3cnfOnf65/PBFj7c0dSlwz1U6
o9wPTQ1SRHLt1Xliqwg8NGRAy5I+x4BPCk8q6BbFfHdNVqcv/uj5p5MK2xuDCC9BYCga+W8XijAK
9nNyVobOUpFT2pUtP0Jp9k4gwXDTI5Ru6sKMQ9u8a6MrermDyyXKfgjL3KfYl3IfojqJW5GeJ7WW
xtuwW5qnUZYJHLLlIyFxRdS+NABdx1nMo31WgQR40UZYYHewUUbK0tkqjImDmQda3Xc+ZMxaOmKM
ucacKLHi95K9VUAHc+WkrwakfHtzbqn/PFwVsj6WJMFDKqvEW4Mmz9hYVUa2iqzMqQj1HQL9DAX4
mllgqRZ7JTU0PzM0beOXxsShNUcKzjzHY1TqobnLa9isEN7y4bEMDHzbtCQ/Rw2Y3PQMgiWq8x0T
J42OFPOOXGOBV38h531vrJoWgeIpkIkIbYJbiK+6L1ZlogUWMprH/WvabKBMWvgS55pPzmo/qF8j
tiUaaN5jZJ3X6yEpxBVV2Ja2dumW+IoEnlDnW/fIPIwSNhmWsmy/Gfrvsgq6PLaT/SgKYiywYw9T
lvuVpsTMtd0V7xLzY97ABGteCAoZj/Hd9qLKGFtSRD+qrT4xVYHActDaW+i7yCaN6bgCIk3FmDL+
ajkebX/QXRRWFNrUAcJvw5a+I0Uz2Ru3SUAsYZgyHyOLfRHJ0vKTeRx9NI8pEuiiZ0uSuKfbsar+
TrgZhjVS6Bu1CCB5qG2Ys0x7JtitNrZOHFCy3Kiw91TZRSZ/MVm1l13KRSPNqxJaXVXR12bIVHg1
ac8j1Ejm7nSkRVG8T69gAjUXiW1h/HZzMOhIWQ3vCmBrx6gKOzRlAm7dfIygDfP8DyZ2h8+Ay4hM
zLH8/tml05jZrz7K0meWRstuApxsAm9j2ff8mWI5UE2vQabMW2IUG4PuLpGhRy30uUcIfJzwhtp4
p4+kAg5fdXneHQAEUjm3ShKEDJok5YUESnUhNNIAB3Kuo14gCc/Dqy7fi1ya3Z+7NAmoafOOv1vl
BSEIclLndyIjZsSAQSka0khYqfdPDZxavvjw8exYs4kDZrydr6maynMUIm+Vmvg4qjlT1fJkQCPF
dQr8UD3ESKd+X29pD1o2o7jetK16CUa234O4BHANy7/mZ/6saZz/3XxF5RP09NuGK7SmlxXoO7x0
06TynEBE499R8+H76YsmyiUw/knmK2tZZzf3tg2Un9Kp484Oj27PVDLOZZjF4n3TneIg2fZXwO01
vUZJjff+F4cqP5Ygj7Xet19DcBi+KRlDx2/996Y1dScQ/O2RKU2BOrPvVGM1Iar7I5SvpzetFhwq
9BAiYeBSiv6Ut6CwshjAUmX0cxpA5wAmNOplwnwZe6cGDXswLQ9yiD6O2Y1dTVFfNLZM49EN61/g
XtEuqUxnpe45KtKm4Ln2A6cVUvbiQ02DUVM0A38xcc2yQ6+Qzah0zo+INccdWANqR4flzOM6NTKd
KgOFeojgkgkNib3/q9TiXZ6TCG5DI+JE08lJgavRem+GEZQGbpfZJkrLi4uh97YC/E7Ejr5oQBBw
QlXd2ekLgyGQA9tj8nmj8vfU2R9wBc0nN/TI/7uULRvUWKkl84XjFACk9qeaRAcKl0Qot22AghJj
gORnh4FZzBwsBz5t+i5/X3DuThqTFUEJog7fMI+7nwPb/04/ahXQfX5axMzyYTQulC1Y9xEWoi5d
96x2/7QjuzO0bbzvIhecS4TMp2RxcZfRSl+5M3XuDnuQ8dQHF6AXshg/4F7Jbr8rXHY8toIumAwy
uj3EzTSbRZRsigyP0UbjQR1TBRyfr1yWyNBjzSqtkswg/tBKW+KZ9FQFcoX/dO4vUzn9PmVb5WCT
D/PAJ7NRnVetLJNYFf1LGt0L5Dp6WUp42/KkhiQfedMSp5O+M49NPEAf8CDvXpWIxhbuTCBmKTAg
sSkehahvVBDi5ZgEaO3LcSOvJZaUooaGDawjoS8522Qy2mpilqTkRb1192vyilO9/ipmnfrUvgKj
OcgL2RVzVI2FqZGxNsOWFj9hnK2TO7zH6xIZ7uyN0TkOvf1hjURwNW4ZKqEm2L0MP7oF4Y/2mlNG
oR9yWE+pU2n8gp7k4AFgp7ykwcFv4a0I+M6vrxFaNz8uglf/486uhZGaityzHwVtzB5A4bpUWjSY
KRMOLCC3qfp1FHER3tzRPOYiBINkiJU+dCm1uDHjIMJbj6+mLKbnNUXIAO3cMYkDu7gD3kpn0oQ8
CeGv6WvfLCGN5eeKNOpo2Kuf6Zllr4Z/5il7YC51JT3j7uXHCMgDVvUcGP3uq0CVBDH6tnb7DZo/
VUZH7bTJg3qa46kRtMgWzsVleGTqv/4Hr7alVMWULgw8IUYcYYLD4if4QbtEwK9OOWKVVsVLpGj8
eWd0Bf+7LzGVxwP++Ymtg96AgAzdSmXcQZlu9mvhjK0tHYeJiLUpqxfBN1SK1GByC+cJc9dat4Ph
fQfdiUCy4GXhR3ll0rCtBT8f/yFUc17OggnwfXDprUoix4t5Ra13kiewR2TUPiw3qRxhvhDmKkNh
rY3VlnMtVa8xK/+N8yB1JwMKEy6eHRvKzB0WF+qMbr7/ggU/BeBX1x5ozFLQfekOxCeWjDc8mWjQ
Nsi8KzyGzmgrzFWoiA4RImrl1jPXCZ2motKlc4hBfG37AzMWpM/whkwkca2BLcf6jD/8JEqLsMkK
ehsK8y6nmPjWeXxm/o6cW8Bl6mIrz6mcZoDLz1SS+5SrwfE/jFo7vR0oWxA12Uuh4EypVUOQXTdX
iwustd8HlXinD/5/KF13NPnkb1XgJyrcPI1uCXCoFwnhjX7hEWrakvM2/wNjUTf/ZQuIKPL5WJpI
0azerlEj5XGrXg9Fy5pfJJjMpd0rvL26qWqx1Sg6M4D+D4y7BVOUrnqGOov/yvKuL9Eu7Ct/+qps
/hPjwVjr3yfTcjqVeBmU9WNiOArl1Lw2QCYwadcdaZ2d2ZzUv1sbDRBGuUapxF05TWqLMJ6oumNp
E9wUgtihtDa90S1P9JXLjzTGfi8rzUe7AjthAZgEKYyE/iocFu2NeHyaeiz8hXrSVmcfoSNWB4zD
dDk3jrydfyE723OZJ8DS6BKClS9z/tdwd9jqOSeGUFnikraqNcetxZSFneEhw9gzSsNmGt+HEtwD
eJM1B578KS2TP5v6Qw6/CdxX6L0btUo1/tLg7/STVakGI3mzaPKZy1g+mSX2IvF2d00+PUVBf6fz
Mz1LUK4yuKKxyr4oQrLBqTROEblagw6Kez9qa/N6anHbwizEg+IjA7qMN03gjMTHscH84HIsSbuC
e7A/k4k+X2Nunv0JSXkEyL9kKBL2OTrmZFrmiEZFNGHHptWQL34AV6+TbKNLBT0iTy+OLh2JapdC
cuWfODCJndOxA0l5KLpwk1Dcb8Zs+jXg+cb1iU8w1CZPfvXcZolrHX/9TmRARxjXFaDm3eTBmnXp
V4zoXl+stS29Wb8Um9yLejsISJbeV+1j9BfxfQoFZ/kqGk+a3WIFkQ53h+hxSef8l93+tlou6yg8
FQ5ScZm3i5PNl0hG9YbbZwa8JCJNvt5uo6WQaU24buSB7tO2RXxq0FtFZPb2Jz7uG//vAUZ1awpo
j6QVc5qjQoKYv1+YCCfgp711g+pWh6yKMJBSO+Z+iXGbYxqFhEO+O29wEcTPGuHcc51CF6AoJuqO
sM5yPcvF6wi/TdV2NlAuiXHgrpABNPGGiuSfbZmbf/TFSOCfgfzgGWSsIsXRBkI8T/4qDLn9sPkp
FPHMb4EmxtPsaETUgApBN/L8qh0D6rgnwDnHN4IY7tFc2yQB1bIn/Gxby8EyYrv6l0hYcYBcQeY+
bbiEhEG1sx6Q12RyCYgAGFHBr4UCP9bFayGgMuBdcvX1fLU3FSUOcdRdoYPESjp22qd0GTs/HOtk
6jBnB4B4tqDFpaugiZL5QNmfybW3sdVTL78ze9fpY7xo1iu6jRZEus7zaxCzfeMIvX9csf3GJK9/
usbn0L6lJlGy/cOAhgWLCuRquXicfTot5ZMB2a/5Q6CbV4iNTUar92WwgdDs704Xek4KERearQuS
fCTs2N+NpOODit5tgz6/LA/KU0KoOS2mSG8SXlxz0dZFddp/yX2+H641CmUR8jmqQPbcY2Otz3XH
CD8sVC5S6xhHkW1I8xXajern5TqbnAVecY+0oc+I9CPdGamSCmYVCKwC45ZEJVd7ly0BcghX2C75
OzDJHFoe4gcmLMQzcIERcgzZIAni7fm7RMoPzvTT1Mgt+fgZ7CanLo1i9sl+l5sEaA6WRr3M2A4+
Jax42nKa2l+94ZpEovqsAGgCZt18+YDWT0brVRP7iV8f+MBOdefPuxLckNiVqC8yTmmrUxoHxYhR
2q4hnMGgtm27Dbx8L2V4JDsWg3G60lPXvh9ZRj9L5iZAiLYM/o8lFWIhwGTfZWnIH2Zy4mRt98cD
/XpYfa5fbbhmyjboVeR0nMe9R6FXCjkUNQgM8p7blBuWs2NHsx8gDvNafHnoY03NKs/Y7Wlf+sfj
z6tLuVIgzpSeegF52YkaMUVfM9Bm7rw9sJ4dtAsGO7XQs2BDQbMz51xsdirVD65VOuIGVZBdL3ZN
st3WuAX3XuJaAW5apvMMkgDiVxZB0jV1NoEjIrLeT516eywg/wXz0rzistvZ5eAebrL88sSOvvyY
XJAQf5xyT0pVqg9HC6JGFj0FWxgpOjcS1V8HUbYu58F7lSaM3luS5QhdZ6IN0V7MQitkCRfIyb5l
7mRN2G1HlypVsAKJx9G/2oEjsWiKsknpkTe40kgriQ4dxkPY1SjVT6EW+hQp3SNVu78JYp4G5l4v
Z5lyvZWfAGKkiw6PgOTZ8tOUtoatzovrGoEaDhBxzvgx/l1WP4iaMi1TFx7INpFsQBDQk3qzGF6T
beSVp9caSAt1lFEZ7S2f19NuPzijmq1Jh2izwJyYxrL+GVynbsut5VhPjpqXi9yiI6aRMkM4dK74
bCk6TvAbgsjQQiV30H84FaqaiF7rkO3L0YLEt5u/Q4sX/9NhPUuvwoiFsBY4xWv0Vxw3vvRWGFlu
jIHhCV0AR3jA60CsJd0UQzCgPthiwIqArzq7YydL2Tr7BwDyDwuUZxpShJ/yTPtmAWUFsOepSEbB
ICsIkzISgZqSyyThdC+i9GhtJVIcd6MKtH5ywDv63YViV0HhpYiA6OUgotWxWkrVYAdwJGaO6X+C
9BHzPzjFl9kqO+ksTEF34bnOJ027QB0UpIARg2JndWUXL20pz/krXEaOqP+vW4Es3VApxpEsnCFE
6ANETRRK8eRUjQmVsoKdBFRqc95r89oWAr2iC3soRhMfDBK4fsqItJnQhBpqd2NUAEOJRu1zLQ24
AHxrSJmVGEO8qTOb5Nao0kkz2i6zzvC3UzeplOAOZ8th8aCmJKHoV+FvuMWMKDhUnZgB8S9K0Xpf
K04wfSFF2IYkbOzrc3Ml30TVsebNZTefT6vEanCph/dirK6hc2XZom57AeRt/qf3R5fVhOCE3mZ4
JBaTaDdINVhjWrO27HqAsGhQ+ZQ45D3+gqr6XST/FfwUH/J22vE9exRmKUs+qcNGErMo5FUGvB/5
vWDXJUJohbbtNei2iz9lWCmhTp2XdEd1r2sD3WsYBqXBlj1t670yN6jYWaRSnlIdlcIQB77bzdgo
RSerz6a0eDrNn6gAygExON/USPi6MjodmsEEzi1tnK4FMz82AgrzfhfzXjNyxGHgU4PjCbKl2Tpc
psuYL8vfXvtvd8VIvX6kwIhbVWZ3TNk0EbZPdk/NOSWgOpbIiKCdIT4yYeGyYidWw0T3h4R46TA6
CbAy1rPBOp2Kppq5BqKffJQSeo0uWcz1yF7ngEyZLCuTzr64CjLiNIJTVXryR0LtPSpBhhSPyWrI
h8ILLtd3C6yzRTzuVyoDsJh1ptpB3f7nV1dXZHIRbxC0uZbpAl6TRWCv2pGA5fX0OstBqMzGgdgS
QRcgEriuALg2THfSmWu2t/hZl4juoNYgjq7zSXyP0QuCpPv/endG+VtNcdkvz3O6odm+Ur6R/51U
O4QpCVqyN/Yumt+d+dq9eFj5YccG/kIGuNlOgkoMf9GdnKyU3+gfTbgVZP8XQmSCeoukiIpCabWY
B8PqJ6zczp0RJ6Kv30I91EFDLn0/DNBhMkBdQ/YUEeZLODgPKtKSU7r4U37gNMLsrRgG9BN1VQtc
OdBZIS3LYWPkW9MdKJmz2nVKdTVpuQ+ANq73IiFtD9fOTYsCzQO+sNbhxaaSD6yUt8FTAkCtCbii
sIMa3HbJy3wJ+RiApQUvzTiDgQYMu6yak+T00NpEPTBAike+ROxWnTnRAq5Afqy+yXnhLptCgrN9
wNjCOnt/FxEblDVc626Q9qBwmRH/Rwybw1husyp0lKyXiNNd2rOJOaVhlSGd0/0PX2Ewf9mDorC3
dNxlsjtLl8pI2GakzkK5aeFuja+fR1/XOr7vRFhhXJ/gK+c4F8juTAk5ieC0Mos8yAwK8JOr0y4T
CTapx7KU5IYrQx2kujkJmQ/jplqSIRh8TsdHmhe/aMiMUIT0BhkUKkIrZPVfNN8Hor80oC7RYSlF
3Z5Jb0WJsdSDhbtOyj1gn2kN3XDkwMyL37p3PyY872+VB3VPoThlNggsk4OT0TQKRqUMsqNBvwGK
zkH2W7fltNvI5d1byWah6erYkP4ZpZocpg0uwHyU5wkwKrAXLkzBiqEcBYrkHGyKcAyvkaVw+skU
+EOpcKG5ehbZB8iW2EDtVW8qYB6AtO/z/W8a0+k3I2zey9REpcVzXdvTU7tNzhJ/33q/bgTnJ5TN
Nerjd9Ucxxd6ZHLBp39VdtPtPSitzEQCl+yAz+rymKUDbkRKHJeKGOYlGYxHYbYKwyfwWurueCLH
WoiXnT6L2LDqVJllMaAIw0Y9VNaLNWYi9tEFOiw8FJgSLutAhRJwYSFv/FuK+4PoVxRufsisd2aj
YehSQaB6OBnOL7NoQ5i/KeDsZ5rWa/RVesSy7fWoHGn/5CzPM2w+FMycn/Ur4158jaqjEfND2o2c
F5v4AsXtPZ+JX59XZVzM5rqDedvYPVewHNUiRKYEwwOsJqHBXKvzaj9zC2I2txAM9J7CYnLE9jky
zGILPzGQizPSLv+LaqWVHvArhrZrIbMJ4kQYXeVX20Vq2M/OVIta7wCfECapB73PiaoGY0KJS8az
WdzBW0AGlTLh/gUJZHp4/VWT2/jCz2XXnNs/NvhqxWnpFJ6N7Ev4P5TMjZFX+rQGoReViCur2NGy
brjLXrd59VAKtYRyV4Gb05XBDrx/MWhqMjaUU2Cvz+cwOTblU7e5k4hh6BwIBErHmkGMJySOWDw6
FSdfQqFpODb9L62brKsmiN54h5+b/e1gQYBC9/e5zVPTDMrF5z47QMbBLjdG6KrqoRL0B12nJ6k3
wr/SmxwpbP0a3FSz+6FBW9osa6de6kwNdHMGLlTi7fbP01gRdMV62Ke5IlkCMfhWda/VeycGkcow
hq2S30jdkIVSTVQZocJJlx09q8kCK9qQDvYiaxwKhRB8ek2niTzmWrsHhKsQjAEu5YOYVP0X6Xsw
HwZV9SZWsNDKc1tifvGhUjNxGC4X8k9qMCr8PoWtFy8abl/NpjhJ1TDm+wUcSIOWFRUtGfZMMFFg
e4gd3slqXjkech4RF/SkrR01PGcOFN58i9TU4fftQequtFHC0IVFfCAQaUz/IARaQXHH1LKIEr9M
QtxqZjSmgeJMaUeCaKJVCjESPfI5x1ttD5tdYy4VwLPN1ORRhgQEiFkM16kb6/Ukjm7Fm/CJA42l
wIUcvtEM30A2Lmw5lq0f7GvUczujF1uEKBCeb5Jx8jGoyqw4UNjSVJyhwHMj4M+Of5iVfwjQdp5X
fbHf0ckh3xiTCsUoD/FWXxAW1eq77BAUjhaaD6QkvvLMYTB6Yv1+G8qPiJvjYkeqR28Vhy82e6nb
vQ8dtYTMSFmOI9i/27hvLjO+SUToMNwhSYmR2oMKGjkq0wzNP7DKsvmO345umFGeCGRhAnez7+D7
pduAXDa6IaMdQwWJDCvAU+DO0f4k8f9tBhQZh5K6sdqGUfhFPETE+XLFPnAwFDFuaWHTCsHF4iBJ
1KIw9xi83XiGoVUKu6saOteVqZHFxjcxHKwHGUGcXlv4ha1ZdTOK9teUzHeQQIDaELykBiU0vcs+
HOFWRmFxuYO5zsiHUPAczS/2gWM/2j2akLt+OcW2BIWrhT3rUBZ6wWIywd/t0SyWxm8Vj2Fu+94h
/IhMg/V2qL/vZ6H7/SVOOmVNH9LdemS4so/BVg6itXhA3Cxs7yoDpbd2wK/pROClEzD98N2GZYUJ
4sVu/JjuNFnVWkcp/xdoyPBchhtwiTk9zrC/3eufzJaWsAnmUJkHfnd0CveHhwbIVlgwRrTvLzkj
mvYC0kN19pBXQk4sgJE2hbskIlw2bcwWcbwLrVJUawilFE4hbBQhBf5PA27m8RfiQlnAzBukdF+V
X8IXYjGBgtkjmQiy8BDbCTBGMBMsjAjbBaokgKi3N0Ql15Y5wHHAkrv7+fh+k8eiAPLAgblgUfe7
ldzwjk7Xa5SzL6XSvGbK7WbbQlZ0xiVDN6+MwfZSOV7tuZeyy+qr3s1XaGydSUVJ0JThctjm9RNn
wywBSYU/eHiZUj/mQU2rnj8lMpgR314VwyA3BioJte5SZmaLEDYC6kuQLTFOCvw5iInAZR9V+QqK
huJfeNS2Cu+7iHvDVeho3RNffi3sUKURrAb5XNoDDFrlHeAix0PDal1/RpFvUEUqa0AKaYGt15Vc
qDFdfENZZQcuylLC/F0ThyEgiwih+Wdv19ja9kEnyqD2JCndCAI989VUkuItxcClNeSYLpIekw53
1Um7Y+xYVN/AgxaKvHAh0ZPFG5mscEK/OLXMMRA5aDEgREbsrlOGhLHuMVqJS8wH3jwP+IukFA61
u10dHWy9RVjk5SVeof9ngIffnsqOXaXPg/blDSN+6Gx6yu2H4vxDciNTpOl+y8tggUxjXh6LZPYb
EjXg/k1N9l7T3lbkq/x+bRMkXpDDgly56k6HjgPSjkXQlxs+QpIlezftH27XWSBbxzVBv1diQxAB
KyO+csSs848wHoaqWDBTWUaX3/In+Hpq/ru5//mCBWQ2dSA/V7FwiFmpMNhd9tpUpfkrcQ0bg07F
LqODwzpDpDPKR8GXIKDSX1wW5ItX+jVgi4wFZnsbQNN2P3njXTEXGBbu9p9UhWiQX45iIio54gIa
ly/avb7fyAo54FNkLXTMVbKKgUL8msBIArndEnXbFA9BL2ETWsi+2O4J60/hzZHwOZBuExUz921z
4UcfQ2UABFgkfFwPQN2xgPK+v/FVpqkq2E04FTjsiJQGr55zM/Nk4Rft51kN7yKDUjSWAhVzQdln
//xKKWw3J4j99aJAtZXmi0xxn8FE0PiIBSAu+WE7GI2mtO/Xyekb0tXl+W7evO6oD39LxFSbSoaf
WkDG9f4vT38uILYNvPYXYowl+t7v58bd6om1fgtaNqgz1W/tPFrNMouYfr1hD/0PiFQTSV2IHA2z
hF5pQxRIvEoClhYDzjFWgE9IY4xl8mKaA/NROrSPtLOnyG/qDqzdiPRhxEqxKL9yOdX5KNQ2gR6q
eyoVBVwVdkPRUdd92rAbsws39kgdcL40/6oFp6/dmFARCT5pk0r7HNpiB7Qj0hjnRCPKZBXfoA0K
Nqs91vECeVnn9cHAY05/SBG2N+ouEWfero5sPw1qjE8ipV5pdvFhDIA84aXQC/GboWF+JcvnP9Ej
QDWZ5ZP7lr47TjRtmjIQBSULnVxizQ107LsrI6LYtoZe4F21xc5iPLtoBUwYb7JATcIRwqIIbaEq
MK9tN8lhQ/8V2d0nHsw9xBgcwl7SbHrqhsn7K2yXhCopN5ADW3zA/iI2j2D8SNM8/SPwi7CNcvbU
y+b4mgq7aYcjHvv8rkYMJBEVuLr3IyeMhcy+XOby1SBf2x0pX56W3IObrUzIfu2pB74u50ZIZ9mb
0C+etfRjCUB4umCVtE4M9wzYDmSXDhg6jVHn9J85qmCxVneKMDbh8uD+UGbaIAOP3Gb2do21XV/b
5ngClx5oavAzV2nr1TlnkPfa6lF8zKptkasa6QvGC2GSc3KlOLM2+GuewVihUelkftIW/mpb2VNm
q4KOoIWBAGmnZSm0ozu9kx3kMZHKJwQHHEmDsI9wim6wz1Oi+1CoAXXqFEBFLWK5kofVGn2EhWf6
CQSLFaZv/sAj2eOaKhra1WybvZwqIrggRbvfKD4RVCetCEFLx5zTmZMj3KM2Jb7tL6LM1YzEHqax
y8w/Ru3ARk2Fv52hnwtmamFleV7bJNnAxSHRnGUmuQKhjlKdewSGxoykpNpH9S4aCbADsNbBAQ0G
ZNrZSSt202g7WIoYSKZL2iRQlEInz0ToK5qpoyNjynIKhgz2aJFOdPDRhH1jjDniKAGWsIVLzfl3
5G9Af+IToeU+yr6m8o/8c9o84Uc4UQaBIWzXgdqsRAgdXeBHvhL7QB6WdMTwXfDvgnFVCNFYuntZ
AqlRicmD72VN9PN39tAeC3z6GPKTM7IFtfWVNsyattRF4c8ozUmQjgqPziWlj77uKTZ9ioAJtiCM
/43r5xd9AAQXq6qwstNB7ttlJAakrOk4B5dSWy/fYucV42RZise1tP0HaAXs1HgffobHtd+Gf2fS
DxfOonhOXFN7FeB1ViWWCsG0QZYKO1NqIctmMEOxd/9Loaz72aY5YMZTtQmMQDkUrv/ZHzDRLKuS
RNzTC9rZCzqQDsrxzweL9D0N8BQ/1GxqEUj/9NDbOrBRBTrKSgkVIa9ClKvObAgDvyhsBtjZ8YAF
qr0751WQ8TxEFtmbWFRxN9X8iCNoMJLAyctApuI05II1X2uk8LqAqbbin/JAkZrx+DK0hN6rnFQY
Qm1ymEt6J6SsMczdxgvX4JjaM8foorl/Xum+lJ7LCn7tVpVcJulJZZYA7ztFaj9zdLtH9TsPFEc0
ygWjnZDevzWSigHx1o6tXxdlZybWmzw9bIMmLZQl2PmVnLuofwn2DbwYwhZQjNDbQq6cvTFV0p9o
iSqudaWl5ZnfTmVsZ67yr18fvG//tESd0p+eyMRTsasC0/GNGBmR4f8IH6tnAUWLmt73aKzuytqA
K04Dy9TURGZQTdTNK2/NXz+loPOL4k9SJhlb18gT5S1n3ftS68bGB/hfLJqKg+36fpqIOpXuSIPj
GD0bifO2pxByBC5QRgBtAtLlKoOIUdkVlNY9T44+ukghGY+pahGtqF5Mdd1wTL+cexlQ195enreq
xjeXXaFRV7suZAKW1CCsH9v7r4Z/qF7PiENuvmqLh/Yo8Ig42Ah9tJlqadFTwBoCOOm0oOpjmXbG
+SoOUKbRVbe4Crge1yPk0HAwACwZUGQQc/ylOUwvSEuCKjVwn0JpIAwLT/dgVmkdzYA+pX8R9oF8
4jL8JevOlp1sPEyikFSppXZVkf4boeZ+e0u07OYgdV77GkUGti1h9MX2rvXm2Ud4HxpB6CnBzoxq
Jcz8qXhGOl4+j7erNr2asaoa3wAJAOwK6Ac2l19hXR7dQSnamV/I/dxwawOoijrAp1b6Fvr3hcSy
1e4ls26/nGmlTmDQm5zsI4oGTeSjNKfuGVFpJ3wj8tcIJyquTtn2kdagD4m3JQW59opKQ9GGVdw9
E8ebO3zGr/rH3TQvA/6bulc77zgxS4P1pE+XZB5eywM3XK0vxrfDizMgIlDXg65JwPpQzHDL7/2v
KTKVybc7J6VWjX3oGLU22AMJQ9zacs3HeYNM3kNaVKoUeX/XpS3wrPPvqQyUSKympgGoOboMgZqO
trOvT5eBC2kGVFxL+luoSx9+WySghTqi1z1jcmQGm7zbLcGqK8n1e4cKMCYrbGQ+VLqO40/HBXCB
8Csaip5wO4MSC9cro57zPP/6Re/+tP7dKOgxHt/wkav/FYkRzX0qca0bRZv1p1aPpuW0O6V2SLAh
6XCqdPRn3m5UJxenvzkiTrPKnzqOD5DNtQDtLInMwvEtPisFf6sbVOT0RzL2tYvsJrxDSz0lAB0G
Yt9H8USxAS4aZIbfc1QL3Q6Fo7C02ZV2ve4dW6WuA7l3n+LyUZ0IuHZLY/72QxWIF52pGssYh2UL
llABXtqS9BVEpUzGBVanMn8kLeoGgwYqUzdx56idswhYLWUPzBL1kBmDbfup6S5IVc2kcHVga2PY
6vkRGQMAXtJAdnMYWQy6XGmveoTpiG+/d5/H4nT5WQtg1Ip/xGZMdgBaVsXeR6MdNnOmfd1IOv5s
1yUBCG/FAiWhnJMTW6a1Y+xIH49LdevKkrHchjOd2gsjki1DMICygRts2GylJuMeYr4W7X3YdZbP
iBV2tIMIogVDHS+k5oQ3CfKN9oTDAYKv0yu2dNo+ei8aSIkCeLv4mbfaR1jdtGTjDWYb1dxY9cpx
F47KGC7GoovjzFFzDMU5UKkfUjmiq0tFSKtcayRDyz6ScIzUxjwjA47/Ur3EipRXBTF/nOzwBtni
9D5iTNEEX47iXv40a3BVpkxkMwM9FrEL/lgJEryOl/7EJSiTyDvXoiVR8FxhxPXkhQ1bi3fCS8Dv
lEdhTRQqM1SzKhboTwI2C3rHVJ0cNZ092SBvf7OKH6XKCMftTCBEnnPDaOGeWgUf3CQITfpAhznU
b+LTJbIc684bvi/mDPxjO1gCm8ABQTCQtPfBFgEnxyVtioYWDLKLeNSyrqzT5AXoDvCzOx5LaAgm
qTGEDkcdsdX/7D6fY7VIkk7PRjU9NeK6sd5xUHafpdoQykr7hQI105JcMzGK1Wf75Unkt/lNlzki
Q4vAZyNPEW7Xt0jVUtK74iailOWwkmYRAIGXXKzkzZ+LvOVB1vXeaMNlWZ5V3qV/qi6VHphfvpOg
PZxR8IaE1JTrRmcgvxGV3rjB2itVQcC4FIQLQTSDh7C75x7zXdpvT+hA8wK7eyd3on+VT6V6ykb0
kzzoYiEaPoCtlZQZOoufwOuzsa0T21O07sR3GivjL4NhIBV+maW4lwP9pUITKOU/Mn86sXa/CNNS
fxEHicsCc/dYhlrW1Gf8HXxnZsfHPBra1Svyj9KN1RaY6Do1OJqmwgKmXfENriY8K7LFyH0Nj7mD
F31i3nqGwRiIijOIxm02qvy/1nmQCCoyhJtSxhWOCsXi1tR9yrp1QaktZCHE7YtG0Xexm/CIroG/
Zytq1PzEsK6dJnGACsWYdwfUDTU7wWTQmkrRqTogwuKmJVIM4mRO3IsmcbZzMBMIMhx2ZEMWE2DZ
8tJ/idr5Fo16bs+WcHgxq4f0DWMbH31qN397Tf8DIv2mEY44kuUi6tY7eE+lP/QLFFRRbLTCFb+Z
VbohcntB/FOHO7Ji1MFQDR6YSAos1NzEswWPlXVNNHlw8oruU6i5lcpiiJybjB+4xDu/CqVFduCd
2gMPtI98O0emyYS2fEc5UYNR4dfLjJA6/sVrzIs9q1tIRT0f9Ko2iPiXZV9Z70Ca8n3kYPzVcOU5
8qzPSb/xbxHmrZOgvLUP3FEgVdcJYulyf8bilSpCdBIAoqfQfoVn3+RbsALiEe+bPuVxTnHXsP5j
w5KCDTS93qNOeKiZKZvQ5ybGTZzBqYuv3mjRnS7+gw3Hth3n7SLmhQIL852/EqHKK65o5M9dOLa7
4zZVz7a+BMAuS1cxIzDrFmwWTqTWN41W92QjL39xpMiPjWPoQo8cCwWPEfNXJvXxXXDbQuJBUJlO
yfiTrrc788Oga4PCMtaDVTHqz7lk7QZeaL+H95Mkw5kuaVLdBT545m7ecBA9zuCL3H1ZHscL8Kvi
LYzXTh4p/Oy1ghhs/ReDjBThEbUhcPmhQXcznXhaSqCxGqZQWogjjyfI0pKU27jXFgca3tUEYXP9
Kj7jrX8w8poyyaFcrqBOYyKMrHkR0SJDH6DtxtmDH+Df2NFGQPhSBZieu/hCF/IxKtu3l7l/n23j
dO+yWTbU6XsEGWwhtpA6PQOX9CG6G5XTzryKh6OILoeBoEgYZuiy6v4gJAfqcJMezwY23VwcTABC
aUlFlWn0iL0E052UQDcX8Yq5y4z9o6YaNEMmsh5tn1vVRovmJTMwbzhqkHDXkyucG3QLvysqZmZN
NF6dLyfuDHPDEXXbbupTPMv9vD4+gNSc/u2Z1oQ4QxKawWUS5uog7PaQZd8+5mHY8fI39Mi9cRg1
9iFm2UhyOoFRF6KXYsiYq9fX/TF/LazmM9nklV9ZwU/IWaXStxZzpuYMU4ZBV4M5np+F+0XwYhxW
JFHKr/KAn9Phvvygy3+aWNmxiFk3fGX1TE6fgoS9tTwwP7DiRbPc7jeo3mf2NV+9U7gi1HY4EyZm
SoMQWoImp9hC8RCzNJ+xgWW83t9FFk1Z7Q3Q6MIxom5WSEXvOJFqAFHBwE316dZwpoAIbRIbT50C
ovdzbOHTJ86PzN9WQjYg5UV+73JEmmPlzMEHhatmQrtxskY5X51Deg6cqetjC+95cZ4IqVPMXWHa
iKV5wEz0/pLRyiaHfyE8IJm8DPLTFZJDJ1GbAiFdNZSqH8QhVwaJ8q4S157yCF7S5yfYVU0aTO4c
qhig6IuQPYnM2M6+hOwcdlHfrxop9uiOcVcLEqRMibPiFOy2qbzX295odIQRSvJYEgxOKiR0ORW+
5lWtvIUr9Y/updbYwykq0SBuoAKyAdY3qHHXXDoYPCjU0/HFXuOvGmaAWa0FV5jC25HdbmTMFyci
UFMi49imigScED2cQeO2HvQAYRIhkDJbuH01wHgg6FRijU1P+8ZrcwHG+GLYFyAGpfOstPtKm2Hw
zkVq1q8O4xuY3/H6TcUAIDqfRBJYyFRrJajQOvzVT9FwMoIcknlisGmKV6CtJB2iwtMQFITtObsI
hYOJmjKfhB3QUtT88th/dGtzF0Tz5QYCBCldKWbBeOFg5ciK8Ym6YIFi/a043LZz1eFCN8yiD5S+
VpxAxdmWt6qx024uu83Ewcw2YEO+oZqbBWBNZQIyiFjyWYNwQ0SD0EcqX1SNLEXRw1X1AFhKV/ph
UTknLXZGtrywgxgGX0FyWJ3VpSOk3jGENdMW/2owLCSfSlhandINgLhzncMrJfQ/GgNfjEs7zGWs
grct3zBxyZVV6R09Iox6u/1Rs7tr3vx6Cwfmkzr1am5qSO//WETyL1Qdk+/ZB/QyFn5aiydYAL59
DhHxZ0RskDzMrMlJwdVl9+iotu9+x6K7xz0msrFJPuMnxD2IrMDiRJ5zqSOweDoF3FNe57wUEiE/
GcpcQE4oem8yBIrKdvuYYLMdsxQTwDb33iVkclURCP1pV7MrLfqLgNEIvdmuaq77u7Emx/AG/J8b
emTUiddd9H8Ix47dFG/5v2xy6PDFpQJJZrP/uLcr1yHryqnpiVrz2nmMU2fgB/1PRPEVHlTxB6y6
2pMxeW1MGURBH/lDaAmoa0hUbmKqz5AXXsqJrBKvlbiYS+Wq06FkdKEy29XZ76322mxgYh2gp4AB
sOUkZVx4WKqZS/iImKHpDxsLL4+lFRp0kRLotR58jw3hhHIqcJj4AayZ//t4NujkboXS9XhLdRU1
RGbSux9RDWiWu317l0sD4g6zJYBwDzyR9JIAWnK/1C6To72a8p4PEA8G6n1A8KdJL3OYltTSVwrG
Si5f2k9sCuoUlURs/QddT3nJxOSr42XGITn/vjctqmAn5k/jWBP/K62SW5HMLXYBs/6h2U3/YnJP
E+ZwHOphns59jA4zlcE+c5MnenKXY0sOykrJGtpyq20D5kRRbOu0CxDQPU8H/qDfkyz3uVbWLjlL
VLT3lzThvgLxgkkFN1rLyUvZi2jO3rBiI4XjOrhGMaVSJ5o0lWJauWYu1qiMYGttNxegD4+CDLK/
IbD4OSIKwprDJWIwZKNATHydjETESVkQkSotO5GdO0uUR2s3s8NXvRHJ5ZyXgbe52n8HHH1yoPaR
CC0MdHAhb96VM3JSEx1uPl1oTQgRN77gghweeyA6H/M6d5g6GYb5fNw3yOtGArDGORPnRmAQtnzz
wsoy4abVm1nzUI+1HkPoxw70vxmN2lPJYkwKlOsfDS31IufImV8eJbClMr3QyOmS2u/70zujbUqn
ocPpmMJsNlrqDk+wyAo30uonxGDd7+asynBEOqwi0XWo1wntTJHu7eISXIHNPxE0r+y2zF0AkGQs
xLONdqzbzp4jlCtzOD0nW+S7DSCq2VpSvZxuGseXg33LB1zf4a88A+K69o5Nskq8OJZer7Mk+qFG
JICN3cUOo5KvrCSxSNDuXTJcQbozThcVYiK6H649LVObLsvrw2X3co68XhHoafeJd4LgBVXIZJUX
HFSdGVdyxuqH+FnX2J7eKB/ZhdGwj9Lu2hol2G/9uEy7nTbDsrDVcDvuFDqk5j+FayEfn2eCnvVa
MBUJpLsM56WmEHYFQ9j1Jj+/USMW6z9jMZrnRVlnRa1zN05xiOwfk2svk6VAxWAsCi1+6nq3j4BK
fP7gbIFpzn+Eh+jlkgXSPfgYXExZU3fT9K+lQYI5bhwC8VWrRJJKASZPwTY8VCchXzhwJ1tuSEX+
1mpflGbDVnbuGC6FjYddBzV6bB8J7fxUcDN6jsvlsx2Y7M0zXz2xTqifWNdzMO3Gkjmnfs9EsikY
SsZLLiE+732DcdmIgwT0344H7lF7XffzZFb/H9G1TWCIjT0CkDG03ccy1n63os1OZylfeeypMUGq
IIWrIyJazuBC07ToCAK9xaXKb1nHvUCuwKaOS7bhxTV20FicyEqLadXHLoCnvBk1QMkz5lmC0e+h
UdRtS4XvsWfR0V5WHXY14TAXnAp+deCG+2CHOFxZ2hDiHbf6gd8YZuoY8/HaF448a01guoM9E4FT
JI7faOBd9+xr8v3r33LotXOhtazpPNwbAHVqvm4lA36QCvdM4dQwwSbMpd7CCbY8UfTYBRbbtCJ6
DR5EShqc4ftNDGz2lHBJ5EFMMl/Tu0sBMWKLIpSV8dthI4SxGjgDAfXSssBGjI7wXkM0vzYesySS
Jc3drrmG7lO1FnSTa1rwTCQu26m/gye1RrhA1eJPjR6GOdyOkjBfghnKW/J39DQbf9TSwjCruNgV
NRcxoTPoNQv/23hOQM1ThO5aJYSM8BXOn1PQ3LsXygreKBxwHl/13ISl7Ubvev4z2eU4PKw4m3Ds
D+j7PAbiDXvPPgwfUuh6G6vcxg/EhbZ2CKm3kgVHmUh7mSNiVU8qDqvqo1ihJFP5AM90yWfRMie2
jPT/wjHLd6Wt8tI86MnqgEsmggt2BOILUDjB90Lsd81e6gUiTTM4fDPojej5F4So8gidwZu0JxkG
yAExya4cC3FGOwEc0ZgHaltRWwce23x6vrBKVkJtVrSO2tKgWm7N5VMGsxP2E2Nq0ich36gBlx4h
2E1slnzdDx2IdsRbSex6UaYNZYMmHA8Ik7e/94M9svVQPv+cxGQyqo6UWXbTFGP3dheThsvRC2gc
Gk/Y7uVNe0wBKrR+cO8bjOlVBW+pNx7P1wk7cXuae9mJ6uKXuftXTHx/e14qkU+o69c2wLdhNeCh
W/9Z2JQWJdSRf0sBIp3284cVlgKz2ijxluJ9k70kJgJ6ociJjM0B+w9JFqaPaDoAJRD7eoo2RbES
DetcSNnAcjmjlE+0LFEGY2fQeLIKyRhtGs4hTimYwGgGjnTcZwWiVllPYdOqidIvsY7g3blgTLMQ
58qMYs3onK6Z6rPXBgpRbA66jsfbdC70fnpSm/WJj6/c0jXxnguNtG0PnqSrw3O0WOUvd+eKdyw7
f+QoM7SauKYRTMBowguj/+6SJhCMMj7pzCPtHca/vvCjHM2zYJq92kdZYDSUHu4sPau9bjq/k0if
irwcrt0X95752Quv2QMpDybwZWuGNkgq/UCPHbQH+N6Te7BOD+Cnr2mHBbSUbPczz9qa8c7IJQGT
1m10UDivpQqx44Ef3YWaAF+poOtzTUmVCyrfrKDVi030KIm7aW9tkDKZw40zZEqV5jKSSKoPmPIo
80b+quTeOUbzUFKez5oD7ocewEGIp684TeHFI6asiihKjOE9aTbNvSi2xMk831lgjKIU5J5I70bu
4sga3RnzRlNjFFpbegKevPDdTNqMcHZOCeX9C/cB5jPJrJiQAxFYo9ov6G4cHl0I3vj12BBY+Chj
X59rF0rK+7hvCh7erds6YLNYzYL5P471Ucv1qFRUy39ykGDFfW4AW1lj2iXZbhf0TdxjC0emiXbc
xQJiaiH1HAoRBVK5P0+dvTZvIrtaisdmL7AlsMjhETSIwuTpsbbRTSezn9hfEIOdG9G8yGokFZOp
rDHywi+tKAWY/GUVmA1uUEtEpBFt4Q0aZWSjhyQXky+bRDt7FlXY322cR6HLzQfgMsSFLTwxi/VA
f2WEu4KvZG+1UyQLFJGa7H07HLYslla/fdI5Z8ZpaLmttSLqVuB5Wg8gUlnTnMWwKln2lLCehvRl
Zpr5nIofFMIR45yizpdzNBt77v2I1PcwXVZOBnXhwAKR51VJFLX1Rdv+NfbeUDnHSlMRZ/B1OBLM
qO84Hp4t4fyWIwjPXfVawThtAOd22MEres8V94d/fbv245LCRn7F6A1nmhTIuRhGru5oGN3Qm1fW
pj4lMeKDowLArVxPJwhaTEDsPjdH5AcLX56DwpMngEjHLHkzkVMVvA80lUyHfXqDSnCxhyUqVTiQ
elmtLPZFnt6GR6JftvC/Xu88Y5Bo2oa51W6JfUjEkuF8VKcd/Nl7ATR21lJuEaswfh1yRHJRV4RQ
WmP0NYTo9V/ejl1kjWGJ88D9oE03GMQ5OTCA9+3mIk/jsI2y8ofn5xFVhGP9E6BhvjWDSk3ZM3Ca
k5vErnqsIRAihlIK5LuF0g/aIuUZETGEp1DNTWfXZIkxeT9b8tNKGZ8dWoUouWnUBPKUflRJjrJw
vw3w78ikDZlq5XBQ3J9Ryg+FzR2BHulVZdeFfWbkGyTwl1amjR3cyXilaFDZOcje9mDMifxgBuIQ
e8MkDghEX9zz5BABmZMuogN7Y4pK0wskCr1Ck6c3reiPjLxfPsEqQ6NeNsV/21KUTCknQMIsC0Zp
rxmYDERJKXdxF5vLtGkndqX1pgQ7PdJJ0UYTgAyePpUIXf7r47v30SNnLynlzcQ+LcsApzTSGUHL
jni1xzQ6CKLpHVaZWdgOySlpavDluPPpiYODSfAKw4AsnHCdQJyOL6I4H1g5ovRJp/Zsv4Fl8G9A
fvRmAj0d//s6KWQB0wv7e8Djz1LfqltxWZg1faZLzK8G18spZqUltIvSpfyu4hd+mwvxjS2YbbZT
lV7biU6eXGG8FNAC+B2Lt0czRo5DKrSTAiop2eQiPf53yqFKJyuaPSRXaPXNOT6u1PtvNJiLPxQL
6ElwfejajqwFpPi4Uzm3a8oAHMyVj0NRajDjjqfuUHuw9DnB2LZx20XKAls+2rHxJ6UXuUbxZlxv
DQEwpVqnDXjWMcUVlUHgGEEpaErtVNeN5Z2nb34RUFVX41cRZoWGpXyInvjm7/n0zLUy9Axj6s5c
1hgsk6xAeyum6Yemw6HMnUljMowGJt833TsoM5VvidwNUCcJBu9hCA0VExkPTF5uJbCetWmMkxr1
fJiwlkwp+Qwg4OvCDp88MLSPxhzamY3n1n2VdC5AmIQExsT3feb1WJVa7HllDip2pVxKKw4blMCa
PVk2i7PHcHXfq7+vf6kJMZhTmeKDNEMZCVWeX04GVPyWM7SZYlROaoqG4EDjdO1nbhoUtEvWYJE1
Y+lx+Bk1BRWse0TGnLJPRCSddk20jZ9Qfoi7yXkdrYz0emCLpM66u0on/fDuO2hGu8Y8Wf7Pl2y3
DDkMO6xHvkApyHQHiVsqpe1akLZznMDNBUYVjEeYSYbQEHpOB9qwGvneojftO3yuK45gp4os72FE
6m9kXRbHiibRSlb8sSKxUcegX47hVPWRl+YuMQ7JfpqctGVv5sUfNItc3gxBq5k/OtFyeH1OMRR6
J8EoUYsKxfHqnhMR16OKmj5J3FFOvQzLYmVspr7K1S5eEtjjSnD0hVy9dhbZ91so2EbExAHeQ44g
y5nAJwlOWyk1Kx+rgtPRUqJ57CfiQC9vFtvZ717gnoc0v1uUuG7o41OS1QwaXeC+SdJIvQQ2rZc1
elOw37NFhBJM6UgY4nB7gszDP/bwXcv0ILx0AXZNLmiHyXJzRXmnrLLP6E0dFlVAcJ+sSgog+ezG
qpEcM85Wh679YniL9NlUPbgVzGkCrxyN6M+XiJ9+BDkBEkDLtM+0w198STknxqicjOeED4Yc5Q5X
2xjXlV+2Saz6sw0xN1pxPwUrbfZqEhj87XmYyjq1YraXfzxvjEw5zQk4piWvM5fH4nwnSj2XltvO
Mgh4ezePVr9opsd/VlX7eNpzehVCTkveUKX8Y9VL3vrts3JMUxpn8k5O1cI9sFQS4iRoqLJCW5pZ
R5zImwQpbfjEK22haqp17Gij2OWmmdIXubyQIsslrKrCecdnRDbowJv0nHoI2OLq5DMDOqHzbMcD
U4aeSYZEJ5D7aoPGkeZRv/OIcaYUTmvIGqehaM3BAxIop3vBwF1kdhTw2zgrsOH8l7BONOzF9TwS
WbUbq86t54G9Pdbl2dQ8UnurFI/m9Ij0RidTSaDIIGGKDY12r6pyIvHbb7Hti4wV2eshJuDz9pRq
k6MSUADJuqn46B+oSGOTLfQ8AvLuGDAnODJJvL1b9Fv6++C/VRP87/hIP75xW5/adiGZxr1F+zWi
8yHJGT0gGVPHxyuFcmZJfJ9SxbZZYpgsZob3ICq/AXdt9u1hThcCbKIfEymdQeUJeqqRURcciSqw
0k0uMrUfPLu9uFBQgShsHdSgn9G1WOdiieSGuqCMCBIVLWXHdBARoFL5afjggdCnvaWppwohbZ8m
gQQEsyCK5IRkO4skLYqInRZK46qR1lkvQkqMbSIXCc548nTtHvdV/vOo66GOWv8XcDzHzuB578KO
jp6GkW0lZJWDWA+7SutkKT2RId4Jm7b+JkffnPGpEbF5pNtHGUIuAm42ONRqWzPgcU+B+D+ZVHxg
Qc54WeEPL95FhvPA+tZBbeMsMSrEqtPGeNM14JNkpSX3PJZDSA9PHkB3/x+yoOsgusdbXZu+PqTy
ZCrhmzQYDlo1vBA17mkjCbNVrjOBzK3iUZ6RKotjXKuvsirUJrYn8O8iPQdg08sScF9c1qrtcCAO
fDlHjtGsI6scHkEYmOfjNTtkbhglpMwQ8AtfoesKsH1G0C36f69wSm9Ahxhs70MCP47ljTNzkg5/
6QA4A291hk+84cLMqKqnh0KIBdRs76fkiW+gkuvyXhIEN++pMF51YatW9ePczbLb/jpKBnhju06h
jnFbqzYcI1BZVYenqrvqJxSx0J2iymJV7B5aWhQYqO+Qb0AG9B+SijLW/AX9wA5BDLGW+DuZSLxj
DQyxRL6s5y0vjaw0JYfVM2OrC1t+JjgnrokQyjHxwaiKQ8xXg4sW1fVUW2DsToMWBTm8XqK9S/te
oCMu/8UsYCYpD2d+UxDsH/zhBSVKoM4F7rX5sLk7yn0O3xGsDwRrfJMyRops4q1wxq+dmtfEodvD
OQTVT/mN1UEaXziJ6dEvuSHHjt7/TuKIRClVFP3ZzlYYJjw8Vv6u+OsCfInmzeNnfYyhBXVvH4dZ
wgbEsAwdGl2sB2vP6+V2LM4RxKLcbaaOl5jB/ZJxS+AruMYUVAv2K3VrcNezTlzucykhMtxyy9rm
t8PXcxeGIRlHnV7RhoXmgqV36Caw+Ib1LB6QsWF4PUDOwwf+6cU9fUvfJ3k9iE3eleTOXm5V6M3x
YbXnpmpNAEDJftyAdzHHY8IMwOLoRytEWUcODNwNyrH5Vzqm0uhtikoqJFB8pFjBdwAI8r6UAwnm
2oUlhlwl4K8c/e5mdBdZlh0TwRIBNbOpSxpeN7wTsgNVGiIDkRCp0EdmpYYKKQDxIbHGDIU+khQx
apJoLGlfV6UQQQtUqoBlcWegCd117Db1LUZcfEaBfDx4Gtf0SKTg6eaU723+yEbMxtwKe3eMJbHC
ykvOif9cqJhWN8hkjAvxaxuQOZuL3WicuSU3s3vwvXfdC8IJYD0fM1gRWoUkotoDiICeowZWX+TW
TpoUIn8fXCOpnvEK0iKRNDx/aZ88ZtOJU88YKXnr53IJqqcVwyrjd8DwcBX5A+SZm0CfbvfZsZNi
p28fl54E+99DCQ/9vlYxTBQEy0DYJV+F+jj/jV9b19Exr7BfeqONl1psDSM0qKzpWBLJN1dltym1
vYv4eGcQoY83mQKye+eMmld9pmsAhWD7uI4TkjOgfLmetxnQUkDDeapMP36uymdT9pNA6yL1s4Em
bB3fzs9clGgjEij+bDB6wCohRsdN+xLh+p0npTcQWSuAp1N5U1W0WrwtJVi+bTqQxnSD+V8ik+jz
+1/Es3uQ8k0FcWMolCh4K2BD0MyGBF3QFCD1zCZDxPyNZywEibUG2614M/ymXqg67qFTffburmu4
besgPVlzDlcPws8neIPz3oFQK14noU4UMUhJiAxuDyNhiCxtQ+792FI2HCefzcN+kU53uDXVKt8g
CNL3jwV7PBiuLFokzOeZwr6SQqUKXjlFPjxDvYAETL49lItRV3RetQFb2fVfbFiqVW/r1e4Oaexn
/WeLSYB/yZPnSgEby5ec/WBes8624UT/ib7SyOQgYeyF2Rous/hwSglx7SiTTAr6WRi5md4pcCAC
IRRs9F0O86xCbNlhFMAYdszNEnwcW6dfMGbc0GQjsWX1p3tJG1YMcMF25Lk59og7ckRYbzgwTZjC
Sks3OtSY1GU64A/8JidRaKRW2SOcjoR7D+8sEvWAWrv8NQsYBXdzueZP7c7kOBtaDPOxeQtfUM8o
FbpF8o1x65LpnmprkfY4F0FLfjcxMJIg+ucOal2obISIfHAMOQT5d4voY9NQzAfkgyB15xNbO1io
X0zyzHi90pUDinGvbtZ5P67JPqofh3dsiAH71/SV7oRcb5k9FjDhw5oJd58ESW8ULsocipgDMVib
JqpukI4NvRY+GNrYnPNBap0qf1HB6sOGBW1hnjfk4DFoIuNQ6+OAbNs2RRBX99hUOxUOQDET0Vos
J2jqFkvGEDqOXdLdpXIwu6zHYG2UlLnoRa+h1+vAGmMyUpsRhc/y5Z0zbwXo1bUpTiglJs9a3Ewm
eTHaLuK3c825MqqmHeLl2OCUBjL69HWjw5hU2lwf1mqvOlnnqfd1bWUiGluPSWXoxSf3FCCLxoo9
0tB8PUsplGMugq6mvXJojvnqR9W4b03+JrKyKQjA0HCpgoq3vxiJNTxcIGN9ASOYS9zl3WxdjY8A
xIFGnFbGv3wIKOvvoLMzgG+B+n8Y5jHHeNeVfP2M/1rafxhK+Or7hbK2wwQns1iyz3BSlrgx22BK
MTdxQ6KNuJFRL5ix/KY+8ozMgTLPzvV5S0Za4k63nVhl9XeVVsbsYHlHR1FPo8dmr4naFd/9+3qF
n8RzClr6pQDWhihnKyqEOHmSYYBp8eLKPRy7Y8w6rlCyaEWHUA0kX+W6T0KoY9rMMyvLiLP8P7Km
5AUFaYeDEDLqpStktqMVAnDOCPe2HEeQXd/LkuKDj+Qb/Tma2k/jVV+bVa4bYM1R6zLFXpxc64gg
BMq9C6t8jgtEg5t1wh13JJcpRD+lZUUKttXj0dv8yOUXHb802gfMMjClMucdB69MOxFrymqIhk1P
db35acD7xNESJCOI3WnG4cSDMew8ZodM4Jmi6itbi555ACXtbSNRJpVhaJHxVk4J/nsEH+o7YtEX
gWKB3OWft+d1InRYTwVS3XlaAS77ScaE3BrKNRABdfAeKRCTu4bxw+KBetq/l1yo5gWgXDhNxlN8
Eg4oSEpv8Ap8ZhNW+xRbfevXufS8uc3asUtPbyvyoJwADxRJtR0GEgC1pUvbFSZZ4v63ezMyKe4K
DQBGPZQ6bfi2TUAKuL4yZSa8C16/jF8eQhZrvGddNLFTWc7dP3vlola+NRwgzxxZ//GiMKaYXLRq
MglpZaBUxaNIk0TXDT6h/Rwp0anIdnMIOMijPGCHiRw2ge6IzJcxVFP0aLW5NKFpOvsGX63RYyW9
rAsT1qG4kUz9i+qy1rU9y7RNZ40xtqtzTqqO5uBdQgiyS7db88DgdxqXYwNqhrY8apItwwtiV56c
b8lKN8kASnGT1ldciKAwC1kpzGrWBDrLciqWVA5EWKGOnQpiUPyVfQH9I7pWJHouePAEwPydmlbm
rNn0H8AohylxLUbqkKNyMq3NsXtPQq9al8C0yzWRjAoIPMXa/kuaylLN8z+m5zDhGqIeu8eHbMZ+
aahNxP8cO/3gvtN42lEJH6ASHWenmeTP8ahy4hRgTpzrH7e+a3NkWy61ZxX82yQe11OsiRn/+He4
IX7fbc5JqK0nFhBMZFiiNidjiJ7ycffeyoJODqfGvyj82kyw218mtUXeiTFuqMc4lsUI9xvYWOyM
3diJRoiFWrXeMPrvkm2SR+76BWIFi586CpprdSfG4MpHyI0TQLu8S1tf4zpnE3ggO6mbogs8G340
xu9DGDXWpaI5XjeJtcCqeA/bHPOPObsS909JZzTHKNpcyZEwarUYD26n41xXWtfR+qBCRGo1mSYk
9imcfH3VvkvCrJpv5yET0Xiat6mPVRvf3UMjLsQ/GfsHoiNMtNsupk+QJq6fEfVEwtFTRE+drjoQ
Djwe840hztrPtJGaMdOR56okR5au1CXl3cLu1M48qi6mMRP7ahhzeI6XcvJvEBrQMF6jH3eZIUg3
Xx3X+1rKbWZYJ1wh3c+ihPbDGm44v6WmU9rvIuJfD1dJYvoF4KOYf6pSGdcu7g2RnqSRhGEQ91o1
bg19D6nETar+rBMW293hJd+x68EFVtVJscBZ7RF9aypr8rF3/3dq9PgtZH+LcPc/9l6P/9ULPliB
txD3lBeWjL8JslmZf2cEZc4UJYvARXHszeNEXFOs9eZdgW5KRta0dTAgj61GbEac3WtJZO4vxZip
lPHz0kgx+CA2GCAOCBsOe3IrMtcIy7RV0CFn+K6cegt7wSkVd443+/s92x6P468gI40xUDSoWDkR
u0fH8SzWwqRb2p1O1+XFjsN98NtWIbZSG5k+qyWx7LgI+u81nyNDOlEZYVJIwdUe2aLkaHFaBJyq
fsNvN+7Ibk2mRiXC3fShBFHrLUhctHAbDhzRrFp1co2qoh82rG2hBPnXQmkxtxeKnm1XBPiuAvca
YFV+vJFHqeZQEF8f6Hyu0jY6vKGA95z3TkxK3vU3FowRhAKtwgnWqIMzGme/Djao0KN221TqV0CD
125E7MYZv39YNuy4XduSVQd7PM7oR2S920uYKC77r22T4/AXuarcgmajKXmVWZnhBwg0JdK/hAk1
T6zkm0XhWp22CvsiX8ro2QCM412gOs6LSMaTDBVBprczWI/Uge7XC0bLCkUwoa4mrGHpnHEcg2RE
EMVSVJmuiOSi7PDawd7pKA/ZFt/EcU6//jgyjJtxebOyuxdmVq83yrWRUvfrjTmqdZWycKfwuSGr
RWGU8YtRizQ0dBpCtL37Pm4X4sgm++zeh8jFKvOUt3VNcXX0FmSMYpKqWogZXP4S0YGNgGyM9WWW
nsi6kQdxPXpZws8FWkZAasFqYNilpDscSG9Dg/vZ6cIkwrJLn/7tNastAiTB6yb3j4EuYH24raeC
WXu9WdQRA2fAf4hlEllsmPADPNOPa4b710Yg/AGcdHKi4jsftBDCAJpFMtwxFeFSLKCn6zDZSHfr
3u/scrBy0j/b0higJn87yGGtLuE8AvCn1095vcD+ePXeN4hdj4ZjRBTbDDdUB5xfywyoiVjd2Vfw
oiUKWWEqHeySbTsWYsjd4orDwIw4U2gdTIpX864Y6oXNc3YgTNeJnUJDLW9XDQEo6N5N7u8vHeFC
o3OqxDfdEdQ6ptWwBYPERbJdAaKAK69PcUZB6VMvIDa4f73SbktK4Ux56RH/4B+0TjfkbPgOnMPe
sPrzNbGOhfryxKNvtXm0/tdKPRDh+mKhCoTEG1GklcQon7dmobIljqo69YE3iMkaLe8qBH+fVDOB
9sMJU+ikIsb4y5i14n2EqrrWS12vRGTMNHbXWtflO3cIQ/kOoVTzHZlOy3BrOXYT/TwYpytHNmaj
J47alsifnvU3OyTpnaib1zlHXS7uuKMgeBGyVfbgbQX6IzodPjPfgtwN+Isxylu7PmzfR11lnVvL
MOjrZmznhgVFeKAP8uUnDc0QA57Z4W0sY9imWfNZHRU8cF7qtWT8dgDuTeMosB8jwu/dtaJdT02n
6j9ZrtM1iEN8TcUDw1MJb2k7o9q6urPL8RRlVk6yTb+x9XIHdr/qdNiJPzq9hVKCTKfMGfjsXpVU
BNXrupY3UKbpXiNLGTZTuoF5uDoAh4CJ/D/HU5W1EbF5O5AVhWUQhdgWtw4FlptkUL9fiXIpTXCf
bOp3gPTc5Fd5J9GeMQVDrIMk4BCbbniVeKY7H1mNsAqhRN3f09rzMGkwZH93aoFE6ZrNTQn449dA
NdY13gTThd0913mq+XBI5dLu6z2j7dap/nTrMViBMmnqMi0Wa+qiPEFDMVSuOUKbMyMNaq1zH2jF
dN/jFnPN/JE8kYVYxNxb3qQWpqdN2PfdBhd3+6EPnYv1gaItimBVqB4MXOBU+aFIr61nsvAxU8tv
sXSb/aoqu0VuKyxlRwsmIMxEAgSqIEP5UKwQ+k37i2I3RJYQzfGei2LWKIFMkI97nJc2CkKRhCB4
B0/5jREOCNiDbT/9GB6lCCz0DDnVKpG6Suna4Uh6S4haFytnY9bcHdMPIPagUPiwLpVK4KDTHAcy
2wP676e/0bZtKM+wmNR9Hd6HJsuNKkIYMdT/PK88loH+qhp6wiHJaeBhXTjRsaHv/4hwnrrrYK+O
ncwwgLlYCwz2tJgsf3RVZSYXzSDBKWseYZp3A2mbZcsqitX9xtJfcebo+0jFY8FsmFrszdZ/UlWr
fi7tnbJiDa6OtNILSTVT85Q7eWR85OaZLQHCguL9FKHVSNtuwh2GU/Px30915tNTpP5awL9oGigK
8tvMFh16lfuaZcLsPmu0qeJmfL1yccJnytz5YGY9KJV0T5/5n2RvzkelhBSurHm+8SCi+TFzpFUB
r4SK0gwAvLy+/Ixh+YKoms++Cn+HtxCKTjleMYKHBv2LGCc5Ry5GzVg4jg9hg75Apk6bjk47x93L
i88aCCUut8N8PuvEYA5BQrMiIm42Qp6wY6ksD38sP89XR5weFZ3SWDinWGLRZgnx4riHYPsREGtW
DTSSJTHZgDIR25ceOnafFngJtgcFoDSmJjfB1GMO/21/CXY0/Yk3I2YDnVabzH22JpMLrqIu5m9a
ENDFSaVCYyvEomwoWH/MAZPaZU0WfurrPNtn8G0vzHlJk822Ht/GVrJJFANuHaI3pOMmTHDtuXrZ
BQYaAyYb0ViyudnIwCaKAQP7zs8OVGrCA8yZQy9vELPuZyRQyYAOw7eIh06PRu0p+ohZEBAnFyWb
ClXXLDoudAA1xvQs9owNlB1jfZkr2ZiggxQsEuC2mSp6Gi1M9om4JCvl9OBwjiDroZ4mepqm8ytz
udETPctlehmuooXeeicAVpr+scx6zDzPPLFHZ6wMR+oHMFEmk6DLiM5aQVdLhMsoRII17WhvzmUe
da/bC/Bu8+sPCwGuHtZlhqx1LGRJPuamCgIYg0YFcVaeFcs4TeTlXK1Qetx13L/16nTWis3HJMaL
nJ4ipK0NtsI/o4MUZn50qjmx47MzPvJDDDqQT01krjBEgYq1nlr7PgqZmx8QurzYWIQYEA5wu6jJ
cBESA1BCSiWMEEwm7Aour1W/Z3RDElomDI77W3n5vUwoP9FbDuTbCD1CbvjSsT+PKqeHVHbDjeXh
NyBlh1PYDwhDty+ATESKvxnEJl+fqJV3ScU8FtmliRm8NXCoWrFKs4HU+6BtArvvYa11wYaKqeye
pffUCWgUQUMJlWDjsyxL055Fn+xzJl/3kmvTEbXagxKs4hGrHMDHx9aJ5jD6iPTC+2FnO7KNiVXB
fpoq6mnozWX+rC+cOjigt8ugXeslmTmOs3JTuLB0i/qf/3TIHfzdg+SHuZDNRLCLylO/sD7x2Rs2
Mw9rMd79+d43+NKYfM+kDnObRSuFVz2Np+sJb2MYpaVoNHe3tsvzXuq4jG7gM8EVaj+nh6wCwqgA
/tFzwQcRDO3bbn5FrQEHLF36/AwcZpGHn1vbA/DZjzQbvsal0hmpOW7PH2o+aIiqSXpElMBPmpyI
e+CaHHHQubMZ6DJvssFeoBkiTdIuv/9v//DX3AQo262wEoWOcFqq8iUqOECkaG8BpGeI3LOaAPvD
4r8zK+LMVDphfU/BO7H9l67uwYKQQpsRS2UQzbclx1JlTRv0jDFtFFWHeL4JxMAb7a9vAXDwJ9hW
LnJ2Qit68c0PE9T5ipO6GIp1CIvA5WjQ7yqEYwMcl+whyfkXGiB74f3Q7+nfUP+j5Lhmyi6GG2GT
sus1jLWN97eqOBJ+/BgKfi0CpCexgJeZgs/Zi2gMAD1/MhK1plzgTMObOzX052lhMkaw7+//ZV1W
tuYOhfdDBBfIy5Pfh4tKivEzExD01hxcRfn0X+QPJOmmObY6HHVevuE8OHg+wHVCBdcqWXQKTIrH
mhC02ua5FB5s041lCrOOeTAWuhHOKgWvhOJ6HoX4HBIpUw/RjGWqAMRZBrc6vd+8SsvHfOtQgPR3
6me5KMrufYSAFANrMv0ZL1UfaE3Ot6DwUR1yee6+2nCjHEMGTxhQmJKJ6pp6D+nEVtbbSNk/VuEP
20dPYN2Rie4c/OJVobSvrW2byVAoKpJck3tsyZS0/WKzDKZb3QUGKkEd/kaCLmdjIebZAKBP9CW3
GOdBz2/z7CodkaLnXLkOGemfj1ZsFzQu+jLkXYh//u9JYRqqjyqMEnT2cvtqw/vvita+wbi3PF+t
En9pKYB3gArj9n/92fx1aqZezo+0CpsX7SvaD4EHA1C+HwMavntSpPHoE3xC36Ckmq6qAA6iRuG2
Yhq2b14S6orYHljTlK/sid9GhtEF6d7QcLtmV3vLjyigd5hU/xset6JjuYJ6xSzGtRzeInbaM3Lr
t+ZwIn7a8WM5JGu3NSdT8pgs0OiXfXHWZ0dr5wK4EMPzh9Mkrd7ZIMUa/vFJ5BtDzu9u4W6N7+Ge
Szt4vNg4Y1XFDPttyMzjtwtvUcR9nNdYHKOgbVOuGwbC0yn/0cm7xaqIYqMORMk4DM99kyDWLkP1
7SBShptlTQp5nWFCMGbX4Vjvboa5OLQpgYwAIq622Tuc1FQ2mv5zk6y/SdYUqfAwvKMqiictPtUm
CZwwZuoz5HHkRN+nMzARKXSTntduZfOSAvLjbutKhULLS101zLnee8LJ2UkfpexbBpkZlkNp8c2N
ba6CWo8CLfUUct04nLZ1QFlScC276rY/f3UV07n6imd8ChTbDUzd+qMdHGW/ZovsoPemmZiPQolF
HY2c7zktVkvcyNVAf1TKBCrGr2OpUQCkYbsMyr3jr7/S028CTZogZ9/nHRPwnN++rL3+oMRNlSWu
22klGtE3MZ/iejyenSaWcpcbzYcYZ+GhS2AlAR0Tz0+IUemqjVxYwk2SuEje412PrGz1jgYEjdzw
sJApgp1YCOQkV3/b5il7a8ub3JbGv0WRi22EJ/gTvh0zf+iD/Ewac8XbWAIlK6OZaMWdrM14QXW3
0SPEFiS/ev86exKVdLx4Rc1nRl2xU725ehzj1fsnYql8lsgkJNe+zU02HCQVJdoeC+Y8Kp1MMNII
swU84aOoQPSV9SJT+I2aFey78AEZXl3ZFBBinxlrRYElBt/xbUCx2OludODMoK6FWq4e7M41/bWI
pZH8UAdXoNvSpROzNVvVfT97dJ05No03mqVjLAIffGjeS3hF9oF7UvauFhCaN5O3vUo7c/pyIAno
+wP5MiecDF4A6p0g3GZ8f2iZDCg4pCF0ZGK6Sheg8f/ssunl++h+UOqKXGGjr9II3dUSuxThdjnZ
AfabzdMuRaGZKeu7nlShN5ryv1Sm9Tkeg3cjzQEgLSkNmMVL625GmOLrNl3+eerUGkcU8CMNyyyA
RQt0H8q5iVS2cRto5ykeURDsJygvWPogo7gSFUEoGnXl6Ib32tkDtepkO7DHaWozzdqWkJ23jILK
RcDqTD0M8x7xoJE6R0X6D5Ivcz/y1HU9g7AmP7EcdI8phvlno738oV0nE3WYEgGRQFYLZQCacowL
74lk0Sfrhs6P4Z+WakDsjpOODbHYWyAlKXtItPLE+3EPQDWfZ1MLzABIKJ0pEVOdrpldpqbVaU5W
JKz9MthA9ZtRANJv3jh6LuyPnw9gEcCbFJaip5xKJ/MJg4U4tXu7E8LeqEOGJmusoDE5YTPK1VzF
dslEU/chpnoEcTyahr6r0KaugloAzr1PKwd2E9xdCzTNNUPRDWv5w+gTUHR/o0IvOVIJ7OIWh1/+
oNTt1JHkbFtmouIyk38OB+19mgsY247to3ZhvvgLcfTwMovrLirC6pr8zKKDGEJX6Fe3e6NH12nJ
QVktFubxpdopmuovDFI8Ml9OYatmFOsLDbRyvzhtbrsPT2eN9yoCaSYp1dmdyB6uB02vFtFYzljX
oAQTdnTx2hDnadUJSWlxcYRYhhBINKcl67qGDjWRdJY8oc1lqGzbvHz6xoE/92zTseKqmbICIMz4
/sYX+JfkliGJGd+V0gDY+AnGhrWra+JnP53aMRUJyoTbpr6nf8oxVntFtZF8qzdJfMI6LE/pPQgQ
KWtMc+fmc23hQSjPuzSHdVcUjo2UieI+5AMJkyVMsMNhFS+k0ZV4GUpax50P8BPCokOSuwjiwjU4
b4Sgmw0ZNAQD4QuslCjM0ZOfEXms9R23LPolTy5kst608GKJdEvlQUgcQUGOc6Vwb+qa+qADFC7U
yt5uy7PMKyeq9SO1PnPOMbL3MckIQI9evjZeD5Bvjr3+olwcbqThYPb5aCbe+5tYVB6jFCFZ7OeX
+38U8TIZHQlImsLNMUYDTNhMRtWFjxXStAUR4+rqRi2vo9Dndiv9O5/igtC6/JtNY/m2CejlYA70
Lc30UEpz9GbbHXaaz11jXwv+VEb1pibcauyleN3VzQXEWvLzHgp1NzcZYa6rungQht+IJKmhq4v6
wO+Cnl6WXqzOLb3KcLZlVCvrrdPQ+LJ90EiNp4ivKak0pGw6yhEw+UOEJeU7UzYe2s/evdwkoH1W
FL/qAttFL3fSa7gAKm7/5Nw/1JuVTvznzf+cysMedVrsw0qqu9LHNcWzsa+30IRRlSKZ/oUQ3dvW
9UJQlOlJMtAJW6u45gvW3F49SkqIAQE7Zne73YxZ844nSEt+9lU+uVIcZeg7vNZc6krnxwW9H+he
6J1vA1k8HXbaKhIkC8CPkRh2l49MiondUl7dp/ABWaDQazGTdqB8pD7cGnm2ZFdaNUHD/AsNHP+Q
uEPijqD9rSPqYVvHYGSPNNiJXCryDuQLjT+7f21tt3GbUhgEfIxkqph/199M66MZBJg3DkKUrDHd
BaVqNPGN1ysyVQ9WX1MynRAzJZefnXXL0lEPkxp/KucKzfe84w4mjrGjTrTQLFTd5gSRXuoPSup9
iM1YBXpvrkdlHMIsS9hZtMUI91bv/3MJFuYAwwfTdUASul4seav+gOI+ptldBULU2L/vXIrIpY/6
IPMnMrUO4nIGm8qnctsuTqB1RrBuVDwKUSqoyEbITkg7MapWnwB2W4QPToiZTykzwUD7b6zKBKPu
VrSQcSe7LyR0A+M4jlkttr1anZUaaziomd/cvVk8DLsqQT4vIFTXVXhZ2pvRfIA9vbbaifl+o0hv
R1Sus3Y5JhJARQBGJEAmwY7MV04tFxbyelcWfmTbMAYw7TJrNcyX35NowsUA0C4ZTA6FfDNFC49O
V9wkP5qUOiNWCdIzYsMrQnLCgRYqCIGE7M/kBT3KxMOzF4HLOMb3ir4Aw4lIPtEUXpijMlKodDem
tkF3VlkZWhzhoyVt1OKkPGgxHw4kArhOrtAen+VXM7EohEKbuX+WqZoWx8ZerRuug821Aa8jDmmo
gUExIhjQ2v3OkAQk1FgfONvlqLQlkm7oiypxzDzZTYUQS8SUvRCVS2eP5Rkz7oqlq6cy5X4voUa8
rMFb6C9TG4LYNYI5NxKBQaukSviOvF2TTWydvM45cKdEj3HzTbbANHHRMcfOY6e+J+LqrKo1/2pT
bDEDhxFY6PQNq4uvPOCD1DyrydDkFXhLQWv6jG7pL8/uNrSydAS1SwBy/zYQmixWibQSKn/ZLoY1
601/PbkGoutz4eKKN7Q2eC3cAnXocYr5ToE2S1wB4viH3s6oxoT3x76n/zVnsUr14a1c74gMPMmq
Qv471cTLr/dkT9/xmDQ937PaIYrB7vcVQuPPpGv2DfD+ESygPufRE2BuAfuBqwf3US7uoT0LrJFG
VFr4ooSpA+h2lcm7x2kQhJpoYZYCSJj9ajBty+V355sQs/EwrzjFDYhyPxKF6teZpNiXRwD1AhK7
XIINAwY1zkcRSug2K+Awo4/AgoFXZGC2l1CQNJfJ0eAKmhIDj1dhK3Jy+BpjzT4YZijWLqzWw5fv
tnAUoft7yEbLMFjMZGTNacRBUS0FIjUXDDQ5dcSEKZmmrL0rVeV+wVBY9X3WZCT2jurmieAYX8qb
PIJ7gQOstjNX32JjWKu1IMnEJNxKVQKrkrOcJTHXm8mt+fwXAyy30M2WJFefcQUyuAn6xMFOrcJP
ePVek6btcbWv99BDnfDu1NizWB5ak++UoVi08EvEClWMenokaYm76kPmTOHRLeF5XDEU/91nUmfp
ZEwPicTnLcALhKO4cw3GLeSffyHBBd+FzQS9DU4rgS5rCrsamudlNmYlEIw30+wse0/B+2DnZTGo
ydMOLsejdQwV9IEg+OyXC3Con6FZA3BEBZmHkVt9DZqbUWqKUDKqE94oc3/CnGw5m+3goeARHqcV
W6FnZySO7zIr7Dk9rq0qoOuppKyC+SHwrTAc+FjLwjIuuHASXifM3bSueiOQcy0lZnGSIsmWYu94
CVlYbCFgLjI4lH1dW3vcyyQWaDsWPDgQvg1t3di3XbRd46iD/nx9vblyAmCqNMVOVp0v1blQfEtO
SAh2QuKYU207FTo7jbapItjwz1a7TGwdl05M7nGNV6DZljjbTRPMOPbld0iVEivvT/oj56u7Hk+O
lSOKQuEy9vtbZJniBROPKs7eICa6zPub+5ZUg8lpX2jOvrPsZrq3S1Q1PG/8P76MLilJFPE+UTSi
KEI+DBPstcznX5uzc4VwgKLr1oPq8tOy6IVU5tjbr1EURsZy/ZFrpitWhPQuo7RcWYAfQReRWZ6S
E+pxMASbW5qUI/K5lyo+Y+z5qGCX9sCjNPiAunzFsFttIfzJd0JeEE806M7jbnc3vgH/jY6LeTRq
vetM+8CH4+2vUspdlYvyl0lVyz19U6cHVaqEl7xCrOfjFXuiZIwQ5E6UG2VSEim8ehkdCrmYvidd
QxLGAK9vQM8bY4Zx9RihIJ0PEAQCfLmx0T5bSyQ0hnoFXkZ0ClnO9X4KE+E7HlLDe3Fx33eJa5Lx
LR/7AV0Biv4/TaVuSfFGsbFi07ps+PjizGfc5xf2cnNNpVFCRVfMjdkoc7nPY/Fyr+7IiBgqANuw
H82U2v1EVHvwGNWWrkjGM40pfEZSxCneVi9uK1f5UBAUoKvGUoVRk38Dcyw4G7C8q7QOYKa+TYuN
ieVmk0j0BkhoFRcewNumVu2zAeIhpraC0mnzxbBXNR2Agd6VV9Z7RUaZES3BAvz/lpD7VuaGctPE
tB6b7eSfM10L0FjLy+PMRCIfpszpBdqsQDrXMUe8Xpizulf+zUq4xKarejWBAvMv5Rq1TvgXmXOz
UM+DFtsKA7LCld57Wvd2RkwY4udObirple9+zk5iGqPuElKvVSeLDhCemUpFfOJj71IM7egYJCj4
yRBXF/5Ay2QWeGfGr2rNV25BgUw4+9PFg3b23FeA7F0TAM5/VfY/YrypmZE457foc6K6iXjjtavU
QUyLaBzmTv9ca6V9+3Fo/uwb+pGzmmo+S9/RvXww5G0ZjqXsaXZH0a9EvpfEfDPo1HzImEiM5Ovl
QTF4VeMa23PsHTb0f9Imc+VL/DGSiHghzn72N4HjiVc3l5brHgkY0oCVA3kBInEauHASYY+lqpsr
BriseLxVJUTy8fXEY+K94fkdhwGNZ9Kjg3sDic+Hvypa0MGgiwt6SY5z5XsjEU2a7xRO4nFqWayv
HMdQG4xNiUwUDAU9+3qsLh6S2FC0yivUs96SMC9RQPWMA4AqAbYRD7u5kmMsXhX1MrZmpY3bV5l0
j9TJZ/8NlAc+q44c7RHuFfaIOPTNyR18jljMTRk/f9rDmzxmj+njilEy1Pz1DqixlsxmOCfThuEB
NaFBDAux/qJzO9jutKWI0fCHkgVfcVDtR+lmH/KbXXN1Z5jNDGk3Y5W8LB3gO6sy1fu2HwlATtjT
qczb6Z0eNUnIgc9Mep60tElTk+zc0Fe9+HaF8sFAO7pxZDH4H0fRYxblMFdvgz8nmQhh3Fm4EpW9
0tjMo8BXRHYWT7gtPQpYYqu60FHkxj/YM9tvdHEFPsnYgA4PPMHYqnanFTOEArxrc3N9u/Kc68kS
MuVfA0TfOwRGO0/1vaTnFAukV7qc5MpcmzoMTdgoTmPJcIwxexYUknmoGB9G3MZ5PWv8XqCMGWg/
YPemDdq5CsZ8klvv0F696G/fXFXDnl0jCvWh4A6IufnFU67buUvHooO+T2m+bGQRfR8lzp5P0GiM
dZaW4gPfffsFF8O35H7PmgaqsbGsvNFRwFvPXs9++Ux6PBwrvkOCNGYqsrGVuAeaPSpfDR5yl96l
gbj4Rdl5qCIJidsOSLL5SJVcGL33MOEhh8aKjXCp4eV9pu3WhqRuhJVmHbDI95qRH/qATs7tPuXs
wndK1Qgc22y5+qLRsG5YFFJHIBuPwZKTr5t7iDyk3MrgxuhqsmxFpWpVCYWgb/xwurhPYELQF7jB
vo565Pr5NQqAmvkhA7Es7wp8EyPvUnHmS+JzJpu7gLgXAB7MqU4+1t583v2qPpj/5Iwt0QIxBmWx
wsxmEdA4GAQdlnmXjZh0eP7HgDDED5TFuDlqhPKDxLllqEFJCtXl8cxTxNG/3FR4h//qjvx/rRg7
h7xj2Nr9o2RQ3/vNroiKFnx0LcLtEmAHsAU7uNAF80zRnPdVFG0KeJ3hEthoFngrc4jMEqrApA7h
r9rf9IVLPNPopuM+gXMyqLyOLgiwj6qYArDOUoh2pATOB7cnP5DU8hM2cSJbHLPeUvyyBRkZgDie
bu7GHGDgyAqo9JAam4Y+hybp+a7e/cwweFSR/KJ8t4SRD6f1PogESPxqWXAqMEdB/H1v2F9jspXT
elVcYKsp7rEqz7LINRnP57CjWX6P3yZ818PjGIeonKZu78iA4tgGjXUrr5kEY2qUXqHbA0jp3Ion
vcJkipg82CxuiLbD6JdtxbCKpMiueqwy+VwEcuzAsWxk25rWfZOGHgsAOpyMYaNVzoBmdLrmGd69
+pLPpAs8Wbv4df/li4hrw83SSPYcXdQ5aArGYCR7Zw53Kiil4aRXkOZ0kXax7IFLBdeXFD9y01WB
3XlrE1s/ybBKuZGUy7ULtoFbgRF6ye59+Rv1yNOYjBhQgmcVuzHH5u4lphemN7gpn8EoaRAEZo8q
4nM/bS2/BIm1TL/nxLxWjU+SN/x9QSdJJ22lSAFesyafKtZsgBnyPYmNIudBpewDCv35lP2sbCy1
Lu/ewye588nSl8fWTXDHwB9W1ENfuciozy8N/o2YBErLJUvjmGxB4Y/XdVGVLc3pF9XnM1Ds0Xb0
eUBCXNQTzyIx/LFZfs8FCYL/rsTzyzMz58IIphRGn2b/+D/mcbz0wv0vps8+Spa9sUX+vW70bJEt
wEZJ+E34d1M6HP0P3n22x81I8nBJIgQFp1ikxdHp2ytD5BTbqU13SzFwazPg4UekS6KIYCqK0lEn
3zQ8vtIfCT7PXLUmZTUY85MypTikKbuXm/aie37QODoykZzhEF7BgIs78DE00I0AQtdwyvw+keyW
E8kD7OV7IIoqssoEjJmFrLyoVy/mM3/+zA72NNQeRXMspnnWvhlDCsRhmZbMdtMca6WYvJeVhZWA
LBJIrzNrZ/jxVppSs0hH+lk0eD82LnWOt8oDcTeLMRC3HFcG2f5+7549U76DkqbNtYQY0ZIYcOGO
7XOPJcFehxBrm7o+OplOp3SdwXdIa4D8cO5yd4YcP5/rTPrTbXuleehaP1AKQsKtpVraMf8Ohniy
jmo06jvMcSR2ufcjsIroN5QatXmDyDr0gQDLIjbgz1VRbCsiDZeUNt0mldzzqlQCSSExo2HFAIgv
J69dXqCuS3ks17jbYkIw8noUBDTxPmrhlvRaBKsy82ZzhO9xj8xGHrR28c24ny1f5SuSPve/yIed
9LXFUCL3lxyRwDMydMaAwX2WGRNEcvjlnEw6bVTHtnRtiAaCLBc7+Di0D3NyY2byUBOcw6cZolmP
VeYc4j7rQtI37x0QsauoT279uo7rSlp1JLo9U1Tq5i5fCFIZ4KCrWUGIZ8h2gS+ADVM1hIy458eO
Xbhq2rGM36bCY4PS/27J+VHE79jk8mJnvgq3PTxWpOkxNhL6MQ3ueVGUiWIQBHzcSOWFgsQ0Betk
VpzwEnkF9zgaKgRonVrLNH0Yh9oCkr4yo0lzcANx9wQ/9NHQwPZywdEd2R08ZnwYaLbFj1Bt5o5E
ALdbT2bIXbC5iVPDGKlPZSfSQrwxDxEwwKR5FX+QCZYHkZi9DepxnyBlRonaE32nPgAHjsnv0X4E
Wfetgrdisw2Rwe//BclwLUcWzKRQns+IEk3K0cSEm1N4Fyd2lXInvkj2EoMAm3LqrzzurvMzOsNK
btJfjzS2krC43CmjJ66tw4mg0Dchg9jHoSLSW/7D2jYbs9mBNitq9zu2KHOHzrJ+AlfaCvaupcnp
3zfC9FH+482+9ZKKIoThm9zXB3KSFKikNu+4hc0mACXWebnDxLIwO4HYZxTubbQdpkafkEHbXyiS
iWTaG1sXkECO3YFanBBt1cVy80VgCDvqOKhZN/MXhsTtVUHj5wQWP6jWxv/O8jlAANqG1+unP2L/
c1Iz5tzgrRf2NYrg59lYJqgTbsLtYV/qI4+24AB2orGVQSVXZXL+Wy3hdMbymztK205ppnfwH6qq
YZjjOaofj+JrWyL7F9lpVFWb5Ns/LlsCZrd8Y7WLgPZOcBGWB6ByvX56WZcK50SKaWFoeDFwynR8
057GvzOWfgHm13zcLboIWrgLccLtXU4SPhl6Yh5nJ8iZChc2Z5hGqVGok2YUCpkAQWreKPC1Ngs+
9coMyBDaxE+65vAPm/AOnVOKv6mUMzmlmX2NkXz1qFBHXqvOG6NLAzVCCLQ4Rqc1d2QnxnVgY+Kh
YrxHszTXKFHhqB24tQW1p0ZdNEA9oHdKPj3IE/n2URE6ldthBGXxH+iWrT2qQdf/GZ4Q0ycaNJPW
fVAlUonqM1HYP3rSSYMS4qCDg6iGF+cusJj8WwTC8jirv8/e4iA4R3tDhXuru3EkafZRxwF5iWvr
J/TtgwdXlM9f/ehaFOsmyPmtxfiGZv3WtskkEJw3wNamJzOmjMEfR7CekOBNkv+oHGdM8tOOp5xi
QAoAeQhA8rf3UigicOpEhzVb7/JbefcTuqpm+uTaeOBxhhgOWMpCT7Hbhk5b+HuwGiqKTA5ksCxZ
G2DKDwDuSVK61b+EjO7LnEmqhSXr9/tCIc2uBBP/I3mi+PdkCWNoM3fWIuFI1Iu1VJXaFPqU6lj4
dTTb4/UtBtQZ3K/aB42d10Zk6AVXE4/J9iBlipvyRbRj87ks1qEuJPCXvhGkAna+JUmq0pgSuUGL
4g6CmENiadJgcV7v4mFUM5odq1LZA6F14fe2Hv5x7xkkHA+aMXEJgyigUqvDtYBhsgdcN5UwiSZK
1SIokaQsikK1e7z1RyOxUjNkyHdPcrQ0BjE3SavLt0z4J64/Xhhg9pfdlDQEj18bB4KWlnDVPCBq
X2Ph0+FCleapbWwkjnjiV8UtkQGcHMneFzaWAkOxF/4Y+owVd6zsAZTLZ5If0AsVACmsE2dAsCWw
WiVTZ56uV32W54UJBXhKfOxKrU9v/eA1pdZ1Y5ikg+wK8C/USYGO7g2YRJvaNRvNMgZS7HaTthxQ
HAUebjJkXMfbp0uDBSmQUruVOzhpVPoGB1vOy4J2Z+O0kUH3IqKxs/Pu4ojmAHXwp9ubmEYW5hAG
WnEvZ3XN1xGb1110UBdjvjKeAop6LLayOF2rhqYpyCy+5315xvSFago6u+RInTewYoKNh/OwlvYT
BqkAzimDieOa889/A54UGbaczaOtw4Iqia08RtNSnrov8nleYgMPf0AWK8oUe5W3E/O+jRPhF+Iw
uh5Mm4KWIXCIkYGw9y/1+AOqvdq1JbKDnnbvQQSAImoGww6Obt0vJgPb92l1XFryypbNleOgwmVV
yhFPQEyInXZf6++aPyB83Td96rsFlMudQzwu3orEOhYIoAw8DkfRrLhH82PbptubQEiOEdlc6xOu
oHHEwOoG818OfAUCyOtCK47JWWDYV+rhrhCwRIZ0TjPJDwuiwtCd5WOpxnvkerbEngmRKF5yeB2x
VxnPzbcEDSvWP5ZazGtvw9ikhrKVIK5C/x1a4sjmRf0uWqXB/JcnYcbmATddE5uGnMRda+rq/jQb
8TuoGftyjCt0G0cif9XRo7e1yNWFGJJ8vSgfvx99ldNu/hHoEKAfaKCQ0EexJUqi0eFO3JrIj1zb
8gGe5yQJqbqLk73Ec+ZfVolPnTCoYXtPqjfXbTol+xaZllh6uKUur1dYJSkACxn8VL9QmU77V7oF
2410TabyMHXeth2+/dcVwP2LPuYodjVWzQanZuTkReIwQmcb9AYvWpdj3JpFjO0x2SiBQsTybbNJ
PAH0Myc+1obukLG35iOXm0BYwn0tSYt8VBErMDlSJaIEZSLa/lEDqEH3pBGkscV06WABRnmoqXKU
V8MwbfL5e5VVj2+s/0SkiunqIMwDZtOCbeJnfUn7Em3AwYhUXyFpW9wlQ3X79VBgTn3iV1jZyzg5
M/dbsXdZwQpvEPT3jQZWYwuizzRbh3uND6uSIQqdbz+qoxH3MkcZzTtbZ6JU7tjyLOL4B+7NLsJx
GGEAs9nIVAf1wt8HgPilM/tZ+uBTdwJHo7kvYFG54tgFgoqtx1RDyL7YaKQ7RHLFT3tC+H43LlPT
NwcQhGaVJ/p3/rRcQwxoeX3A7aVYX4fQG5Wgfn1J4MgxDvvtWxlLgvqhtfPFwewIOY1YF6EjfScT
81nomhzTSY5kg3VZHxrxIZATPEJIBG8CXFQKa+3+d8HtXL42niw7TEMZ3IAqXfM+QtpUXM7Msrrd
sEVFEnpvG7RplJwgWXzDXjFodT6OmtpFdzNwCtomGCGWEm1m95nLT4ft7leX0pCLMG4esdK2o/FP
ADs6ipOj+4oa1JZdvh6VdKfyQNVti2flgqg0brUDyFGKPXUcjHAiIxY2Y0P8N3nhHJE/Hi43IiUd
/2m7PPH4rPtmmTdYuR4POwKXvBho6QGe6vpcF/uZS2KQaZhqn8nskoAFWbsjYuIRHBzdbhL2dsoE
lQTawZufRTNsiNd2+KsFgWqIbglqVyNjgIcZy1kPraOQaqILD6gmoRUXXUtyVMPmCE4Xthmd47Ia
YcPfnBVzKZzYRZ9AD7mxfvCrHCQu45QfECBULxgx3SEtONUUvnTh4i/q8XaYTXNB4iRUJJpxhsYi
x9NvTeY9Oxpzk5BSOKCmWJ2ltNZSw9IAPd1F66G4xNkYP7/JyR/D9CkUdETNj3mM0x1aRsnE2MQ6
Ol3ap2O0sQcFoowJJyIdlJ6mutQmF3XaXabgoL2lR0BAdQ/PdOythqbHyVLbkJkzDRwRsY3nTsR6
3BZrAT/X6GiSTOJ0f/neqKmTvJkaofWBmFM8Wu6PDKAzkhUfJ2VMIuXGeqnbvMtaZqQvyle4gyzo
Dx6QxamYCw5tmRdgw/qWSnjLqUooJ314koHv1j5cAsg9GmcA4Ez/4mUAzSZTSUZ/Ruw2j6q/1jFr
y/6DTjg4sEOP4l2f9byzBSYQMf0H2rXGQCE2NQp/HecaSdVzcVH34up6OdRJsnuD8eSD3lMw1WKo
vlmMBmfTLlz2L+BEoBn8BAeFUijvdjsXeox+NnkVdX0pmL95AndSxlkbSGDH7g4ryy1dkGlz1no6
VKKr2GAeY9aDfTKiUkTwy4Sc6gRyokG09o7czNF/bogRvwKiSbTCUbUgYRuV/nJUS864E9fwiY18
OepEe5ONZGUZWh3UOt6r5S/sd4k/0G3yeT8qU3qkpLXw2+eoNkFe27T2zt+U3opKTM57VorcGAvF
vb1I5cTSw7dwBjiG9e6++dMF0v6l1ysG4GpZSo0ZSwPTqjmdGtshBTP8JIyckSqVAIyAirwA+7bk
n3v3WIojubnUKTMxg1qPQGwRyjuAxRWBh/Z/kVpqmrbGoxKsykTZxyg0z+baN6Tg7NBiI1sZPrL4
l9qUPFnaYmIamP3g7anx+gW8OnxFDknm82usd4J+T2lq3pQ1/szZQvPpEDdudycMLB5Ek4ztS4iU
WcU7tShJfk/Sh/DQArYCYoQ5ZQCB+x4+ob9CAzymJqwSFC/1gS75eeUTfIIsZ11eXfd6XYFyeGhh
jWHqthxp2dQHgW+yvjR1gyNMst6v8uCpM7V1d+QnZ73FoMkR+rvNQzn2bj8HOc9fZ8Mc2dkz3Kdw
+qWiDzKEnP8Bu2TPi9ExO6arppaRWFGfCxZZROLcvf+8RCiCIGD+QnEIKk01EU4ncFyp/8wK1BT3
Fus0w6R8m+Wco1bO2gREZFrhN75kngPloVUv39SKDRVH8yE07YtGtlxLhaHLJMp32/0DA23kHqd7
opTjI4c/u1Latcg/5knsj5Fa9rkVVNPd8afzT3QWVvhlqK3JImpAtFAHQ5xDNpcXFvumdBw/o/+z
YctFm7MDJXWViX6zll6YtzeE3ho3UByijklKSoNXhfw0uPSZGrtBkV4JzekbThu2bQrMdSuu00S+
xWcdsp8Z7qjXiLrnzXkRq5Ggs9pvAhCy01cSiTUdsCUtF6eILnBEOuzhkbtic4eqVp5m6JEiWRNr
pu6l8jYuzCeVPpnguEVctsKXOwZvkwCG64Z18llgVr1ketVaCms/MjffZ4OzUQU3dmJVvMYcAJJs
fPC3GpV18MIFy2UpM1pxO5xpPqMXp+aKU99esCIm2rLxmJ08wuAJj0epWy8w0rjbFuI0OCVhT3US
LanV52KbNdhRQ3zkELlIH4RhkSH57P6aiw6PdAl1ovPZhObLn3pAkVBu2ml9taZVJ8/sVIFpdPmb
yBxnxZD1GMtc6RuCQWdheD9/N6MxCyCb7Q76eboLkbn8Okp4dMXoBWiQk0Y+jkzCRzVjfEDvM8xC
4dDTnOoUIS4iqXDKwufVhyws+QxIYxbXpa6aBMjfAd4j4D5uzGGj93EOsb6k1hbU273rBDoobiK7
maimGkvyHbxHlRwEouVqFpS5vgbSroAI/pGDDcg/7Yn3+2TVSthI+xNKFRJhLNvGBKtvSrzpl8ZV
EzTVPmo8PzWeQNiSFBORfRqkp9VxaWZcbKI8I1qgvT3K7xcNQudW7ldCe+A33pMVeNEDbEDAWGqQ
MVXc9WCSyqnJaRmOu8kXQwBABUvMI2rjp4z8i1YDl9umoW0F7iMIYc3I1PEMIwJVDJTzqkQ3MdPM
U95U9EU8U0ya741EeQzFNkyhgPaOuZQoly8mxigHdJp8GSuQlbEhWJgd+pP6z42iekVaf90jUZMA
ShIb+Q1NyXe7x6BfDkh+DYLA1DTGscbLBebN5+X+IfxU2lFlbXFQOh/0PYwTsUMBDEy7JUamvNzg
ZZnBZ4bsx/6yRveST8ComDVA2HWEYgrzxJ+IgbQbJrRkCcfMH50YBaErB6r4fermOfwIlWVFgMBZ
lcoxB6jzONp2SwCEhyfhiUI1oThnHb95N/Cb/qPK2Wq+M5Ej+VvafFKUD9ai5CzveINpEb6H8tR7
uV1jdX437NXbqaJtG8ufK/G0Gjli4vnbKCw05f+RLaF/zkMqzZclmSRZ6h0g479sjCntE/ikJggO
jRcGh0H+Ry0ZahtcBXgf8yPzMgHb2TvmOx0EI0jPhedcIeCXH7OsPso0MtiHRAcCFcXW02L44Ivz
ql6JyXde1ZffjTh7QdZtleTLhGGWusQHcglFMDE3xS+tcuxzf0XGWcU5QeGM513BJSnZpmHYdIgw
z89pRNkyVZzXdiUdb7PHi+MnGei45hl8bIv5zS8+Kii3MedyGX20S2CeISlK+tAwfxEKc3yGWGDy
CC2TLZAn9HAcnW6/N+nK+RmmvIQE3MFs1AeHqvdcwNf0IXupW4VS7VHovb/X+mkV1Li3bFrtOlOG
FFVwznZzEn335wlSSg2ZkhvtpLagnNuAggvRQBLUF7+Ai9R85R5fGcHfjlN75d1hF76ZqZTxngLP
DHNgfmVuDkbhHX5caoByrY7ProtHXePNirGm72Eu0hJOBs+GSfDK6XkrS6D/A/ViCr0LBqZf3R7e
T4xJosibnGBc9hqBskEOXdPc/eIR8Wx4pYGzcj4o1WJDMtDy0Iu13nzNJFVb2t2O9ZxQk+KTeuSM
tP62qrccf+w6tfmELtJi3sAD3NA646i2OS+NazGDd6I3oK8YniPV/pI6a6aplCbWZ9NDh7Kf1BGx
hXa8tVHlqG0ZxjTKNT4JdmJoCot+2y/a/3r7xl5xPoOzsxHIB+chdSMv6NK8+9QAEfIGxz4XFfl4
guF9JhFSy1GYfIPkZ/fZ8newQt/wHklZgd4N5LEf/KUWhpbnf6QAWYgUcbBC/b7sp9XIq86ERFJS
vfnFLrDj5lolN3LMV+54XlwnMxfxE2rK21ETZbkqwyzXfTzYoIKY+VkySgsgyHIJ/vDbiXSIGNQK
kZhzImmaheHT8cZZc/fWi4hJK9QpuVKozJhxqnpchp5CJuhqdovsOrT4KPtWc5qmMr+R4P+TudWW
ca7MfFv1dJx0qsaqW07zE22hYFXGoXZWDOJXjF8fJgAfnBx9MaffJmJ4KwzMSuLoMA5aZ0QX7Dk4
CZInfNMpTEU0yyEHXWDhSd4IONpVJiq/20I5sv00eDa9AaAxw973pjttzX+RtZNvdxkZmptN7rWS
biGJSJCFb/irr+6cBQdZ7/d895OdJzzu8RHl881f7Ol6ypPMrABAXYpBpLRjtxMPzV3cqQKG1pSL
reQDb0fhEBqfGtCSwxE3VVsOIR5ZYKI+3TCJQOAekT4cfhqc/7J5AloGArX78Pq4CTqfmVf8iIBk
69Xl0t72HZOi3UCnGc1a0lhHk9cQsjUOdpRQE1yB4J8BVOVmdI2rj6JKhV0fZfWSEDxndDfacal4
U+lErwVxdzNSe6/eTvc0st+lcMvtjHotqMZ3/DdbKJy3z7OHONAZ86Po6hq56Q+ubLysWHpt6yWf
e1GOL47ZWgr/RYnjaxfyq9eGVjMQx2cHv5QZp7ERNvPkeRumZf2W0OBFEveVaUaB14d9Zr6cE5mR
JGYdn3hqgSuHvrpK0g+2EPHpakrliQXEmb9VGrGZ3deXzaAJ4ffits0oqs3y0TNt+F6t+aNehVcD
qU9Td9eON8dYQlXH1wC5eI+nWbKKWjahTY8MAY0RclYlZxKQ2kCUzTZ8iOBwhs7Ilvs0PwEl5KHL
bxAN3AgCpCwRGAYEc2wUNXOtSKFO/sv4p17zCFmhOo+A4C+mFGvENZN4Qr/yXo4scygEoAGzGydB
rKRsV0LTSCmhZUFkR6a0w4Oz/kGg18nKRvu4LIwOBDjrKn+ZwlrAlCGihJ1uvg8LdQbFnvUvALDL
sQdnqLcphbN/YRxXzn0MyveIEKDjKc7oGwbbCT8fAsimSUnRJHl4X64dC8y4pOI95xcxceZLlhvD
XVjAK00hY0bAa7F+u0RbatfVEefDWlK/6sK62scrwgWXXYorcZWUCCKgG7a56NbzUTiNNp1E+6zh
CAbAp+UoqIxbsjx8OP6215m8SyLbi0EbMDRfh2UTPUDzkmdVW2J8+OqBY5jv+FqI59pIYLbx9bb4
u976n1dQDkjoLUfH07bd9Z76j0Zhcfhle8cbey0I6PvZeWImEJipG/9OUFWv/oUQAPTpWA3GRhvS
N31OhUdpplzlZJLLu3eT5St93boZpGNJIP/r1tGeLTDDXm9scWJEpin0XF9kbdT6pDalFyOeKg1b
KLruuxxPnEIHl/tfLcJiW7KbZv2iilwrO/eygQMHWBUhqhM90N4SuiXtF/xvcsCiOOw4CFu03hPO
2C3lZS1fOAcLJ4JaLC9L5PiTWdLBH2o2mCKCEXn+cCSzRo51ssOC9sr5D/w+xy9L4vX26oCtoD6I
3C60fIV50mJzoeA+yfZpMeMO3XkjvpmCMXJc8tAufTcWlaRYfTUUipvXjev3oGBcxgXRyGA2EdbU
AZGq7JGOnS0K2HKoXi1pwZUXsplzFU+uflP2ttA8gsNEj8arvo7ot3HP8btig8W3GA9pFsjsRbnV
IvrSeowMK0X0zp/8CeN6+kCCF5Ek1bo9zZiWj7pzdctVJ6IazvnuQIeUIzWkWwopO9KOzaa6kJ6l
0ENkI+Ik4jvqgBge2sNQ8hyFxzmM63aCxEAAqRCFIn1DDQH/zcHweqN+DCA4Pl3jbHLakaj8JRy2
gbBnBpa16sNY/SJVbn06Kv8z7euHaSOxhjnqzNzvKw2dWgp/MuIxWzLQFM5Wfh4FuIa+l8LoaYf4
xDqEw94SzE8AZYjcr4NdAszxVEiA6xmDDP9vDX0mAIfd8GWGFhcRfBsce4DZQcQsYwxcvaSw6VCB
CMsP4bbq2bg2tCE4uxldnRNyYhdRJ9ZmOaSBPun3X/AivpnmdQvZtCqn12n0xwNC63RmDQ8ZaK5M
5r3oo0ru2kQYFboFXStNqtSk7zJC/ffAe3H9WXM6c3h5D59kGdusZGtzrf1cA0yj3Lb0+8x9rYWS
rtmnX2dCsQnZZUMtMXdamwWuRqcL/6q9/+8cYXB/7OugAKtQPwW/31cjiRq967rHNOpaLUYQ9Bvu
3YPf2WE5Aa86c57c8PWCDHqaFVJhPenKf/XxxYmAwZeFxUt7iY9zb3KUYcHGjPT/3IEWJlIxQOrA
rbtXRPzsBX5QQuH4v/akFEv2fWCmLJntaQGrnSBn+h2kBPZxLxLb5fcSKqmRYi/WzPICEj5pX7XI
xiHGFxpMM/XWs2VPIw1qC9LwLwvJi4JQ30fXjtyx+KxFHLpA7P2mJ9XK7vslG2RzHVLj4b+DgID8
q+ZnON782cL/XaH5Bu5vILcOynZJ0aE9AQb8Hjw9cmrnE7Fc/XPwVKU/xuvKg/WY8uMZzZGgttBj
a8tVglyY4/Ctj74unPmcaJe8OV9WeSmDIwpkafKFy3Nb0O2XS0gTmKNoCzvh4bEnRMycu9uj8V4W
NK4NUif0GL/NPaAVRik5Ks7ISh2n9c6L/L7aldaIRoCHysXTkL16J/1rJsoKpEhd9zosr+dVXvuI
LNnivhqiATrokKpKbfKQJT86KmJ6RA0OxuUBad74q1ylPBPwnrVX9aAkkzpsmAujjhKwHhEXvvfL
G8oLEg+Vb7a+K8s3NlA0cYMFB4U3qYN9YMDhH8UCLPxDWmY7LMN6CZ5evovmqhFaTykChrqoWVsr
m2gRgk1MzJbhJR6Sf3NIMSrsk9oSaOw8a+QLd6W/AxxI7JbnEgUS2t/vjaBclFSK4W6XAAo2w+3A
JwfsUGb3u1DjMcQSBj+7sPkkbpDKaYbP/xtd794iRThmWJKd+3LmKaO8zdo1CCNtVQiET5qUyxN1
Px/UbxjTPL/Yje/u9NunWBT9RYbh76lEbM86/3kr+XmETGHjJMXukbEyXByepvPSjkUGjXqXh3R3
VXu15+hfbbLHpLztyUGNTKm1ERirv6ppkge+eJyiUtXzdQHljpfMbiLiGtw61D1S3P+lVeIezkn6
bErDZpIO53Kp5EYru9jAHfCJcHyg/KH9Rl1AeVHihJW4LyGDUJp30Gc4iE0Y4v0ZZHj/r19KGym7
MMcP7dOWW7u6I+bksANcdr2jTgm4zcoTEuadDCh+zdUH+j0HSB9yJhtWZrzJ5vNRg/PcXoNE1mcC
S3y09HDgix15uzzjzyPl/Zf1oXJTldfyVmO09MxAodAdZADFOgJvdI1puB9f9cm0KM2Yxd0oC/LR
OlCr89IC5bzcNx60PmmXIeaXR84V8B5s8j1xU7NP7F/ECSl1k+PudXVSrv5QD/yUG76GW7MIaESE
BFVvXouMOireT4m0zfgwIAmHgzhU1EesKqzVIPQB6UYGl4G5SpLEdvP8cnq+fVCZ42Gc5CRuU3iZ
skqJqWd2++MFOz8iD6XVz+9MlVObrlp70vDIFHNwRU6FyNQ6BWnhqyBkJs4nIAMg2dOrRDzb6ufn
TQnLuy46Fn4ZryuFELwGYEFonnab0g/gg+A9ZSwgj0Tp/tzxr/JycoLySVXU2V1Qd1iCIAYhHMWA
ftdOtrxXADjXCkXAL7jJvVM2DFDq1Kwq3FKN535qGI8JXIZiVlBAuhvnuTigbFw3Ps3+u7o9u8wU
S43/3DC7jXhUoeQ/UAFkl42vgzyP32Pf9kEnWk5eRdTnaR9VUVO1QmbtsJTym2H75ejX+i7vif8G
6nGRQUWojy2gQSNDhW1k1duRhdA+oLm/COaNhrWVurjqJr5Rw+eBHY5hHZB0ICdegvjehQEeXGHx
jnAMV/mC3XNz4DidNSrg+AuuxZk+h9zm1OY9HHLMbylN/AkxZZ6MbduARK1+zSpoGAB/0TmpSFgU
72kelzPjswQSZDqZWl7hgVqju99wVJyjjv2WbdaAMWqX8qRWcQoVs6xeCIjnDhvtcIIHwyEXmeuR
ER88/43/UldLKLxtmHYmVZYxBKQNR7mMcWYO4wodSX/kqEYIiuIvxCIfT5KIilCCwEYPQGiClG8u
D4eQcu/m9lJLBwgdsjlsN5OdRjUzEqxu1EC3PSRxI9p3VmruPnZMwOBCrhMFFIPNNDNYbGx3PbAg
7sHKGIInqqrIe49GF+/w3XyBhHZcRuwONah7uiHQaiJDbcIsKRoTxoZ+LoKE01wfdo7DTVmAGp6r
kvF6u/hdQuD8gPZTAgVBEUVvCR/DqhYgueLZkI1nyEopJOBo+iz5CR0cgqQRMd3jVyt7VfhrncTt
knPfGSesGZlpFktb43CkM6XsJ7wZ1C4T+t68+Uam6uwDm7fyOPASxEPQmtEx/IM3syeOKlzgRo06
tuA7hwxGclmVY/0IcOg6yU/J3AOAzpCERaSMEgc6hiqEJyVqA7bo+rmCt6QCtewbZ0kZNWAWx1qG
a3skI2X8w9tNjmuEOj8Srn4JhojMgLXO7pZu/CZBAsgwJ03GZyS0PLhGzZmC1UroS35sGa10dT0q
k4N6sK2Txal3bdbxnUkVEKCiVJDYTurMDmaLxBsvkCH3Cc+G73DrZpjHL5g564rQYWiR4xy6vSRj
B0f7kE0TFbaJntXJc8gNuWPx7reLsxb/RYpKj+6ES78w2FhKq2PtBuJkDxuOWfOdmWBbLVjz3H5p
UyUqMHEQcED4aWoUYep1U+O9j9SguaVVV5swCoogtMYWzNnyKdYMHDtWUEjqqIwSzo+fks1OGQ9u
vGBGhi7FJ/qm8jEw3YZYBhwqaV7Jq2/629lMZkRqSrPOcwngRWjHsxOyVuKPR/B312dfKABCEkfk
6esYqqfXnHgpx0KLwNaD72n+Z4kcivNBt43wjl78NuP+B9Q9PKjjOVpcxDVZ3a8MnR0v/6rxM+vt
p2H1RqvHcnfM3TrWUmIotmAf9eB3tF4QAYE+5JmWp3lI101caU+IYe4sOraXLucmi7rvKw9qQo5Q
eaFO9q0vmBTnEyihnETYY3g1W7kFoXXafyYgn3d7ClId11Bd800H0FqJQi0LBzUfwjN1mP7tnlSU
BahrPSIphVyjEE6xXHJlq76kuforc1CNJKedkt+Lv82nnm1MVWatVFpAXfwNO5SjXSzKn3fdXehu
KIZ2cBOcdUtOyWf9gD/wbxEUeblPHQj3/6Jg5pKL73lMzsTLqEIo+Fy8Pfqm5TDCmVtQhLiIO68U
L2PJvp7gjPPb2XQt7f5duaD+sAIuaikFxzbAsj6Y6QFaoUPQnL+6B7b+tgZeMwkEOMhKlHbRSJAh
GmsBrPenvA/SdPgCV6d9HHCqj+/6GFpIe2/0pD+/7hIJH9dCJRuDeXRYA38f64mzcE1FOshOge9q
OvAsUnOqwZdvup/C2LJVI2H+CaXVDlv897HxuBVwowXi+r62wUpQWInqRAQqueoyFQU5h/18bue4
npoyK7HQmWvxBeerwWgng+7iTWGqn70s/c9VQqBr68NtuDq/sBjG8EhbI3rENCmyiuGfkkMLm/Ae
YXnRGtyjGL9BuZutFDK0Yn5Wz9vVoq2R9W0tULzHlxMHiQakaomwh9tYa0Nv3s6REHGjdDYwDdgS
8z8WhVv46pvnfoDZiqrDWMjJsVUlYu1r+HC7dIt0R87IgWYAg1CM05dphZ6Pts0e2xlrY8hKpwE+
jsbE+Qxyfm05TQ3cfxorAkAu2lCTBkuiWi+MOBY1GH2QVc/mPP12sJ563LuNZO11B4esTFpJnIAv
yw9WW36k+MEZsqryNUuI6RsmEDQ9x6pddL0DWrtgFUoARLhISCDewClOTFv4wBS0LUPOd5rn4ccC
QzWzuo8ETtaUPqecvrDtSiC7NXYOdUJEPYD2UQWAfsqe33BW95AGWFdHK+UJGqU6hRj+AqLjUWem
j1qDL82bq+xUB48BWKmFzmzuHdZmK2TWTeNfplyj2JVDSAe2Yty6DketxoUWD7HuxVgm/XyotFEr
XMkg+LWAPooFvoECj7yJl1mZlyspN+sQOgsKsgeiW4sS6cpp6paWY+ekBN6ENzV8bBc8+9MQ+/PR
d1LzZ6c1ZmhPD/A2NmBkKZDn6kDOtVgSnHQxvz1NGV2/MatIjzEBJD/cdyOEwg73nEpol4WOMT+t
IZs5tripq1dhGpubKbOWGmR1cOzDQqdgZw+f/01d7zURmOw5sPIxF7Qx2qHk5JBlYZVwBy8Y6C6Y
vLTg3mmyyDFnWxDjacarynldhHkjmeAClMe81qFuBzzvl/o5M41lFcEbwdM7OxTjq++R5snm2vp5
zJn/jxGWeBlJFKcTOKHExlr4EK7ODyRN6FL+ODTZKgI9UOlH4o5DUlSedNlLRebGROWe71cMnbOq
5YQY6ETE3uom3KmHxhPnICZfr1QgD3Bky+yfoBDxMat99iUlXjb/8l6opHQAJ4H69xQg8ifoh35Z
G6aFsW1r/WGnzAIBAnVhdVNY+feZdj7hsFOUDKcx6YPQJppqzNz+CGYMygzkpnPyl7hPRJDlBvuz
u92qCpNSuuM6NdSdOrgnyasxLjxzjjpDl4W0bLtYwkkcuwZrW7etqyWk5IEii9zLzxzaKpkhbLSn
P6s9OFcv26dphw6cKC78doXlwO84mlRI8jmW2aCPbvSGWRsaY6VNnZCymK+T7YfaxfnEFP1PUZSs
WU+AjoRyvh3mkCfs3OoGN0r1O0iOhszgTxJstICFpYFxB/cdu7oRaY5lx5nmmZjVMdAln9h4DHDB
jH8XFUb+/TBmj+BVLoeN9zFLYi0NQwN6Ckd7trziIXiK9ktCcPfPFFVwZvbePpks6FFB8cdtrPNg
j49ImXrcVj6NRlQH7IMbDAffYC4cKLJ7qhsqSicv7IJAaprE5k9yqWxxuuVRVXv+Kymn5kZ8tU39
0phECvvxOw/VO4tuH9fAMYZ6F7TFG+ayREdozxXQMdpCsjCCHGc4r7mCcZfyz5IBCqT4XjZy/Cpv
8mO0cS1SSnXEynS1N7peT/LunjC+7liwDm0ACIh7dDIfNlA/vRjmdLKYT7A8PGWdEazENgrl3okF
4iGa+TDW844ISFQX6Yl3rJqguBCV+BNqG9QxX1Mz5Osjk+PUwthBixiQAXMol5tOUN+SHoe5621j
nkW7hlVppTxVWGT8I12FrL+eU0pfdn9WvZivfXiblwITDE/GNyGmdE6QxQtuHzebNgI54nTp4epF
IW+K06D9y3pyBPsv6DVQxNCSW/CzWLMei+XIcRxX6ew/aiA+HihpayiwBy8Q4YZ/1qwqA1ybpDBT
p6njbr/c7SvOiac7kvLrF21iglzV4aq/shTFObC0lfDUISODsnXaUSPnrM9r82ZOBd/Jd+UEhiT8
krxwOgJofF0kBhCrPFq+Mu+r4LNpGz4bSPAzrcgmDYQT/T6swf5TDoPCtHyETtCsfUOYR/mfHhnq
2L94H4rpysQDEZ57T06sRlpFApz18Nnl6P0AeUQdlAIKwIrjfzMmaQkUwVHIWc9zO7tgAxD60Y7K
F6cqP2L8BjJsDhAEWok4xZoKjZLrGgowBHZ49ZbipThoRSWJmo40S6uy7Ad4+plHkgxOzkZsSRZC
8btk0ssangHbhtzNGF5/ZHE7Ese7RrWb1vQlAfKKmCGQ+KzoKwp622FrnsCwJh17Qugwsr+EhUVL
SO+ZbopSr6BInW41LYkf6ff1CUZD6UjeWDwUWw0nTG701MW1pf3/MkwBSSYKRZooaKUQCBc0p3nZ
FR3ExXw6anJq9KlIRaWOWWde3k4V4EIe3z0fsDNzMLDmPY77HSKb9+x0WLzMqClfQsnG2zkUxl+E
8JxdKOiEMoLO937qwfZa8kP5TrxawfcN/151vfCQvs7//WY4MThm/JEIHrXQSnBOOvVPWkW/Hwcf
j5AkBNY3OVpoYWbww/fkf6bbqINDjr54KobJr+QLcviBEqZ4DzEWjA3BeH3m0ON+lwGfaEhvoYcA
o6zG2bs7hUGrxtOd5QUiDhpvWwhiLPJbtMUvbpzsupftldexxm2UKvJpE+SfXmwkP3ygbUKKFm5u
x4UbIaTlxUSlHi5mthPPR4w3xNDUB+/XXrQ9i7p0FBCjp1thXAy5VFCYKd9gzrEXKUEryjZZkg2w
q01Ra9g0U97R/dt/oaYXYknagFx/zfRNrSAX5vD2wc9/gw7iHwFbC9AMfR52dw33EoIfZJ8/vzH0
WF3BHOqXFTIzD9AzXOXH6swb3N5+cBfy8QtJKlSPQOygMrgjHSzkC9ivcenZ0W3i/M3+JSU+fyv4
geNNq9W8ZCcgn1FMIrPhBH5t9FQG5HyHNr4tcZ8vpBhxiWwGHClRr4yqo+rxSYCd/6gkGD61aTKH
KA8kWeTzAqEqVaNKHzKZOxO8n8+HJQtj39g6SieqWPHtVLyZ0Mx+0AzdN7+IJmSE4tf1oTQMb3Kp
5TO2sOWigHtpE/EHmkiJrlYFWRgsx5eEDdQMVY3H/Xkd1BrmnwNUsFU39+NOk6xl/uhgaGi+/QfV
27ReGru3KzF8uW9RQI9knQwTlyl8bFm1GQAne3EX0fCj3RByorOCvKzE3X5jI99vYayyHN8hUTJp
UMO89fJb4eNxuJgdyWOAmrJqpdcMwRqkt1CfKefUp9X0jsh10zMPwZvS1xKXdbbmiRvHtibQSMJS
igL9uPP+BWHkfPchXI6/qnFvTSeDJ6xFq4LhJ6ULLINj8W3md+GBFNRUJu+zxF+ln++Dh+SQ8Ush
lUEuuXPAfMIE6gj6iwuzycCg1gUEz0eD88+Ai9a3q77vwsoBqOd90x3ffYbTFw0iBMetllW0jP18
zIr9lO566PRvihd2lgkGg4mn/sNDOSAqqEU6U5emvhnhonj2SWcWrw4+y2SuxmedgzJOPeoaFS0l
s+aZrn569/OQ7+NPUoOzEoDazSdaM6ithLAGUiV0bn9Belca1nSAwMGWeh4QLGHTCNT85aHU/oxo
Ak8bp7VKe+RPtjkGQpCxzwvbdKIhzY7RpToCEzQ1v4Ni4CFgpWBu66PifllLbsRwRd+g8pJlaBod
HAIwGrzH7Sn9sLNYwNtwYdQ7gf4Jtl8iXakSBFIhgtXTjCJiQNdWYGBSgorb0m0a3XXMNipXXI0S
MGBlOxRj5UD2yk+yc9uwhF7mKDkOo/RaJW4Flk3Dg3iud31o/wJePVc9UWzDyPLqBczHLYV7+z+x
bBYgaAYsAv+dHf4+0AMXwEslYHb8x82xRl5nBRc0Cj3nY6g1ontmJQtwqbfK6edbqrd3I+fBOTn6
ajD9OG7APxV++IbeOL7fPtdc6sT0TVQD/0663W12tjNA8AionoCI9dlvWcORcdn1OttzjX+O6I+4
luqxIMdNMn3+6DHXvHyT7i7okKRIQiR60nY3ohmudD+DNtbQrfvLuezO70AAPFEg6MKIitI4VxWW
kc1F96pOh50mChGvQe1WuXkUF9BsiOWY6/KIHJuRwERLP9endJRTSccIdVEG0x2cd8DBpyVVBzP6
tYHBOXI3i17BYvEMrjR0Do5TODaw+JQ8KIt5/RWez0h1mJYowVErXDOpElskYvwlZdk/p6DZWS7a
1flK8T8GHtKO5iYZogxYu4czbf9GrmP9NaWXa7axFMxmmHCrOz4X8/nGjKQMp2I8rsQq3WyXVRlR
tiBm+pQR9faAfd+CdjK4c8HMaf6q7WHyFAlxv/pkcawX0kkXqEL4kAUXOCT9+WdYESxz+V2pw4SP
x+JqAc5tC4MV5cMfsSDi/f0MuS86UsXMFT3oZiViMWwBeWKU/Re3BljjB8vxda7ylh0hU+x236q1
1ZRc49HLC+7mvj2gtjt8pwey1Y9qrEydZEWDBZ49yoswwb9qfy4CLUcekPFo2hdckOCchVKt2fXH
4VzWzbDLlRCGHqwUCQ60cmBYNoMUibNnAD2ziWPusCcJGlNJVhWLS24dVVzWvkVkIebhBcWvTYxl
tIOoW2QB4zAwYl9/cZM6eg3VtWQHBZDNAIqphWB93IkwV+H++G+8dM+A/1AW6psNnmouiIEWqVyr
h5R0FTOLg2EaZUwose7dRkfgAqmUc1nHfyg9RKCGjY1dSRCpm9NxfwqWk4qSwlu48bYOMVhjCWez
dC+uV/FOzDZFaGazXI9JcfHgYaDd4C9VBk3LAVwher8ilEQBD6UjuzEvBgaFMckBw99n0UuIGdZq
7zshbn8YL1OvB4bHtrmnp0P12pLZbe3yqp34XIhth2z9vgZm2AByL6oarb7ZgJIlwK2audjsXWnx
99beroFHTrV1uQQ58WeRABP4tE+wCrEopqAcGjmlr3WDXph6d/aBqoxepXRKCpq689jStEzT6ihr
T41qh6DMLg0rSK+0k8cx8ktXsfDnPW/o78Qy9UXGaKr6gMCXiONFifOE9wt3twm00mbAfJv4TYUs
OMy2T5l9an8RmWHcu4qTpTn4alVMbnNCMyYBwDe/yfCMYk4xkRtDd1+nYPAb4rqkAeIEd0tmXA4q
ruSOyhLapCIwx341IrfyFLUZlaUWdBM8Zb+U6Td8yorDU/tw6Qym6Per5GOcEwvzNEiU+CjGnum2
70W2OqATDwBa62ewA6AagrCayEcmCGV5qJKK+wtQcCaF/ayTD5Ws1Yg4+wnvrk5CZo9AGWWY5Vbb
x4NABx5ksc0Mp07xpFVBKILJ+EuSg/qENOSF7kN58+Id7XD63azYfl0ypHXCnzu5KOT0lptNTTTd
uFfsYBNaoA5cbPt3gk1f7yZU9RdW0ieTj85ypP9BfpSb98Ts7L+n5u6vMMDoB88dl7o/hYL/puf8
OE5SKXV+7ISjlOniesCmPTO6ieXb+rDoAtOis/aOXa/pylZ6ZOneB1b2DGTOBBu5OkPEHF7P27r8
4FzHwCAGpv/soCo76+VXHAv3yhL9SECKFFZkbeDNm9zriU8NN+zROsAFlaYgPhYvZDVISRqU0Dqf
Vi2EOszZg/dKFqTxwzkOFFTHBOqpm3lkqPpSxPS6XmgbMPEj5Z49RIddVA1ILkKpeQvpMH5ZJUF4
5tUq5FfPkgmtpmNIkYGLSKplCIUMFMIJRyicCRrMbinofJtN1TwB+jHmld4+AxwG7fMgvyJMa1Ow
mGJ5awkymVxYLTidsADKUFPqUZGQINskKv6DFPA4GZnKD3UKfsuz1ElnNyvNg2Qx+dXGCLcx2P+1
Mod2Yi5cEXe9KlF8DXX4IZ7QZ1YCjuKhVQjnFUCa41LlIyT/dmScbf5amwou0rzBwLeUB4mZjEAf
buSNN4HR4gn5MJ50svwXGI37Fyr+EJCmk7jDkqcC5DS3vEv9rcl2aQJquMgGKS/JxsBMj03W+o5l
Y71QyzzEwHWbNUxkaqyZfSHy/+4GWvpZ0qcpADRtKFN9rB/m0wfA3x8f8YCZYkVcAtZWCUSCoC4b
85nQhIzlWywEAD8xD3fELMPS6qO5KYWxc8BpdWrJQWmt9EdNkwMT9FoW1LKKR6TApzbYH3P8kf/2
6fuDFZIzoTMPbAep9TZGCrFoFQO6QgKFkESs/Vl801YS+1G9JazLlIYSoucaTP9GlKEB4elh94LE
Unc3ONDwOY/R5FaFH8W7uIU1PmCtaJHtxEoBD7T+dsEn1WyalxvgL/B8FMhycKxGmvKbmOTluYae
o4WWpPRBlr7fKppcpvpsoFKwrhWi5LVUhVbx+uzSgCsYQFdHtHFHLCrmQg+GDZ2QyRXxY6DyZqkf
Oy1mHJ5lJpeq2qOol/crlefkVRasIVihyThBkfgFhYXh2Cxt+cLvflyDbPIhIEQ4Mmb1EnGKAqzw
VAlgz+6OJ1fZmH//eO/H+VPDFl9pSa8jRxLrpb3YMSs+oIFK011UgF7tb57S94K7BfiLZZ3rCNMq
r6ubLhYE0P27PgbDQw4Xc3JyJU9xoseKWbK0b2lwyzG8Rb/0n+cxwZYDfPSuz5t14azLlMq9ZJ7P
jHMm6sOaL3NUObYsgaJPaFOsL0YVbkJq5f0NxCSKsea7NCcbn+Sz6FxsQISKwZa+RM5VXPxzvoEK
KGOrlUkDCYd+gscsdZVulh0rlstzrejCq2/vPW2EYnI0ll6aUQJdu9+FzcylwYDG+Tg8wr89sgg7
Up63imccOykiVjiAA6SbOZTl3N/q9bVEXx2o7jqesPOPQrR6nSDfOqRDHrmrXHGkGZIzZAb63hQ3
kBFgGDJdK4KU1/84vaSLbIpyx9t78nMVxZnZJIgzUckaprC7dLApBDxm/Wf36HRDQs+ObB/eXTnf
4tvyPxrfXecNoNhdiBl2BrCFjeEp//c1J14GzKAlbks3brSIFlt0uW+p2cRyiO3Kl/JjbYzVctrZ
35ewA/CD0flFlkiFwxKuaQxOu1GTUBIVPUw2nOIvc0Z5geeZ32G8+k5Q/Uso5R59qRNGcGKbQ7T/
du+glp5K1QPp5CVB0A9v5GJbrSCxiABDeRu0OZdfYHc4tM1hpDTnnre5pTuHi3alSL8BKpASv9Kl
HpH72YlHKeqngv1u5pDdKi3HHgm+cNHQLbHIXmWnOl+pr9Wvux2tC+UUEeajXyfMSbL3n5sJji5g
IMbdV33/BFvvf7vfjVxl86HinXBkbL8C01KmzrkQFtwm4A70pdjBlC7h78+KwRXiVv01JbUZ9zNT
/6eAFQcYXzPG4VSwxDykoENNprP35Z7v/nvKKKs/IVc0Q07vkuQwTuxcHtdPgw4RPfuEOpNDAyVh
0S0cUiq1EZL15M60Irn+plDh/OUxJJ39XkkT7CVDkV3xl/hvsWzXEaeZgFzXA4Tiy/d2kY+0F+Wr
3CcTqFkd97VEJVtAhh/BmALzL0uASafpGe3NfGEpEalY1lDsn7YDCOpqZ98w06/S72vmuEHp1lsB
42uLW4ypgqz/Mvj230SQL4nfIdUpw4O3xV4V5NfH+K636/ZeQvGJYQZwtyX8+e8qb3o/gl6Rh5GA
ED3bLMIlF3v6saWTq8s9EZaNAM9WJiGWHXE4gliXt8LArkPNOXxdXxqebTHEXeViaE3Yqa7bcaJt
zOAN8FSUP9xgKj5yJuNVzB7vWMFQfh51VoHy8pRPDQt0bzuM53B6EnC5zDSmMHy7dDLimI9rrg3O
5phJdoz5gZrAsFH7O3a8jQJfHfyntw/BmwA/8IpgacNAjskstwdi766Brfeerp8MR0a2kv4EWorq
8sEuhO1yll3h1LDIe8xsWkg7R16cObzMdRctiDJeBekiK9IkVlVr+/Bew/WsUKQnVSISCeLkCWjB
PaKZOEiivd6mA1Y3V4fhWyZeMxNj8ppQ6Ad9x2do04+e48h9QkUzlNJgmnYvK95Yj4BLznH6CMmZ
SVDGawacC1iDLG2y+AkwsfpWV5s/fZMslZjiqQXAABTXjjxuoUNIhyK8bnSw0bSQqdto8gF72UWf
pVnPRXS4YQGd+iUO280P6zoZVmnr/wjcv0z03XI5IDfvL6qP23uzvYbjZy4czJK11yF2X6HB2iPe
4SjnjUrd/v9LDmwrafj9ziZyGGVY8uRR+bZBCa5NCpn6nrk53QN5/Ini+qu6No3VAzeA/kCEvmPb
eOaU+kK6b9msmk1lAp5s+f8ffie7ji7Py6PAIGU4L3A5+LPjaPen9EX+7klUcTbfevkdc8UJWasE
9RN41siFVqXXCsk1lot6IHQ0iLRlMECNNm9koAq8fU3xAaKylm2mSMaVaP4TnjucPttT4pqXFm7h
mteDbv5xg+SWltguiROIiJqT27n9gqkBgAnzhAeoekFnAMH7ABOSEt8cNRwePv02P6BqFYYwUSTM
fnzhAcZ8VWg044Ya+2aXZPNsvqoSv7UoFSnEBXoLQj7ffoUdb4RrOjuGEBWfv3Jshk8oTF/gnQ1x
kaND+BzEx7BbQodQY4B7aGC3fyTS61eGlb002AjrrUiAyIz0N9O/mDl9BkXlNO+ME97TUmKGCFaw
LKgw2H2yH7xaD4ZvhSSQdPp/Y7OVoau+X8Ck8OWpuAtTDP3EjXTuEe1opysDR2+SUc5q+MaOK1Ii
VzEjozYcRR3hJctqf7SOrDi+LZNKvJwu71f5iUZ9Smbhq1GniM/xExv+OKgEuP99ciQ7qiLLOkia
FgVO6p3yKlwqao8MPkhCybfh/Ci58Dofatv7lD8DEUfGDPnNWwMq1XAusxnt4YHFNHE+HmBss3su
DLdkjzKO1gRo+NlCTuBpdThjpF5ngZEuLxyW1mLrWYhtR1TpqWFxN0ROomHsTLzBYe04wnWioMeC
A1YSnyO3R5LSFobkSFO9j20QkplhtWlNuM421v78Ai6jQ3Gsac0ZIxP4pqnDwr0omIrhCwNub2Td
2UVEr/zUdl+ZSAkIskH/eAibg4jejHLGEp6TyJIK8HpAcJD+RxfT92/4AMzrDhgI0dM6C4Ol4kX2
ZYQxBV+e9255m5rRTDQQ5BluRBpun97daQxgT7Sjpqbbl31MlymoqBCzuPKDEpfmLbJx8rjWWfAV
P7oem3XBBg6zicS/zChwuPZUzFMh7eZ5vKj5DTjYps7vxUyPqOnbjJOJG8wgou/YoZhQcKxS2AKG
79sjYxVwchlO8tHQ9KbFD3vXKvyFGRZe4ATEkxuD8x92LrWTizCdm88jqzJeMdWak2rYBEGgOkX+
lSHk4gufcTnjmNwVZR6My4kGKsuDUDVxGUraYcyu2a8tg1zuuQ6PIBOVndwv1bcK9ZZJajkYlO0S
UKvT50ZwAUjp0fZmYEpucbWAzYVL/KwG3FGa/pzFEB7ZC6GiXV4GEKAVpv7hlB2k47GsUa3bM0h2
tAqA2o+S7OmfGVMlG3wvhFSY5jSbuWiK+EAEZBY9toU1XuNoo0aqBXhM3ERaEc3fvnIBLpry6Bs0
97GeJ6giqk7YtemfsnmGvPnOHGHf1Koyp72vxtC4HnMuY8vENxKberiI6PQy6obkjhUmhZqUZoD1
UAKjU38tBrqJVaNrrefEEFS3/vqZq5dnoroHaYNIQPbVlxR+7MFZE8CbN8TFeHSnmmcNeZbJmqRL
EwC7/DhsExhT7OFYYTnI5Z5L4sfMBm9as0TGqQSCVE74nGpWOkI7w5T8nomwKUCMAnvifF7qyXGC
quFUK7JCRSMx7l+ZeXtws7pwPbxBOVMqUSjImr0vNPYFe882d9Cgzl4BC8NbX02KV/hMfq5NSQSU
BJktc/6q/DVY5Hc2fgG1mBneFRO8TDfcv8iwhwweGmeMm0mRxomNlH26gVWHhSqaNVt1+mOckIhO
i8HXLdBaF3UhCOX2+yY7HRVUU7FoHaKFMkyBR5ijTeTpPiOCRIS649vS7rT/Mu2q4cJfpxFyxBDQ
vuEaWdhN8cqos78GUF1i7C81XxhaHQkKUhGAXOMlE3YKPiQyRzWw113Ft581sbvOuz1SU5qkMk3c
4doCjdXza7I/1usWDf5X7HP2Hbm7tVPCgOCg8Vtpdd2T/Z+1hyRy81dseGHVopaj6mIBbTCIhQ5q
p9Jjbrcql2V6e9DHlGibEhQTb7M4uY1Kr03J1Bawe5it8JUUOvxderzGqqY4qr/O3YOizP5qZaiN
onAn7jOO+HUhYE0Ya2ZpIlnbhxJCBbkEIhnzEZ4p4G9K7vVt6ndHI+JRtIrCK4HwS4HSy/8CqJm9
Idyj1AO9Mj2gOgYaDBN0Otse4AHx/JvtoXeTvMCmxECnvkK/YvGmB0w51d5G7TjA6e46KSoet0ie
X2R+xgnh6r7bCJ9yquFw+S8q7YSybv0ScKz6pNbt5DSixq7hGQaAApng7Ixj3WLugGOirdsuz0ea
zbcJ99XdCNgyFs4HLfhFCkRVApchJjRJCCVw0DIQsby3Cquvdx3hOOmA+SM6n3cVnz0ptxl2PXGS
xw2sqlwxrm9W3Q8A4ZcOKggHJGs8hJpAwZeE3agVDWIBw1pgUXze3uMLQo9ChSFAyg136EJxCpLY
NJGfx9E2ccr+ycOxMB8mFXNdQrbG4lcJpIlbENltsGSdHTu4bXeq02N/qD4rkUrxxP1OMjyTsLHc
vx+d4gQNp5qEep12ogHFuZjE9QeGjvwiRLLRz334jiMWqf+r5+MSl9K3zee67zIR86WjcqFHpMdo
SS9gNYXfesT/K/5DluMGiaubqV2pgDH9/ynXxe2x6no5O+LKnZ9bLaMaPwQakVGiytAOyrDRrT90
Wwynf2Z93S9m1YPB+QfTk6Tw55Kdf9Wl/PNgt2hwOEn2u7B8cqKRPyT1L1A9MKT9h2aVf59ZKwqw
SGtZbe3ryLnMVkih9oUxZ3gxONawiANnc92BSVu9pwtYyC+HDiZ4PjyjdqOw5MXuEo8BCPnoLkYw
BzFgfbHnnpakLjP5ArZ021Qs9SNuo8F719e/j/+7vy6hKt7N622Su+QTTPktr48+9qArKF5ImH2+
GnSqalc4LdxPeXWwYl55SnellWgWKXtcQR4GJvpTn+SGULO8zB7L2Ni6I8KHzYkauszn4oWIyj7n
cWXRDuCHYpjRoiUVbnFJJF4M26PRduSN9f8smRKLL7a7mya+qAlagRycCK4LnJXpCB4X9pEusuRu
4b0wsByRwoVSo7gBagmztF+bZHZDguf5d1dLJ/lQYYCamGoAj5yfkFCrnTxsE2ltBF+ZEp9aJZHj
q364LTd6JIz4ckKZxmNWy191cSycsJYJKuvFWJ2y06bbS/J7ab5SPFY66PR7rdSKlIEW5iT8Guoz
T9bwAKQvEwZKKwAPykV0WbL/SUkDTZbI/OoT+y/IsMSDRNeWH0a0cpd3MIG//S5rtroMi/20C4d2
KAnrrvDUAH9Fkwgu3JV0NSD+sMXlW0jCkCOV4Y5MApxYBs/UAco+2RBsqBQINGep4SN1Fr93sjuq
WU4QdUiS3LiOrIsySQ2Ld66ucplgFmrzte9MU7SVYgQwpFLO8SqeifEo7vJw3ADZvj86NKqpb90k
yr8k2YeYicEN5jQNfxXvSF9JHvq12lVMQXyk7pjdE6VH1y2f2DeAk+w5pc975v0C58wJ8rzrE3M3
L64I2/AdB/HlQAijxXmFFrLsInCAemc21u5fZ+BFQVMIQ8KXvPfbDxnDIPyCEMKk3fGkcURSTO0J
Oh++7yov+uvsgGGMwqfAOiosom4HHM5hvJXoR11/w50iBOpnzfjVhLfSrDblt55mVOFCmCXDs8CQ
u2o15Q7RSQYsxbndjr/9xla/1KbSA2/SGbbYGq3KjkWFYXX1W0R5TQUT/gPJm0omWWMweTbd9Omu
WwOJLfdmBo0Wx6u7OaKKB6it7dNoE5ZUosqITr23XTAPk82n2b6NiOCDjsM0n0m0Ufp4nqtnKTaV
qbk7f+KlU4RVmU8ADAO464/R34QLRbf+eaUWxE5E2WXdtgz3SUAxJ6wDgqL73s4hCOAzta/gg+XU
/tlrt9mEKLHpsmtud/nLDmztkzKhJfuAVBG12W5STp5QuFoKzF/un2Gn28YQFOVjSGRG+4GWoW+9
HC7IYyUlHD36l7Zau+oVNBTeksYJiyKG0U6unr6rhmmKRvwPQ1NoX0K/uMqNVjFO7DLE1++azsbB
rz5X2hYsVKwGG4V4vZL2Y+6yd4ZtkyrWYwyfHVjILDKuRy/LIXp4eSU9M3ilpKiWeVnGNrluv1ya
pNiHek8gzk15aAkXgU6FAwehivSbnQ6d1HJcnuzx4hENXWgTyROGyxmYCXXI7I7sU3nz9Bf6U/tW
uDZogr+FQK8OL/TNVzsMTP54QP8XVNynO3H4VktKAS89xhn0DI4hsiPAhfUisoA4IdIjOPDea8NF
esyud7Hr17ydXoIAeN5NjdDnEPmLvZQoFo+1wEZ15NJR2at7uz71/HPNuvqB9ZpRk54KvoNKH8p9
l1MCB9msWceJLXrkdhb3TVM5SzvrdZASfehC3nTqVHe7fTgMQghDK/VGjPOKzsS+ChEnqdpq8o3I
mwqxN/TNGRG2HL4YZBrE7bH8cZbGNnNY38phMa656GCmlMDcFrMU52NiVtcVmVv+sKzL7/kyFl7f
ynHc2V8z/AMUn7h0UpRomhq1X3fY+i3/18/Tjr1FLoQod7Yq+oeUWklV2Oqw6erkH2glqZxo3ie7
kXfBbs7UoT18MtFcMo+X+2TI1GfH+pKhM8v0tJAg7BZitHkpwxhqOGLjxC0QHHiOdJkYl2spzVm/
p9F+VDgVq1Jmu9AA0o3el2w1q4Wo8ph7CPr1Y4J8mhVBt3jfWderQ+mw0Tiraw8QeJHsFMtCoMmi
/AtzMMe7snYW13tZ8jzZnN3ZIN3R5YEdldAaRgIAcpUpS4CN0XO7DnQVBfkZ+PxkWTNx2Wgu38P0
h1lRnIqKlHvaGLLHWb9oqJZGe6YJ+vKVUun5hEzmMQIYueDDlUvufsAkeezo66sHIWPDR8svfszZ
CcC1UKBMfoBNd+DSSj2i6uDV2+ytd3Tw6C57ri2QFlZh6WPfUgDxQRJ5ohnpKfH1hNNf7MsJn/f7
G0jh2sSJhjXCvBaJsdkCyARFCUCKLc61a3fuIDEuNUL0cLIGz916JIn3eeTjMb7VCfU6co4ilUq7
AKRNDQ3LquC3wLoCqZUUAV0ndZX8rBfaiRk+4fWElbVDY+pqWlspPSAPIjQb+y3cS96vON1YG5k6
vWRqLZWEQqqgihoxpL4RXMVyjKh8JklMOR3xAktLwb/wIrb6Z0kR2FHv2eAwyviIBkErXMWWvCzn
IaVJh+2xR1+lBwjqSVZav8p1/971b/HKohGIwDq0RynmwK4UT47yPp+S56AUiRLsbkNPjfL9OwHg
4V/iDA0VnErFynL7amJiGWnyhmuOvfM7fc/Rzc3K89r+HjLqwmjUyd164qTz225ctr9H8EIHU1Mi
TCWcNNZpoqw9GjdPGikzEJ00DdGFR8yBJ8qAHgpXnVk6zfytPJHGQhgCd4EhMgOtnRUzjaIbev5d
YgFpv26nTtFqRm16OBP7/T4fy2B7+QyeZ1YxLPaOcSOJS9xVhY2p6WHgkSPW57j8HdDnuMVChs8c
lv99L3q1HdxDMVXIaMo07GQlma3gjQVcMa7eMSIjYhjGCOMer2EpZ6Q8QAaDBObslrStr0g/H4D2
CByKPEIyUuCHjlpTRbiqHHpYW3yB7XtTP7uf0q4zwqgD0wPS8YXTQpwcmVmVAHKr0UWN6AeQP1Cx
N0MVw97MZJrHTH6cXhc5QH1WL/l0y5WfY2apBk/jIs8xU25XjyYVAirTA6P4VpYyfjGYfmt0Jjmh
vfCveQNQbMQklJjb+TInNK7zmtRn7/qfC8sE/ZU/WoYSW1uBI8T29W6dtp2C0aTP0KIWA1lF1GGc
1FilgP00kXZEAzLKKj9EdH4nTvgdX+PECt+NoBcyXfXZS4bYYQMPClVQM2zEkJGTGfUyJ7IKWsVl
yirJIzso6nygM783zwrLMVjQ+jsfzcHqCmVngDFSgt1qyI9PmAMNBnIEaKPpzZaLyLdaU41M/0jz
CBqU7LHADjHFqMABsZ6bgp07Yo8+I5YYWykR9oKOUlHA2xjzivQ3DSoWi9X0xnQ58aM8teZH31Wj
IbsMMoLdJdGELK47f7BoyJ0AF9a/StrFRpUUuDGeMw4i1gd1DLwBqO5QbX91mo0Q3djEwYvLM5Uh
e1pVKRwWBH+iCiXZc9q3tznBIJA/uuXYutB0whfEkQCeqMEMKchgNjufXeOGPsLj9naLHOyP9vk/
iSeQnyGNhAGXCG2hNiHyXVSP8EVrR7nAxNazHbqRq6B68Zi8O2yss7bbYlUJC76WXB16Vkf6Kk8c
2ymdf0XjR6MK4gnVj6sVh28k6zFJwEXgn8E6FlI94IdvvbZkvvD9oE0LrsG+BJycgRkmM+WskPvt
GxfUNUmopEkkZr3ezuz9YslYq0Sv82haligYiP03atQvrH3waDpYdoba3s1AX8Hh6ddmvsx70m7b
XoCuGjr2bU+E7Mg3DClqWX1iluJmmbBuf3M/QtDQyntmCoAGznTiFwqhAOB4ICToxIlozY9W6aOn
WA/eo0Z2EVfUXewNvy41ewIIZl/ZdMjWL4qvLMtEuk2FpiIe+8ZwR+Y14UMohqV88Azp8aAyPQpG
4Bv4UtIehM0ROXv9gfVbGXeH65tdhZ3lIdzpdHbe4npR3AqiKljU+D5sZyj6qGovOHM+b+nUs2o5
4rwOBP7/hAQG6tTRqzUx/JYIula+AiA8NIEu38c58ChcIN46+bTbkyJ5jOOe8jfnezkJrLCXhvkg
TjwyuTCsCSRWl2mnw6Gs7dv3FCVBnr3eXkSAudLaPPgnerI01QZXfsjDrPK/9z9oEJNRFc/X3beT
ogGBdouU4Ot6kaIlkZm/STtVcVB6ZZB2u8eC+QJnDFzuLObmpUKZjA2XLWTIbgsKH50BL97P3Hee
J4vWzF+w5Bia3BLRra/GECH43AOUT0pX7d/WmIu8pgPINJjJubddXDHew5jS9ngDe04wlIT9Ej9k
fqdeTfWi9lVO73zhuwd7KDewBl1PhXy/Am5w8u1qmqcTWlvdzY08RdRROt8llcHo7XnEXd5ORVRF
qXMbgL2R4RZ23DqbAMBNfSk0SbKJ6f0t8hzHdOpmD82Ol35P4lFAOWHtd4vVxKk5Ep3ytcxSUZd2
dLfomQ2hoMN7wzozqDzVZkyRehsADu0kCG3miHH3/JoQzWRF/ASuSmy7slYPRttpePtfW0CKzDJo
hr1Ids7WXIIE1qAsD358w0TiCA0uFivxx3QkxU8FmmJyW7fz/uZRy2KxetlxcvB2mALkXjcACRMZ
Mb19iF2z657S9oH6moEyBoB1xvYVj6JQTA2YBJ2rL3yG1T/rTo8i6FT50luKB6+hoA/2KIWn1vi3
tTj+/Sb2Ds8NJd58A09lKfhYqDlzTy2LRaCAwCYbXsTTaoAT2/9Ks2VEVbo3a4G9mBsclQDVgHAs
vx2gFWggfJ03XzzFezJ/uSS8fhDBFf8BBVtn3fgoqj4wXnbJ3x92Y822fagsPBwkkMPRtrgvROO2
IeE2rXLtMlZ43k/vGQ8AQSMYZOlG92BNzdf05UMbW/x3dosTd85oJbkG9A9XB1P4/Vp9KweG670Z
NgRQapX+zwX7q0C5ZHjb2oVRllh9ya2OJ1/mmi60AUtmQCw70jIb8iMbS2f6TJgwrAuOSX5C99dN
XKWXtCGVt7OzZ/KZ3jVjSbUofNbnfbkF/GX1p1ik6mCuInfVXd9BNzz79dlngcInzs1SA0D2HN7W
+STBG7+veY/kZXBAISzQrMG4qjeVjucpnHVKcgdN2K4pPyWMTSPz6CluWz/UqJwy2JumqSkp6Aew
idEUVPpxmvjqid/ew7KFyVbymAQlBCI5gJESwsO8zhb5H9pfl0hj1ssOy9E4n7bv2YTkMsLVXZZH
emDr0fRTIueKjK6wHyHWYSc0ev0WlGeYK8vGNHdURBTm//mXXS8K+e9Sr2W83XmcNLgqcIafq7VQ
I5hlgcDW6apwidFuOD5e4u5w6CYgPMvB8FaeXPC2fhj87nq0a7n+bGiF1I4VBHIVG+CQ2yYeG2Qh
Om/jeyukF2XmVHtXq2JScPfN2zike+XqSa5rrfigEyrUPKwX2SOdIQMNbyebl/NZ+KEsMXL+r73l
ieZKDnSRYD5Aqtvoz+ohoXDFiizGl2vntjoTyztMb6VWtUtttlbjBTRWfKJrIIzljDl8vsBDnv+6
9Na7buvW6Q+OGGSpz1XqogcX8q4+pYeO/N5+n9NTJtG6ppfWQwJqUID8POPdDvd2JN3Qybdz9hyY
4491ndq4q1r99U0IAfjC/fZTabIav5vOHGdJ5F39MNZch8kPZfzFuXqA+qj+ZpCjd++Wpxu08u7Q
rsWWJtBYKLOYzRVhw6VcwWQ+TLL2H2mYpwQEmBFMvXsLfI7sMSPhpm4Hzz+RIpQxp9trIQBVy4v/
3+otMqFsTar2LoT6wFagnh7GmtOgjKXIVtpuDMVG9jNpkNiyaSIv4YoHlPW98tFPqBScoa8Xmwse
IFfGNxueSzaN7iASGLYz0AV+ETXhOq3uoONsNJXbuw1l3IPbo01oiVk1Q7hSQt/kd0wDryLCsael
xtA2T2LWrIHSvZF6GeEtivtfvUdKzgp3h9Qkj61BHd/2erZj2RYSgbpjkfC4FLm6SIreNXwU4VkJ
k8KoU5WeB2Stuodtm4PHXYMjcIEa5LbFyAHzxskFJ/NCNCYC2SrFk3NLERemOXFfCbwJSJ7+wCN+
oQIoTeS6lOuih4y9p5TY/qYqDYoaKGPCiVjXuwE4QTc6hnOCOlDVlXCvlgfuXcLVmo0boOk3TXuE
pIcP51zoko9Tc5AxMpqOFnGRaL5sLtcAcoXUEKvJ5B+rLhE51IBr5WUAia4DvEXNE3gfdoRyeDbk
ww1/VCog3/2zTHGhyB0kyJujEdFlI1n4YQj46ZMOWN8ZMMA+QWg2NOMfgSxPx/+DzL1g6AL3v/wV
aUlF1XWA547N1dMSMHGerjw9/7pHNOIxT7y2Uwb1vd5YMR3al9G2HrElDOaNcrzsls4IYyaVuDoT
wliKSMyMr597fvpoUffUgYG+aXkvYaHfOqRAueXEMC/ZjHrBHkjcx/pYrHCbXp2P3KkCR0SS5aAC
YDuCXrs7yFn5yJzdecQXfiVTe/9kHVrljFsXKys1+0PaSgQw1zYm3rEWurhkDHS6wzYv+oA7EjTG
qz2iL0nVPN3NKNfod0UrMxhrxkIbwVU51Zgt5DYDpQWzW+Nddy7s+FQtEG3hMlS/qW2PflUUD8Mq
d5iRXH2ftGwF25uavI+Ucax/OOhHEGmFJpDtooSVQ3tRFvzm8H/zKsZkxOzAXTxoQTidRypm9gPz
RW00rKxF2wyszjviMDoBmYcYr5kFhAkHZIk1MedajNRZ+iBVbD4KSOGQnOflo/aLCmO5SVV8so4D
zpREv9h3zdEjG4gjUNlC/1XzehtIke+/f+IhxBqfnxz/KpvnooCHlK5fuOeUmMs6GqkODz4KojT8
k453RkF6YGAWEok32UqGw3isOybaefeJIEaoSP05CKq8VwSF51VxTIs4WfMvZ6aUUi19i95KBL3C
Xrn8B3UG+ETZS6jrMvagRoLPs4HYdNB3FBcQ3Q1vHqEk1SKQo4TE7CY7F4IdZg4FKpF3hZjZkDwe
9l0JVrTdyqBLjlf9ETFrF24iVQe3O82fii6si52ULAqO8GTlJVaf5e1oMD/O9s6Jm57j6TjZlo0f
eqs3faJjrUbskRfIkXwj4WB99KlKUamwIHG4pGW6+S2ObQj3KchSJI+lLFLkfIzZ457fPCtC61/Z
xRY0dplEE4YtUH3Dcfrnf2ke2wFyJXP9AppWMoGH7j/XN5zfmoValDQuhQYcqIbymv6Dm9Kmy7kg
7Nwia52LvwuXr01lMVQChzVdeclZp8Ofn5l0mONDAwI4kop3GAxDoypLf/xM0m23l0MqepWj02rN
nF6XiCtUcZ9S+XIShsTSanBkFNKlb9YunINPe5EsgqNb0fTqTFe00N602citBeod0cmFsjdMtP1V
qcNdnNaYTgtm9aRC6qj/95lvsy/G1WawNm4DdCUUBIhFXlcHkFW9AmB+LVtBoVBFkdfem4nRbSTh
F52UMjIMRFZHEjc6lJOJfV7tS2ZWQafOEMJKTWRK5oc2FE3RreiOegkntkFTJZvJblXALIK5a6xp
4L5w0BX7AaJmUIww+qW02DZsosgSIU2mqfggUR6Ps8Vv6/EYAtq8cQC1qJvUqxfMar66dnqgHOAA
j1oeDv+IV3Oap5kKwML/liAqoMaXSVRbwjyLwrbSIJjXdQY9gtPCdk6hF5XwU6jO78D5Ak2iWw/w
UkrCvhIKekTxvATpvxJfvO5+ZqY09kLd3VWBjfe/I6u4+IBH2Uq7xIbh+M/O/ik6gvryHr0LsgZu
4xwLT6rfY8wRukw7776co/bwogj0DwxqR5ZmGn1SBeZA3mKh/8kdCUHXCOFrml8HCx7Iu+WaKZWp
+N3zMAdzXs95TrKegBTjyVpzUx0gx0BGwpS+3ZovCQuFfz83k6JhOvdLUD+0gNSdNK4aCVHVmclo
zozR4maXtgIj6VR0FOah6ByPfhDqKBam3sbiszM86pKmlE2hI7qeO8kaUFmdaFa8twiM5Ot8kdTN
H2z+mZTEG9NSkUH1q1ED/isX6hKzMGZOqhpIKueLVmsBc7jRaiCCZUgbAMt7KPXVDrPSkjkAppb6
ZycF5IBkfNRXhdg87YwnkwGsK10xmjwg3FSloD5Fbte/WOnOIO2QHcNn/G8in143EasHiCe0f7lW
yDy/Hm53A4123q+1R8c6LfWYUj/z+vY9P1UI0gOLNsq4kxFMPgIhMS/v+uX3BM4jq40LrJwrdlpr
1/NfAH/Sqjj5dQBE4O8eW3BwI/o1Iw3a9N/QKluijxO8KneeYLGMMpSyNSUyXNSmaVsEt0wbkPJk
/nQgz0s8ArWLu2EOmXSRV/Z2f/IerKaH68XoWs8DjjZNcMqz0Ur9yeuAtf+eOG2Cr+jYytQBe53b
jCxVBUyon0OfJqsbHoon8ey3sNS8aCnFZjQcgQK/ryGSvJ571W4R6gEfsfJi0wBDKUVUWRcQ8Q50
kXvm8BE9KmxVmUg9a8oCaq1Ch0rsBmk1CrK3/zLS/VMjejiOWFkUaUhJQ3TOWS77drpDqpuzXZuC
qqVA8Lnn9RFqU5KxjdObhnmW+sG+QqGZOjDJv/Mu8sGqF8Z/uDPhOGcFy6OnmTcGTsqLVDFHz9/r
1zNdM2/5aozA3odDNxGyvGJ4zqgIAEH7MTiwwganrQIG/ShU3w44R+Rx2cr7MsX9ZQ1MiY1fWLdU
tGPBS+OVfi9XDfl5TxyOwEsP4sSwcNEEYTbZpELT/EjqA58PLQWJqwDMc+MvjCzVWN6aYeeYPAOg
ecQTGY6TTOcQLJL0OwDC8Bo1pMsBnz4DTgCxHpidoPyvvdOemujsOVobFQ+RYs9AgpcoEVk7imI+
xlpHSe0iX0lNBY4zbtOdtOTbM86zQdATAY7BfcuZTAJvX3vXv9gRR+LPWXC1adF0ILEF6iCYgZHl
ZkY7A/sBvWx9qEVT2UjYt+oOGrnome2ll0PYQbGT5s5R+nAxbUKL5LuErJCkevlaZlT3DG8O/z08
2bKDDxYo4FJR5504vHDcF/b2M7Jkin7eyXwqvoNA1XR7pomMNUCZApIdzwGGPqrVnktBwAucdTUn
Y6xoN/TubuFGGeDA9o1qiF94AfjIuf+OXPdoi7RWzwHGOl2IoGEfQGNSPE0FU3MuXxk5XaAtB6wC
K5hiRpvAStSO8LwP4EvbwzVygUMhEMijAwv4Ehk2lquOox49EHm2MIgmRPdJD8StK5J08WblMmPH
yynoTn3agnPEijNUQRG1/Pbl9XXWXtrWgm2pTj/RU3coCW/dicoLbQ6ijdiBpkUS1GguzMWIlY0j
ztb42//oyBvQuZ97oSg5NZ6wcv4daoaFMa8aVQNYzxjnMiPzOL5/Z6VTmSX9WPgYvj4FYtc4vaVE
cz8Azdf8z/qQV2bcps7qZ1OMdCd62aXM2+459gy0vjv+cuxk1HyArAIIDLFI4MDXCvyID/mmb9nv
ZC7sAEWuhoQSNH8WyareOCHAuE65991/LBtXs+sr5zgT77vIPPBghcM9Sz9dKLoxWRXGV+KfytO4
yhT7TsFSl0CL1Xd97g9sXlsLtCz2mJ4ykalexDz/U7zcgKSzEg0RXz30lA941UcE2hLxOhXERwJS
N4pBTwe5vQbx2W3ud8PwOPsMKV79Yg96bw272GEaWjRNZ3uQ2JgZ/P7ljHzENJYj53+zFYmYLwtQ
ua+iVT7ys/91RkeEEVrs5zpwVrDkdmWyqpYFNOW27h1kynK4saR2zgsdJCzJIIcgN4Qg7OvhJkjD
Cb0qHI2RHvCNaiKmnyoeaC0wizC/0qFmXjv1wW3fBiLBbrohRGETNtj3EYTN5TU8r/UYZoXLRhuM
tenJMam1nZjpnedmtRpFYFx4sFXpuanudq8QeoDbmi35nHKFSSomUI6c4QCIfK+OcCAKufLrwvPc
/0j1kBSOheU2cbkLfdVMsMNE62akIONUHO0W5K8bsg8EjxupvBwNN/478Szmy0EQdk4aFz0fyLE+
gLiVbFJujyfyOmDGq+5tjBDUP769AZlRCNBnFm4wBWI9FO7APzO9UVj67z02yiHEPII3qExxxj4l
x1V3jPcEcWHHXkUR1OZH5i8xuHUKN5ZWGP1aiJ2PhHuODJNYiua2r55Esqzc6jLeNdWEYZVOr8Eb
/Lq2kL4QM31Y+EJfYwgZ37WFoY+Ck9DawG0NOs6gzMW0TtpbOUnKvGX5sWg+w6RrtgltbpZAcQEI
V2A12+/dAGtMvwMEbnp+5RYXYuYrzqK8JX8ClpZ+nTRdhrDVrKaYLBg/te/tD2jeBL11Yg+mF56Q
qbpGveTaKNhwR7QEIJeoYIWNfnFlL33bWYqJBpn0PLwUC3nRGbpLWhWVrTkwdrjBJdkrz5REIGGi
twClEXpkNDd0pVzQU/Pp9zdGlgyTZxfTvgXujRZ4DHOmtc3XCmaWmOI7y2fv0DrzSLQsKk+f+jZK
kobzhvgG4PSAhBU3uq/oc3kKpvZhzunQvw2JtdEfzDQ+mRLVgZ/aBIExN8f+iYjc5zGhuIhalaKJ
Q6F0DNDlKbCVNNSrM69W70L0VDqYdlCxWLCgARE++P+YQ+Dw8doOZclxE9egTbt1F/DFTLNFIdke
U/Mfm3RcTHi69fBIM47xaFCzu6PJQxaXbTMqKa6XkzS+lsnXPmjOTW2KFBVQMCZ4Cvmn6I4GVYoP
Q323tVJaCNvROZ3ko3oroduEgT51yX/ls5qMRe/4j8JW8pQzvRGKU3zTzg8BbWpFsA2/QerfrEJk
t1pISTJ+vwb25LCV0RsELgSRN04goOGMPVmCU9aVgjvq0RRoo8Ny//F5is4+VxaUT9vOA6o39jZ9
hGDN6yQfQqYe9m55EAQ/FIMoxhOtSBhco3G5JpcCe4pluqCrXFiwx35iQvT4jTwJ1nH5wRVnmFe7
hjz/qhg6IbrnhSx4g9XDZB/4KIzJHvAAuMiJP06LdH+7e9a4LDG6kPvBLroUxKbMqtGahIGw0EEq
IhmOANGHtwn6mGFt0MuO9ptBVMMie3uCvWqSXiRKOvNZbRYAb1ozHthtAv3+SA2fWMQCleVaAvEu
w9J/0LIQKRjhDmlxuN7u9rm2PM3X+5u4rsbIOp87Wu3Yo5sAiKuW4oEJUxbG/ToMOPJrerhk5iqb
nzNeLGaW4ZtGmnOWZFPNUC6zZxES+QCZQx6wGv20CBnqBh8ubgfflDBNsjbFN11hcDgFmysN22go
2DbfqSpo3oo6jpErzo96nXX0T3xr9bpUZv5jXTUcpBsVnOc9yaJDxuvYyDmtCt5dIYmKZbVV8maQ
tfuDUTW8HOaNC6m7AQZwI8V9+OzAawOGNYZt6nny3ULut4OxwKIw1L5Ru4zNCS31OLH9yssyGagp
20HrYcgeWiyRVZyp/poEsQDUi/CeloYYOu84/RQyhljbuIWw4KSodYnrcEHmR4AHVdwrs4f4kyb3
xa5hcGvyk4OkBSHGUKnnUVecEsuXYqmVrnCfWIhvJTn12JBlXC+SofASGZdKX/pNleqGa1xPfI7l
ShsA9L/MamR6DnDsAlSv123jNsODJ121jj6lXXkeqIeo/LglECayH9Yb7wAWUv9fdbJToVUnVs4a
AJBP6Jm1EM9y7LuANot3HvrkW5ZwgeXmxRa36aK66X9/z+hTth4ByAqgGowkZu3g4bVoMH6gOfT1
7dP9A0dIcqawqx3iFcmGg2iNDM1X6tyBOmCxQQfdj9HOkWsncgto7WzehFt833pDx/fAvvIeYYWU
WjgDV5ho47MxihKUQh40++fYVLd5i34B1y/lYGFDRu689HE/ZavhngxQDy3l541XtGoC27XOXGmc
/HuynfvZrcq7tSHZRgBKunWKDj67WeeWgob7mk3d2v1BgmP9D3ZBSD/ZrI7bbYqGT+1HJYEgPxlL
0XkH25PzOSqqnj3UUaAP/43ynhlPL9mBamWvXcTj5OM5raWzKaF6b/v7kr2WZzPOcq5o7LasO00L
NeIi5k8jArSSz7KorR83mYWajOzJ2mPa6/WH0GmNRWUvKZ0Ea2/RMXowVicspb7jNgNxBAH+FKBZ
VzL/t+VXjPnNKjfmu4g0SkASgWx4F+OLo748yarbAd6JaM1TTnbeFktcnz3YuN657Kwa1lPc2Mvj
GgPrgd/SfWK7qUgxYtDHkjhEsPFWCBqebgJvJ8LsUJqcrdEW9KlA4het8bHKh5UCvt2LOklaO6V7
po+bJM1hjiiYwUNWBLkyWP8dKiqAaee33Fd0C6bnNM1WLL5elk8LxjZzU2A72w47wS3g4djSNvP6
tpF2NhmF9wMQ8f9AGC92b4Zfm/4vQItLx3XXb1xa3bCr12wHS5G6YE1NiUNzavy3KJTUlt/t3pSo
dZQTaoywRjCIHLJbvmY0PARLKp0qmZeSHBq+lBI/7T0SWVuUN8BwNFLLN1DArqNqZiDIGzKhp8iT
mY7tnp6xl70sMeZRkfjr/+Cuxn+NgRj2ForaDE3zQilFbftx65YlZxQSGH3/lc1X1aEfGg+d68Nh
ldxBO4CCTsiqcmmdPXvUEzxKp77eMe6MyrAFUJom1Har+yF3qbFmpOIi5GWEno1A1BGxacvzuian
JQXfaX+ugnUHJ5untJ/g0LwhGY9a1EZtzKvP5x6XKnvDHtIxkK2z2HzvHlJ/oNm02FpeO9+oWoZm
XDZ4d6kSh5krpEUxYHL9r4CePtB769ILpPpIDAZdA2npeP9xafsRPdyb+QUjbZPiUPUadOpgqX/M
7izeCADbimhsaDABcifK4XcjN6t9f82GZjDgkBb0TwJZSxAekp0WMpMLaXN6K0nwjGoN+mOjqil8
OUuXTT2dEFw3dOkZmzeAvRi42XBHqdMPKTJZEcg6rO1bN6lnI0qR/mI8tINte6iVUx0BAdPJCbDZ
P/FkKpa3cAkCYKymWX9XCqrkLcEzSqnDwPMdsTNXRY2vOGG4a9VlHMpA5f4aNS3BC+SOOwiTy7bt
+gL4JZViC3cMVkJqnozerz6TqCfHRaQHsnyvaRJMSnVaMLsBXacGtM1XeajHo4L+RWA3brATbulb
D/W0sUnRiyaDwKjfTLBOiURysbVlJBedI3kgk7n8TmTPDnYDGm86oLyeTkMydcUTC6JsuD7K5gsk
NFMnbLyQTWRd670gqFSi1D4yZclFytf6Hq5/OFz7qpsHxciRUrlHwJq1yqqJxg3ZJr3tc3B4nUKo
oyjv2JHkZsMiE2qx26MPvwx/o/ZRsM/mYqUerpzc3Be7qsORfX0IB2VioQWrwJOMChAxhAPdHfRV
m/Ah5VR3uEYmVB0O4b/8LmZaL5lbH7fcKUz3EsP6WSyYPzQBBlfzt74XzZEEvPmlXxUC8Uj0ILU9
MbPHmXR0uvBerg1StoZ+xbZO3COsypiwPhF0MXgYGD+Aly8IFJQCoSDyKZ6wvsskXOXZVamXZMIu
v1TiK8Qj3ZPBcHZQSGB1bz72qgvNHfDl2fk+8IValS02saGl1JNsRpGuy2LkDWkjvX1iUtxREiL+
M8eOasGPRKTfI30OehStHfCKRIFcQ/COsT8njsvQ7TroocVDSb1gbXQlVRcMyeRicNMDFj7ncAS/
YhpRS9lXxEKDCcnq+y0tOvj6pZnUjOh7VSBZt3alIgP4Dcbp3vS9L/JOTc8sA9fiO7gYFxuKIl3y
m3qG2VD/4eK73prx4V5I6G6MCjiMDfzxYQGpXEfKxaCqAZ/tWbPf2WW6KOzlLXAos/Qjpex2pS1G
8ohKQ8jmjNZ6zvtPLLl7be4SM+Ky9viPHT3kjfAyJ0zxiYQzFX3bFY/mUXuaMODVfSh9EhsQogmK
CIWQjTpNdhmsucwou4/jdrL9s8gbRtvJOm+0V+ffcPAn/xgDu2HqM4DD8dyL3p/gYz8wm1ozteAu
RTUE00/KRkQr5YoKeeV1G+eo4KxCA0YkMN1gAFzWmxdF75jgBUe4jL9EAXFFECkzCORWceGD9wWs
LdWzi4P1r0dCeelKuRJoyT7xGt7fxBlOZtW4Vd/LsUHhAJMlFJc31o9zkcVMhUT1hmGNrnZI1wYX
jfp7iRsezyN48+eSaqahGOVPgJii63pSI+lopxQRzCPoFfnBoGp4sZEhIsKpL62kaHONMRqQQ1F2
CC+wU/7X4JGRuxNUwTpGSqan/u6koJNIlVaYV9yKlUnbHDct96ZJYa98rvgsHsObFJXtKRYJIG/t
UC2tIVSti2kPKR1NhJzyMYqpfS71xB9Cjkg9YrMHK6NuMJh6yfnZIAQoLVTgYpniKXk/3VZSGqev
2rthTdPWj53LlC723oIVkCY8PbpmzOhL1O/8gOu0lfjGIt54inqBozpA1zGdnZplUnCzBL8sVaEj
dsidGPapHuF4KMFS/vuc+FsZ/pzpnwkcx1MSnBzooJVsL4ZQf7+0v0cU4NnBrObL4zqgZBPOV74S
0lVIp/nkXqNm6ymzcYKyzcz9fPAyX0tlqMY8F0gCs2OL4nzcQmI/fFgDFmZNmgj6FwkkkuKqKMJy
9Wu3NNb8Ic0XciwJ3y8NmomfmB7ot3euz+7iBDpku8EXkfgWYR91/UNmKsBi0B3jmX1kKBEMKwGQ
6JPWB+98OJ7eg5LWglp7/fOUqYY9TG+r4mssq4DvQIU92QHZl7xlFiKlqlqOp6wZH4jQ8fV9qPcV
rxP6OYGARbK++uTJhHAGbG5DjaPvFz+k/MuU6Joayd+YMA98M/m8Pq3NDY5fzmfUcJJEHln8Cy1l
vsWuC4ySjitm+qR13tYjNmLO/UL9Eku8kDNGatPCJ7Q1H1NoxuLcABMkURwri5naTkt0XG0iRlG3
cALsDxcfThNGJ3KTSfP6A2D0VrSbOpu3WLJFFw/SsNcTL4vT86NWTVVWyueFvnP20j5WFK1/mjUt
lkU6m3nOjcgex8z/6pFwAIphvne9S3snYQ7hTrbHCzf7TUepE0tPyAI3JB47hIhzGTgm19TrTSt/
SsJRa7V/IXDKiqHURY50X7KGyRNVW5EFs0TYiuz8SEJK1/hkNz6EkHkzrqMwc1OHmcQKmnMjggpJ
bZt4mTL1IXZoeh0v8RarHIO/VYXoGfMoKlRRiUu5xB4Gcu5Ck6XApa1DCva3wd5mSGZqpLsh06uB
HLpLEKYwiri8Bcb7f9iY0Wwuflk7m+LRzSYMN6AHcsrGSOTgpVMKiyO3G5dwsNaHA8HONbWv1iSX
iB2g+EYv6jCvgg0llMwkijpjOueSqdOs5LlcaB55lnwyKVzBj1ABos0P2CWPUvBWLA30Egg+A1ok
7NT5vapRfOZjjd+0zkY+sHMqJjXliIFmikj0LWPCeILdP7Jx/SD+8MTkZxkmkf4etDrmRwYGE+La
ORB0AL5CfXr5MobWUsmMo0njQx6FM6rylqVQtQeBFJw+zDQ0vEA8Z6Z/m8bdLoCu/Zd2whoJxJ29
GJP5H6+EWvVTly5t1ZodgJ8BCrSfrwftGHFpiJsvtFGw70FsOfiI/r3sjK2GzcQn3wc4CKShtJYx
WAL/T5UQkA/6cpIkHhgliLMTlkRDg5wcOvkMzP7qY99JnHT+9jGlXPIixeuEeFwQ7szFEsF/5z3y
vooegqIbCIkocTlBUn6Ri+9IpAeUk/Z8h2/61u5zXKOboBQF78T38SkhA4V6hhl8n7opDytxaUeu
H13cfi3nU99wC1W69L9B2bOtI4C9UnGQuwMkugtLW7ymq2pK0wKXBWmpjlYlFazcOgONJkT3RS30
6bpBGcyxXn2v+sK57n7Vg1hLWfupzG0S9nUU+QrenqQd9oTqi5g5SLSMNEW5kQg+x8VRiwjw+M19
SL1wTGzzocTK/hAiIRdFC+rneyAVm9B9HJSHyOjy96bHBgfhxqzJRK/5CWf7ITcy//BJaZmuJUHI
GtyV0aTWZxsyQLBsfn3SgVDWB3lDfaIctjISdxpt9Z0oUh5C+Z/Out4EUL+FoIzJt6zF5ovy1XeR
ObfUNmkPbmGTozmOyy9BoLCtNVMGmwh0t3wwq+rczBuucvcTvrC0L8mWvcBhTW+28a2hq13xX4OP
wc9oz1iug83ExOKKFMUGBfN4CvwDXyVGWrUJEEpRj4gXsMPl37+lyvSOt05khhQuQnyq1SFJyOko
7VatO9HNgoAa3RKCqi2cQk9+xr3fwWUV2mCLBIRLcfBrY1d4N8LxwqVjxMG55k+jibCshZSJIzYU
vG9AkH9faWEJOY8D6xJzWT3hU2LFfJZB52c7AZBk93XkkDBTdOhkz1DLJDPp7uu+GYcAbW3Ihvyj
0OmrUoruWkz9C4DbHQpyX2kNqg1vZ3YQHT93iyXTSp7T/YvncbnczjazlX0L6MHPKZlCjRrHDoWh
ADuixBSysKKRTSFF79BWj2S6ZeKM7qZ6K4wy+0vfQSxyohXmCY4SF8kAJi/iuSazCA1kYdiei55t
DNpEwIb7DcfouUzQwKGP788bZp2pyxbLehtF8oupI8wVTXzUuqA7TcOHaVEluO+pgB2xWPYRhLTt
UygF/wN463H2smaHvGLzsBf2N89e8gLmt/sR84Thi+P49Kn2o2wZiU0i2MO7Q5zAaGf5s3WpnZyk
UUkonp2TNgND1n0426qLvFJOw7v/NylEoqdVHsEFjJ4LmVClFsEAoXTnH4iY0dm3dqnEAOdUoJ3x
cQ2BadiN/+kCFVGc1nsDS+vA4Jwapvh72xgsmfLEF1IzCR84a/6OQfUNPnsysajGxKPz3/x+I8IO
AuC6ZznJ6KxVa5/s11T/pL9lo26JzQ0qbDLZqWdlf8PUltMgiPCByTzn790Qw+eiGMdUfhtJNjKg
FjenTVPZlz5Yhs4ncXX8ZZbIxaS82Y+fruZda6OgxKvXA5reaMqs7CSOZchhCsFI9mTceGJHUs3s
kKElSvGBG4r1+KqsOOoroDKDObGLZyPH2J9a4OJEpL7g/g5mOyD7aNP3iBEdjm87sJ5n7/I70hZn
7/qtWmjkpfb1TJgcRsRYOPoK4WSZl5SKjv3zIq7APbA9VZMYd4v6ViD511w5139+mE6VnNdvwP8J
0NYxxVWUYIUJ1Y9QbSZEFp98/hrVocIpeWeTu0Tx0ayeVfvrSrTn4BWqajXuCtbOV5a5VQ25reFd
QGg9AviTgaB8KpGDRQ8frjyTcMZwyPzSJtNO2iOcOFS6i42ScC1BSx0qa0D/WQuR3uyvUVlYOyhF
CxyFmnRVVZZEh5VqGxYmTr69LQWUybdZSRUvUSaMhW7GoiHte1bbdrOz50R5MkmdU78WbTbiuMqa
UyYatcY0wyPR3xG7CJ+sep+ZlSYQjiukNyD7qe7WnLz0gOfAjD/WouXbNMPT55Q6ojo9843/R5g0
cghTSd4PB0pmoxvIjolxmilyDgRVI/sZ7+MSHr9DksOg179Tr8MdsQc49iaOU2t9BuiU2GaD52WP
j7zNJOqZKCmJ2ypK0H48n6kcTXvp+JsaMFtcVRsn2Ol/9uvhs1nLqu4hnRHPj/sq6wbGduUNemW9
KpssW3CFBhRsNz3qOVy6VziDd9cTldlm/78mZgQURJzPcpRZB7GAeajEgrqgHCjhhkwAKtkaBecc
85g5c87tlSTbP3rR9izLxcIe8YSJtQnUDucBjPh2P64RZvi8Uaybs1R2bYtL7/irQPec+hc8B10e
goKPtOmMbgIkcoxlKorRj3f/lXNxEA9F8I1o8Zi3sVcq/CeTaeIh8VSMax3BGTrS0C+1qNr7v3yf
qVAokquxgkUpgRF+M2dncq5iBEojOVpA+6F1uybdlyY+BvuFFot2hJDmzvaH9Jk8w/4ob6YVifIX
Tq3yczk9UcKx5DOf1NoQgZwTMEx9Tma2fFkPuBRpfJVD768OVAT+JUMxPyCINjlRd7tz8EUv5CZU
pOict0+ArvgC72fs8DcjCdXryqJeX/DgzQDTr8OeBjLKz5sTtrD8L0uIpCLpHjUza3hUAWPz11aJ
yBVTZ1bTsXbq2yEmP0u4Fl59E+qzjjpa9w4CFg1oXbWCLzVyHraGQvEybhCB2x0AAH7fICJAe8dc
ywEBE6VzMRCFZ8r5y4j+Js9HMcHg96tiVgUPrAsJKeWx5qKNXm8RhSBiGruhpef8vRConI1Nn7jG
fi9Qq/BRaUIRBvbc9jvNx2IkifR69VEcDtSleE5fwRlNgKx8oMPs7cO38Y7FLfXzS8LvmMsQG+Pr
EjWq96oNTRoHbSzS6CyL3peKwe8Q1M2A3PY8LYN/kZ7511nJ0srTZQB4CUuAM1t5Goh+Wm56ibG+
oyYoaxpb8iUTnkRlH3WtXXho3LafZ187uqC9no/U806aQpZcwSWe2jfPxlXVXA8V+C9KhFF0WZhX
0+Al3yOO2pLeRNEyqDdOOdhJ04wt2d5uo5PLlJ7efx8Jz0Vs6DhJONmPtIcA0lbNYtfYOt1JrLyQ
4bM5CmM1QYWvPd1lRZiUo+K8uwggKX5kL3YNwzDEkc9qXeU+fiJqivd1WBdktqQckPhnKN3bXYAa
gXiK4cyxKOaeizJJOhJjYLrTaBxyt3B85RVBmoRqTx1ypxjO0q1nrCvy0HlxJcOPD4K146mSgWWh
3kDT4AmAGcHJwO3SMnL33KgeLBoJ95TtIzYSNk5tip91hQqoFDypXmp6AKj//NYuARgb0QSZoTSO
iwbc3XUXf21dC3wulOiX+JmzubgkNtO5sOu55mZPUj5+weEH9dczmmw+54zGJ2ZqSa3gaFJ5b1Ti
C3rP/Z87p3TnhHolTg3wnjVy3OKeVsUGbY/YBv67XTJQnKAH7LyArVTZ5bwf95NhQ77M66fW3cSZ
CKZYp9pOsL2II1rfxlsyyCc+efPV4dpA442Lvyh2tknKl2qsUXmkueeebdt6gGUa7UzlG2awq7VG
KvL84VGZlutkl3IeXddBumSQWCL2yD5BsiVWx6IzwPwSIUUCCTk28zqCRPqg72MjUdbMt03anlPc
x99MWtZkoY8hKnNvz9pd1iOzr8Mo+hwETINgNOasMHCfzN4h+eQ9oRB0STJZ+x8O+Zv7lhp9BC5O
5gx+uGuLP4j/a9Okw4JE7aqP1ScMZBQFIsLXN1xqdeiEmxVWrPnG+hpB6ohBFgrRsngB9mTox3oR
WE+BlB/IIocWfWh/sPf4z+GJGKKOiMbBFjeRfnl4HSQW7uf+dOTfllNFA/Bw+Dusq7zJ9gjgQeWo
MWPCXJy8CYomS1jWG3ikNJCzbH4ml22gdtcT1x5UcRlneg4U9v7rE/jd8CefBkyKQHG/S46HUgyt
mbGhjKL1XoJZuZZqHTsEkL0NdsZ4L3Ub4WcLqBRFLRqEfaot2LiOHwb9lEb0Nk5WV3MeFKN/0tBE
2w4+Eft2cIjL5gjqnWMeCPpYHkvDjGfTlzk3HdDHwoMiegT4VObQk4Ky7pT3zFg/Ezm2LGB4XCXw
yhFQUVnSjrjMqqvJ0JH2ayj5kkSlVstUWh+z/H2neoUxW8EEDVtVymrUx9jkl7B0KjNuSyxwyo5K
K8op5mw9dwvuMHw5r/oPX2MJJ2ZU+x5k1vTenz0Xv6QTMifNZCELDMddtqg6hQluaW7uLUz3JiGs
kwXxzhzehZ16Po/IMtA9VNFErved33SQtGe+m/dddkX3ZGtGjq8urMyPl4D734RH0muNBDMdK12k
JcWRXjklBMZwHmvwJbMIhSWBvR/CzVqMD7YGMD0uMURhZUKx7Vpe/BSzm+9QqcjKWnPhmKVScbHR
+taO0ZyndsxVXnAtpFZclz5CmFqMtNOBEvfe4RunnFWbebC/kUKRBEFr0g4ZVVZlnsic3VozuUQv
8RCquTzQ537IZkKslxJpSrMpHzZuj4HNGTBwr+KPZHPQ6W2wtIsDY9J6/ROVrhKj1GdOEEqPe+ik
EvMGZ6tU+F1QDfzpfnyQLqxoJVfGKPBvoCDUe9p0OlWJEf+XYYOM718MsYr9OSr1VZ8mYYBhB4g6
uDv9OdbHcN5SKLlC2hlNvttspMaflj0AYGAGmEdZ/or03JWwhyys8WH2Pb1tqNfo3oE7QlLO3dey
H6SRpKhFI7owh+qbnScTvBH3Cxw69rG92K0mmiyQ7MkWSLD29byLzUDUCe83mLzEAT6rh+U9W+OS
HwOw4GkpBWb1gHI2UOo+KKU0aY1TZPEzS/yGd8Vo4op9y4KE0TLvlHWRKGUAay75NvEsBfvf+FGk
oLFAViyKhoXAJsckjq9VlyE7NeUluaN6awYa3nfXjL2TruqhBSgjyjdm0sv5qQZqv/RmqjgBaFWS
p53mm1xonEKXHdm1WgAqfSERmlhLlq4+seFBfndGMaTrar7h5xuKqmdl+mqMErX9P0Vy4Ge+/Ok4
OLJv1AwF0P/GTiBcLnRrxy3AJe++nXH5dDoPCmmqyO4vK9enLEXBsBycaMY6ixD9c5ZIIXsucaLv
a3BES0Rlcl6UuOo2rYbr7TFrBdYQIefbReLWlc1qyecB+7DOUbskSe/V7e+pqg5ePcQ7Ima9tMv3
01PbJRZmT8yzvgvODFp3YW4XOqP2ZsISkUHfrHehEC++hDVF/2aQZ1zVoJM4cQvEwjpXn5h0D9E+
ej18yx/Y18GCiU4HfTj/fsE2Cf3DY57U3gXIQTrfs6co/I4rkMVuYr89bOc7TC1eqRVuLMN5KbwR
zJlZ3BfLGFT4woWUW18ypuA9S75bIjtcew/wfgVaLM3Q5BzEItOfbS8BpPkjhfbagcrd1HIQLkKK
VPE9raAf5Jmr08Hv3Ecky0au9j5AL+avTDOFNYdSowYgBfkU+gMSpmShCbInfJLWwtbF+u4897he
0y35lPLZufH5UPzAddjyVRDjyFC79b3PFFuVjNpzDnzPfJ61TikOhTgdAtG1PqdbhIA1yMNMXal4
d7uGYYMiOUDkL7k9Yab7EiRC//z2XzbVuWvgaj7y3kSGdyQqusGAzNdpzbPRiq7JypDXrawZL8kR
ix8BbF6X2pnNlNyAVPgae8lznMK12yC9LhK+wYO8XVzcznIr/T5R4mVAFbqdFuGY4N5td6X1BSNY
1VGFUTpPfiH/wjQXXc/ReCoyvr8dyPwcTWMXsmLOHln/qFnXX+JkWvMeW4rbC8+aFSKekfINEk3W
q0NTnacex2Vkcr4bV+fGu2+lTFLSr7LMrmSxQdQEbWwU14zbkH6xlhC8Hi8IpvXele31TaXLf9u7
EAe/JRSAbqIJiq9MS2ZDLQYMiRP9TlHWRqdZnSUQQr0+fCnKYD8igyE3w+W3UWhi38SQ2NU6TEXH
McoCsW1NyoGrnWnKuYsRNH4xFzIWQ397Rox33OQ1G63f6OWKUA+CFz/927TskDIbxChvKFCRsw9o
zzx4JveuzAzyavNu9qFOWK3FMtdwveseIhKQIGZCbM2RtC3HRMp8/5wsJY/iAG8gjJoKfJGiY2DD
/vyUDVdxotRD0eZ10k+IlVTXxSfz/ysj/1i3oELTFvo0j2454r3R3cxWmIqvQU0iSWEqcjkCCHBZ
xw1Amg6x+pnwA3fgFzyclJ0/3fIvlMZjno1OOSKXVQPiF4SGniJHw0xEt2v+lFOuAajrZhsarxEn
o+yJMFBsPWnxk3f5GNJ4UAn7UIqh21qQMptTBBMlpRsaBW6Ex2/9t1OkxzCBE/aoUt179ePnVSWa
XqmPM9DIe7pt/M0DfozFIauZbkg4+ZpmOyX1tJzDJ5ZzGAZFEV38tlLBwTtxk/gJFGdHfTZPDd4F
HE5tXoBr07xsaKJkCoM5jOIGAt0iZRRBUP5TBnrVP45l1uUW0Bx++lldwJnXb3CAHGyG3hxd2HPv
OVFpl0XAadavsXB4GLKR6I6KhXhXvchkPftBz4DixSBGovXjhG67RomRR0UuBknuBpyt2BaD8IK0
MCvLYvdEFbuY8a0nv75RL+JnuGDJIhC5kFcOWFWGr0b0vVfq0VYPyhTSZqWyMyGtyowm2W+7qw72
gbxxS/jL4nPCEfMmQH8GoZAZykUOFpjaCVqH/zG6n7nhqWnOvaDuUcGYbyohZfFVYZG7+oZBFduP
4ztTPZRE6wAGCk/E32iyWfhb7BHA/NwVQIvNOduJ9sgALJrUj2pXds0MknXAJsJms3l3T+2Ovu8I
GcbT1OXg/EU1lyHQErSTABkYsvhVLw3YpIqu/yrIJA7XWV2wBHfnNMMi7syJStX8eexwnWRhVouT
sAi6ObuzQDWcqWa+xO0r9dRuAy8d8ugjK+lXH4Dz6uZr3HlfzfT5xiJpCVo34EMhbhrORwLrQlUA
Zq8oUGBSDa8LJlDrmxWvsmj9RGpwqq7foyFmvz3qqxHgU2y1ot5RpVEwfWhbVVbdeav0bajtdOsu
ty+kgW030jaY/pAnMpj3N9rXo/VGOcSRDpk7tJOYMzG2J9J2Dzx+v0aHqyyZyBKMgphshJmMuNSJ
LmTCv5kmPXaErQLCcUDJl350EBr7moPjZphDbdJV/EGHpj5jy4zh/MCLMKKNuEJGMsZu7DFp0/d+
2t5bC+9Fr87ifkjUY/kLPCud4JAmGBEvukaF23RX18j+bIdxbn28MuxfjsJU3HUVWcNZZtVQ0Llv
8r6CHdIpoLJ5H6C682SWC5Q4ozb2x580Xaw0u/5bNxyXdyyfB9qRrOuGT50inbfk14ZQilFlUxcs
WLzRAHzLGc8vXnMKBa9VdZ5pBVPdRiQckelDQ+oapDXaN6PGJgBwghlH8m5yeMNrliYYowWAUTRx
I5CFwpqAR/uPyd5cE53oirUWY3OKprhuqUJ/sYGm2zEmCnXJryrJDPNbONLyjN3hAM3Ii/A5dnXT
vAMMfcaSCa4KRtGz7iJFva+wvj8SArLAR9lhtHukyvlFH6a+AyYEcx6QvkFlOPpSLzYX0H9NSqHK
lPp3IHDo+FtwFQzqJpTXpNy8Jv/L19YmKBanRedat03mFgGpP+yl7Mk9QqgpUTsyGeaPkJONeSXJ
5k6rNGTsn1jBz16soQ82G76CPyem7EoETBHjxBZO12bBXoa74rufxusjCcG/VyP6FSH46PGtwNTW
2V7mzz/UBNXzHdsFvHlRMTUKhDQRzyoq/+eH450s2I9BZfzvwgk0itpqfWVrP+LgC6/WKlhQT7cI
rhVGUW0c3mghHbRTPJ+25f8SjNEQ8U8/GrpbMy2YO5xdI6ODqaEsOfW0wc0FVmva7v5rVs7gjdQz
iWV51clX3eIxUac14f/fOlg+MDNz8gGTGw7RDJL/wIFQIAq6WNoVK5dU5I0Eg0LXDs6kXrj+K34k
eDPyOF2kpslUuJ76FRlxUEsE3WdHA0s1NRXEjSg3uVkYQSBexz/Zypll8cuOc7VuXoSQEL3DQv9+
bd374tKn73jNfmIQR5rQ9Ih2Tl9PDZCmY6ijjxWje62WYKMDY2Xp9QgzkH8aX4Ptpl4QtyxhWnuu
2IP6JvIXfJ6CdZJtbcNxFM9mhaXsMjKHSpsyf7vr0MzBzrva5teQTsXvVp50cCC5p/fZvfZRGWZR
ziPZsQqSnGFt7qqV4YcJhZ7QwGi3+6sVxFvGr2t7yJQnXmTgQNx3akMy3pqx/AAgUpn8L9DdkW3X
4LHkOcwgzYtzwHMiVaIVr4RpmEA5YGZrTuqGIh9BuEeveXhVmHg2ktlPWLuim8MWw/QGMDxVBsWm
7C2wZiTggNrzkRCgbQmoAsCowN8AVdEWFZ2LT7LpCmcacR5uWNrsJE/1/tBe/B+mjh2v17Lq9ouL
OGb7438fd3FA/NPXY1WAYdAFc3GEGFalNfWk66X6DgyITb7rg6+NP1Riv2rTRXQ8J43NhbIBOC8c
tSyG+LcEMxoQFZnonTuKtgLwUH2INEbmQFfFGQATw+ZGVQr4Kk3WLq8d+C0vGQjh/NVX/6yVckzi
BsS3da2QelHnet9EVFsvLlGNMa3WNeDLxwAbKNdTMNBtQt/7H2ytsA0wcgAk3cDTYWG53r6rN/Ln
+MDOKXIgo68HidNhtoE9xBND/KIFXvI8wV8A2QbxifUjf8AmaFu0K4tKeFUXg0dyzXV/lzx/MjC0
7s/ETqVTyrhVvIMbhtO0gS2P+l4dwWlOZZdQTmd97V0lX10BnJFwh86DW2Ghn5Owam6iyMrMEiMa
gA9UE4dUFQ2e+jvRTuE9dEI6n77BZ+xBH+noMkrsDivz+VXljD+yc/mXNp/s00mnfi884RbVE5xI
pDTcJKMQpSr/EZYKeWopVkjMkHVbFmWPgq34JNJTBT4LsxA7sRw32IGx+Snhicr+ag0TGAUdbk2y
6Wb0LfDkMzKIqAItmOEVhxqhqmHURM//9bCqDbYNqbmDQxcsXbPMW9JGghC45wu4TJ9TuSEEktQi
FvUsd+WW8IIRKx854FDII/HEoMIlxFHEbItuEYKPSkO7Uj1zMfyl7DmbJarYY/KLWr7InhC2jIR7
bncy/My8QI5fc1jyhUNyknKrpJ3f0QhtPDCBfxuBXQaJDKHjLxpJcGcgQGrM8B/weEvz2oAjlkTQ
2Gtozgw6dA+eIbFmDtW/ukc7d8u6QAyeuUDjdUe9cWvVg759vQ2BnVPa5tCjL8FpLMl1Jl7jiEJq
6WVRuIA7xh5SCDWp5qb+mlRasn8Mhba+W4z/NNRAhsr8jC3KfK2G5Va+7/8ghfhihhLdUzpWwJOU
SZn07Y1hl0od3cqQRPNzJFkQkvsx7Ve2WPtGjjWNdv5tTNNHKRtaZsaC5dKLn1nzByxrBVLQP7Pc
bh4qqNpNa/3LwXCBc1+L3RosF+0BfDgxdKh6u507wPFsVb/91o0eueHt1RP8LJW4ylTElBTsLL+X
oJJ3S/daMxHwlj03JuAWUSOjdqp2h0sff0hTpqe5F9s2sZ8cv1dYt5kbxwrZ4QcWF6Bs18ENmM5E
PHGFuYvUGGBpPcFfZdQMyfXU9t4LmOuHRTw/OO9DeiIkXUOXgDLo5hy/juR87nbeVzeFx8KodpZo
VYM+tGzeCC0tkDU0y4JdRac4Qa1l9tDehPqighXFv9Cbm8KbsLnFD/mULwgquNSfR4Q8xTsVh3E7
lduKz3Fuj7lXqbQKn5xklRuojne9mEhWVg46XwPRBM7Blv4nC/kVZgVxEwrbIR/pPDYHeryzjQWe
pfntd+YccOjqs1/y7qxgFtL13cP9Sw00fvcQPdBTRdGKaieVzoYWnTKZ93dopuzyEDn3i/LfXBqR
l2bIi2/Q6CC1VhLyLauTfO3/ZldjZjTvTrf2UQc7Z1MDYVt626pavXAgpDwllbVp9pfpcgr8xa19
ZXkubTUKIb1KoZ4tIQXzf8RkHgenfMJz3hCKQsISM89mb5lWuJdVvyQcjO2EA2Z4PdYBVDE0H+RD
ew1axUtr2WrPelX08XXJMCRtb+vtZXV9LJBP7XfnQKtbhzbj4Pc9yqHm1WF1X4PuLu/VX3VLOvrR
uK1kDfjyNdgpfZuGL3jCEkuqGAJ1OhTHC/RfcwDhj1IT5y1cHEOBQpKIUlQt5nD/g9cvHFEt4Lm5
y9b2Syb2HlUJ/u3p1oE0cMeFwUAEsHM2gQOpETBmTSnBX/iiBkdBtdwMa5qWX1oxbcEj36+5kQx9
Hd0sBeuKXXjgqECdVnljg5FP6fBOdLfsOFUNDE7ZKm61qMEJh9mTI1zxKkm4iZnW3awHf8i7u8Zv
KlrAv6rnWFnDd7P8Wf3v71nJznSIcNYY9JsR6aEncm444i6NNEBUNet1S05cJ3t+0ckdp9D2baBS
qWIJyQcG90mzqddBUYZxukUORgU1i5XOkR3LIO1iv+7tc3xVprr+MYq6nuFh5hbfAGv/bZFKw85V
LRfzExEY1XB6w3t9nZoNA66GTjA21qB+XJUfAnwZAq+0FzN2joKFtF/EHrtMkXcWACG9HRNj68g2
ofY35EkKCPJCDcEUIVOX9DXpR5Di/zVeRxRQv69enAHQg8KG7WCzfo5ILQHuyEEcQ8q5nrlmuyqd
rmspCPfE4EC13XE9pIEjle1oOV7EETOsld9UzvRgTdrsQFnsMp+RgJ5tHqJ0XAdMGk64XoiVTeKF
PExqUB1UstlPFoo470VEMLYyxghdgmrPhpgfdG2+agxGP3bAyNIOCMGVDqBHs4JUodz1G5POSq2A
3SofRIWzo8mtz1V3fHdH6ts03WGLraRO1adRInZoCOx9RSsSSewjIJeTQaiGn3wR4Gx/x8u/OkuI
Qr2ldbIkGC2TOoBtd3KGDBPIME9l+bMVlzPh+Dl0pqSlM+rSuHPb0OkE7G7Qyb/mN/M9ijZSAHto
9SNYWhe57iMy7Cs79si1PpibXC/ne2SviRP9kAQaLbdKseeN8estT8VrzVA24GmX1C3dt9pcihgF
Z28U/o74DgHEQPjep4JAoIOWeOZAvyvZL3+8z5YL3FAG2M3cGpiuWe29+lG08IDIB3XN922flEFz
+H0Q4qiFEKSc73PapeHh61/cCvF7QZGd/y+VsbeiBajmdJbC9drnYtVK1ixR3i+GcPWjxuxGmPPS
1PZ1uIoJ3bRRG6urkzbcKlsRUjgP1oP90HjdyJdwSRdTte4aANqMfq1ivi9DZJ0O5th4Axyj4KL7
q2bNwMbMnjzdHv+0GSgMUSzzCfxzmoJPnRJpw2YKb+YSk2exGFpZxqgNdEd9uihxwhig1F9e1A6b
sRFh5gR29MckvcUNw83f0KXGL+FFKDJvRqYHjHFn8Nk1gWIVcG8fK6imOF7m0CWSLmZg7z8IwL/o
Nnhi3omp/40YJ0K5AadPmM88pWJvNto0hUue2tsxh5/J7TSs60LmVQ1Fb8LEw3oMO7Wywbpcvju0
Wgvpa1y8CGyXRAB1OCIePBQ4RFAmE4Ck9fKLPBsp9Nvw9IkQ51xPLL38oYE/2wetgBgfGviilZVb
vBE4IrEntrrdMqlqHqtsI/G5x/GZDikqJsJxzIjR6AZrfWHyM6Y6DnkqwxpuXT2CW1SUARWnvo4p
mxP/TNSO6SxoDnYyMrhi+4UWdxhpM+TANZV8Lh5sYCKtCkl7Bo58dYn3DpaLpNMudbU6QVLOA03w
VmcGZX1yEVwX9Y3vynuxXSBE3XEFkfyWZRlRHpTRTYQkeXwUO/5y+9vQiS2+VW43XrnW2fpyz3o+
EUtvKzSAanAiJZbQRGdeLO0pUX4/orhCPZTgod/fIxykJx3MqD4GRBWoTKAjwpMNGAC5yLoyiRGT
8eEfQrMsNngkCsUXeTTwnew9pkGkErhfJ7izDgL2FD30btPdEi25IzjVUa45THPcE8srm3xIU6ey
tunnaebWrbsbZJj12qO/DIObkOlkstaaJcg2/wp4MEUVD6wLaion072NtLVZQniBSW8aswyOrz2s
SMMblGQHp9r2POv9DAUlZSrHkxoCmRX6r7+4jdqpoIxTv40Rx2H2W4t+lP6Y5a0BgsUN3/0jZ2Ik
r5ZqPkn33TPUQd3egwpawQx0j4IGR1XtygTpBzfrYwi921VKsZpVM0j/sdi43tPgEe9NnCBtKGrv
wzOYIlk5aRyAlyETbV2HdIDJmzg3HL5XOk3vTHX+C1/M+VxqOeFO1ZLMvBacHyllfOLQlXyGO85R
Ittuo9yQojeX6kBdkZivFa7s0m9KWHy53Tr1DtZ+PNn+iVqbMIQII9x1RhgNFDJli5QyGrDA8OMc
862uMlvWgggcm7lq7xQA9Ly5CRYEgLlGLSyj2AXaIETR6yQz719mi2BCDPGbakhs6zwvhjSxNdNv
AUZJL0Dvxz9pTlQSKf/u4l8G4KYjN0H/zUuUZoU9wiWEV3qeB2wWSuRhrW55pSE9KtxordUIaGqe
QZ9DwWE/iSMcj1c87uuW8Xf8RIurVeYHEhfV+ygIizJCDeK5SjAgV573VfbFzY9VAMCP66Bv+933
30W5KKGP9GG6VyAEHwHrTIUvCuwaAis7es2mXz03A6/fwaDf4WTZjtfzxTiEdmOMqV94p1l9NunE
O73HXGDUk9MJN/e/cYm1kVE5bedYtEw2x2j0kI5bk/L0tYA/dCrf5rS0a+HoTTTMPoKps1YtH8QP
XiREhr1cAPUJQn/UgFE85LUFur47z3YFTR3h2w3vIe3hrqp+ZoS7nqRsBtt02RVezvwc2XtLHbAY
20Fcbyh+LR0RBDvatko8w7g0KAOWXu0ww2qclmNVITXIKlFEdgb5IyQjwnwy0c7Os+Ouf954DvAE
fPBJn8syNlFLvhYopPH7aQ3tsVUbEr/R7PGrgtURgvhW+t19mJSnq8mE4PBdX7UGW6EVXKC/ky6b
JXAdU/2EwYYixz4fepnojFIWtryIw+0huEmn6ZuREgNCqfw0GAwW3lNgbv5TsAErDHToEDpbu0jF
5geV4gFs09287Pd+RU21gMnAPjZda89n9xqRQUVjRiRMg4xiYAymawC0bQulw48ApTTlj+szxn6u
CQRK1IakzRIKpwlnkwlleQ/SyB9ivTdHdvYeJzh4PEKxlUdiDnn9fdpfdaT027QM+VmdRSX4MufY
GxmUerU7Y9tDj8JDgr4CmY9TBeuI8O0CdS9fXS/irfhLrFqkw26CVnhNUDzTQcOUyP3zHtlcQcn2
RWhRkUQxfD2ngWiXgIXkT8dSW3b5H7ITr+64qB6OBDSTSB07W+qvJmTu5agJKXjhpVPSotiGiPn0
hsPFuZnyGBhos/8rnFULm7U80WcEJLPCehyiXL7Pu+mYNiwb3Il0p0geu6wbLHHPsTm2olJo3ysw
xXBVYf3NyJAg2V6lb3B0hozhurkF8HRQjgYNZSsqdi3LwK5sW3YFEiLLfpqWO113h4SxMQ7PKLnp
xf/YxxaaI+gAGDKocwxmcKoJTCPY44a4OMGO2Sto1rqlwJmTZTlf1UmvRyZpHrJLR4y8nfI0JE78
6r2WLbPj06fWCfJfk8a9oHPc2tN6KZUptHS47Bqgkbr77E/tOxFvFULpkVAI7sRLHu1WWCUFnCJu
zBKcQ4bj6wm4H3691PCTDcSxahm7mqsViiL07Ey1DYGz1aD6icGyCYs/rIbDUV0eA1MnBiEqIpyI
lShYJDlxfDpbOgnfifkh9wKn1Bwo3unrdy3TYKtv3L5ikN0/Xub/1RkhXcJzJANNZrRt/woQVAPn
wWaZaIcs6/extOF1SiEsd+Jyu2VyZoEDVMUovVpicMQ5TusF+SSdjDYp/nlKfQPyRoGxGBgEEXYv
UWpJyc04ek1Ck2JmgINWxyrPG9D6HcaREXXaCi0e0aZy40Nx20fVbmcXyXBGPN3b40S18dyzE/aA
RzF+i5QpPVc/I+44g5gdvEPoS74NjrycjMqHih5LVHsdccTOPOgO1Gr5iqnLzn72bWTMtCzPFlE1
AyuduRF1lEoPkLqN7WFySLwZPdzw2CZNjrKy+dnjGuPuymcrVe97e9nIP302y0SgJaeW4frdsRho
ZGaD9z3s+WZ15FOaEAHuc03inw2ZekpAsju1tHsNEU0JeTveO3EdfgSxvgApDCuhK5YqogZkedxC
ceBP+dKvuNj9T6uMNNw01yd0fkUIsoU173fxDvDA/Zu1+xfPN8r3Fb+JwPcbJjDUmVz4HO/7xjgx
47oAAZzQTetuF/q9Rd3axbI4hbfr1SmvjcdHTkCUWCCZdDWZps0zL4EY9UhxPSQj7enA+VRormO2
ic+FSBUR5lR1PT9f4+nD/OKQZ1tlynzmkXdUzWFiOhTTN7NiH8sSjHLkzZMFhshR5blvnmZCrjnN
eyldbngWRyb1TFQttKOtzRjfxkui4TtXNZsyMY9iOgKv2pedx2rwLSm0j3hvs/Tk4/Ymrwi71qkQ
SBMw92rdZi21w1jlpv8iQJ1B+sG3fi30xFuQY3/u/SSBlCas7JbMn6v6SgGt7ho/juo/X4Td+R6b
DMhAFIBDgaStMAAp0dk8qN9/hGDzOeiRbSX5kH/VlXz2F4hRMN7on8cgrl0lDzYaw6c9KMNMYrSu
ZSvD4jioRM+5mbDKAllk5KfidL4VkcgTdNGkDsVBVzN8a3JmCimia9O4JwxLTSTkv3zM/GV0kQgf
H934AquNuOU0RMV2Cokyzo5p6f9n85Xdzi0REtUM6Xql5jTr50Q2gou6bDCQPDOjKvVtJM/FUHl6
UClbv+lnitLq8SYtWOB7l0VCh2rpgBa/a4IJtTe3hUn3dQBSqxX/vGdGJwKUTG/204HuhbMAIJYR
RjQ5cMJfWzRk5KWi25qzMg3Ip+pSgrAWBPDp/DOAxB4kc3eJwAdXdtMNRSaOimcdlhbXGd7/qF7Y
IIokPUuqKd+XYXp3W1QyHsr8U0UCjEkW2ul3bFlSl38VbrwS7dcHqA6K0Jbm+r3fnpk2mIMgI3VJ
fyLUa7P03g4tEcKrP6qxWJJ9oGbpNNExJCsjf7Gre+P7sJRAV5Qih+xJa18LUB3WzOPXuEcw7nRr
UPDCJoooPbd90ANJDd4Av3NvmDcLjKKfLI4C2IgG2hZyUuGURGfJhy4RFzPF8WAwwLs4hglF+VHX
rzSgwzMY0S+qmmMlktuMQR4/etaMd2mC7geycBLoCW9DfKXxGBJpxM4P3rUA6LO0tbIfNRDMVfWo
X7dorjq16EsP+REbdax7uOK3wUQlu+s+X9TqITVTopxYjeDhci41BwW3r20wwPtKj9Fq2RiRZUsy
W5cRKEvu6ZUxjURf520VCaJ2xDSnKBB9e+eViAHpB22WxDrTd5/V7mJ37/07+8Lg+LmKdQMJXjWa
93p9HCTWG04XQTX5H4kC4P7j6habHF0iLKEX3ymLIkoBcw2PX8ui3pdXxHVE/06zCEU6jjmuO1lc
UVk/wz8cNtxdTrBW+2f0Xghh28FtgKbNJmcpgKbBX7bzRBI/QdzXMFGshWfjP/IHpB5CtmTVi1ti
7Fi46sXIP+yS4d2z+041mE6wSLtnI4JpYxoFWPA53S7CV5HNkCzidl3UZFIXdD+CaG0JiQOlgtsC
0Y/DO4JzTqi2aUuYlrVUamzv4CHO3QUtwU17POgc+qACOH+VGD69ddSkwAW6xYK+VnzGj3FqdEJp
zdTd1TpTNuy+Hw3QRE6IvEzapz/zhTYuYvnhdYKEAZeNEKerUpcGoiM0A6JAumqELyv+GzXEpv1z
R+eT46yBp8oxnBzO/ujAQZxo08HKmqfs9VDcjg66/JiLhAggP+Xt0C+KzI/VZ6u1+EyIXQ63/HU/
AynhluSVLIbxGj1PjJabvLcHgoVALUDqGR7Yx1Wotby49cqbA20s6l1ylJHtEbbtNNsz01xKSFKH
qBmuD7LKfS8UYmebKTAGt3+UncafkprX85uJLi10/a7nvOwMNkEreh9pFVlLRlbg+zh+UnloLDTf
vKDu/mBhJ7aNp0xbnwrK3hG23aDSo3oJtuFPBVPNjBwumUXLoJZDSzpGqGTfqUDUYo8hskqwGYpa
1//F3u8JTg/XOPiQpjvIKdAzn+ucPoapXJvO+efpQmO40SpiJaU4tnt/xqp2aYP/1GoX35FPlMmu
f+aFtZToKR2MOyVlcKSkOgkMXHQtJACxmxFpL/X7hJbfPZjH8tTi5NElgjACm3+ztd9dOiQx5lCB
Qkev9LzXv0CqA+rx7SqLTRVhPuX4SdnL3gbulj8NGCHHWGcMxh5fbZTJ5v72mbjyQXYMEiqvR6Di
9nqFAKUpa0CoM6+e5b9B/Ccs70u2ygdop82AJ4zyTVGi7ffzwWHRhIO7D2VYK22vvy/DeiOhaHyt
uxQ00aKF1akMms6jDACQu9Pl83LPGXFVaNFiaZ1/qn4BdLa4k1ewDc4DzkW5Bgrai8hB4wDcL1L+
MLQ8ia7U09PbjFjbHrdP1hMvER7OJNlqAa8eMvOjSIAFc6ZB3+pI0jMeE18SSdOxeZIdREQlF7dz
CZApYzXoOuptarm49Ycw8YRC59zQi1vNvBFRZHCUjDgL+ZwSXs2WjZjLV5029A2TjoStisiqV6bF
JXjFLrKXpM2hvwf6mWlK395IS9S7LVt++ZHuZwGKkcyxS69skOTRPV8geR8pe0BrWyINY+Ij351W
8PSVRY1UjSTcVUDv0Lw1fVA4n6I7Zg3Tp79KtskF3TM4LIiI1BoP8aSVjp9mH3X5hcEXVehi+z4U
cpY3HlITj5I2MzTfjq86NHut2X4ASbKd9/hG/DHn4XPIEIB4wb5NjTV9tVZOgoA7DhYWotPVEzOp
gslMPig3Hrr+NtWMhii9vd3d+9al/64D3w5FelN9IIcgEfmR70oIv4gRpEpo2DxCEDfTF8hcm13a
A9ka40zrT/GWdiypLQIkG4BNIkM3B6siJnnegq78DZHTaNpzy0m1p3VSrMoPZsGx8bJeP39kNw9j
sJNhoCTio1kbt+ESp5n8zTu/+7Uqko4rbxqM9cpk8OFTFcCmHYZdY36pq+DADP/D9MJFU8tmnXNk
3X461GC926PehqUFxAZywmG0ZmkFJBbbEya/FPHa+t6SfWOu01RnuWj+XgWwRaGBR28l4zEpxfpP
s5GK5Hui3X9ZQrixblPr1WAUe3aG7YqLolq2k7+DZDDW4z6Rc+gDGTSHoHn1TiCWefbiD6XwnNYe
nhO0eFlXDIrCvwsW6jXSZi88lYpPqsUQqo5vTHoMCdZFSZhrP2/2gfenhMWFO+y3FVL4csRSlfqh
AVfyz0hmW+7HU7yJ/n7X1OgEpo4iLbKjN4FfuRVQmMUj1HuZvDaWHDJD9T6qmryFzQovjfnLGRdy
0yrNmUdf+6IMpQnoS2lfwyxAdwcyZTaPdBVKLtg2NqAQxuqSjn8YwRx6IzQsLUzU0Io/REQsOUCp
UFzBK0t/IM3usB53o9bwr/J6LGWaYPdfMfzFsulSSxvA5xzJgoPegb+fNUtWPo7LtTfGlb+G1MeF
5h0raGOdae8BIdKlRsjZhdl1eAzO9ODYhDNRsctCh3QM0asxX7e36MQiJiws+lYTYy4nEpxC/LcX
o18lEN7Bz2vVJHe1EsKAxD3iJzsSe/QVzh6bmwe+sde8vtzdkN+QoNMFSU8hTG3jIdunl2HabZp6
NiY7o9fdXOgOfUUPcP3Eypu40bjjV3KxSSRB8JLqPmTNvJ3BaeK74BUyiSLmgolkzELnsijJc6pT
DZ5uYv+1wb1jlJXHnvOEdrZnKoEY/rnQlkLqoR7Io8xmvg+x9GKaeipzW4KSlYUAiD2QbIQguFFw
UEOZ1rOrOF6qXPyP07peF9uKp2a+zRfbIpweW6v1JF1MB99Pd/47bCWkbTpfsz/XRDp27IPKKJ/R
Xyw+ZeW79x5Uvvb/ldlDylg1R0QlyUpq+7O/dWeTTCx/M/uF8LrirnDBMnmw1NtPPFNaBzRKmuoN
K0qm8HCmJ2GyVeUqMO5vOoG8+cHKBq9HbgQ9GeYdar1ORlDUZ92nOIkAlpmMASCiYqxAfTHBGL4z
JXAlH186SANSxMXhQ5yZ5wJqXFOTV0mxtuwHFtibxJSrtfKZwpRo/o0cWJWRmWtpKCGaMr0f8F/Q
+fZ5pcV+oUvSaY1in9AiILbbNvu0GOxLQs0Th2O4WQFkV7eicvR/YwVVuEm/84lHuuPyigxeOzqb
v5373HVmJ08Uq43zk3z5aiIs9Dm0CqBPJKZ3X+YjV+3c1mHUKj40jX3V7ZBcndbDkplU0o0ZL5PG
tQEyGf2vJ+iXsFVyg6p8qhsrLIictZgcTfrfK6q1RxtrrtArI5Hg2PnJhQNCZuxHw44AfZQEYPs4
4hFF88giVYF35moJxJ9bkRbuL8aF38tdVFVmAtR0N95AIYoMlBva812Tvj7kgClKjnGIXNI/1VKr
K1F7RJcOasAvyT9kf2rO9aSgFOKaRLEmK4SHi6Vws61g8vWdQaRlH2TZjSwI0J3vgxeuqMLXjZPF
9GNrGJOTuFehdwTNDVcCI7X2Zqp0jf/jte8dY0L1XQE/1RgHNMhFhMN+O1IWCZrKbbqWIASifbVV
Ol6GuJEHTZdGDmyWWI/Ajw9n8LKV7LoexFFFE8YEMJHtX5LijZQfGcOBU2E0yenz4j+c2VETO/76
6kirCmhCkw58+Klak+tBqhSIELnvHiUksM5KtBcw3QQx+nTEfBOotxfQSRgG+uvfkYSxnrJA2NGc
hzLpNr145DTW/ZpRSneHGnFC+2RuQF/tluKlTEN7G3KR/NeeWtP/7ubebgTkrIluvY3BO/gmfxUB
jaWF0cuoH07Q+wjvgp23zd/wVCAtz62AYiiRNFpQpXNdCkiO3XUqNDoKQs9xY+5KGGV0nARL+dPx
Gh8OSZRKiRGzjL22FfhCBrHnXrn+ZDrvCvFdlBPaG4A/ly2aMCY/BjnP6IQf/7dTb4RqFuUvG5W8
MxnGCU4mE4K4jutFLMgziGkPtdaX6cpSct00kt3h3pzJehjMIP+hEdwE4y13HrhtRecoMs3vZAP+
yZfPguBDA9ZK/JNJSYS6wcMlbiNCQY/MRWe+NLYUNwzSwOEX7GwmFC4hycS5hnGSMBixk5hAun9E
aoS3eQADn9lPmFzA2y8zWuRW1Mz8LgWooM8bcxU+9nh5NLzrDToV6bVcd8oqLOWnt2BfwPwl4ftc
1rroXVANtBYyxkei+lbxqzYkpiVR7+Lgpw/dDDCmbYvthzCWGBJez9pw9jw4m6/d3pliPfSLwNY8
hpF/iMC9B4SRj7BudCP/FN7TmwEX1OaLI08ZJTCBBY6vq5lYWT7F1BLb4O4+Tmt671fltG1ZYygs
Qd/5XG/p6zYEJMXlERkL28hpcEDi5QhgW3Mw9UVRBE8jaeifjhEy5piX7ff0ygADGkitcyYlYDqD
2BSjrT4fHx+iD5yDaZrY6xWFX30obkchZuTsyvk8e4tu/rjCcFFCVSGBdhsKK7AJWhN+NwYeYwOZ
9DgrpBcHUCQoeRwSIyANJ1hXX0lr+m9kgjcO2320k8oxQ3ctGGTyHcVp64tX0xuZ2dcYFK/8UbG7
aiZ5VuPp5naQTOY2XrgQzbjm1O2ZIiYwFMrV9pIBjPZhVTk0CVNQ8I0w6ps0Rp2G10lXEssWAyUP
CDFnvqnRRKkhBEdini0kJyHPGpmtNRym/YOzxW/u4pz7SYTqWFMnImHf5/XjJiBBmBZweFXh2WRA
986fjpZkx6AJaqiNrjBxZWcfgb9AFa6QZGzb085QHsOjl15axcxYO9Rm7bGQwNRMBP2FBQEQYRJV
rYBTdEeAl3hP8skhcVXOPaT0SLQI+L5E1t14UArdyrOfw8DL9tM850tMhEZreKOiY1EMiUcp4arT
z+KQf5sjAWbq316I3dtTvooIRrAaR7v93szZ6JAu0BecYgUwfMhQIiH26yeQFXb3rUZtRJz6b9wL
WsACiQ5kJQlFUXX278BM/wLSQkMtIm0SrFxbPjLsQ/q0mDqUzgvEGAV9b4YhpztSthrYil+Q8+q9
73i4w2W6JFavz+kFFp4gxWRnUMtiiI5yohiNRRfKlEKWhq4m+ZaqmU+h+b8+47JQKU7mZX/aUJ0S
1JqeypJmczdB34FbLR2X/cSYCmpawYLV82oVHfY7N1BSULLdVdfXKJdGelM+SPW3NistkBM1VObI
rwL+VfWrmen97gfIIOsZuRMMddMgYQdoWIr7kZjGXPADMQwrkbLTjvywIitr6wkluaQIQMFVo0g4
9EHxJ9ZMQih4UQM0YoaOeD8zIMcfn6R21uVIlMzlfmRZG3CmgcfEjzAvPDJ0pjic+0K3FuxZv3NW
NKIPg4/2+PG4UWlKf0WmTQxSQL7jEvj0NfH23Msl3dJoLsg5keJcRo5HG73+vkinsvUM5V24Avf6
BsqKfizHZxcMJShEuXniGUnj1fVfN1ZbijuB92x6dq9nzodzY/eobJo8urQ1tTCQ11jiVq6OrW6Q
wCJKx+iPlML4hr5XkC9hrhakJczY2+h1mmUL85mUaBsGaplSsdjzGtRWtcKa68oMleVuVnVLUgAL
C7wHz+ARgdz6nUGVxO/QpBKzZglqNdRTyl29o9y7dqhBXeJ7iV0YkHF4ia9lgCHd/77npRqPWt1r
BHI+5HMHGfxxJ0z6LLRqES1UnHZDK87X+2eFt1Hla/uKXQRnbL0IxWOHuUPEPiYH2h+O/1YNmu8n
+K9iFXiOTMG5+ojk8WTOZ21P6ugEsxWvClc7UT/rikZ3eeQ8UR4gFBRfs14iGY/rErqbxKfgk1g8
f9fA5ANb8Zx4/YQHifp/TLRHM1iTEnHiSm2fUfr43me2Xn2v3mKeaxpHw6bNRwY9YkcGOmhEnTEo
+igZ+Hj+wSIgjIBdHIig3h7sUMI0IhVS0gnWbQljSQenij1vUHELF7h9fygiaoP+o+csUOnlP6sw
JiUZ6vgxsWjGLlalnHlyEptwSVlMcaWg2wgpCjnINnbZDXnTVYpXsNV2N8nbzwTOAixuZ0FzD0Ee
ZWDMUYQzgEhMGsWNAruzYGWHhbYTRTqAn4TZ26uPoXQzI9yb+2ZUulkFUBf4fMBWSDwIkvL0ln2u
B3ZO9Koy0kgOR6SLA8gX0VtfctSfPe1wi6rE3fQ6B0e8ISFZw7UCZFwUO1ddsvppm8JaQL7GCd2T
tQn7S9/uCga/EhZwkXte5VQwfAiML6aaEI+R822ijcEMKV3yd5qO/wiyeQujmTcoSvwubbH1nyAX
AAIlStB20Bxr1wyLtRT5cioHJYJsXxLCqDO35RRK96MRW7jXOOS6loJFL61PI5jzthJ+En5lzqPH
uSlnVz/lAQogJkSr2c7bsebNxEPlNQd6WrFfm0kSqNgPZQqa0PplHCmxo2DnneSe+QNOZXHg+/nr
L7v1OlKyMN7ITquUdNOZZCpxDi5PVmpj4RMNsBmyiA71G7KXz2yNMhx4qJ/FAqnTh8lvvNswt6XG
+1rsVveMcfE61gBWdEKAA2X91i2kFLIW5kOM6BjVo5JUIqZwR7myNoAXIgGSbS0NXDF7f+jNbqq4
SV5rVWeQvUW705FV1DsBuMP/TaN3Ud9JLTTw0hkPCJHFmYJGjxvx/+71p9m8wL4aE5edzVMtorJ3
YsUcd00diLqvDRRAa922YnIlnOrfEKJ2Z7aJfe3wMDObzNZgXwuat0QInL4e7jRBFtsKRnmswe8p
bexmCTTYfynULREZHPgI6cmNrlFQ0AKcAFBCTTiYuuM2/eyJaz15xmPZ5HqwbEb7hS8qGVQJNi49
liPREyidVm1JXox0JAT+fLBNbeN5O5cGiuqBBPuyaYFqIZSltS/BDrpr8v7FJEnDkZgPALItMVa7
24ESnIOLpGOxBKSrYLC/4YLqEcUTPxKoT5I1hZtmu3sgEBCIJJCxX081/5ixU16QJnWPd556Qy3h
5cMZR6YLNln9kzQVEPPSs9nM5fMESWVmLoXkdlNyqBS39qbSc9i0pp/7Y+JjE5I5ZsH+ai3bmnSa
XesrZ1rtxzIeNJO9dWY27KPOxJqule96bXTanvBgGGW41rI1InV33ny6gpz/wILigTtzhsBVBpdv
tjie54nc0WEiS4M4t7ogVLy4DEHj1tj6UtTGmzVX7M6C04QPpV2ctOyXpZVdd/IRVhnh3YZDGE3p
Af5ePzG1m9UdIDYH2FLqpM+pkW0s9lkrJxHq5A/SyC+8ZO/xcPxLzSZoyyltPiH90NO+y/SkEnDQ
/I5TPLfJFtgu8sOkJxkaopkk+MpNCj2qYq1Et3LT1xUb68kZ88X35ZmSkTxdP5Bg1HarpV1gLoKt
HgO674CTfDKxhpAEXcniPK+ZGHTtix0u2b5wIm0panRqRMfW2KbpcKbe9rC6xGmDr4tWWeAD5WF1
WYFtGheu8JI+0dI2uaEU8MfRgh+ouAptkKcGrcpG/njZRZY0Ta8Gj+CNMeU71C8BGg5TNrNP1a+r
bRfZ3GF64VUD7skMIiuaMF/HImXpPSpxMeOcwpiVMs6Ad2Chsr/orMMC96WwXiP9NkbV4qo4c51Z
DJt5pqtdO1RygyB+jXvPF1IQatdVzBWQvvs8NMg+xZYNFg8/fSPmu0Yr6aLttpYFzyu4r7gG3bl+
jgIViSXfvU6pJ+pLt8JCZmo1hdkyILtCk4KlMdU4rOtc3Kh9Tca5gqkRRiIfPy+xOqd/HrfWOA5P
vYme4uxD2fCXCrtouWmUPKeZ51LBxmVIN0KoDzI2XyygMYoWnz21Q5qbgjPSM0cvdz6G/QEvVvMN
aynAWAH/vFc099/8w055UhDvx3MKoXPlxu42gFwsMV/KzwPUciBea6y3omoJXAdcJ1MZWwkHR5QF
WqfERZy3QSDH4VX+0BP61KXGrGi257V5/8NkzXsFBKOQXmBFLjvoYdYAFe1Qc89ECw8LDvhQhWZU
3HJ1C9cFXA+BPV4Ra+6H1c1WroPIeO/Z66Gc2+DmtGOzna9J29sNIUQGDfQrvInqipHD5QXFmK8W
7X4N/i9XMiI9xuSB3sY7dHgVyco1wcotLPdsyPVQ0aJYVqpcDiEjcM+ymFDXFNutPRgwStG9fDJp
tert8DWNELiqwQmx9XMB0xkl8ueyhRX4SJ179+CuCOJRbWoi5J8TtUOiVEAcTqMD8D8ZD65Shvh5
6A45Di237C0y1V3YDOUwdCpn3YMb+zqUUQrs4RAj+obtahWK8b8xwmSgxCxGGD3gVo957Dj5fsD+
U1osvtCAM5F0/GitZwlhz6BSaSCq1N1KKR3jTUS+3giaJxu48tiLEYaDbslHKoUWJ9FprWZnlJOl
jt3Lvl81/l68m2TJdcSSrQQ5ceqAddlmfY8hv9wdsT/KJzp9/aGwudU0C1jJJD1vTqMqLukuFNHa
eKjKdbpBrUqp7sCG77GeZ9bTRN6lscbJQ2G2g79F6HA8W4B0fJ96UPO/dtB7GN0Mzo24o6wI6Pe3
nMMOCiiQpEWvafRyXFUJmbRyuSbtprsdYwMD1DZ3Xn6QvzW+j24aYd7alMb8epKJdNlxAua4wDok
LhY0FrGJCHgV9gcco6OneE0yb31Jwi52NGOzH/7lfSTK9UgRW2S8wvYLGC4uRfqSAiSYzhY/mkLa
e2zoToGhyMTdqeoFzq5lf/ZKQ+dj3FXQpZGScPyO4ooNxWUvqhvquD/cXeU/JrSKfxT4haGMwmED
CADzFtpcGqKLDQ6qcmUvenTWN2+kDp5lGrMnjghhWTknCYTFxnC9V1SLqLDgPqofSsuz2ec2nBNA
w8ojEGWG0SIEyEUMmFI9tSBXGaqrcfoSQlEtaHMaELgcWmo7IXljR1BLFIs/OwHZj6rOf8Kx6162
TaTva0Jj8OT9qjkfLAmL73pXUhKwWgH3iG2gSKspcPCbCp4SlRaHflHFNF9VDheSZKoZZbiUDson
eV/tRaV2JXjyXKzBaWQixY4TymGdru4oysPcws/nuCuTSFHnFnUF24eYnXM1XgLWGNxvc5XhqY8O
JCGqwUrOMZPEelGE8pBYGWSECU3/TAwlIjgVGN9+dT3dIjQBMXKMY2JWkdO2OuTbO1tv0zYflyq6
dBoBT2TnsoxMeO4BcP5OsKnxxF7pIG9gx/8A7SBsynuaDI6C0S01uTYWPaLh/BkzVDUuup40Ts1/
8OTUFmWcZ/xWAIP71hhWYoqZLlj/ncRQ35mwBcqk6VKqiJyAWBeOamD1d89xTmOrvGAWkDt02RsB
tL1qCQPAWpWN9jeVlAqfi5fbTrtbk7TBx0/T9hqEwCyEZrrN82X9kY/12vbaGBO2x3ejdBIGEm4O
/g6jfrPHg94wDRRJxNw0mRZ+3bkfq1lb1FSV5P7EGpmmY/RS/2p70xvn1ryuugfdaDZlB5aTWR94
zGSsAXhV3FincOHSIJK0V6l1epfjyuYAD7lw3fVkjEQuQGQy8DqBQEl+bZNVb8FrW/JSiNcoyqRS
aLemGrFVZSW64u9M2/J/V8eHR21zGjEFoSs3a4+3cySjUVMnninuW5tF/6qI4C9fz8eqtvfFBjom
rNstqujt+6V+0stF4kjsAB12etw2EL6Hf/CLHEArh5UAANnGBSmJqir5+i5yLcXnj+DkX6MMclPh
KVMkcwgQob7aKlhNFuRaU7TrG8ImbymsnJWSitBEdWsmJf8yY6+GEzis+epGTfmBLZCJhxYcJD7h
zZNBpy16UhkYlD/DQtSujXhtAF6jccaA6p5pzP7hIAwesBvGcXB9kjf4Ns+Cznli4snrD2uJxOGg
TSGDbHU5iSy3NGBbllvwhVixTGXBzFI8KojfSI1NGQ323mfbQe7zCedHuY6BwI+51bhr3jFY2Rvu
H6h+nwVOWgfFZBhxIlEDcat/J7KF4aqpXY/m0LNPzpNCqO9wDD63v9pZkYeajR4had/d7IIn/rjP
Lguc9F3c2D6NU4KucHTExACvkWyGtWr95BHY0HoRGrEhY3P3mxoygbn6MVxrZBvDu0vAL7GY5zIH
gImnHVdpaL9wBBMk0bEyW0eW+Jkoe+QbdJDWFgEOyW91GjejBQ6SFzDUNxqRV6a8L0OHiRwJ/s9i
BlqYv5DgVQqERX2oRq7Si565kArGbHO9NgADuK+x0e9kF5STQ1o7vgActXLkLYgJ52H4OFVPK4Ab
RhgaLD/jOXfsOE1XNciYzmjqfwqnhsNEQG2JMiVuiYvhJq99bV3n34Gfvn7sVh9M6CAcK4Lzj/Zu
EoGcM5fRNqHJHrm3SijxiO7o2RXg8EcT+g/rLgbw0E4JZSkKYYwvcy2qTyekmlzsNIpmw9Q1Rdkl
2h4dtHRq55pqK/ppC2kYx5hPAEhfJi/qadNZnFz76SCUg9p/WY4sDfcI3SumdD/4NekUCCH+0klm
p2XRMmGwc6CLm+Pd4uuxIjALo+OmnyyyC9vy/fCb10bga4BwHGSf8XNQtiX4eEx05An2BbWyFJ/R
aIIRdvYOXACEyK16jcp6WbJEw3I7knXsAj2BPRDwe1MOO2B04kMwrcHVlaaLLQYfpaQPA2Mlc06m
GKkAX6Ye3UKLQQjD1CPP85HOtpm5kM0y4NYEmtb0IzoscS/25FtrepxaSME5X1w1EKapfdge5MoO
2VgZgVlIYj65mYFHcAcjua/tunK+ZY1+4VSsyxv3wolrjooFQig8sNVVz93t/ciXrqK55NygcNq0
5UtcpNw/NlY7YuuRLPS51YTw+TpP2Iwzv4Bwry+otzOoGBqH0P8tByzqd/0TtJcnQpBvGdzAdeNL
j92xRUkuAEz3IWqzRKHA4RLbs8vhnrdPQckg9fM2BWyhk7fksHhvleiTP6wf5buw4JD0WT0aw46q
QB6CjFP+hjVYgjiTwYvaVassAjVEi9Gr+zsCGOU5IZn3UtzR8YFO9sAgSd7MpT+fbXA6nJeTVkDL
8dzW8OHFbO762KusxUtMQsp/uNz+F6+ASuIRUYeGTYbjNb30r8TH8cG1LeZRdsh8PrL6T927wN1b
uzToD/bwpbnjBsMT66mIiJeRUhLgH23lNH8+ld6rj+r0l2vrLZ3tTPvi5AsTJ7NKmqUWM3bbiyen
c4C3pSLfLtB1Hk4zv4TOqgF+ZPWKV7+3HKhJihNxw6u1ZTG4XwDDAl03SRwEQba1Uhtmoz21XYNB
wF3YMEL1JeggbeKyhPHQ1tYLP5A0OFW+gjPtbIvG57X2sBVMdXWMqYNJs5j0a2ttbFphsDv+12oS
LT5Z1qsK4Qah5/4GNgsGJt6fh73WEpjRPszjgZJvzsYeNIljN2Zi9Cq/TXcGrJ6y889AQrj8Edua
8ujq9OTRj+ewcJybT7shv6Rc7J9Ry2w6y07+CGWn6sD04yZkKbfA3NbwPTkdGMufMMbEjjnoyAZr
qrN6IT2pauJZkl1ciwTjDbjQefgDrWb4Pixc9ct8qgUtOXuG5PrVvTLNExPKoihuBAP3Dh/0iqBN
DfncmKSKYGEzQfTUEgNkQHqId+tIo+oFhPKP+gxD+B3PuKzgISxb4BBSm4h/zIhrVFCVenEHs0Ig
lcKeoHCN2YFAFLCWQ1Efw9s3IJNIrl7FfhWZJ7bsh/dP3/CpoLCP0PTpT0TNfYsDNo/8R1qTw1Dg
m/a/Hj2k8APWc+EOAsHypBOfp0uUCqNQe3LhsK/UB4J35bzkQ2Bgy/h82oR25P1ARuijyKWfIjzH
Q6/as6xrCEu8lvy3El0WIwRLIp0SBqbsabAkuSnD3wSHtuzo3vxGwebf7fuuADNySsjb6yDucOAR
8r0vrrWX3Bix50eBkiZP/g23kppPLD4DnUJPoVh2spOxwcyMoHp7oSCn4bRWPXX8bpm5V4Q7l5nj
RY8gWv+R1+Qg4f8W2tuop9DoZ6qiFeEbz1AJ08kWPxoUdydiUI86C9YO+/6id5vbiuDUj3f+Afla
qSy1g8IrMeqmgAiBT2JmVrvjK4+sTLan4tQYnkerXYQg15iF5zX4ceNSI19FLtXIonvInr9AOalR
nlMa+IyrZMh++oJmJ44+KwSUZh0UOKFmBpZiJ58zl06FZ6Y9A7x205rBXeqZhR/rXaEAIVlPMqTt
USO/ZKbPPfpp0+w5z2mAdbiMYCbRG8nKRHvEAZpapCa96qD3giJ2Hg2koQdIDCoSDFUMQPe9SZSP
qTPm3i/hfhEdF3pDbgcPK2pdR70ZzNAC9d0+onmrAe7Gai4WxJatn8wg641jQCSMw9TrjdKF2f8y
uoxjBcoD35AARI1bu1c9OLuS7uKQ+SEwJk16GjqvCVAh6NEdlfWkwx7J3k65EYQkO2x3XkveKuMk
OIhixLhIZY39Cqz5/gqGroGS7PdHEMMtzKzMBkbig445M1xenV1+rtd5INGh59sQ19iYVWOiLD94
SOH+81rRCZIGxjP86uaNbsSyXBssAVpYtfaW9KLQEw+X3csVR6Jy48/59gRNLcOR/5AsbaU73TDP
sYKac3yFOXlAnS7dUzpMcp0rCu1eFokMe4qp4nQO7d1O32eDLrtK/vFukEw38civj+90Q+CoLrK9
i+pRdDKIVZ0CCvoGONK2uaQZLYvtfermq6SkViaBOfrDSrEqTHXwl6/j5ykDuCTn/0VOhEkZ0Lal
DpaRxq/1vuS6RMoqGAfi9d9XEXVDEbjHSasHtnpCpsnleKt7L4Ouj0A+AiWticfGvljauZLq3le1
TxvDaPKu0d5BCQSW683R+HD4/Px+R4xmuNtiduK3Nl0gMoFnf/5MQ1E+hhM2ao/63IT3mYYSc+ut
fyAej/3RxUA+cqPDN6ZmtS6ztWEJm0GmxY5izuZ0+WsJLPRq2VhVtpC1nf8QT0RP1f2bY22PQcfC
k+byrM+3pwXgMllHXzCEeNXtWg/Vp5fMg2J251/10gpltUCwK6IqnkU4vEEY8Dsr31SA6mynbcsp
vbOSscxn/2jHePximPBKB72c/WEwVPfIBMoRK3IdyM31nwAIzSslFBgkVoaPfbxpo3Juupt5Iyyp
zmjdGGbuVGIWHY5gfX5Nl0fVWwPbLbTwj1cMf1wVTpw8tN8oTgRqeJKz4Na9jfqhwIx+HwdBKHwD
ndjTHG34SRwOFYpMMBCjdOdgHBITfPT+U+J+n9IlxpaxFm1R/mhIJtQiW5AJZRNoZosL/gfmq4DY
3R6Up66HxAhVZYCk+sOXJod1UYWdOa5QzwzPM0AAPz/DS7WriecGcfazG2BLHqd8gI+tJZOTi85S
68z+pFgP7mYTP+1O6tWH1hYGJMdOnBQMOs6UH/WZ9mpZtcE3+wUydh5bdJ1t/Ly0kW3NvJtiG6T4
es1EiiVF/7+BNwl3m1t+3acLIZpiCWHxSPKEd649IR4c8jLljyvgB1FYa1Ex7Ju502kKAkd6CR26
XyODesSZlf/sWIvi9ptkcxUweqTxojA13o4cdW1ZKxB4y4vXsTsjkoHOh1nUOcXz/uq/sV8DWWdt
9kjSYJpMJ24aTtMCG0jb24jt8p+AZehrbMfTJOLXulu2ZF+z5Y4cYLV/wLwqF8bsuJieJUSDdnob
Dk8dkRow1qx4XCqm3GkOFbwblgmPpKeF6CD6gAtZGPHAdMl/tprCdClmy2kYn4fIYpNcyoISnzZS
bElDYgUYl4gITQJQ0h5f9z2Y9na4qhxNGMXoIQuZi3OSC9vVVUUtOQcWRQf6r9NbU6x9/SwJzAMV
x3q5UqVpiIOoSK0tqHgexK2QzysWW6SA1zyB0cVeo3y0/Dy1rkNhquEjtoek1fa9pp47TlT+NXU6
sH96QhD1HdSSKAHuTsN/l+ni16EmaBbQKC0QUlzBbVTLmMVjQjDhgq3xz4ccjQIGwBT2jL8ulAku
lDYHqTgjPtw4LFSIFC0f1xxegUaVz6gvqXdmY7OLUZOjxbmumNeSf93Vt/enXuz7vplSGlXxlEn8
CdKVi3/GYyd20KEc+r/Tm51RWuAlZVMdL2D9ck+hL6ld5S5xB8ugghTtpemAInEUto2ciVaWa5ks
Lc2cbcrW0GGW9JJWaTjcJpnDSCGSWFZ09++pJqKfJOPEI4KJ3v6z2gYWkVsvY+FdF51zp3F0WHuX
AwZbE1v1SLAjIlOdsvroFsCmYTPxHMehitIGqddvJO41JQCDyZDylhI0s0FNSYsWA/Lqm4qTA7gA
7rGyvzLxaC8peZCroZ41xO3HFGgaS1GVuFiMfyrVCGGsLJqyge3iy9EWitSDbwRguB2IiVoONWWL
xsOwhOMhVc7t7BHh1YB1UdKxORTNekEYevJOKnmaQTOsIYbXpS6sZrft80zi9nwqY/XQWozN05w3
qi+s07tetbs6/srxiP3OM/f0Is5wHx3xU0NsE7i4U2VioaGV6ADaA3OpN8PdpIfKbIMtL6gUcx8j
uDwSp2wPM8A2/zA0HBIOyLHaiYSDlc1N11I0gdxEF0AGHUl04fYvLHOOzDxXvUdyOHgQDmZqXaQO
S4a+BVs8VGM9Qi1y9BXgkcnoQTvPTXo+3qG9CrnvSvdO1jTLP4hVmbn9k2gf4Mj2hO7ygAVCsboX
23sLlqOD1wVDBaS8HZHe3J8wiqq/W4qTWHPbaKItpbArNtmvBM3NrKhd3QMvxqT4NKIzpPjWC4RC
Dl8CU3Sl0V9GC7KB5sTuCiCKaCCU1YruJDbMwyPgyQi2duNZftpO6+DE0b1B24z2ht085oGzjidi
vnEIU2WWrmL2ZlQwSlNujU9FMKrCKHtSfyObodULavpMyJf/Uz6q35+89bCmjH/B91/MjHXA4lmo
I7Jx3ctW4bl8Qogt5jSNT45TfS6M2MbrLffNMNY7yXx1LsyPK/kf9UocyB814eG0Kpa4O3PIZn09
5mvBCcyt7De9jgoL/ttjC5X/kNG6ig81HH+HQ82XQ++8NlTGj51siDPB5eF5D1lZgkvHi6EQLEoJ
akTXm7ZdVd5PZ6+5N6/hWnp/AajhpDSyDruVC8Rhfv7soDxzgshFs+zb2Uov9U1kVXc7mWAu7zQ+
sOi7OIxupUKOfYQsPbhl9/GdBZ/qaYGB1CbT690eQmiY2k7gKh7xRGHSI8R8AKYv3YHJYF/MZ0Og
XCFkdZVnlWMv5GlvriSWqzmCU1pDpFFcNk5qdzttDEgqXRFfIEK+yrS8kBVepngDGsIL/j9E0Umk
/n+6YNnYOTu8a6PIOiU4Uu3zFdYRV/zR9Sihou/p1QyrJj0Rob0fbZjoVy1QsrYgxtnov9dJeAnw
8CTBeMw/YeTDvDy7N0fr3DYA9iqo64RbZlI25raXrJA3CdtFeZuv75v4ejUd6673Hlw9vr+iAaAf
GDPgp/V3fjvrSK+2w0pf7WyW6ETI0RaPgQ1eKxNEQ0Hdo6B93odZ6D3ZYh+dDoIJzS+iwUroSZvC
1HnXWb4NvVGkbroyYvCnPMCLp7Jx5t99Kyx3Zx7NTnczXy6ytDRdgF+fI9gh7mNQViwftPc47fxh
X9cmP9tg2jrrxtuYI3bGZbfGjfGGuIUGgqS2nVXpTq0y8isnr30Dw+scsWmq+D8Lm9Kyooohn+L/
UVa0ueD0pEnwUUW4VaTpP5EkG8C0RZFNj46eRqQMBdDF73Zx0zSSCziyF6q5y0a0lPVJJFoXU1Ih
J33UrZuTeD+akPWpYT9GOfRajyC2rzblDMvdIX1SUsttj1hh9YPeEKMD6WR5yScxnuuzXZ6NDVsk
EeaLxeDNe2lyp0Cig/TgiYobY4qjcTtQc1HvYURqiLRv17kgvuWsgBKTsfNENBMfRFCE0kK391uu
YDAvdy28rGnT6N0hwsVS83dE/5DIK/92CjpnaVEVJOZYmxtfSElTg3iz/+TSPn5IUMpb5avkCMEn
GzNCT8P0F51rRdt6jP8lOE+edPFBerIJozpjOBIqKBV8ZCOf6KxjPFhyYaeHx6XmbIxJNv3bUY1u
kBrlyJB1Xd6Yvi9MAfLnb6Vo5r11Ss7ByZHhkQgvSZpqFOaCdp/6nTZiRHIwk0YvaCTE+jAOBLae
vCK3i9u4e9C6+61QWzWouypwK/x/ZW/GrbQJEt/pU6RAR1UgahfZdu14JWf1eg6ylsfdn7qsKUee
s3yGpp82oZsELoM2S9ZM7P/VVDj3o7/TEEFqHmn1l82HGwDab2FD4FTbqFZTmBpPJguhPK1zdLCm
uJhDYnnRKTnolHLP+KKYs0syGEQ38nrUkB+VUt9rAHANDxZKHQiFJwM16/Mk2VsWAZeBvw6MgNoe
sKDK1MLi/S2w+XW3QrdAADsCRjdphXr7qr16CfAt4PtpX1v0dn2P7E6aiQRpo8qrZ6emQS3wFzLb
a45L60f7f1sWz2rqsOJHKr7mjHk2rKK0ww8qCMurwOlZf9xYtVeaUuqlzfc2bGusMR9Wp1MKI0JC
bqpjYhqhp27mwiz6rRc7b64Yqnk59lj2QokSLrLHtO8197OSFTd9bz9IngPlR9hEUDCFyV1ZVPiB
2f0mzVPSoIN5NZp91XCDiV7pwUCuw9SsmVmcUh3YCX3QCnkpT1dlNDR1fAhddbE+4cpnHGAkAI9r
+ydJvffglVmcvKiGoRpPE5c2B0cf8KFDX/ECKZYdwlQWdZYqn/eE34P9cs68AbjUgnSK33UXsmSL
3wqHhBOoUYPKcCSKZzVvfXt18sNyCBTxTrvz7+yRsUouvKPYU2CVPpG+0Im1QA6DmI57ZCgtPck2
koFVwE4LG+V5oZDZaMATaxnCu7OqmKiReov9PHwsdusXDkQgDTs0Fvm8pFCzQPlbIuHZWasu3obO
GlQ9QD98y3fq7TPaRFfCshnrwFVd2mIG9tUBgT6rGURw6nsyxRSd+Rx/3P5ldcsIFwLO3oLWHcqY
FPSvdFOvgJbsX1z0qrhjJ3pmI6D7uafqdFv8b5aVvAbJPpsDkWKjIf4X5y4RuJfXjVaim/qzl8cg
Ay/8VK3yJIALnxd1eFLKtCPA2gQgIjgn6J0oVHWaI/wpPrshwH6XEHePKpuFD8fVh4ULLbgxe9hu
iaTtbLcCl0/MRttUNnC4/IMSCaLG+OMrU1c9N+A887JfAoT8SPTcU/nZ1TNtlJcSUnsJRJWLJ9Kb
t2QkYj8JI46Rn85olLFYaSAgltkrh+DlNK5f0tlSlCfJpEMkovypFVXRBuvdLK+n4p5oN/a7dmnt
fz4DnvDTQOz/qus77bjpLJF/4yExgVY12FqkSyuvfoPTF96ouk/qyHJH9aZdPyzCc/qiYN6pOd4C
BidCnXraQpWQQHhkVw6ShEOK5X8yzsLjr5yk4C2tw/ssPxCF9VgeAfuTYlFC37by0/yLuVM4y8ot
csRxyRM3yWFys8DFX/+4x/oEB4M5oOT4D02mbiYXKdzuvEK6z6bBfX+/SOPNHi5leHFlcwM1y0lg
78EEPgTv6Ia8IRhdl47jBTvT5xHaRVF/2YzB9FYVQtxjZ5mbyQOPIn+TSLP1sUHy2Mhf+T1tz5oO
I714fyhMLZBRPlD1y2l5dMJy4/9zd9dDA4ZlCjH3SM9s1zbQzgNCIEl7OmvnYVBLR9u1PpZeJDCH
UgyE1yc4GLGRO3TAt8Gd4aAIbtoTUJH7B6O7ts/vKfQBwis/cVZ5hdmWFV6xYdfPMB+Zh0Sx0CeJ
/IR/6ncZjRhRyDjY3td5VdlDHyi6X91Lr/K1iR17B4/TO/73AVQOdD01YDiyvTu9LAX8f4cE92kZ
Iv66CEv4ZehvUTotW5B/FMiJstr7xjBDXhNZgcmgVlMy9kAhWF93FVDWRMX3njyTYs9e3h87y9JK
50fkWt+38pjnl4gtC0Ag5Wrbg86/AaELyuSwirpeZiz/sb8fqmTzHWOve4S6rFVeDEm4F+cLcZEx
YB5Xj3EvXxaFs9hG9l7nEOiyBEVjGLwT07I1mf7AZUrHT+glRS8Q+PTHT6UWnK8Z6wY+/XS9pH2q
150O5eP4MVAcox8WIIxmz3c3UzHQKcuG/h3u/qjbSP8lDcja2TsR++GLlCEeCsKQuY8KqqGIUZun
f+zgQTh+maHQtPPzFvqAy4ixVxuLbvj4D0inOqjAdfeTmApNrc4oTMk91D1zLfxIkMTMd61hfs0k
B/qfltIvqDErzmi53qS4QhoFsevliDztsp6qDjcOQ0zqCn/EKK3TJNK6iAT1U61lhDCyiphbYorQ
3n2DElcm+2oav12H2cJGFiiYE+V2qaa6I4dHra+KbsUJM2sxjnAFo/0+DbB3iHHGcLVmTEBmoGD7
85owIRkMrMegaCnMntgchy2ICtYaVgDCrAuA8omli8YEut2OpYZ0yzbQq/HrIbXIZ4o7KiPareQM
xM+sicoIzGKtFwhtIQpIUQHps9ESdENExi8Q433XCiov1bsW8FvCORepa9Tmy8e0TA2VfA+uAt1H
HTvD7HRa90FcTEyhJ552Q5TNxSuqj2GOn7+W33Hp+SYJ5DeyP108sHuw0vcoi3bTwM5fqrPPLkgF
++6r/h/po87/NPqg+/nYpT+5BZB462RaStqQ3V71DvMTPqDizLbXT19C8F3EX2KF/NXR2Cwjog3/
KUrFMPicjN7C5chd9hA2HfocU09SoxcGaRk0KY/XjKsWGG2hKxMtTEJEfwXJ+5fszqJrIDXnXZle
Xqqb+oS2sCf9fdslwvlEbuuQnYhIx+Emmj+VRa3aEQfiN49auRfT8c5dYV1fh0c9RkMO9dXloSjV
inEsm4usZ4zqxwGHLD4J5X2tyDuBGxY0eB5wnXvTNBYKr9Sbme2+vRStsuyAUtiKslJeq5h9HncJ
58JgoMVo+YuOooU/PsUzYo3peDnLb4ycCoa9IqNTFiZ8Q8KJia6Dwk0KeF9F9toGZwyL/EzM99Rp
Z5r4uW76mg8cCi3ubp3oXudPbgTwlEO1SSWVclLujRODhzIKcKPWrqWkFoNvSrHt7eL3oZAF5KLD
GsNOK5HeKt+bEmem7hyiuCTmQ8KnG+5S1V1daDZ+/eTDFPX9ohP8LqeF/weaJH0N1aNR0t9xXN3c
VNR2RgEfLdUVL7DykESjyaLi+yoNEQ+shBb3Pqls0SNz2RnOl7YgXdOB08A4Ymtg1i1MOQ2xlSb7
7c3GqPiTV1ZvDkENRzA50ZyK9Rb9Xq6V6Xtpl6Wq1j+/MxAIlR35VaJjEpn5E0EEVG8kJHODzpBc
jY88AlINKt3DhELtuvxZJ73CVnRkLjIHfOwY8/Ob9tqFFdDH1KGH2UdRi3rjXCzKlgEwe6JcRVIP
CV5dW51ldCVSGYmvds9RoLfH43jJgeXgF0DBVxiys9XVXO5rhTSYPW+7EqN/Wb/IlwxOKwm72yBw
l3AHUVGaPU1rwwlqgfBGoovHGTbcNjL7xDj/9eV6bF6/82t7wkuNBt4N66k3c9WeXkc21GvFc5ym
BTIYu/yO5IogZVJxlI9q9AhEDTtbyXJCgKFaCnIaDg8eidnqz6NG5cmX7jYwDUzAapIXm6upFQRW
a+aG1JszEu0vTt+Wxg3+k1lZGlTS42cIUYpZ4ZUMVrcb3gaaENCyule/C0J4YF0o8w9txfLmHES/
h8pQffGnuJc5JheYs0T1t7dBfk6jAqlaQh8jnMkb1Uz/VzYSzS4g5gGN6C8ztHCb4C5fRLeEcjRU
JwPFblNfNMY7eiSX7QaT8T2VArmFjEKEbHh9uArvjDN/7xaT8dA1NdtgVPGRyDbBjwL61OJ2KpzC
UiAadY7wqajVbDXrRZaGXEaVQvobtoBQIGOcyIpO1GvvdJJ9CrTvMSjrZPJo9JB/aJfAzNvcWlZI
ZKDInK0KaJcRAaAgDVNSLVpjGYqTmKLtpqqF4eJRBgfiCmjileQKNhoLLygNhBs1gLsCpKqwiu0H
ogV1hMcvWaaf8eYVvHG2dSBn4eGm7q+2rM5t4T57wb8Gbkh3FJ3+zBqll0JHeBNx855nsy8xcf7r
S777bl46QABsSsCoTrJkghJyIHz/pQwIYeg6dg7ZWuxmOb9degR3sT4wb0F5QmXZY2wQhPnvuJcz
PqFWJKKtMOt5YgpwpIRzZfxherSZv668HVZqGh+6mjsz5exKuCAzDEJi0P9zM2KAsyI/JPg++/tW
TPiZvT+sno4oEQG3HfPCXLKbh3Ke8M9xS1Y+OgD2xOoLzl518OcCcrk/JOiIxov2c0CnYU717tX8
oJM/IS6F9Yyh5t/xt0RHEwYX4ZCOObAdM72jBIFgpE+y7CTs4A6lhHfqc03aTuDecdktFEpNbcyk
34p0PqYM3kuhifv+KKAca5vuC5X7I7KQH2EFMsnJwPRr95DsrzX2T346s3DwWw7u8kQ81TaPMxX+
ckwQeKIeqGRLdQ+o6srHOg39iujsvrlqQkBe4OQOuPkEJMBCdKIRd9W5oCl2G6WqiCQlb3vxu208
5Unrx4P16MF4MEhsz69vamzQbrwLcVpaeE2PphO0uNnJybRCVcUVAlAV54HY0YP+tNFJR8WlsPIE
bnO6Pknt/9bMB7r4cdG/hoJFYedcFJrHW1g9AzzeuFIwef+4qVKmRJl0Gfsa8P9W7tafUtWGb13G
T+PDPY2hHu2hYdI2arttzh1YX0q16EIUzTWRzPkTeSyTKscxPCF0wkDql8lwB7yu53EDMtk4IRfF
vNS81j6TJu8zgXWRVpMiKJK9L/nzvh5hNoQDzaKfg8V86QtNMDbbTM7+EM4WpBDJp2IsNZnqsIGd
vLFGZutQcupwtwNQZ/0BIOj1lOObIQz4vTIFCoi3rrM0rThO2dVwlOq7Ck0z0u2/akzw2RQgPQ36
sLklgka77Rxlv48ebm+sSpYh7fdFxFEOygnmRRCsHAT5KnY96VJX1K4nSeSp2sUehdGFxd0Mm2Sw
9eOzjuBXpwkHg4OJZBaZQlP3iM/eC8xrMBUoHM6WI4T9o69dW6zS9YhnrgY//rQm4S2ZFWDoDjYk
vvmmroLDXYQovLoV+x5dYOs/8+PVNrZv2h6hgteXS6prHFZ0TCsn3z7Dyk8QIbVV8OaIiGs8srNt
a3cMRituutUPKTGzhaZaA980I2DzNGdcwSgRHctycuUaV9dg2dyBl5I/l0aoeohahdpWSwEsCJWQ
ob7e7xt2QqgZHccrVX696isQMMdaylhbdCIZj7NMQEbeNw4EVYCvtB9E86mHVpUEFORhzhsgez6S
ShChky6b05HJLHplQZiGEAr0iIi4AdaBx1LIkpLlvUbfXXPf5ueGJchSk/WBy58cJu28KM9wBZZj
J4CSpzas4x1vd3mdEnh8sw2kK3PbFOG14YEaCb451KEq8eFf1rcLzVKagE38XOjEBuQVoKf52C/d
76kO0qq9uLPCn4teP6P9QxvS5Kg88iS/xUGQ/oqvHdUBorQX6Y7tPwZAmRJoHfKRYsGFObtNMN46
DZ/Z37BbMgishfkaSVr8t9PbX0XMp0CqMarDrNgy9M8Db0rv3fwe/JHfynJDlwSOJAgW4cNpo17J
d5LheldfkrZu0wWMu7aX6+PTxi3ivtLx/U/Yw8fZNsRqvkk5n49ihyocvvpzYrs4XQcCe6Hi1Zmn
EUKwdKmf994oBq0JpjfUrLs104nMCiLd0yLb4ervcGiJp7lm8JM81PPBGtxTsr4D4yF/2BF4rk7W
jPiXVsXTaTreWPqKOOPVndcK0SmMt2xE4AqSwoC8ED85dLYKnzSew46a8Xo4uzvli7cSgo9y0CO5
H2ItxKZjhlw/ximpNGx9um2dcuxicphOdDrfFcUCJuFvNF4JdOc5SRqWzrJlUvg1C0CMJaAM6Ds6
yr/POV4CUt1SzctypC1P0baF6cWfsPG2ATVHqpAT1CqGQ9VeKGko7joO6QwJoT2fwH4ORyUC/JjK
Dc+/+n1LwGlJOlJfOwbBWvBzb9UGgM3GVNQgeOKPR4+w7y3xnRYrbwIWf41rcLV6pVTJIpYzXVrA
LWiujXSzG9FWzP0p736xwFvqaURhUkTccKDNA8MX7L7FTFB4vvJ6SaASINunCSGOEVlzlH6hncta
fiNikGgjV5kwIYBcbTtcStTs0NcVYjlIIfVtP2W2qIG8QwlVaCQuVz1XRVyJN7Fo4P/HC50WpVIq
F9kdhCS5ixn8xapxPQhDPlq9eTTP15tBWwYqsDlgJXhJxqpZTU3CY3XbloD/CHKBgrwlHrE99YQh
WZNmXJ5FV/+Fzsz7u/Elap4pZfV9nTSw5qlDhGnA+fgrJ7OQ4hCBkegopLdHT4D9gyhcimSI6yZz
vwjTeR8FdlY11FZH4A6KeuCp4to3GoOAzoV7aqbDhi6tvBug52HbO26oJqU3w/zWhxucKVLKzwvV
JfbK/XhVmYtjwX6dJMaNnelQgmGMZ5Ftb6SvJUGr3THNwiPKi6itQlEBaqgPNAOeqeQl3MW0d67t
8zoS93Cwnq55N1ix+BTH19zwKvKkc4pFZG8vNxqa0Dz2L7OgAhvNBchsjOknbHr9K5TsgcQHvGBk
+Ee4Mg6xk6cz+yCA9ymFpPq//8njXk5VYqNjUUN6jf/USTsyQA6KsMxC691LwWheOKMVTzNbkIsl
w8le32gZ0Dw/fpBxwjYVwq6u9L+SMx0W90KExm7r+5lauuOw9vMvj7egNQj+Pg1FdWpqp+4Ofe25
IFVL6Fq5pEWzngGpGt7n8m1pIBAgYFfxzt4ciRst0vakJNonxnPUe+CQy6gT44A6z5quCmUxTsf3
jUwqvJ8MHkG2IFyUWiE9HfadNBBluP7pcAaqtk4JVSsq8wljymXn7xVGK4Y5DTNENBC9GqY1exT6
BA6Ul/IorsFfauLYNtnRHM5cd2xuVhk/pYpXTB0/VNHLAt7nYMeWrXUhG+DMgYzYrNRqVZduKoV1
DiTI0GG7E2T4YiuTiKHixWjlhlc057T254qyxdP0Gj9TtUClCKp5GiNSZ5R4N1LhwDbvuuYeVBsw
Cp9L+EbXQtrvyt+iecS4uwCGnm1Cq+qUFMrpDYXZxV5XgNmczs+RNNvh+EPc4HIprMEAgSV6CRf5
axq+lgF7S2VJumSkH+x6q4gvtLqmyeEhEnDB9s4J47fpVzY1/c8l/bB+DHEhFP3YQI9k/6O5lJEH
/fQBnt2KJoRTFv4j98FfhoRZXi6XYgYFeLyA9ZoIfEkSYMeTqvR2IJf2jm9xCWPIrhw10BoKkRf6
61cyfAEx6a/PKEW+EPse7aArR0jORi/4b2+NBvtxesLLmmd+lf2sqXeSLZfoqibGbqZ0geNEhs8a
lJ9WXdAQ8oWxEX36OcWgh8osP2y1xNGHOqkWtdHQAjvHw90ypyqReFMP7QZmqjlE+1Lgt7ImVINa
yy1luri9tESK2TPy4+q6Y2A68tI6Rj0holNH1RvdImijhHDxe4MiZm3Y28kr6x0UjjeLN2mjwds2
bFnmbMr+yZKikcPLrMmsgBgkOrshtLg+t65hz5zuCRpD4nuLockl/dB4+woGaEoC43Q/YCWrNHLs
AjlR/kjjoxV1l30DfiUn1xRMv3bKevYsW+81Ch6FtJzN4TbssAL9/P1tT9MgqhUqDD1kx0rk4wGO
wrGRycYkb7UWAYhnvS7xKOqM01gNQOaKWhZx0pvhdAqT/41i/0x0g9wIa7sANLyKMWe6vqvDaHV5
fVzaUrKG/7b//jagg+7+NmMowusUY4zniV9JDQIGL5XocrDoOCivOFLz1lJ7M6CZqBd8eDjXq1Fq
bB/fg3m23IwWyA03PhHLKlUWP2x1bB3bSWUbNPNxaAAh3QDygMSo/pz+wBNPp2HDWcd+hLEVxj/G
5MGQk396MRHm9Dc8G6LJwrmgV1grgwwjPvhQkjNzXFSnBHAm3Ne/NFyPhrYzTpDLudLcXA+eQ6Vg
z762kQaU8/QP50B5RhmVY7w/yT3SWSm1/MScMdS3LQohnwVKEPc4o8D2f/7G0K5p4dokIr28NNb/
/MRfqXhfkInk3cJhhiJJYXYiHAZWSnQlDh5sKelKASiByFXag4Do/UWzVbosBNTlXDYIgtFTUZsX
gXRUudseLvt+bD+luEvA5zFmiqI3418Ap9NkkW108Ne9ip6k29gkardtWlzSQOO+5BVKlZVmsM+w
6XcwocRzKdQE6ity9NuIOXu6LrNOYwhRJTBM4IrOnFKpfLAiYHJNSjSDWM75pd9PrrUVElyB5xOB
q1Frb6kgWykJkjG64IE1AG1vGin1j7gpcxTYdBnf3e4wXJDmVN9tYq3Z4FXWFSC2NKG9eKG++54S
Wva8AjEC0uOV/80thhG/UmpT6Q4cqMHTQMfm+VHNXi/b7qf0aJ8SdHylo3eS5/2ZWn64VS08bO1H
XS6Xx/OrvcwdeqPi/B5swlQ4fFJnXMjFF2oCciw+agN4tZnuvOelz+OmiJQ6aMmmgB/UzgZq4/qH
et8BzSvs/dFcAzblsPkUhfqrL5/pCAdgGKei5ndohpis+rG7TIKSIPAIra6zi/kU7sBfFoLgyI0e
rPH5tK2tQ5/NDVsMPn9rf1lQRqxOoEYu+sn3WziKFFdJ9HKyYaLvLbMn7ZzTXvT71Jjkqpp/Swr2
HPVCaBWo2US2qAEKlTjlcnr4dAREg8vkOm7WO+K07IYgQZFIjrOAz2X0p8YjJevuOCpaBzPeORHa
efH9xJXYNx0INuGa7qY70/FRBe4jQs3H5IK4niCzBHKYMHSrRHS9Ak3dRDCCkBmDN8rwZywg31Ce
bSHlKONz165/Z6RFpMi27LvakpFAxNeZs2p8OPzC1OYf+nu2nZGdzZ8gaZimZ6i0FfVpbG0kkCi6
7CNs4rfeedjWKZeGkx8y7oE0963lzuiGi5jSFAkugawMQTQpyM0vWAAjmC5gnFcKml/Ovtj4zrZZ
q8uULZPAEY5k2Ppz+bHx6Gz+qZwnoTD6qpFRH3Ssc/PGFwI9o/T6BgAQB6gy8judXGtWaHpcBd+H
Kb5xcbuKCaA4EMmSNWmV7TNqVaDB6vj3hRunBH6Dyfx73tNNNfSaPmVN+3vAgfDr/s+DD3iYV1NH
d/VO8STz1nSQshnc9l8Qhtp9freVksQRC6nnrsDm8JBwYrbGxPXz/WxdkWjI1XzaZObhKwIkwAYA
z9m8IIzomihFVGJwWlbvchES1aUiS7YH5kL08jMzXNshLk7I+osPDXUYaDp0kOsjpoIFoEvtBHb6
ujD3Y6iC/hbftrClH3vVf5GK8aLYvSx7bqKcivh6RziJ3L14UNlgmkVM+rSXuGfrMZGmrQ3f8WXa
+TGS17Lsq6gmGSyxsGcu5KbgE7z67kEjToZF04Xetw6z2uCjqbQMQ9RblaOu7wqqgWZCALsWXkdD
Yn/lr8/xwjCl05SPv8xbGXyXHtyyArlIUUJsXLJ9DWaYSEmmDNVE8DQJpeVjdegtjFHrhi0y822S
c9xrN5MNGq5R1Je86Bqe4v/UVrfzvhN3Aw4/2C6/toQYG/qAPMtA9l5K8CZBpbXnN1VfpRlgiKGH
ed0PZbz/J5X+ospcGORPqa+CZGXR/O/dY1bjr/HDwkQFuxZGIk4Lqm7KREf+xzhelXt4eWK2ssPK
++zicul+zWfxa86CjeVFFHWEf/QpbduorkfibKk8B6cl6HX8gI8VjO6tErwlHeGkX59KVVw4TDE4
7LP91r578s7u0xTdetTMSiXRD/NaGOmj2pXOZwE8jh+ZHdBU3c7Cwz059RGz9yc9vyZaKeIKUXcV
3woN2EflJnGvSgAIvAFyrNwencJknrvLCc5444lbHcFOz7M45PKJGRbhBVsTihaC0cLW+WjVrKdq
PKWQjHgg3JpvKJHj+m8nQlT62Bz6m98VOZfJa3WY5l5/U9URXD6s++TsTSGLNOCEynTIHXmhbDsu
QA44EWPUfUc6cZIbQhci2fr/+wUUkU2zDpcdUDrSspbJNMm7fT8+xr8oO5XOCCk5xwrXy8BIJw6k
VJ0bQwyfLIWePnCuw/e17hKktQm5BswWOIikWiITae/Zk8hoSd1d+sYy8C6ZSngS9LE6e9Q/i+ig
KfppJggpH4mK/l8Wn/BrxHheSXwuovSTLfV8i6JMYp0D1s1+tZErV3+J5VcuNhJlzHwWaLeTfRyP
/fwOdRxP27ITu2DDVr1B5qncPNqu8zEmiH4KQM4LbEwC/9gXKgX6D0UNFNmYi7z2rPhaG3EJefkn
7vB0WgbHq8WZ50K0OBXjwqW0OWLKDaxSEnmiSlYEC7oePfEotWN1imp1pJpi/KzZH/ZLM8q6XUzi
LiKNmiuZCMiMR+sfbpXjcIGg0cv4G3EBxUcyJ+glxn8/hW2QGNEWveX2y5x1ddst8dDD8PK1h7Pf
WaFVtNNlBRClU1KZtXzFIcM0HpgDko0z86gEt+OcbdDm1yebuUJoCaxUoc4h9mru6VPDW3ZMt9wP
kzu/z0+uzTZ5wMM9vmVBHIsMpCHztY1aK1s5SFNhdigqlbita9dZ8lTCn5gAINbU7LayrwTPrfZt
S/JidxHjX81vTqDVlmADsIdSE/r5JNmfkjMyUk0mBCVtW+q8lS80XQ+ASCBtvvO/ptS2nN6h1Qfb
LGy/oE9obiLMI4qYBU+OaNA9iKdXcbuL66or0ObT6cGrh3Cw+bLw5pSOmF6cS0SEiGMWDGtuauiL
bdfmYGwsSPfh/I6GTFJTJxLlLMarYTkMIeCSWS87dEQWNmayeFsm1sjmjvNdeO6g+J24YpwDKMD2
qb1+TjpaEKBis1rb3CwvaaqybtfdfhvV0RDFFRoNXr3NixPwh7CavzdqZRfj1/+DB9eAhX/62MUd
v8sebgBSVsY+2SYIzdYC15GYbuH9xUqNvRDST8bV9aMtFyN4cMxfYmIvSKVCqQn56qxnoQMqfYGT
hjTdJ6nSmZ5TlShF3CWN3vi87k94zyB7lQhn94MOeqL/G+54t3CLcPtN9SQPmK6px2WYNOc3mniS
u5w0rRc6E8aewECyrsKXkUjo7dVn8pgc9t4BGA5IixV50wpzekLspMMYCg0G1aM9B5FhX7qjU41v
dmsQTP71VTm6us7KUKe8CsAqHbyIRVyY1I5s5Fhef3w/5WYZTkPIzWMyZSDMRFRkmrWEMnlCG7ix
SgO6r+s7ymlWfiroHg5HRY7/uzWagniCLnJvVImsh6MIJAEhIFUt7iWG7togMwCWIIKQ2qDDOqyD
N+PGQhFgnTqDDf06D1vC72eORlr9amsjlCW7D/tJaXD+2bALvMZtydQUSPXw2vjxljvl4ASFOIF3
mWiKVtWtKpRilQ3W1SkKXZ5ggV2nbQpNAUBQMvWal9i67DuOaPpaTausjVW96m0nsQ7uAydv8tSc
Pekd6Ndg+WSWBkbgonx9s3JnXYjXpgTrNy57YJkWNkQG6hB+C3ViFYcdespRp4s5/OyvydrAU1Be
FNJvD6/s71BRyQ2e+4/37ycuSbJyfdIvWmnE7cZCVi++8mncl7Tz0l0Ai9+aIC++eQvc76BX5bxu
y28VzfrqtB1WZ6elMfTOW1B+9+wnxx8a9y/ikkZYVDFkEzD73i+8J83uW15aUoGIC4NCKkGMbNbZ
yJEqJ4jqC9fI9nVuAYRSHVVbmUpl96vlRb3fBBHO611PeBG6FAmGRjXdPMqfd2x1NGvPdDYLmmfH
BBV+WZ/obKAIsEtNa94bgHybr95v/CD1NP1+Y8WlL1SLLonDBw+Gwc2vJHDf2f2OtT3t0xEpbLKC
8R9eGfB9wcyHbvejsMeGuf7Zp+SR80fq+9oYamkFKg1aSummx8FnF4gONRbARfP6tXiFHcFGCULE
SOTw7LLY+PucmZ6sCx1f3EG4WEHjeI18RB1BvMSO/zT8vVNkS7AGudn1G1fc1EyL/uWNt6o1XUk8
EFl6X8p4/iZdrm5jXRxmXFHk2MPBgmptlt+TnPlP19mUp/x/Kqg2SsqYJm7yoRy/1L5wkdbt5dRg
RjPeeT17RVOhTYzpfhcVH1Z4TElfVaxhSG6hZ82Gnp7/e6lr3MqaSdxLg6Q1DvfucElyCPJRiX6t
wHRAQ2BOM+d8H4yAbSl/RakA/pet6WXLlQtUBgrisTkrNYR9cVTLHx79PSNy3jiz0gpvefRdU8hJ
o8d6vf5NaRDf/rxp35mrvII3gBYUwysSE64qQXSSHhZukrpvQQJRI7ulNPZP/GuGkGf/XNtTj47O
krRfoR+EZUKyhnu/Uh1MJ4DaWaP4KOadREexNz7ZNfJzrJ6tdbozRcPhazXyEacihkam49cO6QyH
voaAMYfuJU7D8I0w9Zen9adOCrJkhgT5dEipBRtmftvXzZxG+RJaSXEGZbmn5ZKDdBekyr77YOCm
1QJzXI7g6EthZf5aidpUVJ7oXAAA8p82z6CjhOkHBCtgPcn19shSWYKCVSzL13dJzFBeiP6n5+oR
/eLul/Tvdw00o+TOgB+VzE4VjlUiU98FSgR2tsIRZpXKWIEPIzeuenNsZWzBJb0mIPEUNv/pW2fr
XghfcKS13IAUWcrA9zMiZ5nnYSNRjvxOa0+NHvMbOlBeRE44T4SelnX7LGh9AkfZkcMSzba8+63q
EUcfFkcmxbqFUlGx1kSJbFW0n67Mluy1w5AIsNJLNzeqP77KvuEBpJ6JUeHqLuAX7A6SfiovSxh1
7zWWPlJu89aT0O1w0lmcse4GhgNHtc45erQyKYgFXGUMnKSvLwkCjWQv+vB5sWp2dAAgDf5lOgCR
yrIin0ONntsDpaMNXQ4SyGOjdN7bwFAhn0dZxJ2dbLUuH/3BRVUNRJ9cnR042C4c/hJmiLGqo5rQ
pCaMy1kZRJxFgr8P10NhEGWmzgNAVwpK2xzG5Ielzx8rlBp6S15YtZ3BqIotSoe8/QYwynUA3uz4
BjEUBqu6FVcR4aT2eyRJ2pGuDA131yN2gJVoBprxe8G6oX6eMmsYj//sPVr5YqZg2CbZFnwLUSiS
qUsJ/jX6fhhMJb+1W1G/CHC24bXhEFQaxXXOdnns8vtMns77tWf7Ql/SFJpjIaH0bivx9ne/WJ98
F4S/jB37uNAVUlJEDCQXtRW1xzZzmPhJgKmpyBV2hnZxk8kpMwoUwE4jEJcnmV0g+222thzxB47F
HNmDmppXqxYn6moG662aKL61T1wVKFVtsQVz8WW5QZKFqXQxsuRLPUAPLZpN2z7edHNVUNH2KTZB
fmhWcxjQxQuPi5QirGRRELUrmK1IddoChLiN3YP1VJxTU9ewwOhn28t1zMAuGZxRwpG43J8P4ttH
c1PqSMO9XpvT+/VGyFc/W2OB+h3iMlywUPJ3ExfJ5HRH9/QH4+S/LOBaoUHRtAwEsWWT85xL5BBx
bRjXvvEXLieDuMUJZj5a2XVhtUw46DYe6mQ02PFH5tFVncJJfFZHzqNykLxff1oXc8uxgz3A4PcG
083CPuoxOdSODfCdHuyd9/SuLqyyx2tUoI40aTwuSi5M6P6Qb4YIQhc22qC7J5Zh5ZyOYnPyiLQb
soVZ608tJCCnAJtEfcyMOd7FQa4C8g8p0biKvJit0dXZ+QoIaJhWk95JuLYInq8dSFNK2xMgl5Qx
Xo7xLQEKmI3H0Gs992oQAtlYmXkDQT1BBZ/c7O04ND9b4mt8AxZEfJlEGATJgFI1udAnICXwoQ2y
iKAF4+8Hl1wjIowMbFcpbLg7o3NWI7MgX9mB0ZkHP9A5AUmgh2JEf3IqnJlm5ZXWGF0MBapQFUH9
to8W7uk1gwEeKx2MliSnFVgnMkwnrfqQKZWXSGnA2SzZUKgp5ib7G2ZCEFTNo+G3FRuuztWyjaM2
SIa5sfGFXOc1js8VWKDWmNx6DCU1TfXJgrB2ljYSNvhhEMZxc0RYN39Gkbh8Ouh+H8uL5JainU1v
CHrcXO8haSP37qLqBJVnPMJTlxshiU0F81eYStaHNzZ15P/uWdWxTm1w9OK/ex4HYBFmHSL7FlY5
C135fGPrl344Z+pc5/FEo2zGS5qJDdMj6g5Umir6otW8Ki+vgWkR+sIeNuqgqoTH6fzYYm24++kR
Ev7y9omOr8bO5f1OtEsn9EpO3aWF/h9h76Vlw0BwSLzLmmgQoqb4AMBj6thyP3DfZSzy3WnBY/RE
qg6P6AJp8Xqi1cjEC+W3A5xFp+DvExN+LbGf4URd0/XMdEakyneFHTxvMBu4v/UmYhSrvPFHf2Xw
BQ32WL+X0QTWeIUv9ob12HP9S6KXU+9TkG2+Xrq9GfJ4qJtj3IhpXYQzwQ+ESWVgyDFfSwPUV0TF
XcUaaoT+teDg1InwpPNE3w6SkA9wTn1k1BvYYdSCY/HgbRXN9hHAKLEShnDNNAGZZ1/gNgWLYn2z
LNPhzmeIBeBKVkLQGe/IJ48ZFyOD43nOKZShkKI07BSeI/qqYdWasCRFtuxI8WXxMWF8Ik/w9us0
PKtLOFNEwQ8B+p9Y35upMEXNjqbIbbifzOH5TQU0M5HsLCLC8okCvsh/xhkbtVltH6oMefzqcM8f
awmiz/qkxTbOIYxUt86HyLX5SaW6421+2fbr9N1SV6MysNmGqjiAnG7aCh85mgYVjtO6ptVWmQwu
iFOd/m4EDVaa3oaBXs0ZPjdDpNkif5sOphgIyXniorkJgiGpvNXxos/ZIYao2RLtXC8hUgeTNgiE
FlL/0OjZdYfuCTiWuov2W2SngY11Gexx4orccnCBTuJBtVkPRvuQypITYNIkkPXJQaAbt9Fu0Way
UbgKRtx0WpaZyYHR1FnSY0zCrJRgWKilt2BF8OT/SZNuHI7VWSziJtim1uQgFfXyP1lvA63Pcgyz
qD2Tz39+j2xx+CV0MFkUFUVsflL1VTJ5pdvja8kQPBOYsdUK9u7642ls/MVOdQ/89N3rgXKyHR9d
xhEVaQ5UMu7TKrxodD35rQc1I1rTxYsYxX1nsHzMUGs7kzmX6200B6XIHMLyQ7QXEeMK1opqetNE
jgK8/tMHe+rbzyPVzYQLUEVHTGr4ow4qWmmOmoVUp8wgUdXi4ZLziABw/mPyclswj2kDncC28fu6
L674OBAnDq2vRDY1zWRUIew20W/qbUlCmA1EiJxUWa5Kx2pq0SgTlEASPTVU3CxcU7Am2ilFDiyD
gkOU0kWqU2eIaoFXmtjFZLir+fBsWRtIiLMu9ZeoOY3pZiPJobthGN/AlpzAIo6KDqklQr5iHjxQ
ijU7yxs6EqbdxOkWcInSDKDlXICYejCUughmC1UJkiX/juAPHmjtmT/nwfOjjqMyNNJtwFPVtFRf
l8SO24OIYCeIGHOLtwXMa4M+JJMeCDpHU9b4QqkN1CjbG+i5P9Y8alrPf/OYMYuecMyOXGp+tb1e
g5X3DNeEJC89ETtByfLC+WamiBPQRX+YzHVrckLt4asiNcVvUQPZK3cdqXEUOsBXz6VCi2Z/LSQE
aJRATs55Azz2nDMfXkepJ2s6PJpJQcEVZkE/FZmQvYZv1hX+LsjYMUiVByXF7N1yhkulRn28gXG2
hjBsalBt2DLWnWsgpEGZHB9r/nRFrERJDYPr04wuah2eeiI7EPYOB064E89PSzf4i+Xkz7xu7Uuv
VSVb3gP52CcSfhktYh3XS5UyKEZ3Y/sKEsQi63VuRXiUFmZax6JTwRb50RZifGYFgSPMyvTeAj68
/Yi3C3J3YEdJQyTp3HH3PzuIQnuuAOGwjLHY/ePZyoHB8F4i07Imk2LKej1QsO6KbQmdiQKVM3eZ
6VTG8n3LSpWomegn1XdlzB0b/AhfneyPGIJwt88Y5kmPoDaiSTElJhR9NLFDTC9Di/Y2c9t6lhXf
H3jrNx3FvqazukFDqBR+y3hq/svDpBwb2GbGJ2X1wVrxiGaV0lzLw1wl9SS0/+AQi45qhcJxaZDt
tCVv02v/XRvthBXd86TmnNYnCJAeut9wOco0cwtWT7KI1KARgVcx6meFs0CczmKiN3j+TdC1Gmdu
p6g2OPB4HUd7g+BYsJuXxFx3DSdXQ/WLryDNx/VaTTWWYR3vvIAi/0Y7DHXiTqrpsLbDV7BHGBwG
CZK/FuBT76E9rQVbwnQFP6SIswROa1Ng+6JmTYNqb5j5sX1MkmUwkNP/E0MgpPL2ipZZvJ0CCeJU
zUtR8cXpt2sZIitFPihx2u90XbS5mTtGfsVttHU592ffeMesT0fSNGrL8IFkxdmVdW9tEg0SiO1c
J1qBJa0XT6k/TeZ+cXmVNv2FO8w79FetnEANtt08R8gZst5F65cQtJvrCQG9iH1ZNRqTfR5dStrP
yUdcloa9foj9Fg4n/sXHcWJR7IhKdHTeQthxa7/CYRGcQ8YihkWSUc+JlkMKqIjCj2dMoB68ayko
2hdC8btJ3sUR/FJgF+ZBWj/uFM+XhYxG3t44ZONr3FTHPHEilGTijt27IEVnaeyt8wbbdvNCH34n
2iCSdxeCJL8zaOGKX0F98qMeuUa02SeJJCVI4e9DHfJUP9Lw7hFI32CUxLhvOk0foB87XZwcx9qk
FwTpuC0Xw/zM7dol2EkF3Hkj86d8J+CMwaO2W3NDb56wXpWlsYDDeZLLLG+v2nVrdva6/aOyxyHk
ZQhePuhV3GpP/QyeUcZnri7MRSUDuHLD+N/1nf6Gyuors0u5ohWcm3J4qaR3fQ3cubZFvBQMpt+K
kky5Ww998sWMiIa2DgG0ANknJ3gV4wOg3CekRyiHGVPGvPEp1UQW73OGiatvCzhFWNRFr6qJ56yc
ZY0M6KXGrpnn6tfdb8QW/wix/JSDQtRfx6YAsmMo3+hS7Jy71SgLUKq5jYteVqgJO3I6oNCFawBf
F1iqn6YUwxixzB4iAt7W5wxdaT2dlD5wTh+S8YpjNXAM0iTeLzohGpVhi8KtMv/XCW/AaL12nH4D
1M8DbgSZpwtql7r2XcYc7+gW1wF/OTFZwaNgd5SgsMmwru+uRpDVlswOKOZcZ49Oqmk+ZuDd4hOa
LOmilXyGqwOEE9ylVqzMYkGvT0pI+nF2HVXJpUrgptFBcJsI7SSjZiw846e7ningpuJTI0ZSefv3
bzi3hhPy+rSbql5VuJVZTZOUGeZG0mjon3e9HWIMxKMfbqatNlCmU+GztxGVXoS7pFhzhwf7x7RX
wyA7M5TxYNXmXFszIr2HMDK7Cll5SwGivm+eDSI9zNMeDRwiGEYyL8IIymEl6wKeEuy8ehtZZMck
wA8OhfFZAL0wcCdl59266V6s1srldMJ/7XQhBWNES1hkdi5wA0se9hLBpDCLWTaXnt4jyR/z54uC
GR3hnVHU4/GmiiZl2pAG0Sv3veYTEklDH9+WHuTaAqk0wkeFK06BnKxaeNJ1FgkcI9ase3hG96PR
f42CX27jjI26XoUYrKxtnuL5YHL8IstzSHDGV4b1bwbdH70rxX9SBJohfK2x60/gnjpZjYjuvtEs
/M+quTAqRRfG75eGyT18lvPnnXmMR4y1F3z0zUuhiZV6ZPipkDrc0yS81SggQUGL28v6x8vh6TTe
gcpKvhbXLXRZ9kNXu1gLruJblAxzTQIpZ3ykmV43sDWkZFR+xPxY90RN/SIMpdUSs+L89M/DucOj
3T3Cchp4YRB04u53moHpA4Wwe/G6PE+RQOyo0sVZf5z8DdXZ4LIPflucypNt4Ktp++3COEAlHH5B
CSgJMvca+XYoUgYykZatTRu7k+gMJkZq0L3zzJilXyRLe5Kt1hoVRl/CZfegDi8ZfhTF/Wp3rotT
aY/MjwyzhayBb89MSyttxpt4Hauush1ZeAawsUarRPyDT+Row5Ft4Ieyc+BOSJnEU9QHJ2bxi+Pm
lzNt2TTbIxYYSGJagLn6YRmM3RC/QkbvtkUJCRTMxmhQ9eMCq5gUgWgzUZxp+9L9ay+1M3EJ85Vp
FAk9aCGluwxcyMsCWkq+h0Y1WX7LQPOxPWF9oaNzWh13wqj1pxeupEViwVBSMUQp/GTgVthPOr6k
gH0+zIbllLT0yPWOmuvN59FQt8i4AWriDaUtXAYB+MmMXPLj2dEG9lg1R0+CtwywirOU5vqynzCl
d7NlPuBFZRmga7M6SO2sf4SbIorF4Ry103R+e4XfBRx7Ygc6S4xmLePvbZ96KGZ3OPYYTF6nrsoz
O7vX9esmIaSZcY9n9ysFPO16Vxyah03vAHuhnivQBeZfSbUesQUcMs4vLDMT84r4Sa9jpXxDldhX
jfv7rz2SPZuUleZco3RI2MIKrWOuv+vr9j/cthn8pTpHHOI0/aPc3P9zF4ppuytiFTy6t7Igoui0
98O85ngE6UjWCwKxi788MEn1ql3BqHx23qDodgeGQcMHzXB7xBiFTrnUj3ylm+r5kGv2XJnciC41
NuxvbemGU0aA2yMGlyM6OLQv6gyLKcqBUv8Pm/B6gVZ9ve85CshoEFNQ/cr75O8cwHA9qGaqSKQz
acUjcjJ1pKBymGKF5uBXfUBFTN3cOmx2kyxfLNgPgOCscQ9wqj+qMupkGe7fDyqdrcfFYSWkmQRf
qYkGErHLssJkyVE8vctj+BqnKBa3X7iyvgBAWipaKx3L0B+xIxoKbp54CjBcpy9YovVxgQsc1XKK
51NEe3MAHNCHcnJSDwDYbJYMeuCNxDYz3ihdkuIrlgNkPcR/GdRJsVfiiLLnHhT8ARkXEwDzUIpE
/pInTfqYwwu34C0jmkEnCAGEUNdgjyMOkMLSHROjahsqZggdM70KcJRqM1bsenCvGDpCZmKl32lf
hujPf4VLF2J+WxmYYHnBELUWaYahsVyMrD06QrjmdlgYgIzKn0aSwKja/poADF9+KAVdTtAu+vbJ
M+1+gTmReYfULhUzEaU2oCnxaJ6JDchC+9/+ji+g7WMEvBQ9lBZTHfdbnMNA6QLNqv9dSqEID9zr
BM/itzLO+ckiXWZniSwhDLxQ/wr9tUn1ovSOVlxRvUvK3XmqXbl/daSH3VoHPyBHA5b/D+Eo1spl
mV9sPFmOE/a09vRx14k9f2qyckE03iYyLkP22WoopzMo4d3/e5jPej3H6f4pjnGQbLwR0sJEfzlV
byUjOQZQFphNKCH2Ni/ZmzK+BxUFAs0NnN1W1n6GtxUY6vbVAZt+XbLyKLAtdqhVavzN18BiVfKm
47Gg4KDhDBVAlaKfCN7aXJTmH1FQ6zRpktD3jRhxndi8S/iBbLNovYyc0pGt6PpfLBEdq/xZX/Kj
ttU8Yi/QbkfQBvnEC+e8kiIELUK6EFMjo7BDGtyx35/TIsO2xKwY/M972SB28hYxhT9kpXT3k1Sp
CXQLSkABSPgs+61RrUc1z6zi49bB+E2X33p5H1vONkY8codERa1NXcmH04N9XlS9xsrkrPc2pScc
goSFGYjGt7eLvG+JgA1oJYVoUtRN30tFKTgyc4W7g1hMtrW9t2Tw//zSOlW23FM1sPBgkZhQBXAg
lWvsUEnNSCPoaH1AQyMm30zKwNPAacjmOXy40vYo1D+8DNYb0E1ZIJ8Y7lfG3+pttO6QycePKDse
I90aLkYBLUp9k6KwFT6jEPxxoxUHF5NpHmfr22w38/NGyNXEM45yyFJKpvnyqySU60WH31i287t3
rBOgWi+nUhG8kOTGP6qu7LJwt9sfNIietMazXcXd6BL7m3nHYOaqgwPQj5X7h+DooJShqUJJmODG
p/UhLGXURPnac6xFq1Cn+si7JS0Oc/xE254Gq7FjCYgicn4vV3se19dG9jwCtRHWR5MOpG9oOT6Q
S+6vm/eKOaqr/tmY7c6apWixWFAAAtinYLXglLr6+vEsvlssQQYOncAJjRBbBVxpLIKI0T1AdUun
NiE55P5UFLOCgkUIrQi2TVQZU/Ddwm4buo4nw9QNr0Md/Z1Z0705lkf/h3nvYYce1AWAlQKMwXkg
3sACBzrT+JhEUsyv07RxP3nbvlddANh/zsh+LxXgMCEGKIDMrSTRKr0erqlKwQOkFhCvFG6H04WW
BQZ1tAoY/5MZVoCK7Y5AmscxDuxk+BUV8ebfIjoAZt0uctWAajpCm2I8Qn/KNa+DoBUO1dE8oYP7
+fV8xGbsn6Kt89qK1RKto88sM2d8zSXRtvLv37MF5ZVctRXnSfmf/VMHxHaYyLjq4LPWw3yFlVaT
tQLn54nqpSfWplhBM99bdpzsBQK/uYHHehVhPOtBFUDgcHpD0uIZCWvhAilNH+sLlxIoO3CkhBUX
kiMcOtb4Kgxt82ny+ojW6MqgMMxTJaiNlZLf2z+jlWwEFIajk8smtagpwe8GMqk1J3AhAMeD+edj
2XR8GxrlxRFDgvYOdmRsYrnyXrQUk+TCm3SGWDUpNHKYN1xbWhCzQxxp6kMn2qG5YINViX9JzYv/
3DxKhV92efgsPE6kROME5i85IwnIoFuiLIYxLSjgiRO3a9t6l67zkHjHg0RUigRNktUhMM1zOsqh
68xg8jU9f7uQc02dyqFtaVc6lmcdBqqKhy2WorEitPk5YFwmauBPjN6ucYQE+6pEraPoXfzs1wyP
Ox3agkaPhMW/NWcaCJ+jjjkmjZNTfTASFWHKRcRA4/QdEA7+X2SkcH1YVKQxBbqp1PDCBc/Mn5q/
TbICxMmUubuzCLBhWLmDbBLnl4qarc10qPdQ1PROU9gVltVZcCSZGGSqTDZdDZ0zPkLv79Dix4Vc
DVUbIvi9zr+Rb7zvtczesM+Y3keGssZ5mE/gxiwgz6R+1LOf5+JO6v47zsilxlStHssgbSURruEm
Ym1b7l5lRFjpmy4yk8uHXck0s5Defs+DCl+gWzeew8GPFftq4z6l24CoGYCDOL5Z1tUp73BZI8t6
dO5F9s+VUMqvGRZ3y6UmVofXxpFiGcLOjwsQsy8L8GT5foyD3JmXZGddGIMTxUKPZ3QXAeoUXS3I
sc94rviB5NUB9gWG6mPivddea2FWaBEptcBVvp8uXf0thhGrAh4uax8AFAroBJV0TCg+CmirbZVO
d9XEok5f9LzxEv7+H7jkI8rEJXIh/h6xgsCiWMXo2AWfD0/VvFW8JlQdRhdoHf/tUnhcEvWGJmlQ
ydHAdHL04FmB8QEeEV8F7Xq73uLymvREEpG7L8iXvIh6MdgIq2WdxxcHz3lC0B+oVwFKUTwOxW82
8y8GnDHIdXi/rE9WePuc7WK5tVfRM79laWaxvdXEsTXT54ppjaUmh0+QBun/6E0nyGdnHwiwdJRI
aOE0Y4UkFwtEWyIIQa9AoXEJ+zJxrtdzqt/gzk3hj7Z2PJOgW6G+0ub2Oi2rDiLKjIyTPp3hiMQb
QTXTNdbpw+/aZa+1OY5HSvyawBakpLhNpG/j9qnZ6LOHXw6THatEuDouIPoqsggEqHoEPTDz0Xz6
cguZedZKSVahDKgQRrHDT/iNfBIQflbv2oggqLJSuNMmhbq2dfwB/m9GFBY+zNAbB2Uj5E7WLlJW
cDDDthmghmDDe4qqt3cIPPvYi8bmXOgBHRb5TX3TGRd6YYlIzWIFSvLF/JjhyG8V0H/2r2z9FM8x
EAR52YCLaj6EnKlrVmmcOo6ARY/8c6r8NXCMPJTsGBBgUGSTjKT1V7sLgbW8Or21Iqnml07nTYqW
gBIkMUcjxrszMSBBLvEynnJuDNu/LcUqalZQRL62Ua1XKuJsxS19yc3s5gDKm1K2Yx04kC988D+z
JGL0bbhf6S4S2TGK98MMJ2nDDqln4F24B611tlU0thsZ3C58LTNNzbUUs1TRRJWTAZ/cHfXxHpEc
axqBT6OclXYzP2nm9vzL7VfDCrYTowfbatPYSzBNgUVOdZQwCFq6Xo/JR44seVAVAmtgNxTkEY2X
aDp23qokE/1f+yqINDRbb+QOtNWK8mwpoWASa4cD64uwRKWt9Z6pbpI/cwACaQRCvAv10iZifnrN
FCaSD/PDCHL9CqQHbEPAvY/fV/OABNy3l0+jXF7u13oxGDEtr7xsrwhPq8rbTV/OluuFiiBnuMBn
tbAuuWJ5hEoj5k1F2Lnu5iBXo50Dd9XlEhFm0Ib5DlGozKEhu6FKzDVIcLWBGOAZ3UUtKHlFgog/
D0ZS9M4cnJc/dbHRQogIe1goKibN7wSEoJQbR8Yhdk8ZcRUcqR5J0qjWbG+FQFQW6HAAfpJfqWnn
GH9fPNG3f3gVk+Wp1EAymtAzmpx89XC3oFQpP7GDYRjgaDJbojYMQTpQSUnl6L+aLOXkDDh5Zcrq
Ay9dt1M4bX1QM9jN0PCOTgJGXeaGKStAN3NjcVh+BbwFa3mdbC1FSzsIJQAMXk4zo07x7SBgK7A0
BjcxFQTR7Qb47YYdJZUhDXEKZXlMEMp/ngqcKPXheSYF9+9HBaoADcqBVOWzEYNLIPia6zB2+hve
JBpkVmN5yjUxy6c9jvy5mLafcp+liDYYikL1tdUlI0sEnI05pto71aEmon3tvDOEucQ/vanpK0ow
RwAzRwlTPEn8Rbw6vIogKOb3ZLwbraL8DnqKhNtPgOFLhOCxifcYvN2l24i75wkZL4scg0mgJFAR
yKrMMiPq2m8q+MeAuP2VRSREjaMRnYDsxiTZ3rrrPRiBmBvIMsd3oOzjys6dRI/3WrXzHhZ/fLIX
iCKh0WIa2T06UbtyEQtPbK4pi0a1QfR86ZB8tZqFYpnkZ6O+pXpBgVA/4RZb8FNik4fnoHgjU5rE
4SMKSkztXaIcIQcB22NGb1SHd3uL48TceMz/s9NsonXOitx2esNgCtdhINMPr7uSQNgW5grphpAw
rrr2cfqm6uKf7/JfMMc35PTb1gsDW/IWCYASd5d6iP31KLDBSjFq/32IY2YARuMkCev/OKwjOABP
xv7YTT9LVZBrPV011P5C8yvf0DQOXyIXjqau8RAlhOTOlhsECtIIHStWGez1KLs7kVnutG/3Kug/
gLj0ZHOknP7aAKrMSiZxGiG1GPl997wZj72c8S0yWFuxwXAFBnrYyHls8mTGqkO+WFHnheF9GHo5
rYNGPxGiLx6ofgcLr1jc3H3SOprJvNeloBCqZ5vne2Xi72BKD+jPgd9+YEkGcTbWtoegMPxfefPR
fMG8YR1epAGCmLSG2JFhbM/GrOJ58NDQ3tibLhNxV1aH9TwaIfC4uHE+KgpOaw/BXxwH7fiwFIIg
MF1vuEPonQh6wRVfUPsFdaJejcVNuy9J/BShSDvxFfJdvVeuY6ipKNJXyozyVEfsGSfVlTfQqskg
Pixhm1+7x4VXjFMy8YRnPOOM86j2/e0jn/ZNJIUUHgwmhc5eqawdfvst24iToRn6Q33u2IZ4Xc0X
16MNv2e4nUQOtOSFhQ/2VYKVrhhmWHEJuBN1lTl+9zNVFIh5oXsPiOJUF98RyOMNeZ2bd5sdJVY1
+s1r5LqomhQ1bIC6UdCChCdoNC87FvEpWi1LkG9U5QuPyNW6nlKMQp59tHFvY1zHUZPgea0qyQ2c
Idys3kI5uoAwa4IFuto4/Pg1rbtlWgwXYlDyT/CIBCnMvjaAjRSWb8JuBFQegkqPP6PqqreYpI3t
4cBUpsshMY9wBstOQ9ih/gUQk5qJqLfknSZnaD27TD3FgD7ewFzQ8a4pfy4WfZxED1MIMF8aKM8Z
9Em8hEBnl0JBlXO08WrpAab0dRjE3FxIXzUqL2B7FnTurbAz1eA+jrXxghHrLlIVwrky7eCkT/y+
Z3fYiFeD3y7zIkbRxSuZrBBg9k83XPHqrS5ElcF0DXBFw+xibg62s/ZpLKYAdBkDOg/0bn7IyV8f
5ZpH1yFI18I2FB18okHXiq+wygD2G47oIypx1EqGkv0KosyBPr/aWkvmoRL2qkmOTBuNDOJ4V5z1
Y9cbU+Dtbfa0erZzqNJHj+DjS/e1A1ZvtaoiTx7tgQDBr2+ZP8XHwYhZqx4XixsLOxVIoYYmwOG6
8eM/o7+zmaS+7WFZCgfJgT2yY+OLC893A2HbN1a1ZG15bfPmImfCLtKBNKpeTEkr+GiI7avVLtRn
8POYIfh784dTRH26VBJx7mNnDxAmNOmUUMsGtJ3MP0Qst09nBD5dDh1pVS35o5kYlQpBQLOkKI0a
FfARtY9gUMhY3k0FP36tA1Baod73Ln+fziHSkW9JMHki3EM/hTznCDTrZtQoyeuwU/h+T9SJ+mit
+HpXFOsR3V3Eh2rNEwnQZylRCU7iHnodNBCBJvwxf4u9y4CyJ0uT5/jvyF2/gWYd/L5dIIK9W+Kf
MdkTkLjPyr9doXVIdEXwrZvRgls2G9pM34Am3vWh0ODm149upDCaPW2N3iZ6UYMHR1oib63wMIZ4
2LiNDUBEyIDho/SYAIuoVFr3nDuvzHifiu0yn1mBAk3hfS2hvGcalXdTeZfY05IsQZsPmJSVa8Wm
hlsdKNvwFOsyZGcjKl7w188nIeBZJI99zbgW417U7lkVkykVmRA5fosVEhqKyduqTPuGnWIO/o5A
l1Jo8tYOvD3eK7zFUAnlMCe7PUJAipDrByVAHmKV24JFc/0fl8y9aRpTqJEA+uyluTMNGHSQTpjh
C/NBK2uN4HQJoCkutaEFYoklucOuYv1mQusmSDb4/9uMeEZ0ZSIiJfQL6zJcesZtQ4VS6ZWpJkXY
fyhf8qL0sor1RgjgxfBFlUE6piGbnGfZjtZyhHIyQxng6uc/M5L/Xgo8hQQ/hUh0esZ1vnB1ut9Z
1aF3xqL+hfxuvGdhyN73fGTH02EvfyF8WaC5UIukw2rnnkbhrOnKASiGJoTtpaQkdANH0Xv2ghUn
R8YNGzpOZ71BL0qsG+XYNPz9Clz/DL3l/PYKPGZKcqISU+07D4vBniqwRQ0IFvIkHisQCZWIUsup
aVu65Bv1X9J5SH7PG7zmpWuAOd2W2Ce+HSXjfxdsJ1H33U5MRAjyhPUYlrx8MSvhFZp0Om42S1L3
ANPSxBoBg8c6euYCYqRu7fHe0QrH+Cl+H4t06yF5Ryd/SYIPKcbxt4E9b1OOaByfHurD28vz2jES
1ZQF6Z9VeBwph4PwpVZlMlIFzU6vSC+F4I+CD74E/Y4NMNvKbGQov5MQmBWIKlE2dsPMRnT0T5fc
dE12HcwD2tHsJ82Rt0MvQemFzae5lgIRKkqxBstD0PQLuMiL4CSGtkFR2+nV8kLaf6GPjJ1C+fLE
MUa8WNhhzwnG8nCIYTCR3NpV90HsMk8/q/iHl+l/kKoORhmilDtc1m/VlwOlW/DY5zlH7m/B1uNR
TZSlAjyU1kXNTEi9Fh77OOPsuhN9vkULhBtBBFWi+5fdYn+bACzgv6tfS25yOyKqM2KsWBNo7qv7
8RP1a7ZGcNDx9yqZKpLgiWVcOPUFSuOkSz2q6Cn0HfTsA91NnLgv8QCGjaOKOsp6jMQyyr3XU72V
KzsqrSI1BXJrzBw8sS6/OYqjO3VW/ME6/3p0g20iBzdM7Oa4ciq55zY9YCs7s9wDRMpIqsTepAw+
d7lYxcjkT3Yg9D6sIPdyPAoiymqI8EEoJBNT2SI9h9NejxmKaeF3tHN22/HfNVrFeGvxmkqpD7BF
w1TyI7nYjHId8PKyVO6ri6cG8h3eixtIY7OkHrensgttV6jg0Pru4ozuYy5cak/jGtMf+zP631k/
Z7edruZlbnd9Qt9Lv54gBaxy12uRCcAJUr7AtS2QeMpd77oXT5ouUuswcf7ppXDy0lf6NTb4hqON
4e6f9Zo5uUnASAIXPzeISmrAovY6vTNFSDWicK0ki9EC7yqlGYdfQbHIijWphh40a3uorB7hl6kH
nn1FbOz4VerXNJdPzm4G+akV1K+J1q66ACoVxYRdDcT45s/zu345drNOlxJOVaz4dSQYs4KGVXvd
rJ3S2Vyio7w4oHBega7XcmYFxeWPyAKM8A7iyliWQ3B3cg+dtHEssk28tLpHzU+EGuK57syrx/2I
jY3baxWYw7VtEopI7ZBJAq/5OoZse22UAXKyNPSusBCkBnn0vpI/NKFTB0/Z3zovxvh8OANFY9Qi
iY1IHTt8NhmECCmiyJcHQ7FH1BGQ4slFJ0MKyUxlU+bT9Tc6QoSwD5bjddCzw0W2qml5GCEDo2QZ
/uT3zxEUCsmfhOXoHPJcChBQDsP1GLnXqTdXCdcl2ZBrkIdl8NPdZeYLFnmQTK1Ayx6W6zoXh1w+
5Rj2eptHSGCJERof4m8A7W7Si6C1+FLzZ0TZdrNOnDj3L1KTbbgUg/A4uGKKG9U8bn4YRX2ebWJV
Iy09OCOE3ze8QNEOsPrmb6Ut9iXvm5JVDG2uvZnR7wU+v2eRCLahk4iMyCSczlCIpKC+dy5Z41i+
37qSdeNsRbPrgBxjlpOFqmgATas+e8gUOzluiAHG9jK5KdxqzYkkwJK4gtPE/GwgR1tdwxAmM++8
ouRQMGSVFvToGFjXxj7VoX+MydE9LONLFyKlFfn2QArZsEVKx3zap5YURZUmW4210NIcObhcq3zY
CZxUs+nrIFGCBgZe9IVYCEhhAZFjPQiVjYJka5MQmMtvCTeFVZHqac4n91Wl3zH4Fvu/fQAbzBag
ZC0PGoVrAJ0on3+QcBz7gyEdAnYAtN15jj22/iyEGXuuKxX9zq01I8wwugkrNlKZQQurMK8RHmKC
BH7R/Xi8yKExNvRC2vpb4kgweeas52jmAzxM/8LRItG1o5vgkaC9uT2uVds7Dd0WgpwbMj26nO6q
/uo4j1voasU0b7zO8B5kUDEiJ6OUZsy4uFMXVkIWFFEl5WzIeuEGoKmVhQBAs5EDdhP7Hzx+wgzY
SgY001whEvtCC5Dhy3uew9QNmvTwDvaOS9biipI5ElEpJi4BaxTbuy6+3vsOiQHGkJwqF1gGDYfw
FqPAAUK2DsZhO26+I1IoLMFVsriTD3rG080uvqTg48SWWSChPS87SJiOqYN/x1/zU5hPyvJuiJXG
Mate3RIGjhQ8H5IFoBv/rGvR43zF+gUHALT4VNavtPvQH6bjbXn8bfo2e7nOe126u8UL4Jxba2Gf
UGFJfh0DU9sc9U+ADp3RlgBt298XJO+Srg0m7AG1/NVAMfQNT4tvLwQAZ/BWjvlm2XHMS/cGNzb6
Z67hUqTWKDvyy4ZVXgkvJYL7LtSvpfAA7Lj7tcYhvjkBxCIcxeomiPgFWOSjjEAiA9AsJihScOTW
blwqFkAvuRjxeP3L07ETakUJNjH1MrM+oiIKMiv8AKndzbBO/Gw3jQMWC+y5YJPIPFIhK6sLdLfg
SUzien01C5d0acjKLB/lgFxvLk92YtyhLXYLh/zy4D76RIKifGx1HvBu1YDYFlw7qk+t96leOHmK
GxMIk/o6KG/cUK9/gzEWh2h/SgmmDKIru5Be3brwNkZuXfnWfgaVGMxoMgbSmJ8OcTQ5gP0fQ1Lk
TJmHNOohtUZggWh7cz97j3nKlfQFYRMhmjF8kfvKUN+boS35hC4ZGXUs+Pjhl2rrqo0hDb69li2m
ZrG2Ts3dwJsxdzFzy5zrHUpvLdeQZLMJF+eLra72QT4T4rcVew468oi3jUaYVMiBDxkVkAVAgCxY
v5/BuiW7zsNtBr8vBQ6BwQIu2JlrOTLwBpmOyMkCp39nLOC/KwK97s1qsdX1bUivZGeeTHq+Xt/4
qFNAYATCvOLneUL6o9bCQarcpw14XPl8koMA2WOk3TlBlC+D0RTxAIx7m4Rukex3V7KbpiwGGiPk
ym/+Q/KoJnYA0bCJRpDKl72Wv5veH6AM2DktqN6glgabujWZlc4rHIFfzzwR5ERQ23zrVDlerD2O
8mTxhw631qsiFjFAdyDCpsaoqvD66bWBiaffo4vuPkIlkqh/VzOxvAL/o7X3tzEdi+wXGOTvLLnm
10MesYNlevyNx0uPEyPGM0a0jnTf52qRTTuK+10Ofc8HD/K+i3bNBHEky0US96wPtET2JGpASjc3
bsdn80twq49bflcp2ZGhWNHGkrPw/JuKn0QDwegkDubDlaXAMmqEcvbzduZ/Mvxoh1eQ3783DebA
jynwwweh7KdhEleIKL0SznZ6G0V4Tbfus5HMRU1vqm9eMjBA1jGhK0aAzIldShZom/YfYeDDgChG
s2aEtpkg10MEbUmLoU75w0WtS/db/sYzaY/rJJFhVBRTDRp+DCdNtxoTQLhhnu43Ommfvqy+2ZL9
sVj2+T9aX5kJsuxgQUYZ77NBMyP052z7NYd9m10xyCkL3/z/IsJ+K3zlnRJbhyLYZ6VGgJRvhnr2
9LPDk/wDtC5SxD4SJ0fp04KXjF5D8/iwUVd+QXeKKTV2I7nb7kCaSXZgPIVHjgaeCRI0sfgPcvs4
1U66fnw+hoeJLajV28bmRWocA1WX9SRU+9rwJJ9R9a5tyvM7vv0rk11MQv/BGVcVZFGLPObGDtkD
xLkJx8R/mnWU/N5qQ/pjhQDX99f12AJ8mvsy7DvQ6VPPHt43OywhqceQ79h6DENKrB4DdDJSSfe7
Ygl5CEJo83208eanFihlmFpUhBbKb46ysqIAIdLEbzv00gX4Wltew/SN34rwkEiQ8d+kkqR+o5o0
1hcdCmZajOihfZKSRUbP+QsAwzLYJrsXdx3GXOsVItOWWk3Q9IHb9//HcvmZXIoBapMybNcPzKKn
cyTGJ1Ca8iJC1FVe9hBE2i//FlPhwf6iT1kiTnUD2Vmwt0xZANbYB0koUMz/cHR7UhL+Raai7sUB
AH3978YU6YbJtku4WzESB4vBDyfk2XGwnsu7MAqgIGiQve4WZMY+TXdzXbxBiZ7D3oezmHJagHc0
OjFO6bupMhQ+RQ/p51Eu5pv0S0PRjaiTrH31h+p3HP9rmNSx3rTVfJhkF1PZhVf6xpJJDp1DOXad
lQ6VzzcgQoPWBqe1vGZYT3CRYyYd/2s5dD0tAq+4WL5clYVg/Qhc4CodLKQ3CxQe79yYHWpJGzBz
iKANrJdb6snBNLXqXpxeU7GbNG/x5BM078DFESotA/C9iLsEoktAai2aSRBzs0NaK5n78GFYOM/E
vlhcKvqEmf8BC6QYyTBWBv08+EBoUpsjZlY1Vs9B95v/b7YTtpNkGCaf5K84oTXvEaQdj0uhpli6
yka2dbi5fqDMJv7T0hATY1GSmgFbDmjUG4/aKv+8k6Qt/RDfYJ1pIAWzigisfiX7cJr4vk3kpfWW
BR3FIL+Q4ylHtR/bZLIO4m5XeE3Hny6TONiK9xxwJElfLiCH0cRnutQimNVxg8NOSfJv5DeitmlX
LfSn5ah5QQ08HYomEca3HNh6Y6+iszicDhTXpnB3VhlTu8dbhuCYO+I0dykOZXdD77XChbkxpT0w
J3OXOzkU0THGy+b+6QjO7MggWl+Z4Ag44/vMuVW+gT25mdzhUPoFj9+txhwf/FWm/p++3BMPNJK2
pqOkkCLBoXmqb9Dk08Nt+7BZUAVWfaApLJibtg5Sb8HEOYcOBug4UTfKPQE9TyLKFcRZAtaoDZU5
+g/Yb+rrJdqhmlB9Ajnnh2xoKzQ2vGtXC677Gt0PcE4NWyqdCqPFIv8P92WI6TcKVNmZ+XBueEf1
D89soXYAxzMj4WATtcX+U4IsfJ+oL24d0e792HVgXpE+4fgrpzLsufUvw88xOWVf2q0oqdWN0/5Z
Dqh9gWbDYXvuiVsUF9KdUsyHR/wCdfYJtJCFSYlVV3SKFzdUH9rZ8S+PuM4XLDrxgvAZ+AK7GQyb
kDJol8ZJnlvo9T8KnXK1HmVpB3V6m1QHzJo9++QFnm+mOR2Pab2VXKFevsSTWheNcO1mWi7yYz3y
5BhAuppDohPsI+aKC8Wp6iNsx34yMVCKs9SFSnImqyMCav0oR7cwWGbSLy5hC4rjfOtHToDuQFy1
4c3ua+ykeahESs0JYUtlfHDUfDl0p+M6ytKl8yV+YyYhfFtwezzxl13KXXYmq50EOIAWOCBil8+i
jUkvAVc6zEx77xXO8XA3B4av/1P6t4w7saHHBTjAEgeHLtxeipWam6nKYdHAzeDVFCR+j3JarONl
upMlIJdswVLbRIowtqL6DYa5nTVo4xbHNmN7qykFpuoXlv28bQkar8oIh6FrTQgy/WgjyFTu+Oin
6wZRme1JVxrnX0+Bh/kKvJB6GmZ+M/MnVKMkpMKvG3/qs6J5sTKUjFUObHxfAPgONmti7UkV7snH
3NZZ/3YEBjQF5+KHSgCGu0QCAb77BnwcI6v9VZBVvNqOs/JBTqptfTpKurRql3J/ixe5uAgULHvN
9pLNvnF+vjWzjtcPBIZReyj43ZOw1KP5TJUt0VWbadc+W9hSg5ixhRbejxYFmwztPDn2MEU88cWU
RFnM4DiAJknSXiRtUagnsByF8b1HAxoSDzZLBBxXSW5BnNR6tfEoraBmzcWa7js4Ld2oc8CMgg2+
7J7cfkHY93nAX86tuS8Nw1DNftSI8DShUWTxUPSSNw36EwnLbYqLmY7HMRqFJIzu0GcDXVk9YJRj
YbGszZ4NRet/zg4bJwYOWdI6/bdw56NMQy65SjqtKpiUPf5dgMjaZAadYy8Vd+JqU+PK8WZbo+l1
L+ZMGi5n1eZsaglgqJviUyy1JNVwz37R+gBrgS0RBlX68EQAiKorDlFwzJdpTcvfiTF7+ZWWyftY
VdGeYvS22jfNdYRWxFX3Wv8zkozO7I+M+njvfSBA6bTuyCzzQVpqyNdIpFiiDeOXZItSShlhE/2i
u2OVYFHFXVZqjKqHSKFdiVe6fXuuqojrNXHS6EIfJ24bYNHsEZu321lb7om0YO4pZ4X6pD9f2g3o
TlZjQoAcjqy6V+MFpflwHxVPhDDN9UbQl/TjIrLwEVvnLnehY65+UuJQwoFIUaf7v/gy+u2xcVAb
ARqeBDQ5oLgGBAnGhLKj7pa08EUb2wswCI//ekC0xYnwspf2tjubMqVX/4BPW/nKN0939JgillJ4
+kd8tQqIfQ0KgNWJoh6YPOCsVWblbXhYzqSqA8PnwTh4uVfbrl5XHMwAS8NmaqePjZeCCzRweMQQ
7YFryak5e7xQ6aSyBPAGWotAbwES5iuNGbw1H3Lr8w8ikGx8kLNHvxU6PqodEWSbFb9Sl1mtfJD0
dJcOXFXjmJDLjTI5NPQBizGlIrP1e1c7U0Lqc/G7AsEzASgtk+C7KTCRXK8F/8T7IHRYDESv5Aip
E7hmRv20YrNaXiXHal39U4j3qfkEj/tuOOD/DpHjjdsFjOPuKxtoVF7FK1wb6/jHiJTOYTZkYlpV
CsxTUPLD4ENSYuegU89C+nw5QK7MABNdBIDBDG5u4sHtV8qBCgDKEDPC78l01jdY6HQ1ZO3L0qe+
enB09Ox7/tf9u6rFMKqKapKoz7al7rfVii8pUAvSd7TVBOf76PLalOiXAMwqae5N5lXARVW28Bw8
dPhx/4QqFSzj9YIMLlYXKHN8UHrpIVM+e+MYzdJGYXYSvFeCOJ2Ng7f7cuIb/+DCk57nGx/VJ+b4
hHfIut5nAdvGexYn4jW9J9OjKWkyQFZDXhcv0+EiGoLjifjxrP6BcHHjhW5xJuLZZHZxHZgXaZUO
At/cKuqBOgzs1GsmDmArMPb73I08Y+V9Oe/X0lJ4S7+gRV5jhrqssBaoOvxhTdOWsIRkCbRAns6F
fXQKa++AJac7c7uh98IZf6LDQ0CqfTEiUhNJxwi/dI+EsoWbvcoM1oysxKzUt3VxiXwTt7dLCIOI
0MSfcX9jIUrAxkCoPX9DTAHsnQN9uN9HrQH+xMqVpoZvRHXB2lXTvRLlKakhjQOkPun5c9jBcwVj
FIQq/vWhWKxT+OuVXxJA1kKLcdRG1G+tZ6NNFtU/wab076PYHOPq8nE+7K5YqTXZX/aP/vKloqVt
wHZZdYqOnIXWIPLE/BSzqEQOeMT8HfaG+p0b+aq1EL8jyEXyJMCE4Gr3vd9VKcI8jWLw11pSaW3E
JY9c/cZ6PB+8NG5dAc3aLKmIQ1oK6imwDyy4bMe5aX/5L5Ug1cVA/2tmecMiu+cJ1j+BQGcG/rAF
ENRL0A/7HHXXaI4ef7Ki3s3fRlWfWQUFIUOx5+VMHFC1yeg8DW5ZD43dCBiz09U+nUTfsvJtChew
NtxeK2XHSuXPzq+9/CzrJjBRqgPaEbwsiwU8OMRlTarHx6cLQn6FcVjEQXrZ/GQwX566NgPleVuU
y76grT25TgxrTZs/GD2mwIedgatuCLsV58gfnNTUtVgvqAteY4+rTJ+DjBo0vJhBhCqmahO7DB3L
luKQtGn/doqk64yrm3fg4fFIkSK2gZAVll9Nk00TEZjBm0G/BDSFRFu2Uo4Rpk3nUA3zy/gCYJzT
VE5p+KzBDhG5nkQ8B0Un2aDmw94h9LCgT9Nl8c5rCudglPgKZAzxj6Y7I5bpExOI3dCBifPlBgot
Ba7TJPgbr16FvlPSrgbYaNES0nUHYAIucBiXH7ASDV6ClsL1WQ+cEJO+kpmzf7zGsCS4aw4LXGys
oiF9t0Ant3hWFJjYfeVOk/PkbJOJoo2JfYwmDKWK2Jqkr4C+PUKL897a3Vx623IScPc29AEnTJNZ
6eyV0AXBzexzHjhn8aqNtsLSbp0VKSEjoo0Yf0y+mBYwIWoiNFlUZBleZp8WKHmwFoS1mk3faL6p
cPChvmdkN5NRplqguimJ/a50Uusaj3gYuV0r5sd4qffW2XCJEr3FnslFsJTdAl/9oZflE39ykicR
h3p81Il7kkom4EwFaW4TlCnuptnj5iqMNnklsBOO/VRaoDqIj3SV1xrPrswVjRzOlWcCa5r5ndf3
Vy/9qk5KYoIDBizmISBK0PrNMlYCp4MeB0Ubv9fAf16VUq5hPgr6HsSg0lHS5Z0HhLlIZLGAyoo4
eGlOfNLXOFYSmGldbOM77vtsgQy9EnkXf5VNEQqmQEgYL4GYL1eDoBh4wYI7Ie5IB2UYFSymuOjT
AO7WYW4WUoqsdmEefz8P98LGz/r/C/8o5aC1VHjLy4gvQuzgseRMbH3mqNjWBcMM/oEGh/6BRGsI
k4CIh3ng87+wTfjlCRzaF7pbwiz+lEaLCXz6tsakvyC31ow1u9H9O6S5ZU2LkFnHcFLGAcqoR+LV
vcj3tZw1RLnXzBbtvvCUzb07zyDV2OEYzlLPQMHptt2nBOABByZv4KYbYGy1PUugVAxHYpPZLuLR
PbkU1+R+8JwRt4gddIRjBRRbj10IPK+h0C3f13MpH0eC55dyTm8Xzt9GXVFdYrnolUUMGiUbyoVc
PJBlojCC0MZNXNSpRPVp05HBl/LmDo/aBt/jrOnZVrysxh1CQdG1TvlnTTNRWYHeSMrqCxLBnK0Q
jVHqGYFryiRmevoBnr5CGBzSSRj+A2pp0mOPZ7kpKn8qc76a4qdMvnPIERYgDg6BGFhfADO+7qSf
kwXHDRUhR258SSJMw1t/cF7OrAVOymZstnXadyoU0gQe+oAhmh8i9AFMEEFkpt44nvkrCHKd+0Xf
vovGDyhmq9QmU0w++WMCazIK8QolXlNwZVKB2g6MgzHPFRtCwsTDtNs4Am9iAMupjy+GBOM4gXEP
lITCumVtVcZUZLXnvKo+HNqBZaR7vr0hZW5LX3VqESJSBXX3rCny0UiBiRxpmuLp/lOTOtTvdZqZ
mYDKoqC6SqRd4dGdLs/nZzjh0oUy27IH8YVFxMQBo3KKDFKHInf/nBeKWIoOvZJXbp0mD/esiex9
b6ldI1VIFjInw55GThZyVWJV+/H5uQQyv9Q9pXj3L8DjTTOzWI+8eG0bBbXsXd3X4chggzhwl1a+
athcLRjIK/DkNpclEMXZvKb1UUk+gNLdNgae3o2L7wB1Pyvsx/wX8SAq7Z7jPytJVBWi9LGHffAA
5Zb9b3eHNdLAlqpqsOuJuxTZUsh/QwSKD74ZaOkAm1uZze8/cCeK+2ImUn9DiVoj1l3MlCqy8FFD
TgEkgvY5dNBiAMmgn6/TZIRCrjrbWc9e1VwPSAxp1ifw8GdUQi7A+SOz5YLI9SLxRGl4SfZ3xns0
UEtdcooGrDBdoF10M6cvJI45hODufEU7xuYehbrm/khfi+kMgRwz1Ef0QyLcw4pkpDc1v5pL1k8v
OXtU2OzbEDO/A8xz/5uiJkMmVnvelf0AThjEE00kqUeoBHL+v9DzoVxKv73H42LdCeTY8MZ+3oiM
qbc9tjQZPWGDA9qBsS4oHGRUyFfhXmfZ8NsspE7kwvA70tFuZtKrITTNY9aURsk00JNQ/77L69nJ
qfe7HZAbaRcxp8+ubNEqnGbmtuJIytxmqkC009+VbPF9wKykSNpfUOc0KlSpP5pnXIBrDtIjJ+xM
SopJVQdineDPHU5smkEZYaEa8ppYXACnrWz1D6s5ALSMbPs359kxNGrOwznIx+moUzNppG+7Kvss
5xwBRJAMc0znWDEvG7+jblJPNuX0BlwOjvIE4N9M3DSNdfZRPAtbjWZ4IX/S5rb8gKGErIwlyjBs
42BmM/WBqy3aQzhk0RkHhj0CLAxNksx9KYKuqXfOt6RlSU5D43jW0poYN6SsgBUTo/01j+E8+niy
6h7cdAvryTVcrorjJw+X24EVGIJKqlvgQI2twNAQln2dMnVeedIbnADohf+1/bRXV6T0b9X/G890
yxGc006roLRel/Vvo9rOqEHie/rM/n+lNCGvhEZnEpkTyVtpieUUk6v0tjWtCpEvc0BT+Pi4/bd9
bgDuQGmLT+WNpBeUrD1nvq0qh3vG8Yju0bFO0ar7FefxE7ZCoLKnMX8Yxcvhme++JsDzXSNi+fmh
1CJsjq+Mb05h5WH/4wtJfbOMkMbKMNlbrlcov5NchHucVWYHvZ25Nes1Q5gUOBg++HET5tkZcoxH
jZOr+3XT24iMG9+bRunb1BpMTJRmTMDQXwSPuru5+eLNQiNRQFgJNIvRZAMOuz1UTFV4az6F1bIY
SOfWNhayux54x0OEypQrogZsKWNSrsYbKO9Lbt+BSpv+8hLedrbN734Oe53R4MkJp1AXA7Ua5fOk
gC50I1zYuVq0wE2XefvKhT39eAUPhBstc/lZCBmyG5sWcclkEeYWYqwgfeuwLvxfbWNwH4aajonw
++KqgnWPEqldAgPf7Nl9o3uNrEw4QKzjJ1b1XoOYD4KJElJ24eF2ATgjd8maVniE79/a0GK62+EY
jInNw9jHpxPFdBuRpzf/liIpkBluWpuEOgLVmmCA376tjxd5YX/LnXSnMxcc33prw26IDMCu2Sr2
FV3LKd5zmm75NTy6A59EmjcdCdVxY/qKoMv6q9u3f6MWPYdBoIZCHX/8s5B2fOpnvHFXZ3eA74Gz
9zTFkPMhmAYf6vHu5uwLncxkBecgYxyrxNaJB//EWGqWlB0UzM1oKWw7jEAg7RomhOjzM0hooaUg
pzYqRN65DF8BaWLmBekvVD7UwqrrCzAh14OZeNvK3HuMfEF7fU5qrIxIeYZEH4UGAoZ0cn2XfxAv
2y1RLA6nsBgIyuz/9VzB6IACnlYXHSHXF4c/NojA6mA+M8ggM5y3minijJ618zV4M/LD8sKwzU64
wjQVtN/DXjF4tNAWngphh3zSEGgsLQ3EjKYeLS/s+3IUYJALRgzFGh7jiK9wmiu01eQoaTHx8IJ3
41uauN7qq6AgUbOMY5K5WsK/qY+Y7XdKcK59eF8SIG/nHVXqFVs6G+s1fS27gBdNH771A+TYygxK
RWRPz13PnuW4OMfy9oTG+q6SVZoQ29D7rQSDZBqxmAQO6HAKrmcfTsGZDfUfu/Wx5zK7OqKpJowe
Yze98g0tSUY0h4njxaxcqAWZE9sXWl6k5J9qACjuCjiZKmUHVzXE4Nj2d1zHAyYDZuDvbabD24V6
NucfSWRXs3giX1+JRy6paFoqHn4k1JIgo+JvoZ5cWgHsLetyOVEmnsCLaC0x7rgPS+ZOGkeLdN7w
1S/2FYv+kJ3Dp22MZhJtb+XbR0UixT/Jh4u1TImJqkavjrd0pW9PIINaQ79wlLz5TmMjTXGJhI5B
9RdgkUoPh1pB0Yw1FrLIiAbHhYJK7ceyBDdgcHfjlcgZgbWHEQ02n4RidvBrEUEJmapzRRPjE7dH
s8BHZY1Lx9eLbTNoL/Ph68CIceHkTXu1R1ROtT6hkrof8TDO+elI3z3dzpRhK9IeB1CoW3rKqh4O
x4FnhRxh7GQhQm0/xgx1Y45tP3adAHdwj+IW5lQuW78GiClKE08qtHPV0tq82YpNjF/XakTq+9k/
qH+jTchKEQriEq27CvxGCGyN5w3voR5+tCmIFEERMzqbixgYJ+ToXbCdwQH6ka1LvH4y8cWqD5O9
VrmfCV/OBcHO1GhGO7659MnE1igmpWNBGo/W8oVMn2r1HlyKoNQiXWcke22XIM0oB8zSBwwb3zrK
ZqY08YNG1RzzNs4nxGVCsxlbROnCN1pvZkbeJjRoGY97S3eJfLq1qinY0ZBvxi+o+DksbYEv8BLL
uLs1ZDUMaUzdVpkQoGFzSE0wL3ZDXJlJ3vNdQYDhrSTiAZmH9yExFW2mweCzE7uEnhYn8Bp0chVK
cQyTnrrSZ/OvCxdCNTvEljw0nLnHyn9Gc5PSHT6Sc5myb8hwPTYcS03PxheshEuBpAgmboFp9ukK
1xIopDKu2NmwGyvJDdtPANF3whUOwuaoeWIn/UWtvciioK9mpDmNelwT+Y824+pQYtD0rkJYxDI2
HMghk2eLN8D1Ngznlh2hlWZd1Zg3s9JCcFHFDCtIG6Re8ugsCEgaa8RX2lPylQeyGuRuY7HsmWBZ
PDt0P6ua1i8JEhVDCX1LztKfHzmWMOw1XSjbg63hJeSHpEgfj9M49qPJ/vD/o7n44Nq6zSD0Giqv
JwMAjdZlVYt1E0mF7TRyGD4RtEAjqEpd/9LJ+3lbHnUMLUGLBQ0IL+5ZEbSos9n0yNJAp9nVt5xK
NcWxLUZUc25GcbXGY1h16RotKXCBQ+u8xtiMNBGQA3enioIWMesnMXX9diqNrZatWLVUMMqj8xzY
RIr57Xb+UHW+LGM6VyJ6NY0fAMomc6K9CEBAUtqaBQ5tQofjAakPthnf7fXKSKJ2QiWkj/ThHaB/
ZdTfuqiFxVa3mU50EuFeUqL5KFw+ydtw11g6KrkqUJKfj3qbpBTkhv5+PSAgE970JnsQ2BN/pO2T
gMrCdDv8zoD14tvGZQI6uIki5lG8T1F8WrIhICYuaC13Ch7RDLDb5+BUcY1KrIaKshLLL0BDf3lP
lKtkjpMbD2xZ+lQGD7MLO4DwxjFEGBBcpe1SLqUTJQEAQeOfmdZbdWXnFJUV3TxH5ddnrKgjPe51
0lPzb7tYq4YxlXJ1wmMw2YpP0t2yKo9K2QpZZadY9V9Nmhva6z1vR99hp4snCoEw3EhvZfGpLXJe
qu1Md+7ErcgITD8+YfhCOE43qKF7nnUYmHjFhDdxGKhCJS2IiR+velF11JFsT8vVZezxH/RunrV5
N5PSOFBl1/u0rc4hsOFoQQ8bSNWV0IX9pAciH737Mf5CLRmVKLoFTiZriubOiC4zMAHdsaZBDjls
rb+ek79/ybl0luNaKAtZSim6ZG82B+59QJgn3ruENdcnckf8p01vf6rsI6NkNOphK5yKw7MbXDhF
3WoKtGM0OvZ+ko5HC+q25B1/zUGWj+C/Wm/qLDf2hK3ixNynRQS2cxjAz6IuvrW6UXL6Z4BlrGf9
e5iLF5DutF9HF9by/SLF5FE5RRtHx4UcmYXTTiXwgpDrIB18SKzyzQCMxVFuMiCQpFdoXsjBMwna
MGJyPqzl1zJ5neUMK8K2m4tsxCVpmnSVv0DEHeSUltpe7eNigujpBnpSFZmiO1zhUf9yCuN2l7mS
J99MUW2y1zAhzds5ek5xYi7+2KHMJ9M3kccTX17E7Au5L3/SkOBhqR1W86FgOrgx2/i/UUnmN/g9
d5wyNSY3rdRf2w6S+8Z/mo59ZiwLl9ldUHqFAtoC1H9luxDnMcPKAMjcZAEPhuC0P1bWc70j8ZKD
seFeEUXIYwS1YGHDaH+62iaWKaVhEYiCGnjMuy53O6W6Xo6UVlfOS1J5EJ12Yz0CuS9vLV9tUmny
1S+OMj3DDifIf9nfQZMFUcl1e/Nr/BNyXrCDaEL3PvkXeCqBi1SJCks8nNaEmzO6ElxwfFbF4r92
rxSN+IJ/+COmRO5+KkrIX5aetin2iGoSUnRc69QtUaf7CodsCl8zOHGMoMMQ1Y6D95tPjT2UuV69
saTvSqgpU55HE7DFht4RHzgJYk13NzKssVhwCd2vTafT17M5heGU2gpVmfV1ckqBTfYTT0JxFG55
D/AaLHlMikxNibW4xBFnuBmRCD/2W7hEH72J1+JcXWkHn+wa7visfEblQkf/Pc2rAosZoemthSPI
XT8TmwS3mYqLAG65ck9TCBCAZ47xtkkK6hEEgr1/uyIcdfXWHG4Qtd0GkQKpk6O9+aUQfPVDJKZF
YXdGItAsCrPqAdBbw32aKB+zc2m0vmymVbEU4hXX//kT2tRAWYhMJfkeVC3JzVAadCj4BIfdvZTw
ZY8COGfdllrvJXzchNak09eg02a7/kQmwyRY1bCImsbpJTk//2PiVWK84uBvpcroCpKgNUIfq2Zc
ALlD6GXe4Ifs0tTAAG6I8PEhir5CXxxLjwe+b9SHsFI293EPPAahG1pUrTfZIg5yC4irustjCOk9
rVdJU5ThoHwMMUuEC5J+jQQVS/JaIHelr2Ex8jXuCEftm4CU9j402DjEDbsLJxwTz4fTr5pqJNue
HKO2gPYL5TYGQD66nJGkyt9qItK0z/yDgp9eMvsPuamNiO+9QZRXvx66G2d8dSihhh15PNkH4Xk4
lEX5PTD2fOOe3q2zTCcKGPDCPKlcDJB6h1FD9uxjHF11qWF7ameN3PDaqY4baOy7nat3RkIsdfuo
+bVM84XqpKqrhTYE6XcnPR6S6cOTe4flt0j/ieblq8KAbGOF/nMYgWTKwu0VQLCLYDdSglVbZJgT
PFB53ey0conjc1hl0YFySXv+rgh4HnHsgj+iYNXqJm6LapPHwgfYY12+t3oqTGncTp56fqN30Yd7
cPB704K9FANvqT/oszNFlbTVJ7bpv1LOrN7Vrs/2X0DbZz+leI0wxYVlISvH5oJ7xsaUiKmOeZWl
7KbVrEBJYld3Pk3ghtFLQmivIOoPxu6NTXwYGXlx2LXwaWkyfEo3Ykr0fTHyAx1myeckOWnFSx6E
DjApjIwjQabvesIojgrSRF5j6f25E+ZvJvrRFZAI6cg70Qi6j/ML8bUnEYvE8mdA4GhDZivJTMKv
R4/SrwIeett/cscrF/Fp4BoWHrpuw7RzIakkKB2NRLCh+MJzhUT+0XZQ0u5O4XVMrDl7ceik11pL
369uzud+KWek/MkYXDRTm3OJuixwA0kMBwDtfrbnsa6Cq3H/7YNEMoxzhQkhqFB672DnbA6N5U6z
84VoJpV5iqNkVOUgDx+L5VYKGYfvlsrMDbMmEIlabkrTFGf5LoN/E757ecIhVyCizEIbnb7GGh0C
ZLzq8s8sFXWvBN8oPOZBhhhYodSiaa/ZfoFDdi9UD+CDO3st+/f886aioK55iPFzyQomtbuBQ2lT
l8iZLTDVXCuy+taYSNNzzPqxzM5o/1RBq+03qo0BA6guDq8YbbsiZBZWn+npPIvUl/Sw8F8MkFo8
AHVE9yEuiaXqevBL21cULZGNmEKh4nOMIdPBrKcQAyYm9YGyVCrX6S4CtI88E299LfWpBOyvs7TC
86UM9VSn05SXgqAsh/F0W09kTCZMn30oC3b50NFYdHEf9eiV2qim2ZXbqCN113ruV9ftQYhy0ijT
MicYo+5QjRJGR3WsZK7Xz1ILl94XTX4XPE5F8284oQqeB/8Xp5OUDHHJbirw7gJIQ3DPoXEEopXR
j1/7tYVase0T1tvlV5KCxbS+/p19Z1UJDElZ1VXRgB3BiyU1vs+S1VO3kr1jMET9f012Q9xEdJY9
WoJoQNxxKqI4HE00mkpuYIXGT2IjH4In3W1oUFWjHHJ65tjZFNoh0t/mHBfH/lNHomey69dA+NKf
MPrvUQz1WfQp4kC9tEs43gCJ9J4hJrxh4a/uUzhAWYYK4HTGNjLHKv9mlAX1ERzr5QdLW9dP2h58
eB1BMJN3moZsv3NIMVEudRKgmwuJPft4x+X3OwuL6fOjzcVhgiQtljS7VIgohGevR3EcNKo+BZ5h
z/stfAOq3/cYnvc3vFRH8xSA/6QSUkwF2mKLJe3bEbLt+2pdqAVsJlBZzVBKCA1par2Gd4HhFDax
myoTeV5zpbsUb57NtjWmEYVc5ECJEdzDmzKTpjfljbEKZ2JArjRRQ+9d0FFcorlsOEly6tqsnevQ
YPahPsp5zXTfk+AqqL7ro2bTT17g93MLj0OoTuTp0w92qQ6oHHT7TTZX9k60V1u14sMAN4yEy8cs
rG+T7KMoDfR1lmzst6j2NOiGn3y5hKeKL5Gx2gFAY5KAKfJtT5RCrcBEoTZYS+TLHOfxeUvk/4yT
GU2nb0Yg9lhtP0XnySLf66a9QUbzXDD5HSrArkF6iwsm4JJR5UAR/g+Y2LvE9BgOWdnF7UR3hjB5
tC3yuOspYMKzhiEzAZiqzsbSxq+NeK0bEf8mmHFf5L7wxpBr8NQa65VTSlFweZtxr+kg1ELc+nOi
m4rTZu8FKUHhwAMKjss5kD6MM7lEgJv7r+YwmC0rcLAdYl8lvXZ1EpDegZUI73Q3zXVe6q07fkjO
/VKxtZuMZH+Tk6WkDOdJfaO96Pw8q6KnG6GIpt8RhQfe/eRPcmI5PsXEsaUOCqI4J45PB9rkV1RZ
4IQ/yyilZD2+qBaVc5QiyCQ0jbYDxhoiEXtVLcfxGdP39/IXlFaezEZdLQvp542AlyiGiIq4DD9F
s7wb6ig0DPdK+XWRo1rRrwhCYxJiUO4UYEqe+VmTHuIIMM5onfrlt5ygd8nphqX4n0KmDcA5AuD3
j6UY+W4zIWKPf8QsHeL+UB1D1P8vgkaQB2FwyAF0JxOHlFatZkbeElSe6pMLreWuNdynisKbRI8D
gpBuTDqbKbX5ook7FCuf7NpWs1qpEaif5dBjvZZINCeYbAL/f/x+MsUy1Ml9F8qe5qE3x5S6C9Bl
mZYdIN0crwrd2/E8hUf+b4odUzvx6sxSTiJPhJaqI1Cn8f2d3AX50MIjiF9vgAbQjL7UhsC7YoK2
8HjChDW2ofV77arT2wytAO95D4Ro7n+dg2V8ZEA804KKPdMJcS51IPxbEGgmFEH5Sm0GExJwVKHo
VHkHz1gKcrAmZ5AOXpZ1mO7btagesmHMw/tnJGp4c6/l2W2Qvk+r/eXcMVWZI3UdL5fj0F9EBflY
MGMGFH0Mqjgiwhzfg/up1ZYVvbieO7VUpZIz84TVlwUlN/zQPJZWW4calnXX9Qik4zlEY/Jj8MV4
ToClF2phraXPwogYZp3vykoJl7nLRAxNf2mUa6F/Zwj5s+AiaCNbJ61pRV9AKuIgyL5/suv0Blvv
1U4e06BdwWnOIXBBkZ8jj2Sb88eDOuts2MqJAK2cczWR1Ug2gliqtq9RmHkIhV1w6QllchdsBNmD
2LZg4nZVRlkzPMRd4oWPsvV2Hl44F0yBr8bzSiVI5EvhhXKZYtjmotXyVjHXo+pUK6ToIIW75QAg
zfNxsnSWhA/EzCulbHMl1zJm3+An8zJd46a0beeRmaCmAp7mmOm1ifccvf2U1pOcEWfG2+CtG9jw
Udrtpiz9zf71tOmYh1rjQpIv+ulJU+Ijklm0tUHi+7OYpMB4fJfue8hDVw2sQiEhFx5nGmKZwJ1W
4S3BV7AdkIwn9ba12SA6Hb4FLK+pvQBALCx+ULWFpNqaqDZo5hKec/QUoTQi/h9QoJyvqs9E7BVW
033JUdD6+a/78zWSrMMRJu2PyxkUssqwhgWwOm+S03OECmxW2qUduiChPZv3UlNVUgJDE2KV1drl
TQy/Lbk/t4CbZKthCVl5EF7v39XmAj/ntNsgd/k5Yc4p1Y7CEf2YIIGf/U8hPYU0fv+u/JQGOjvB
pdB3hw3NkTzW5rbGqYhlnrmrQR3dJFkSKjSSsS3UG85mhHfNoNgIhAPOLW4ZzVfwDL/iSZDJ9UQN
ktoMra7YUxkuXKpHMb7WHSzMpAsWMIcZlQudc23ShvRNLlVjyIaNrT2ICoWki72ri7fQ5WD+Ajlz
8GhZlgW01q1XAzP79AdRYGgwqtY5QixDE8s9BQAQTSXWStuBG4eMWe65UbEVcGlcv/9Z5y2L874E
OxWJ2GCCCZ/ybCFCqGq8+McpCpZYKKOh354b8opY5JUl8dpno+Ku+bQ40+Q5PBMmOsviTSMksAGh
45A116x3Px+C8DdNIfnTWJ2lGEnY3ex4Ug/5OcylzgMPuELLCPmgaS7kfeZ7tjFUfR8ufm64EGgY
H/JrX7kQiPkYOSlny0dDjV9mWL+3CObBlsBTkBpPO9JDaffzZNqD19BDAFqrkHyvZCFVkrlPmZ1+
+jvMQwQVN1LF+ojqkO/sKWL2WXE3G1F4yERVqwU3yGe8CostowxGRS/iZ1jh8qTMWDPG6RKrYeoV
3CVAUFDOZ5MRkxNveHrNnEXjN4antSFtxurcAYrHfdKGv6zRtLWIw5GzMGJf0+3zqy8cCUF8MVjM
1Bz61l/YMt52gkG8GAEW8peAazFlotsyN4FTDaD6f1d0NuiDUCONfPJfa98iMUpfxAfEXM95oOxT
5usrfZMD0iYaoZbvS+QcRW7pymmBSLEXNLKtZMljdy1CacTlA4bep5FW8J/ig9+LpX0V+di2eob4
oYgrwB5iJ+/CeVR+hZkiDp1CCcbVaayxFGNbVyyGdxcH1G5bqhDFthkwjt10GcB7FoL8CqTtjbVM
/PZS1uiKnFRG2HjZHZWHHAE563QjExBIef8rNHMuakjRycVGuShu1vufKStRPI5/zT7q5nhwdgE9
nTIOc0Ow6t2kOuEVXe3wW88etW6TxSxpNyWPMKbL/WI/3IgW3FiQKBfxM+Wv2vTRymRUvk6yf2jS
n37Cn9ZTuSVbWiselcJr/A2o241324gVmQAXr48ANHePYeveoFAjEEzJ/U+cr/kxnmyTaazKAtb0
RjlF00064FqqxTtec9lacnmKLY0K8HLA5rXURuBEXsuhFF2nDHxLhv0ZAP9g+q/gXfzcTkGeg9L+
VckT4F6eftgdR/qVmsIH4wTqhxP2Uu4ys/JVRNNMJQXj9RjpSxSKFC1+n0HSqs5HVHEdc2Yu7HNA
Ppf1+kChgJN/kJB0LD02RHG7qzKLHw8+tV0V0ULU+9sNbMDq8dRnxOtP3lUm8ErLng1M96AhtgmD
i6FIqkLGGVko/Kic0Km5NyaU2zZUZHyu5rgQ8MVBkuwcdCWfdXPY6ZoMvKSV0CTC9b7IIgGl1ePZ
4F0QngCYHdbHDtEUzVIvrIN1DlLIwMjfki+liDNhI5C1rKKWKlJSs2UliQkHDh+g5L3dfebG6xqJ
5O25nrrGh5bTuXlXY5WxZO71wE72KsMqUHaHOgcunnsE42ZZQ9sGGHe0lCm9lMT0qIH/MgRou8YI
z9N3CbbvOvpyZSyaYHhzqHopemFIgInZERapRgtf2kfvYMJsVOX10OmwWbBpEjqod3sHvReh8V8s
DyzQ0bvPrEdcImEiKfLqwspvOXuDiGrKlR7Qd5TOfnlgogwshMX57BM3rCOZdGoTabhc8LMAn0/S
OqD0daH2CvJeQ4XytLhoN/QL9r//u9+puVKJRssDbkn+bXrU6ia7pIndMldlqOkWBb0lGarrxy0R
rwwkxlSNk0lO0k8nrbuuFVXEaSoQc5uGN/QSZbnr9cxovjjzPeWBy803oYvZS7EjJeBElyVW0/fn
NrQInEVTpkc2k6pPzPQ+7JbFYgM1JXIzrukwTLsvyiaeYxuoov3pPdDX9u952dBidZ0bAIUKdHF5
2gGdcWmHa6KkFN+wtIFETBCK0bKFG/Xnd/UCsfcodxBdQcs4Ow9iqv4B5PEH6xZ6GbVTMql3TgwX
EADrMcrmQ5vBsJpGYum5uuU8MDJjDWR9z205sbHdiK6zmaUYX1Ngx40FtqDgOWwDtD4Y2lbmGum2
bynG9U8pngfV/hHp6wIXqfMFXFDyMDNxtLG6lDGhgibadzHtjpa/GeUVB0Mer9GY/y1TfKLCbkrU
rDz3SI4Gj5vHrtoY7rSVdzsfP/io0an5WL2aOw/6EbBx6jvsdEmIzXpUZ8JLetm0ILfBByBIeYDa
TDny8BDZVjWR8BMkgeCJBas4TkNPHsFqTT2rtMb2Iz1q6d3dMfR1l6+I2GZGKCVbsjMZAJ/3C5S3
L7WygIo6yyqxZBK7iMZ0nr9Mp6ve6Lq2Bam3HNsH5H8tP9dbwjIpIgkrUjyK3X7xaElRuSfJMXap
CIjVB4qyS6ribuEonQR82oKGpT70CR2VKKek075VOf73v760Vx6W5Ok0SlIPSI2oj5GaA/fDtc6N
RBr8Ih3st+gDntUlKHit5OWDWh5+maDFKjnu8Xvz0k1y0pYtvOl+kspQCO/zvpEyZJrB4Zt/d03g
nPAY/pPtnjSrwtU6/o16CXDSdfi5AqV9yD30Kp5ltzUjPo0Vm+a/LjROHGLfh0hKLwF60gBhWqvl
PT0xg04jMOE0aj+jWqhox13mKNubiEoluvjTiQF2GofOBGqrSc3Ta64pE0zxfmZKdDdObTeoV9Xi
tZ2MJ4Oq9O4EuBO+z41Br54aPqN+PbZ1KgAGTAmU3d5v5V6ap+NhJjvrBP7paDBqQ2m2QGLCnu42
niwylqf9xxSggLnkec/+VxJ0FXAOztGF/pLdbocZV7st+HILPaTklWQW3aa+fTOWAFjQyWpe/9oD
Vtvf/5APo9w6t4KHNh6oukRfgJ7wq/ZGhevEcPr5lAhzvFFS1GoUP5C2OeDVQabvKuegi27ePSEw
egfK/6x/K4gqT/M4oFkJkxz6LPoikWDk/oGPblp9OoQ2JDerWuAE0jz1iKIAQE3/0+2degmcCb+W
Kw9VIwcZX2kAaNeXLpgnyo9HuFGxLLJYqvpUiTJJkjs1uTCC8+aENmLJ9T2bgtHqkwT2ba96iwHX
P0yZWBbJ+TlCXSOnUE34xtiHFJ5GmdJHAo6fllPp8omqZXPWjkpN0ITeWU32UYTLeJZJ23Z4FmB4
z8c+GMal5oHQCbjOdornkF81LZxWwrG7yqiUBEYC8ef/GuI9hlkTRfdhai4MqBZ65PhH1Twgu89r
NHiYR4vtJ4FnDMVv2LJgTsq5D89Y7dG11lCT1mJME9YOu7Xv7Z/oPimpEQoamYiS+vfvAsKiwVGO
fe1A9/F/GGavvdyO4fAtMQO/ezAPOHhaVVOu+gyS6sPJ4GT53qN7ZML9eQaT0czJhuGWh8MB5eaq
RxvJ1uhiGiPp6Sd2RLvbwnxC7yFMwTswFDXRpBuE7XFa3vHRBOFbXsyJM8SRwCvoi+oQnSRgidyV
xQCbzKmiMhFbteJuutIdSF9NqEOQjPv9EqVHvNdKADIKc9XHricKT5YTHcvQF12UKU+j1aJujpnn
reJiB2i56FoU3PQ52OQAEKJiXgrg57NkdvDMlLXSHSI4wiEYCxeAKa6K7S72Nd/tEhZEtuVeXL8b
r+oVPQr+pZJezGxPOleX58VBa+OjfYMTzo6hcsN4J+gQtGR7CQfA5K6uq838KoPRoEtW9cQyP5tv
S2dY+6PGtm3VXzxp/7Krttc8a2xCkCeVl2pbqGBBJSSYF8XMnAn7dsEO0EoZVc2b8yMOnnppzMvh
ED1p0OoE1DdkMTKfkqfRDf+J8JPWb9q9sS7TdvRMW8DN+Wi5VqB/6x4CJpr5e+UBrKCo/ml2ydt+
77AdF879/ZED6RQrSmRI+nfQIsUx1XKj/RoAnnMEN7j5/ESquz1gD+GVTIMdjGPiP7Tzabr1f/1c
jcHuzUf4bzd81UHCG7oYW+wymqXSA+ca04rIFl5Qr3554PSm1Y1k9VqamZN23rAYsbJO5sahA9QM
ZEA0ckDXBmVWson3Z4La4H3n3eknHf8ZAjcaycY8F2/xIPYHxxQNHTHe1spkTqHYEhqX1vSmkZ+c
00E9JvsdF9rs5UeHFNhFwe9KkGpMIMCvg+waCRgQt4iTkAFb2xSNIfOCKi6yz//xXstJlIcT9k/l
A5zVMv/SvYTMyyrWOn+vIcffp2ztmFdGUbgE8k5Q84A7lTPDQ7EhuThsp4jMKFXwM3exyHbcE6b8
HtKD+HK9whsKXsMZNtLSHiPinhGJy1iXUz8mOkBu3xT1EajInRkzv7nZ6YAbqBbBZ5/RhlYIEpTD
ZBqCqVeXTBdmAe7khAI3faquIcs0C78ENe7dJ/fZ4AsXT2235gRKEOvZZsTuPCil/fTrpABmUxT4
r/UFzO4brAaxdEQy8A7QokyIAPVzMvzwR5MtZKM2sAqWvts3M4UVGJ1PZAzpIec0rP3AD+V1ekKq
jDZa7DidGSmfXBqzCil2alW4H1IDs+9yONjtaTlDYgOFXKBjr/ehOhaAPOjN1MliAS60i0AIATTx
usXxftCZbulE8fFsQGr0kDtwWKCExfXjlxGxuauwdXPtegcr+sjY5Y4FZPt7hoEIkDf1YBEHkljz
YLn9q4+e+zXI2/A8Fjig/1sOyb54y6SRhZFIzpuwGTs6VBNPl1kmHbyU4AvuRXfeT+ngUUMWCf/b
Gj1ht9GdFItJrY3wioHdAZI0pz64pPbakjpHJEFrzJFlQKBirdVZj7T9KQuwqYTJioKT7zTS8hhQ
rmem+xaZM46wyuUymoA0wQAPARoWQimPNsENk2Aaho0lmo30FH1kCLeBDt5nmC674PSTd4Ms4+/C
LctN0twIZGkhR31GUiTdnt4itj09OR3Wvgu6SPZ0xfwUumamTdMQFYqriM0+KftHIypfUrm93wpy
UfH21i+AZ6IedZCaDlXjQ0WFUFtZGpO4Ie4fAX+peEtSe2MGeHnTGfEXFD9Ht4cqxFa2mTnBNlGz
5HeWo6gVBuZfBadCGyjrQLkisVHqitV7P2mLhMaqkJbvUB0V5a3I+MIwVZ48etR/SYWzhiv//JM8
PzVVE52nyT/pHJ4JSeBD1f2ObE2Ywzq8KndUfEfKZ6F6XCaK5KKO228EafSRNt+Th5A9I5k12o+/
+GLRDV81em2U3Z5GiVX2wENKPqUe2G8GDEmkFP2u1TYVvgArBk2GxZGubf7ZeuAvlO2WTv2cOS3R
rEVlaoX9jU61zOvRnE25uMpLeJ2iJwcDHOak+RGasAmpUnjlfy++/hTl0qXMAIO5zrSvZRKrmafq
mFZ9zVWvJ3gFblVUEqKs66cIjw/tLvwcAUFD0WNLD3HR9zRtTkqgEWmTB6kdWXFz5uWsvBmDqwaL
Plruv84T1PELsc2d97Ek9wh1sKvpcxzov7T+iIO18hr7ddf2buKwspP9SmKFKJsXMk6e7doAzPfu
4OdrBu2BNrzyb0+5FnjlGeVgdGNGb2fE7eh8QMnPh1CorkLnp6OBEtdpwXMm4RCvwGujwPv0j19E
ynuN51d8/yjVumX8VqlVUSRp4sXC3ID1LrcyBetXtAadBa0j7Dv46xtVVW/arm0r++WK8/xMElny
3xSAUnjP51lUwDl9TlY8fkb0/vfYPZ4t6aZ9ByykM4sX/iGsyT6s5wvgtX+okS2MlRyOb+ROEs1b
EQEs42R46fRd4AuaKIPZEVOGi7iy5WPnt3XhCgcYp7lSQGX93N3nhEdZr0RFaeJch8DyKsYXBt5C
N0G9m2vkrbsY2RiAgMKI3DjTehTyXXmIdeOrKxRSd0j7C1ZiSMfIgO/3+Nfi14vGmjTfMKr1G0At
CvHfCZ3fUWG40DhWKmTQB7yV/wd+4mEA+Q+JNtTAQvJHP5noqhpOq2NXzYkTNYonf7RXYNnoEYeu
9nqq8015YtHiewtqpdZnHpEZMdxxieKMC4ZcfZOgVjHJYd5p9jv/rgMBrG23ou5mYEeCGediQgy3
ig1QQTknLWmmZo2K1+iRbnEb4K6ipkgQuPsVvnT1uSG2BFnivsGuaPt6+8bo25F9RvTELvGsKByW
CdSwtLlmJ64uCmOE6R3rpET/oAZdRW/+G0IIsBfNQVW6CduAfI+QUKa9E/byTLpaugRBrUMRaXQ4
4VJ30pTUAHLcCjeGRkjnjb6IwsYf71qUuHy4nsePfp2QrZ5eMKP5s4am6wdeV1MuzKWDP0ivOdyY
s169VObBDAU/3Ige0WQuaYVKSmoSayIk8gyydDnT5Pxv+yA7jTPzS8dJAdgCKs+3T+UoOsC8yEa8
VI95L08bTPMseo0XGLaMzQ36L1N6baKjGOQ/Ki40/UOfbiOm7iQXt07mWFnAFv84DWs4mUWDBWXE
nhCD6lK7xdzwK/wmUW7CkWHMDpZDrltQhLyJejH2tBG2/0ydMJaphF/SOWCI4Aarwlfha6MAuIct
cgPqtFksQh6CEUDfM2xlnuD6PI7s8MJe1Y0uGuEenMOz4R5mHIceBwQ8wwcsRXJwbFWQWEghuHmh
M3K+XdosfB7/TLwNciEaVYzcTeA7WWISSAhNA171vRYmhgk61qKie/0C3V/Agz0jndIYEl4JRe0V
cEVeypn9DDE6cnzYRYQMRuopvZKyMuUfgPZbJz18twEvBa6PU4ah0rMoYQ8URCUosD82x3quHmsL
qK4HHh1c0x4eMnayrd4sxLGWayLi6wH1qY1pyAjDFvI0nLL/DXAIx2yc7s/r/OBB27Uf0LQLM+3E
WJ2DgmywmfB37z0YMaIEPVTLRQJhl9MFFML936+F3zoNZCJRlN7Iyl4EI7mjMXHIR0JyYIaQ5UiX
g16/EoWH6enEEU0/5nGmqe1FlEbmJv1pBJ9FXuUSHcw0axsHC5QaOoo0YH4XErBUvN3x3W23GKWC
v3VK0epFK7woDz0auNVv+kqr7+ZAlArUxJuccbhCoXsDzw5oVUmd9Yp/KnGuGSurvbCeONY79A1n
WYf63KjwUYSYwf0MHInzb+meGE/6Y9oNf6GETZLk+L5OS5IkQGxOPaF83UTuqkNyM9k2Sa9CXIJo
JUjUw24ftJWAzRxVio+/OaWQrBgotpZxa+De6o7FSjv+L/O7FIXg29vAiYe4eT2nW9SGvg3vOQ7/
++B/++cqyWWlT08WYDneD5lKWcxwwZ2hhj+Dkfng3DrJIzzllieRI0LUfft+vYwZxB5UypnXkf2S
7yoN1meEzGgSK0E4QWGMPv2UHzADgemmUmq9TTMLHx2PcYgUIUACok8KVg8FO3xAKjdC/xARgICH
oBXDLiI5WLjlRF2AvmgQYlNgoEwkVPFgVXnI8m41sWjT3upmIt+H8nCn5tKRj0IKX94iTdKF2iEq
fN5iseRVpFEyv2Uu/C/V4HZd8wqLYln+FZ/4vFjSPHcZUNClJdK3l2w9UiLJ96V0/G6ClyrTwxSS
huGbyQKuUpRjA9neHC3VXnQDHV4kNHFk1q92+0pR3lnBjKW79Vnyieaqrs/ItTCMlKZJtx8alp4Q
FJV4inyPt0Ep5+zSSClpVPzwzFGSAlYn2ro4s3c5zWURXMZNUW7YM3AVj0fWxGC6K3ASSsQIr4DR
Y6HZ4b3HsPjjZxuUX2Rt7UYBoLeEgXFN18nqWYxAnq37dwpxMbxFQQQpMzsSe0U3LRKnCv94xiQY
oZgViA1LRehcx/TImburYZCoddcHlllJZt+92X0BZQRoiTMNN0tBKgJ4hLkb5FkKoewRaJT/69oW
WoYHywTOjVozS/IsB/DzAh7tNPViw/NYTcAq6aI0u2npWfO0wDsTerZdB14NDVQn5gRPx5P1U5mJ
5k1vqaHUYa3AvSwI8sV/IecZIjo4L/ZLc8SKDOBsl2Dqjvx1sjsVF+JpTKtau/Qpb//cFx3OUSqd
dd6xozD+yPx+k13FVuIkYKOe940s4dN8O02sRClrwARsuWsrP+L+b3Sjc3CWlpEMuncllKsN8Hv+
XK5FEJeEmYYD06yaP6wjFd6dBS7wv1NA9ttSe4S0ZXBJD+GJp/JQcK+/J+1teQUSErmjppe1H+W+
OoMATKVX25w4i4n3JDZ2rgJqtunl6TkUTHzE4wcuGQs/LUcFuks3MN7arG0VZfTiPTrUWzt5oN8/
pkNAe7jobCBe+FXXElzl/NQoNGwPbl6tvCOYR+Utq+YKUtMTNbrECSN7e2vXqkWpWXxoFG4tpqbY
b2bsBUxgvZaLKDgz+aDQou/TsPWeyVsGNZmDzzxe/mXwIe151ADigr0jp1cnTjd/cp5pRYXzDvML
lRZwbhxGm4E3ryhdfU8232kOut9Ani+Fq5oNdbBQfVgH71st2RcUVZyjw8WJZIZ8JfzLl/lRPqSS
aguyqBEbxIFj5OxkMMWXW/l1Hc1pCYcPmZECGn515qZjQIw0nox+VdCX1c00mFOUhIFdEles2iXZ
RakrzFEVWjXFNy8GrQAJu4EOhPM/aFYRrjo8nTwHLync4OYCv6s+ER8SxP/TEnxqPbk05Ez/7KJF
gLoGpramXPC373v8L9mx7vY206nRorveZQf3poiZljTciN+xarBAXO7miT24gvQELzWbWEFdjRs+
M12U5UcI9M6kAu5IRANdp1dgK9glCQHNWbprad2gfZeQbO/OI/eYnKUIgyquvQrq26zgJPYM3GiZ
OjymrPqMV3GJb7rboHmEw8JaklrTCv1dRIBILQPcrWMUFt7TRIuuNV0ltNT3veNCfSclUvefNhfY
GhctEr3yfJ1tGTVq1q9cObUjblfEtWVvpr3/llSmnN2Ndikv7slr0S87jL980Hj4WaDUMcMFh6Bj
tK1r+ptGnoUPhWmi5uWyWiWvXCBDJBHsGt9z72ORXx1hOGgeopYsnpt0jlhjzdTGyTw4nUA2w/5W
t1aWq1Z7qtsETL6sAMROjniqT1ORklq42M36atz4GSsUn2ZIDIunALJGSs3XvZfh5hRKyT5TF6pP
xczffglGQrQXIhZIw1/JmpOhqRaLkKnAAFVU3v4TX8NNw1ePVZVDGL2Ze4VsRqDGreb01h1B/J4U
t54laTD3vCSt3apIW9xKnOkX9xYzDSWXoAoVoreB84KclyH9wRrGxDndhw1rnGysbfNr0sQPwaFN
DYN1KaZXoYHpYoCTFjejQmEwuY+u3mNefbntq+/+hKJiIvONNbc3CCyspM0Hcd88d5tmQlwB3lic
mutgufQ0KVXmjiZfLkIRs8cxX/uc0lp6Lja5+Zfi8uqLJK3kbyHQGCaZlp/xJ6YPnsf6JgPWFYyr
1pMouPgKbL+buUb6bemEjxLI2XXoJP+OvP66yjFgErmi8/DbwLs9bwccL7aDOr40bZbWrPZ9kv0d
gv/wqoi3O3JXH6E8fjjBr1xnk0c41ygIvBthzExlCcjNGx5oH/AN020sQ4n5xip6XPXyaPh0NCFI
zwiL6pEQZzIDx9duYL+kE/A2vngl7CQSRq8vy8t7UajT8f+hDQPbqLcp35UEofwDjnk5PcvxtjNb
1taa5nrqU32RwdVny612GLzBIbqr7/ecpFGztkc7ENwCCGbiBdP/ggjosvYt7xe5w0yTpemadn67
P9F8Ee9zIvaC4JG/CiSE8NztDrYssxFEOVww37dCvZhYjSrMrFjFfrd+KlN5pKRRNkIzNOUIuPhv
+dHUck4y822DTOR4hafMI+5yaeN1KeKMkdpxxooJCLfGkrWZVruIGNEA1a39A0xMSuQCuiv7ZgoD
noZong/QvGKSYdDYcsHvwD/mE/gT66YktHpaGgwScDgGAwzSVZTlvgs3qim5KNYMGhQah5O0UgnG
7zC/43WpTXs9+m8YX2rLytXJWunfdDNitQCza04WCJ7QCW1SbSl5XAxZ/i7k9lSPbQb5Ayrk7GPt
ob16AXnoEC0swqyjkk+ExfUMzxrqWqgvnQ9Z4uHtWgEVA0hLBnWuZ/F2fhflJHO0f9b6i2KDQ6SP
Gj76BkdzCfSFkgkzKmGO6GsTUO3Cf6VaD+F7GSCgAt8hR4ItTbXE6qOyl5U5HiUPCHtcrgYKkyX4
1s+fxFiFG0KNkJkr/VuKgUxTvhEYBVwTgzOzaEZc0xfylV0qAb1btMFvAseeE/vfYUxTnZyTvSyL
yk8eCq1LF5zvzpx3LJNjoDmGhheah64M1umSbqR21kZZaFk5yfHSpGl1KGSNRCfDB06ph51lUUFd
J2PHsdEEZaB53ofJ1Sa18p7LPo77QvuFV9K0ikWdx9RYy7A/fKJYNeSwy84anE6i+ajrjzCXMLoy
uhipX9wjDiLe8Xh8kt02eiYhl2iBiT/02uJ9teUYdxg9iWqwtJFTYCYT4e5RkYZmof3eXE2SOsjO
oKqCPp7k8P9oB1M+S6QRsCIqFL8qMzJOIO1IW+VXnMAZZeOUP12VV300NU77zHw9fvGhv6HrWLzo
zV0oSiyeqGIweY7OUJO+/PBNNjfCpAln0bceTtPb/PQYUo2gBKffhprs+g7GguMy6drc1tE8t1dU
LQ3Y8xoinvxJLoeu8mfu3Y4wnoWvAL0X8YrmP+jpG9vRVZCpjvNMBpb0B8s4RGLi8ojBXcimV8CW
5QUR4v/fEHoYX9xvsTMzFe5yBsPEXuJSURWLM6xa6OZpeK66DiTktsQjuTVCrC84R1pnuwczJJLd
cIvQTSuI8ewm2wjpow2J7Hl7SUmJQGMvTa5jTddqErUMkxKkKC5S+6OVOaDs2IRWYEC7ns3XaIiq
u78lbzjIwUW7KHPcHQJam3Pk/qBH58ntHpxOYDI+qWV1EzMf7OV8FDRiR+w6SSXfm/5o900knJaJ
2EqwZ/r6/0AL264GCMRZSwPcEYXEbU9KQuc0MiZq/ZmHIhftM2WuOMAA31EeNpnVYIs9HUCcL3Ww
wK1XE85k8WPDgAys+jY59WUWa6Z4EWLczPzGCfTQqBWn1ooWXNSCsQJipC4GqunPazDGwsK+8UKW
jDz7Eay+yTrtJc9BOFoaFdWH7kU2lNqcEEKbGKAoiDfhdopjRUfNrqZhcvCTj8QcTVsjbsa8C4ge
oFTTtVKW9hWzoJ3mzZiyC9oUxoGY49yPM0IUE0uLgwh0qu8KywCmY4ZOD6BKNRxupfGs2dANL4aw
XYGPFghPOch1z9qROTlznN3Z8IgfFWBN4tsCenAIC/HZlhKKZ6liLVBLQN3Tvk1grP2Neiz1XIUx
DeeshCt2D0nN3STYu9usJzg6r0ST+aVS0wBDIBYuBGvvP3X+lUEo59V3HQwcZWr0EOOH1sFHfLit
Z2dckVbQrkttgsREJ2IcAv173xsZ+S81cid/rO2wyCF/2QbgNHn3DBesT5A3RIrtXwG4pJvKR7Fd
GH4+oAutvUsmF0btO89F7Bs3FXp6Dmki/FP3VcWm70QCnya9xGoJfU1A7bltbkxllCv8S/ZHFMBM
ZM+7hW21EQsNO1Q6GrjAagzmBWuF4kc+ebJBXlXs6y9zQmEkdzOb8Lfm2SnFgUP0tduJprN2q6BR
8psDsBko+vI8fgmg+CJSO864Krsk0Z9zd8gsTG+pIMbSXxsENNjCFVYrIKEgv1T6ihHx/cwmw83w
aFmW7x3zE4tOMUaCQtf3/OKTnYCGxvWp5A3s/zft1v4+H0836TMcug2uP1A7pXaMFYerXNM5jtAk
xsW+9tDqPkuXJG30J/FWtWkeqfWsS318R2tdLfk0bPA/EXkMEJCWUmgK95kUwvc9JCAhmNj0P/QT
PsEGpo/aUdrDrbXuDGy0/ufhP530LfL06SQgbzA/qWDfOPzpgSOuRTM4+4dDXE+P1sOjHTJk+f71
FVOjYlvlzlsKVP+fVr7Wog/q8briNAlFR9X3+Stfd+Vd6qbCuuOPc77g0R3MBThmyYZ4qi7QRI8h
wUz2uU/RGPHHxFSxS8Dg49MTucNH1Gq3vXlsv9oOMCIaNWWBTj9kaRHEvl9qN88+c0/G//QsVcze
0mGqSCqfTVlYwRxglnsnMny6C+ho8msvaI7EITiGRSGnuCQqncSVq/wuOsGMC6q+Te0rNWrMebP+
eAxJyyS0EZUwMUxHRPM9VVEsBTJXqC4Oi2Xs4IwelTP3rP8O4XU0FNcG6YRW67ZlQWPldtCkblVH
i9zGjCgwBztcFuilsNP1HVXEvtoyzH4KgFhN7wNGrUOTigkeZJaOGJHTlbIzeKmIAUAmXCiHF9RZ
0hCmLd+NbVEN7+xTYNzDKFsmiW4/78P3ybAmlR+SVsxNukkr/Ax7+JzMmklP/fTKw4XSQf5p5gz9
iAwM1gZhq3XpEnoTp8MxX1gI1rtWcGKHGtBRONs+ltH+hDM9uxaeYYZ1POo19AT3f7lNUF1pXDmw
uVsDxlkJJzoIqdDwy+lfhL1ZzY4o2eGVvns+y1Tt23BQasmaOythrcwfe6n/2o7vj/092+em2FUC
YqEVYPfPCoPJ/ZNenEPBMWifleNEUmkVhkPi1qHL7SseXQrPRdqpUvzFHD+mhkT50IpgMogljbkc
W+hDDPtNm0JPJxdqAdKf+uT7zc8mQzYTSushsWCSPTxaeRufxgGshH6Rvdz3EP3OTP88XcG1n5Au
zO0LzYedT8pfGLRr0Dn+kzjdOPZyH+C55jyBBauldOQKMCF6KwU9UNpY9/bBg38tgRYMZUxME2OI
j+205uplrWUI+STyeqdzT83XeKirBnErlA9YfpzCWZC27xhyX3RK49WRkIfxb6rBge2z+hz5u4zF
Vj1ho43IxyF4NNxHPZbmcwnC1SNyrDRPMJFyrrUqj4EtzZT71cxROcsoSeC7DkUPP7pfp+XHQore
9v9skyeQVPeocBUzK1kxv3OKvMcFviOE73vNB5hellYE9zYNLr5/qnb35XyLQvDfSkGEOwCzIAq6
O74Os75i2is27osDzCOzGegvvl9jJeDVIGkMT403UZ3H7mTbparlMNJ3316wlMR/7a3B4t03YJ1V
jL7/pRdlFqjzFKF3kmzMSMG6krTaUg4qpzB4WiOZE+LkoQdd/3/6NSpJc8l5EOvsx2wynFPLUakq
mG/iiO1QPdTapppF4YR/116G+YjpaWkHkxgHVYltQd1TD+S/+87h4OVu5ZPr5tf7kF4OTOi2Epl6
pEJFxbJKgH28E22aNcmcZspB6Kpddw9r2rLgl5w68+SyHR7skpkNBXofT7X3NhrDDv87m4PON/3Z
H/nrfDkLCUT6hP9iALR71UvtGyqm7f6fC4EdfURu+1yODeqc5vrDUdz1Vuhfw7c2khMg422d+rZL
sY4wV91KeWa7JzK7e7Jj22FpYhdI16MFjTZVMiR1TzOgh5ryvaeWY20g+0b9I9GkFlZS/5sbqqbi
NcLWdNe+rcaMvB9IN6ZwRPGj3qbfSQH1NXbp+ngPTPJ+1ayaBIAYAI49gHXGg0F7Ks476i5BKIff
DMUjT81CUyuP5xG72ifPUysl32z4ahaC49TIyLgGxX9wpxIft2qxn8FBLlBdi8o9rh8wuQ7jrXMn
ahDGKpafzhYsVPHRKKyvOvuOUddyaLjT7ER0dXKOu9iqJHK6KMqXTevj8krjrY1Kj+aXGF4Cakw9
co5TLyADQFZDOU/QBW2Y5ulh4J2/RSZGQQ+slcMVAfxTgL0xoDrgk3Nb/S+CiKvbgFQRv3VKrWV4
OeFVFovzg0phX9Qdu1Vef7nhV+kHlY9DKLi+xkwqy18CpWX3Rts5Oj7vG+c+dGa7zTd7P0uS8T6v
t4/+rU9AtWUgJ1/O5OOrKVvWlmu/ROHB4g608TG5BwLteopxNRSBO17rWHi+7H/CNbxRXSOKJTEY
qqJ1UF3WykpMKQ+RULNhnE28zOSao66lkilvpz0x50TePFdHLSOPjhQPhnv33SHyHizTPxdYQ3O2
JTnbLwX5MtGMgrVg8QSNl21uQXOLVX1Aa0PifYU3gGuoY+x8tiGzOh2TxddODlNrHYdLB3y7wVvr
2q1r+qbH3yFAOuWVE0iWJzx9Za7mGdVgn2kcb1Fk1IP8jM9BatMv5Ctur+e5wDet4/oZvkLpfgzS
1MVMiXg1upFZL9pkOIEsi6xFrYBy1PRkoDEjndgaBz+IzUEJJOxZH4y/h72UYLbxJV4zaoyUPb8t
FG4+KlYyeogfGcBKULBBDISlCJbxmp2OKoKXdKD0W7UI4JbUGwHcWrfca1oN3o0rHintIgrYceFz
irJ5OAYJDxIRXIBN3pzeBvMXXDfL2tMZ9afEegAWE9JHDeJfTNeTizAncNBecg1hsdHvEhVc5p1t
WZmDumDedh169kLzgJKdI3vYLoA03gaS+glVyc5GvB2cD3C+lS3WzN+wrTZY8brYOsHtoSVZCPIO
hC/8zXfGKbywPpRHE8JlGP6eKK8oz9m963HUyBdF++ztdH1DhWtpw9pY8PmL2KYOxGun42ArZZZ1
H13dppjj6QsHmkL+j4cEGsWilH1S6hmmd+oN/ELAmoruhuRAxKboTso4/O1REtOzqTavcUPB0vz3
jOpTfR9vviP/U95uLUSlFug/xsiULebzceEkHN6/z8w+KR2X/scEVTLcbEHOL+2jxAvQ9Zu+ekvE
5PeGweLkkwHLwLlz2yGfNmB3iWyYmFEIQKSeCoFtGMKGi6LbZItNBuxPlvRNR37x+RU+f1BDgo0K
IXgu5aB/1bsmBdo3hMcLB724rxICwZniShfpv783GyKBFiroTybC50k9MpgGNkdFRpSK0Ztb3nJQ
ydHjiVIlskDKThnMKliKD50TnlDdl0+ywvaGAGpncvPbKsX6XvMoDfayiPO6FvX5/bQUqE8eQBVb
cF/GIV+szokfL9vhDyPjsJRnfX9LNUIiH02BVhfk6Ud7Hq8IiR2fuFOFfR5dE5C4wXL6iRmTBoMq
uwb6GN1KsbVI90aC41tMSBS7zia1FtFh0xAWfIHZb5xUmX5UcnFLmSvcrh3qOo8+nnOyikg0gK0T
NT5xdxfs18wBO/AFSjrFk920v+O1SeWetiqeXP2OrQ7+ja9FHeqUYImTRRvQynNZAGoD32ZiHNcP
P9Y3gco702V6tScfP+8vik+kTHVD53wrwKIrbIAor4U2DopqhhV+X8WKaAqrVyw8piIAgrEcHSEa
77ESocu5L3s4WrcTnXtJ1clPl13rcPatZy3kiLZxzR+/7nrHriob/ac9KaKNG4zto7G6um/11NM1
yo81eIoFXsrz6ieI2NTrxRIziBE4cHjGvt+1xS5oLsmn676EhLszDHE+7bXdva4wuG2BGrmxL8OY
5pkwtMGaZAT6ZCmAnwM9Pbi3Pvhynbfg8odSKDPphGGI1e7mKYbhfvJGOg5sYk0+rtVJFIWVX7WG
cM1gqVf3RiU2fonPA4SryjfX6jhDY6WLtWwC81DolPAvF3Mdh27yKFPVukvdWNDAt8rUTnnMUn/B
JS2faWZ9BLP0caLFAC2hAOzvXUvyIZ7+T0uZcGYhzfH6ZdKWM65z+ZXWhwkAHBIEVSWZmSxGoqmv
VYdxX9qxNDtyhhwLAfckYOrZtOrtCiySnttmiu2wlEcEIk1V+ZG0tp5HV1278hG/uyf8+e69foiH
gjMI6uHOCPhxpDFL4BzXvQErkrAdfkX0yX8xUUZNdtFpCVjVXb9At7ZgbSGcoPOIvIlc1kbwb8/D
PKe2KmND6Hg9+6LbddnC0ACZZ8F8EuA+A3TLqC053KgzofASkAlUScUMEYu7ULfvQy4FVBYaoL6H
msXAC0oJRHonZgUzmx89BLcbNaCYnPL8i3K1VWEulT8mpt51I91FPC/5C5fGZLykf+7iuHLhsMT3
TRNL1i0Kx4GDqOqiWoLL8GzrTpfpsh375s4qDc4t5SJkolLMYPEpiTxij6AgbML2nq/ozHdp/auK
mGoMnsqeg5WIgAZ/sPxdrnmcFXdozucNaQDLdZ7NXZsvEzELC/u3x7YsR7KA+6/ax7G2xzaaMwkm
UaQamVJI6YeYH4rC3Wrn64OVhHVyL7V/O+Mr0b5c5PYnhRm/wQqlTAOEq8NuaIJP4ZCBPM8MQBmq
ssdi5Oi1HZdK1iaRZB6igVt096456QElqiyfcv6GqBzNS4+KR8oM9D+ZAURL4I0QBQBc0QFrvmWr
Wckw5bm1QiJmfFybs03qhNq0ypqQ6LaW7SPc8fpGZ0OXLBSHfxyManSxThqUVqoomFU6OjZF0pLm
oay2J5FkukjlC5Z9irGiVCvys1uSEBMkOGMSQOZE58JGDUGXLeng6eUB+QlNoeDSdJZWPSEWq8RN
zmYnyXW9DQuILitYep2mUcE4itDuDDXyt70NnmQIm5KYz7EGYcRCDClyzXpsiLUCbi69jpGzNChs
bJEqUtope6izBD0y/wUGK3b5la/jIoXQBj1oYaD2uQ5+yfM/bU3uGLLw4WgVRH+KP8Qz/wtRZCrw
Hunns1ZTkm8f55xHD6SFHVS4nrZvaY5yzCu1y1QMiKhwSFVr0leVcWnJq/rmOSuOHrerdtycKd1C
GV1yJxrVNzQpWMgYEjMcUhzdigYPH8Z3GS2CsZGyZc/9WeitWy8WdLue6WV6ZeUUgeSPT8HWjogi
7pZLXSh7MjsyUcTNFACOY+p6OJpibrCpuQlDCiFvNtdvadKwvnMoFatPg4dONpnH6L6ahUjMMiNq
rzHruR0s6lSnOOJX7dSoaDUvZus9HPaxNyOt81nlyWyNCo04rgiDJHTWEFS+koB2eoxGqasuIMvd
Rq1xnrsL7D4eSDeycrrYQN7K+XWsgKA8moZXSIV972ZgXomMJ/0GIBfabGnNcmZIK1/jbg9kV+oE
WolW+rxD63oPjKInW8WP2AJF1XnHSJs8hfqDJya2gVG39NmxzDVRAqZe6CE8oxwUpqGiPSnsSOby
8VLNeVPxsjR6GWgOnqUdhfD9oDCm77LNXZ4/WGhyS753+HA3C8lj4vU0i+Cc8QBZqtBvjKJxmEdy
WKKEZWW7X2sXQ9Ex07smcNk93phCJ+ykDTx8rlIKEtfrg9gQiAUYzf94MubFqvYit4fwtU6pEosA
SfFEhHR/FQErG5zduxPuAm/GxaLAUCJ/+e6J8aKgymmefQpo79BD0JhZxqSofoUBTz0/Gbxs+fsL
Ky1evqCw4GZogkcoAHfcjxjpWT/hb3qlgoN5UqJ4GRMZ4cBReIzztdouOUeFqso830dslemypVHf
i2HzdP6dhg6hAnOOo9opC9jL2+ivjlrerMfYCaCRCSgysow6jkhiT4LztmUbuRvm0IPWx/wOw9/Q
WH2hr8caGTpOKKvxZeXrC87EusuNVxJFT5BnI5Cu9b1Vynwr+xi1Vh8/YsCiJJHueNowOIvYc2nq
UCEO964yUxGPg+w9E/z6cm1aMZllZgEbZWS70muz8LQZs+w411F6Yze44ZKP66J+LUv6QTKqOKBQ
C0DeqvZkD3/c5ry1t7P0+G5UWGpiXXRi9xB4rGat1lNOU/jgrXPqApKg5Es0tL73KhNinqgR1PP0
vWXKW3+f2G8tclMO4SMEWanwLo6/ou+4YhG8QeixkBf9C+wPPVHVo+/xchdpn26BNegaTm93fx3k
LgXqxo7d6/vktujpReYoUglBP8pRvP+xm4nO3USeufm1xWrVLawk9opbvBlpMvH68+WO70994SH2
G0yY65vKCTNjn2TU2Yh+tEZzlaHu6W6i1Mcce5qTLDtf+q5wzLjN1dLUS0TofY7zB4u6Vhzez2bp
nXk6sQ8VFFxzOx4muLDBH9R7jpdKJQeJthXwOEr9Fgkc9o1y/iYloImmzLCpCzmHCSTjHeIjkxbQ
G8PVQKgRC8NgKS+z+knfIDIwx9XmdDB0Vvrwj2fU3PDOD4tIuuuLsRBzecb5+D3xHWOggg3tZKv6
yNQOxMwhV277ARckShZhOw1fn0/AEtbt0tghh2AP4Bn/tb536HT7hWAtD5KEB07arPFGPDI5Ptc+
0NFUxoc/ezcwahD5NsTDzmCjXRXFhcBRx60vMJe36F5i/oMrO1wNNlYJh8klaP6sOgnMZ0xdvcfp
DXiNNJgCS4YChMZ+PNvM2fdcQUPbFw6qXPALv1S8qCNteS6ds5XSs28gWQDv4um8sBXxR1nbai3B
PlkvGTXM7BpdMt9uAUeII0vio8FnXdMXoYh5eB5aLdslNyck+Sw4mzh5L/wHwVrBhkIriueBQ7a3
eH3CMiuwDTWpZhQXwANFCI7toQlMJBdve5YLWGet+0WuhvjrNMl2dofzctXyxxRVkQVoIegzNtlw
vR0hKMTjEoOYtxmROSEZ2OIngs+wyVcs+9+B+FSdAhixeAnsJGgFlCICWr5F35jUVc03npYsWjOh
kP6WlZ8r3AaBh4LCvdUglKKvIzyyrRob4YJrKMO9zDI01AlIyvC80IRf5m92LGcMB8yw27RF8W4Y
NxiyeKmWSXt4CjndXQ8IwUf2OvrnW96MdPE7rLzrpeP1l7uHOxk2L/Qua/uWVx53pr21lPM7b0yq
Sre4LLlyAZOc4Ryx7+ExAXWiFQzNmO5Feo/LoyxxF9BEDE5iUsJjCSn6oXX/S0p0ZrfI7Bh7Efse
8LNkX7UcPp438Q1q5R1uuIr1u9y6+5uli0IIlAxCsLyOMIvdvEhYpCv0vUDvLFYqO8ArSipItjHV
/k6ZC/p5a/RuIbeJRulQc9Z+lL5ww10lXlwjs550jV85XfHGzVr/F2i/81sMUqXp6bwp2pT8awmV
JWlrl9ZNTB0ibk2cDxa9adm/k8N72ZyZ9Ii2bv0iTArwqLIKA0/i+0aXX9x3mcSSFo34r4dkYWYQ
Va+1GgELtqATidABzUf43prMsGwZSCuB+LTQZPEqgw1RNFIoNE+/2LARzSAiIoN2K3aNTTrOmzGI
gcsVMigK4mL0MOmbmYkOavbMzndcIFo5bSFNoI4rnrvtdnu1awko+oq/WKtvg/0rWa+uyt6l7TX4
qvkIufUaAf0JqIsRLyuXue0DzdlwhR2mh7krK/fSxlTowzAjGfBn7NabtZ5JHTtClUy8HZeAFMTv
f3QEph4cwtUd81Y5dRRFPKzJL9MT+oTSbFAIYCn/HpFvebZJDz2ctJXjQsELsFTHAk2nTT9W6Ufo
Bfm8i73K9dAC2womQorraxr3TvFXxz0TNAJI0iiBCHbxi3BbmrMITnTBNjMjLcEjnWcaBsZSJYnQ
fgroTOZU7190GHsL6anYVYr79Mm6Vmz4Ne6E3xWIY3eunBimlSF87GaULoDwWE2mlsfIeJ9+2RDy
/IjnXcKsmgWF9VzLqk3NdYOUJb5rv5twgDjK8qI06cPKxxkW4jTKNGLKPo3YPEVx8rRdARyGfm/o
SBbB6BGiDAvO/kOebH4LytFanZHzc/2bEJkQHVeXrAC6S1qsRglo2gWP/0T5PfHqKuEGub/q/RBq
E6mcapPxkaESLnTlhTB9youk8/zE0V9308HH/wwlmDQ1JuQtpgAjSc+jZChS1snmrF5/kro2YWO6
msq6XxMrZnqIoYRQ13XlLnQs8zCsnfeyP3jDoZ1y0SsxT/X/RiMmEJ/UyIRaV3/2g70gQ3ZXw3TJ
oEhbP7Z3qeAa6ABSCi46cmRENEqON0LT+SsdCoc2pJASzHNwMC5sgztgVltTqClh7+rdZT5D1CKQ
qtmKAwLe0c3fFQCz2TbpoY+u7Hm3kt+vIGC32RpzWI0e0ZqYFVVximoyz/QjArhbg+R+FIpcpmHt
HIAyjnyVs5yTDDtJ+zAoEbf1IfbuqEeo9bxTyotbi7q7LxPhT8moKr/2fVzzPP9lmi0gBEp7HsU5
aGbWNsm0bbwq7d/5x6/wvEex6uGnPL6FVALVWczpikHVfv7El/PsgCq1GmNlXsIFUHtW6ilfb0C0
iqkt3ac4fXzhk734o0/1bagPZlD0N/wGtkDmthkXHVxguPFly0D3aKQsiYU3EihhihF9faZ+BeGP
mXa0/mAd4IX0UBQWmLZE1FXO5rOoL1JNrfqcOZJdsukfV6kFQnGCzGM+Kp+uemkJuI+PSznxK8x1
DL7ZZuZrWoFTrBYRsPrOLX00c+qo+hW9xVdonE1msm9N7bLt3Uks8ZuMwNKtEchSRyebprTwhEnp
sOoZeWOhrnjEeKiOboPGckEfT4A5MrgyBAl9S1YQS/QzMib3fEgfUvhsU9/YvVvNlE1Vu3FZQ4MN
9D+U/LBtiG1KVPZ79QAjo1VHvj2Vnn7kH8k/hlB0LbcHozzYZ4wNfIKWoqzbJylnEjPqGy6Hz5FY
vuSCgbwPVrCe7kXJaMDOeulQJZ4vrUHSmIiH2CCWH9HDhGWRqT4rzkr/hXaFS9nhEvsV6VphldRb
PVbkEeyLRGxiCLdu2lg8ofNtxOVQod2IlCTMkDChHmQQaIMUiNKPYg/DdBStflr04DNU2QUlVbXy
yZAxku2iRkEVrjVdFYugXQ5QRqMdJ7AgKM9hN3RY+Q5l9fF7DyQiLdmNpeM6iAnzLnk6y1uKq72L
W28bRtQJMSPyj97egbgLAWjk6HldYLgobDzAZQdadXtKcsu0N4D2ZgxDLlLTxn1QDySvYsiSn1hu
dHHN7jvkcoV9X+8b484a6jETZcpPu3+brDaCD9NHl++Ry70zLTEkEvbAjoEfc0Ow/tuleC4SI+iN
jHUwkccg41u2trTuP1PRoUDc0Z2DOMSMv5DKk96Gqsx8wyK7+gkJJxRpHMhLOA73jWhJdSm9FKuS
a7qLaV2VsDI5UoWd+bv5uilBZFOc/kpLJ6X6BuR9wnMYV9+8IsR679mbV8YsmFYiFD8UCJLH9DwC
M/92Cdki8GQ5bnZHt0xwIK77PVRbNj3l++DrmO/QVBkQ75hq5eXPuO4kU1QoZXtf7I1yqUH42KKo
8nsgCzUBMLPzz7VhB/X9ZrDgjlp/UlVZTERfGrmpKWLTStHNdMDe/CKweCCmSPyCbo+MSxH4BtnQ
h2WX+2tnlUeGcTKLHK/dDq/M2dc2N6gpl1yXajBAs4/kJu74sRQ1ZK8T2JEbEuUcUNHMtrHM8F+Y
KhD9FpRmqtk9KUQMoB3yH1coLqp9WqbwqJzVAVMWQ+mNNJR6AU9DrlFuh+qpjpALqKoxTpkbRM72
JUpHQNwoRvSNVAi/udQcR/AVd3LYkebvbfEgtkQGQmoAXoeCHyyRa2Pchumdda52PIFQl10Kyocg
ByKrkr1VyamBP3pcoYgSd6ZZUmDR1cY8qy+2zhPG8o0d9LViYInegiFjK/Texk1j4339eKZFS1xv
7RuDBRViI9/exgzLrhtEmfuQff7AAPsZis6pFHzQzBLVKpKX3Kk0Pm8APedez+Y9HlrKiHkkqjWQ
N6IGN0TmLJHdT3QeKxV+t9RnDTLgkoIBXMXwA4Qlq6oBgTE34hCquU3SJ+L3K1Ps4RENATo5X0kp
Yl2WanBlFN6ci/LK74bZjmqGztQkV0jRu/4Pw0PkUtBAHdDLWwLFQdXDg5Q53QfsIEZbGrr0vYzI
hl8QVtFuK2TThq3uDxz1Ub/0nyjGS8WC/dXwupGU0CldhiVxKA6e3YH3amDv5dwycY8OG8nGIxPB
OYT9/1Wl4U3QUKZ/71u0P8bdEP2dWDKiM+cQE2bJ/+XGQEiUCJm6b0BHb7l6d6XO21dhbHWZIxIt
EvggpUla++jQXENKQ20cKUCnP9qeq25f0cSlvPZf2g9bPmuYgqGu8chjNESRIBgESj4YLk7Ft2Bh
MfZx8L3fNTWkPIBgJ9UWECLExp6dT3Z/iCU+L4/WHY8IWBjGXMWyPaYzX5SEcH1bmtlHn7ku7sKM
h7d1rT7cT4G6MLDyJafoq4oBZFWKSVoGd3X252g70b82I2eKwrfoGduLtuwYcjnpiBpmOFkUQ/YF
8SuSMVxHckNPhb9XEXfJ9ao32NHzFz/TGfKfQ35Q/213IuRB8EKF6tWtQzzrLgr5+GN7t9c6X/oO
yog/4HCmwygYusgrWXJt1LmGDUZGC2psgP3gm5IkNNf+N8E2KNCVEatoYy8jUHVP/Zr7gJmRbMoU
MhUijRP1BDBbEdfv4yulT9nXnRhIw8uCTN1N7guKr6kEzSCZ8z/kndT2sxvfpDx2WPIo033JbEM9
efgUw7yN5kzna+n6Ox5sBXxPsd9WWJOskgs/Jw7tFAHmgqp8zlUbxO5he4XrdmEAz+/gNIcv9hx7
oUY3bHA/xsGwR36Cc+kNFJD1HbuqMl6qwLbX6wrB1OVlhacF1hxJRGjYnMK49dplfxu5eS/7BAAM
Ngu23A6bunwIEiLmwvB+hAxmEeotzOYVoSPDxFc95Dn6b8mfir8pkIlYER9qzbn1c+ZdqAmk9oli
8L1/D/2aBcufTplLdOYv8G1w+Wts3ZlAptrfT9nvRY2vnTnXykC5NM8iRclfnGwY0pEC/uZLkoea
+A/WLB8N/lL9epTki07dMpGZF99k35FiIZwRcsVazUwZhpXCW1pAfd9zjqbPCZO+fgJgz8T7kl3w
H0vYkSsYRyfcbAOnvhdg4t5TweASfdksU7TIKBuRlWDwLDquzo6R8nzgE3uVUAKYtDaVXtHJWlA+
ARTc7pJArAY0ArOoC5IVEyV+RkfR6rBN9Fmr7hAhTAFjFqVgM9QbJKuhkBgka1gtUKnO7RWRN2Ft
CWNsO51Ha4rdYhtmwKP0N2hezSe7ourTieV+3ME/v2pQY8SQ5hjGbU67m8gFixKHCNDcBR8dRh5u
uLyizqOkcUg3o1dhSIzV5g1bWYUB4JxTAyVOgk0i8x9M7Olg9zgDSD9i0TmAXMGg/3EqkgGMQEhn
vNHMEyQpT5BEBtKF+00NY/6jXLtErUwB6paNYZJARZR8t7F+tG2ydGgOw3nRbiEXwje4gmTrl7CK
a24BwSwszl6MrG/vnNz9cdhUgUx8C7c5U+3Ssi4+1pSDpnPXzvvzFvkcNPmS318HWYJGJDrBemwe
mAzD65Dy5MUbCY6yiCgphdFHCyF+PMEiXt6yLMgCzrNKB2IrWwabj4JNa/1UgszO7koTt5FYF+6E
FiQzpL0YZLdQI0O5z0xms08MvB28pOmERQ0dxqrkRD0bL9xHMk0nNhlnVhxSVlCHSbknWMQwngeJ
Qz2Grq7OfA0lC2d+RQgv5MoTAOy8SUwzwbdyWsd9ilPJweLo62JmnknfvI37NXZx9CEYyHX3J+Jx
y3QYzakP4uFncNHwOhibIunLJ2O1kff14LqyiOE3gyM7xV85UPTlfh9dZxb3m+YxNdt+C6Db3IDT
7Gvvq0GjQVRc37H1o/Wq22bSR5fpAnFVxz0i1U1B4b8Ig8PqApDtLCp81jmYclveLjqDogA/aQ+m
YQX1ir3T7BzentZajtPAD6gQPW/dg3KgtyryGcFy9+otXd7PRjDY+pK8Iv+CC6wOWhEE6ADalj8G
ibaaCrcsHnWGom+3AIX177lu71pStVsCywXGN2MPmDl/RXmQWvmmIeM9jfEuFsx5DTk19o5TCdPC
mbgnJ3rcP00HPhIyTNd+g3L4iqyLWI3t5wjH1x89AGdErEomLfpun/HaRbojIDjP2t1JXtfFibO8
Bn9A2OIgcHCfY9hnNKXpr5Roqj8NU8FDp7A/miijssw/kvdg2R+xKv/wkavCTrYbca1TfmPxHoJ3
loUZ+GrFKkBjrtZZ9TapfucYS5NWXSE08vyxRVHpORBWmbFcnYBBnHh9PzWM/czDylV8Nvx4FQuN
bykgfjXKESq8nkrgAnBXdrfaJOMc+2jum8yPslDGfhMqOYPIcWt9DKmJ0vsb8RFlFLfrl8yXP9pH
nJb6JvyIpTXXxBpRfn6dU0fUqLn+ygkn/Pk7j/kBOpH+hfscFOvRZ7q958Hja21I8FMtHZmiloWF
+fOExBkzIXGb9pa2LDcUvTJJNzX+tyh/adlbeLBoOOUwcSieC95feh/SecXpE0a2dHU6hI+O3eOX
y/9VUesWK4OH0U1CkGeYBSBJW17YPqknWRLkr/GQFmCcKv5Emu3UI1yeOXmBJhVzEDddyvEwCOda
Z+Dq2QniST1+OXuEv4ds7rwdplfgN9GP+Gt1tN4C4TR2YWDQhmaWFdqPxcQmdKEFkXGGnAIGiCdw
xeNsIH+NCmDO4aJ8qbLc+btAqywuGxeauAwY6dyLrp9PYazdYsFJdv5PZf7ifcW8p2Vzci7vGDjd
cmLTPOVQHhFjE7zlpjl5hR84rIGiHbPkkwWPjvGrNnF0dVHisQF5DAZHzCHzvYOrUH9X2mfEs8ZS
8JLJRY3kR59WUa76qqASBOmmDb8dTK7R9NskcoQJeH1UxvlGr6C7xy1c1T0ck0iWVFQmMJpTEX5Z
JQiVaZeLnubCyV7P9DLNbky4pt5VHs4aZg74ApQ55vSLvJEB+nazQ1qMwmATIby3LbvOxYCknu4/
sep648NZ8wcjL5v/YQTbG4q+RZg/A6JdyU/OzZZcqX3q9qiaj87NFGjYet6sYeOv7iX+mePj6/96
yuRYmuLksZ2qG8jMR02/aXLOe4a6toKoKFh3xIchMxkJmWz58fYTgatBVX6MqGkJrZmi7ia450lW
iijQgTGZxpVVmQ0sJMlaLYLFFn/gmZjHSEdnkClDmoSnGjUkNuq0hoWKEXwx4xcTwYSfdpSsT5VS
AYvOcrK8LUVBuM5lY+53JsVhAXfgr7E9evO5oM6O1MEzBajg5xyg9gygYYfkz3KgDNVO1UZh2i0V
7Bc9B3BYCgsfiwiMhyBTI4ooo3qvSfrAwzkXEOPTr1Kc1zEvpbYpFoQkvX/UaLYo5K+99+NeA03e
yFVvUlJzkK/p9JOrnVPm6mPBzN++ikTHMqWzcbwum23OnTF0j+QzItYHzLMR2XrGWRZegQOH055K
jLgIsd8hTQEUJ1Fbr3r80J7hP8oFr/3+aDh9PXs5albvbj8wZBtJaKyZtreswyMUjEryhW2Gom5k
gheiKFRtP6eP2TZ8oGw1nmCPXOkZKxFjA5uYTktP/n2HeWBH1f6/Vsmm+tzoid4sJz60b0CJoKYa
+DuouTczWjBpoIhzSA1RICbcVHZw8ichix0OcDEp53uqeiFYvMF3LidW6xqijQCTIPioQppZEjor
1wTHyMERvSNPfPLV/dw1BhkpkSDpzODH3wWywY0/2GMlDDZWfFMm2TsTal6HK3t3xqsa9CGewVnZ
tE41NKvwkb3290osGw/It/EDzeK0X7E9phdWS+8zledNMANQsbuNrQApnOhDVMXs+NLZZsjrSPEj
+7MS9c0lQiLvWB4yzAeaH4RyxYfTdO0ZIFl+tCf5RN1AUVYWnD2j3rc0HKbQdraQkmpvZo5DfLvj
9sRWwWLMZ2WpeJ2b7GhoNtrLhKy8FZ4v3EX0m8GbxzCGGN4T3uJ3mZo1wCsoDxY45FWWxbouI3He
Sd9GD8HsPtyELEu4fSO8WN3m6rgYh+L+ZnFUJOqBEba8/n9RiXzZRGYnb2VdyWHFTECRc5sezoUY
heJgnpPDnoCvcXQf8qBqOi28lS7fBN0OBsMQrTiuVWmyQSreJE/78gR1jlUR3hCNmeof3RyvLt9E
+bbHQlIBVK1eU/UI3SNoR2qcc+GKgxrWNI20mUhdWv5wIW8t596W2+PrGJU0oxDNpFsSOkCRRVVB
Mk78fGHCCNy0elSrmFkSAbPAFRZvVkoxo2J70ujw6zn5TVLkm60tnhZpcmbYnaOgBz2jttlQ+7xm
bc65Wofhbe8gEfjncWNGGHIzSBsTXhVhURFUQPxWCCMCgQIp4CpOHh/1IZi5GAp6zMP96ZxtreJw
R7Fe71cPC01hy+jBas0Iq6Auwg8KQs6/5uj1QcSx1m63A+Z3//oDzIRojtt7MK0GF+wleAtQyYtM
XZoiZdQypMgmaUyctzAWR0G0ggOa2GFrA32soLt2MYGLMq/JumkDw/QQ0F6dqJSOrZyqm4Mk5K5q
/8mB5CBbrNdEePm/rwx/mMKiL6ylSW/pAAzJqhGDnUVvJcdRaHzzMG0bCFPqaHORWup+vtjWKAgU
JEp69U25Vj2XHgK0eyOeFtgcxziUK4T6Secf0VfFJGnUV7aDdCOPzs+hBisTumNRRfg8G5zEr5C1
g8G3YwIGEQiVzzN0Uv0FaFs28z36/xlA8IZrPp8miTWCYt3HZkFNQH9ejKcBsJur8UHqoiLX2khQ
GpACxI1QnSRxzlEHqoiBEmRoKggrOzwKEzFK4CvRJKl6PkRgKq0wMpYGgcka2lFbuP9WSrlvSlhd
bFuY4raHxSZNpMgxiF1gDg9HZd1EUT18ETF9Ph6LwnCSXGeADxfeaJSh7sTBZEXdDznMYEVCFNs1
Tmnocy8v/Mng5cT3eqMM1zSNQdYg5pP82hZdc4rxgKc6oJoC0x1Cet7vKmq68i0Y6OGTNJpTsCyk
yQxjEYgjn+I5+s9S7zL7I5GWUqTO+99NAZ3x2RiKA1z8XGCmZv5nj9NNmbfhARHSXSjq+KlgeyHa
Tisc72axdwS/gH6MHdHyTHWQdbFuViotvDa+ZbAHai1EOvOBKudJh4m7cSN2Yr5WilzkUgStxPV7
4YjrbTaDOHlr0Jc2AecCRwf7BENXeGqlLEhgE2F4BnKZBiDwhkuQNVi6IioJYU92ef/NNvFOJJTU
Ekg8jt8nRqZeK4IH9VsYHFGnUxNxsgIPwPQIB1pEYEdHwBsUAVgjibBcqbVRConVs6qtyj7Hn61c
APQcIDziNMq3ZxYkjpTalBsdMTE7VK68CPZObsgAj7HbtbnKmQxVkSU5AcmB7ctUEdrOo355lTvg
grhQXixIt35Sv0z7ZUD4jvwqxGG/W1547CVEEXPR4z+ikB/Ud2OWUbUCtopVdo4sgGf1IT5+pUc5
Kqs1WJ5dBdxzQwSDU9vW99Ecj5pPhHk1SX3tauE8UEu2UabXtoQsDWe0ZRW/VkpO+w7CSedqUnXJ
n2yb/HjgI8khtVC7LTYJ3JMAzf/rq+YPPYPtRvbojEP7VQOI1v9IUhkQgO3ThNqXUjIeruHfbahR
KXhBoKYI56OkBpPMemUOwGTWcXtufWGHPJCQb41MaHqcZ09X3ZfqV1Wk9u1LWKERuwY5G9pAsNYg
jQMwYll3ztN77IvToX5K47O0I+i464pKGwjAK3qg5wVWgl16IAKb5OwpwuVxiSns/VbGwrGkSOUb
NW11fmWoALbvA/G3r+AknellqXuXggoabbZxoxYUxbZkjd39TuNX+zf4d8/cP6SfXD915r3G3ByM
UGBxTyZhq5+FjbmK/M92HU7UNkYbbJbjbolgvOg+g23YtFVhsdDNOLxsMQUTRlX9eKuVvdjuZOlS
NzWOb0xI0AXFsRCwNgOzfrWRjs2NC1XEs7XXNxZMuKqEQGRBuvFUJf4iwPuSLhwzAZl6bt1gq5SQ
NtkI9W4mLlRxpc8tdDtu8dImPgr7r06biNiMkkqh1yZJ2Z3dXNBs6HYR4DSypjeZlezUPw48gQxi
/gtwyWn46w3j+pDLgXjZPNOoC7IyvnCuP7TqPhFRPO4e9Wc0oGJ52KvmQVZQH8cD+E6Vo8u6ln+J
5dULc0zNQn9M9qHUyTveD2Kr+orlPbqQQk38civikuy645FELNBiLyLfzj6Q4OpbwbWSSnknwxEt
ANpl0+Hv+bdOM5yPFrN5Lc0gOcrnEb5ZPc5rj8jpLsGxYSSA7JnfVWjkd6BWH2ADwT/jMb4Q3PEL
JXTSekQwiuuw5pwqPHQPkLBhmSidRdDo+s5kRihFWlncOi3RMmQqcJJGytvT0mDfmvEToE7dpwHI
OyQzTTvTSDv77vH0T5IYW9L0GBFm4YfyDMYpAMIslFGdYP69NaGqqaOWedFX85FybXbZqTwGAGUR
tOubXLyTiHU5UgBUMIje5DZQ8Lc7/hCGUmrTwfnQzHHsDA8XxsHNtIZGANCzIz0tPsFOouTHf6pY
hrIB7n3KlVEexONlE1vmxIzNoukmip0ybE04baQSwRZ8g/Ueygn/b2OBjLYKZ2vYem1rMEG0ThzH
bfEBzDgvxkdJE+zxmaNZVFTz8i8KyqpSOi3g5h5fMnpRRlKlDRYyGKC/tMyRIGFK+CyKbwDEpLLz
X8jW2ADqyErC+io9xbBiE3kZKV5mgTrnQjFMd7yVLcaDZM8czf97TEFU1r6IDiTtHAc0oW5Ge3Lm
jW+Qj+nr56L7LQLF0qS173AazByQAc6V/OhQkdeR1qJXaTYRafy5H86bYPx3dLY1kI+VX/Z6GHsO
GVP5mkPrpveVUYn3XcaQpQ6bNC4ht/xs1vKkDvU6vxpvkYEPGJMM9B/3w4o5Fvg/foTe4feS620w
Jn/z9DswlUTxGZ7bIOJ93PA/x9CuRgXQxERLQJVGyfmvI3OtAzbnaQnZxKWSmm9YvK2azTf92dKO
ivzygs83vGmVdKcDBFukEus4GvuXkxeVF+xkWRsE6J6wN5/vnT//CdHOc9UxD6If78j/oosplBuy
4CvrF+hclCbVZy29ZoIvUo+GVGDMQ9/05UDNyT9iZDzH343fNJd1iVpejYa5UWy7qCgfWQhq6mSp
vPlBhqgw9RxJDTFqZo/pxX4xZFXH1YVQl2DljGXdtfYnzsKCFzIpEbM4l8WzMApLMoLic/GoHPab
0apuZZZQ8yP/0eT0biaxXeCq5PVfpV0I8X9XLzxR2XnE3XjLp0eQD95XoUfNUcOOK+w/B0uz9KUo
SU+t+hTWCg5tWDs6wkC+6CKGtOdaZj6Ng+ojjLUd81pdnLhYcAXbq+rcNQhfAsIVmelRlZZkkPNR
ar+LVnuIT4lW8QT7iiWCG8VmxBCyJ4JEebz2DysG+QolA7A0dqisOp/H/6nle92ShXWDDrCxzDg5
rGngemu2fDUk4t9qJSKfTmxPOya7fURyh73PXyejxUgQIqRqMNUaCxBRlkKDeCDKe35k9owrrQxA
REi9fFiTNEVyKGVhJP26NWbC+zoFaai33hyXsz+JIcbwc8lFDEV6TBg9XBZhsKfHqKz2jN6c1lsb
KXl34/N/dUdN85Rs/mzVk2Bc4xykJNnIbUi7a2mPJMAZ52pRUHNrZ82MHPJ2ObwhvsQXxINQ3Jql
gzCtPfvMPKKPvBfxKVa9SLPvhq42Nbefne5Rc2i+ZtzdobnEyjU8fWmC0Wjly8N1xxvJaXNp8QRc
mEbR35H6bSGwyeKajKlE8Yn/0N4f2Rl+J92NaD4Edrdu7PhG2jYDCI9SBdtIIkmOuWPSuwNcoms8
q7c3g/vMVeRWUPOE0qFUFHqCk0mq1lcx6JHLK7Hx5XFirn6BiKavp7bhO3XdhE/ACzNIApO3CUqu
d6Jg3Vm3vERlmToMgWAMss2AQXsH5U66KnH/8K2Wx0NdWtdZOpWEAuhuJqYo69jJ1H5JlErKV20m
3uqi1dQ/uqs+Ic1O9jAwGrF9GqQNu5iaX3UubkXgsMONFUks5ZAwJT5cyNNZ7YD8kGp/4aosDotq
1x+0iQW0P6vb49ksm2N7NpdwvSCAxR5tfOKzWopK5q3XZU91JWXENIa/q8OD+WXovKWbLDYedEjs
Z2JimVozcVckSvXrRp6v1uk4bW33DLvq7xplM2mwy7YBFtEEQvkmraYPwAvUCvJjSDon4+6e3U/C
OclAs1c1XjEcY0j0YWEmtxejfKmTJD0QOqbhFfW9z3GJZ+/4R+Lus0imgf6J+9tcApOxjTIsEOUe
IJZqPn1kNxbVWQ6IwoZTiIxjl5jBuQtrJQkD6GUClQQZ3xlzxWf1Wt8I/hKqydytGfNOkL1zrXy5
x7uo3oPgiuLINzMsGwu/mmnu238K36L8N14cnKPp0fM6iN2i7DWmQnIt4++MSSn/oDMlpRyHantu
nXFhHDpR0d7aZGtapvfT+KWSccaxY0AjCzORZbIwpCwvFmIvo1/2DKrtp8tzbf8bW7Fq5q5tDzVi
PyPM+DTKQ60v+X3zSa1gxjdGdq1fNQfwOh1Olp4ssMCULvvwsw04gJqJEGAwexnZsBTHVkFBp0e2
TEEW/pI1/1i9IjaBIIN9AnCoqT8UQlrrSQghl5nko6pp2dQ+y3eQhy3nmAn+X2ZEoXuj4QMO+VxU
am/AS5gDO1t5xReYd3QT7A2nxgqH+wW6Swum+3VM127+FcZJpDhV9mQs/TuN1bfZf15D13lRGWSU
iKRLW0WIwNm+WVf02JTzjHtClKy2AhRmtQ6IretysfeGZ+WLrXRbXYBgiBgBSIc0A8PqO2E5TTIH
E/mj9Jfb8CQZZyPlEnJfQnwuvh/E/SS0nHkOQ7dSXkFI21ixAGLx0izJ55Zjhul7rFuVPKuYKo5o
jHO0X7/YrFZWlzEwfe9qdKXX3p6fgSGc1tE+Nr7QQQqEF07pJBB1fCEaNWQidoJZYI7k9fhuUS5c
3CtbpXj+VkZ6Pbe5KP1GRqfj+mIBaShWmnxgI/ipBdP/CkWklGClhSH5s+CcYCxAtU1CHwwu6K4K
Q8RzEXvJsOQiALH6WvlupoFSxV25ZEX3kcC4lKh5mheemzldwgapRe7r9WatYhq9yGnxg9BTXUV4
FSU4epZ8gGqxcVNY2yXwNBVil/ayfUFr9o7hxGqbQHa1gbdCOzDE4TacIzhepujtYXMuuzkhLWjM
0D8Rl9EqZpdeQ8kCKpHj7NW22RRgjo4Unediv8zFJ4lw59eM8X9qCHSwmvj03M88GM31BBFs3JXF
k4cafnuL2tOSQbzmD5Jd7XMtC3zt31lCrCRG3VjY+qXJkPhnrJb+Z46aYJX/ghsoJj0zrYjP8qxY
85JfZYb3NXwyKYJVLwX7ijx0wq4VgDcZqLDoPqhPVoEg5ynDs7VFuHyqygVTr4jey8bh3lnUsqDN
5+34P19DfPZ2L2HL3qJc9DPKSpeVWY9ddEixbxVy4OvjRdeacZYa4lLU6+XVA67jAbfBXkExktqb
e5W4kTMHgKFHGZijhJDYleqs6ZX1GZAXq7KylQ2RqKECQazVLpj9usOlqxldMk1sjx5/UjzbBwxS
avV1ooK+JifaL5cRfxbqvZXuiOCWDwC3hVxqJyKk0pRUzJEcxAsKNd5/E63XEv+RDLu3DJ0/3Jmx
8ybFYKHnTXmiRTpmgHdAzJ+BOI2dn+GtKNkpaLacmJKqF2bJDCfBU+s8CJN9LA/0ONOyBlhoBIiK
A9+JcEzPIiSkXZwOWHDk/SoA9frLH4Vvp1ornjMtehiFSCQcS+7XC8B2vFx4yrggihBaKVVNSRHo
mKq8oZrnutZAWMx3OO0Gb/nojptTO3sG/eHsGku+yl3RKWXYYLWujMZKyAm5YTrkpsO5Z+uCCqQE
LbWHntm1ZF/fYTwPoL+Mh64rU7TkgvJvojxnj05uDylGD6zi7AWinl49fpv4yiSUq5GwiGrPPkIJ
iz8yO0bH3e6cJuORbdaiR/XD3P6TDfOrvPMgGlXc2qg+DheuW6ePVUOUIYQadtbt7sY+ktDZjJaP
Ttohnl1sgfOHMb27lz3J0GHeJurMArSjVRTSqlZYjZCP6K18D01RPRcUvTac5Yl807t82huFqr8b
0jpK4ZeVEdDQf1RLWux+mz2sOC7XQECcUvHkBYHvg+8tRVn7lMTz3J77bVAvc5GerEg4fYb+ql2P
9ZgyJiycQXPQF28zOeWT7hyLrGMJgvppbjiH2ZSEwn8ZSMECjLTRj7C+pZyU54y0CMmtUkiFosIZ
+MnrsrPrt/KvvxHgv8M/LhxnCRdz0WVNSzwKhqgQHlQBy99uFM2Zgd5J85pHYy8MFgw5xyBPTPNS
M3o/v42WpmbAf+fEIPBfv4tGzLsy7VnYReT/xz5yZ7VmQ3HXHlq8sP5blGG69NaMMu0oT1GTWYO4
MNAJjW/KW60fDdN2dA2P0TIIhoGkNbWhEnBvf6rKsyEru97/GaYcjPBW2nR+iJqga3zfrpIeYUuO
yiYlQ4WvNs1FbzQVP7inpcHSimeric6EcR6QvrlqRqFipDxAh8pGtH+sZffOdgSZdIRI2uLpuZHS
afkZ3ua1jCb8zDWjsiNk+WpxTY0+eNzXbMWG6dpBw4cwddxzhOwh+rK8+J1RyyJ3ztspPEZD2ZyB
PyAcUuRDz/RgBB/HculHcUq9vOfna72TItZL2CCqubeWpJTnLN92jPUEkaVtMfJmkOl13dkqw/fS
acaihgQyP60UXtax2SytMBIJ+zdHahlwwsf4ZbkOtWPNYvA+knifOTxBnsqY19ZH3AjQrqK1mw6w
THk8uHw3EFbZejl3hjM0ZCUjqg72xavnGgVoHv93k0DTM3LlEm3d6TGG+ZP4PKg0xNtfJN+nRra8
qIsYBW5S2PId8Duw32iW5FXL8yPkCkZohxG0SJ7rTjjbzPXry/s+UXtBAaFsNCUE4+pSZ6/jOA/e
zPsPNIpLrTiNK1kpqIPRtoeEx7S/lmzdbmwlG5jGfuTyBMamm9JltIGoIIMVeirVfpo6QRQBBZSj
Et+uUcjLw4YMzIZyduwBVKE1xUjWZUwLTpPw4V8QLBtLPYKlV6HOjO5+EI+mx/+q+nz5uVPcnwTN
uFUdBu/O+0dQTdKHIjS7qLXFXzgeEvV7prGP2v0Jk1Zs/APmwUU/GiVpSS2uSHyM7NSO7124EjPM
iDy2rIhEnfJcgV3hK8xZeDfQ+8DJ/u1MvpaNJdT1pzqM7qk0w0gi+e+6Ogtbu4Wb3DRmpJKPBNEX
9KuD6EFPL0SOUQEXxWNoCxbJKkElMAcFvyTX/iLXm/V3gBO7EQ+GP5jEMkfq3EivqS5DKtY/dWPR
pzgJGjp42/3biGg3f/PwhjzMVTEiiqE1ijWmunF8QY9BFMXCFZLIAQz4kgAu0OURAJfIfog4xg8a
8anTlFxh8rJ5Z4Xz83UUnpCiuwmiGjokzp7nQSEy/mBJSLRMOnFRhElfFzSkdlnWex9rsk7Mvp2A
FSAkakjXVXpNaDga3hnvqsNdJdX27L06cfaTRUA2ghPvjrlNFxlJ0X5BI5tjeWP53Cx4tmsouF/9
EnhwVfCFaeTzO4amj9AYJcBnkM0NkfdCEUgKPHOGOn9Z7RN6Jrb7ZYFmzVt+U47VmQ6xxjGJZpc3
Bw1d/4R04Lpu5b3RvT3PsvPqTDYTmUa/O2Sl+qa0XDqAFqFIG+Is5Lg5JbG4EWM2R30Cci6t7J/v
QdxTHNfIa/j5qG387uuS5WAnHOcx8+Gb0VZ3IpBhR/yGGlnZ/Vg7/iSWrTIFuHj0j2HAJyvZ7Bw8
qwrXV2QCA9bsfzPnFJX0Ic8CqsWV9MdVur9P7VBjmEsEBjI23u09zdrkghAi1D80cH5CE7o7H4Gb
M6VI8GgA7Xmw/OTQ41FG6knvEdGCbF85hX1Y2RXceRzHdT2nd8TL7PdXjLlMCd2+lHvO89UCdhNo
xYKkJViR8mj1HMYKKrcq5SIudVpGGU4xNE4cE0nPKyBqcm1XsC/6ECSsSPDONqeRcbGIT6yVhVVx
Ie7uW0csVans7KHGKGf9zJeYsHxZeFxct9RdRMMFfjZwatJOad53MJkg3U86TxDlRYiIsuGoEePY
MtqLvlsTkxQj0CSYXR43NOmof3ioUWkedQWDOc8av0BTYlbbbHCRpfOnm++NMpJKubGyYSfUaxvm
drAi1cM9eWXOnXOnkJ8tuHf61nzPZ8LFy7UJ+iC0v4NM8x/euQRuG4+bYBWYgwPApI6cfqfLyaum
UHZurDVJQWrqenMRc+xVywmIA8Jj/meMjquNWH4YyLA0k+UGTvUlwIX6SQlPeqD8IGmu/7qaRmZV
v3DcIZX7Bd1CN4dr7POTrwzES62X1LEMNM5fUfQGktvKg4bnFD3dlbVH1nTmN6hCItGFl+czhJIZ
EQqjH3eoqUTt63dpCETzAYKBaNEHU7VIjZBac3tj55WReR2QyfBctRB05DS9h4qFvDX7z7abIp8P
Hv7Or3vYeRdqoMdGb1yBEwlJ0AFRheFF4Bqjyu6rMmekeLR3N76IKWTLq39KzxYxPqoUdPq1B8LK
IvrUm5feHM7pFy3pTp1jg7zvCyzvhH3fDPDYkiQKSc74X8ybnHsUjpaGbdaB4reLckW/WUx0aHzK
1ZOK0bUAF2YP4KklrIsRzCb53jZX9gdF8geQx2MdJojbLWXzbrcDap3xPRac/5XkE3CVB/fa5WTr
xyqV0Jkq7ukFvxZ7sTvfE9XCtzg589HODvw9rl30s75qPcIDL1DR5QoNfUWDuoheYofV7oXijjow
jyuA9EIKOoqF6+GCE05aDM7RJzbg1v1FjWpOKL6YgfxEkdf69cYa4rxbaTOznh17xRK6QS0qczS2
dy2AzV31d4hecSELjiigM+w4xVoUwLYOMtLuh4fW0kyZygtcexe6fTMzg2P5wroHHzioXEGyqsaW
keVSlroLES6X2YJxe+rw4R3LjWqZiOAc5l5vm7ZboLODLdBgU8tZID1sasZD5qK2uCHAiyVe/KBZ
t38Q2scbRuAhyBHl+hrMJeTwMNI9oO6pA6ruwENUMuJo2Y/MqVCfziQe2PkNcjeyYZeLFSIioufk
PzOE2WavkCrnJBZ4iYgJNqO5TEShIru7MM1vIsFOyXGRuCm70lMJd/Z0KSyCiBeFhFBPngMVI9zk
EypO3VrwnEO66rN1KGhxZV30M+FQIq5TcWzwVm5pG0Xfhvuii39VhUmykOcTWsNCMG0Od+ffSFXV
BbJ2ijNaUfo2oZLjgPA//UQ+JCwjEKqoVpDL5SQfnIHbZPBh5MO4+dHgx7cYMlYrvQFb3s/+7cEU
WQeMqHXDu356ohvylqRTEHmZ7FGPXJ5KbcgLAXWBDAt8b+S48Bb5GY20q3zSphQPOHpEHRjf+4lS
jUU73QyHWCd1OSrXxRkyTda++NC5LCdW0GFXghQeq484KWYwct/VfS0X9NRzFCeAQMKwWh3KP537
JOwz5vppaIx8GmYhtraUIlepX8RLp0P78hcm6Scs1YWbkrkYIZApoWtsqX3XczvOn9FWyHlFAMy8
ZC3I2UIhqXVFFay4bu2UIERnP0o9laguqEyT5OXBD10thxYODV4yM7A2iwXXWtPETLSMU+8QLnie
y1awh8MaQkySohUlQwPEecPhFIX8Fc1g1FDk8/jLXA31oHcB72rlrnJm71MrUj5Xgm/gRL08sOXy
GwR6oxfxcyZbwS3ijzjlk5qnupTy5EyL6aEwsPiFPllQcFyNPW6MyhbKVSJzsBXjDJIBOJRbEID3
WyoI88DNc0KRbSkLHoS2Kgwie7NNZESg+/+Uwn/xPmXNFaiQ0AsMsQ3yEDoqbYNz6VcReJkCr0ms
SwzhEvmwgF8slN3QL3TWXC/hz8Wy8a4Y8NW3hE0O06BrSjywCx3rnxV0ARU2HNeZVv8BNh/XKfBX
vAEaNYWYdEX8YlSHF0pec6bW8ug25xUaixQI28bsAjXt/D+9dKH/M8ARoW5Z85/NB48ct19CcGhi
m1/hU1dC3oRK4Gha1rt5pQozqMTmWwclRbgddecjmVkZzFMkLT/MiVpkZvLHKGj0J1xC9jhY6CsG
bwEOkIONhdFtb4bxTDZ9LCwawS02br0tIuAhXPs79Yy7rGRfEMHI/BnggNdVpC8LYaH3FQalC012
LTGpEpYQWu4K5ozi+ecHlPVFGwlXOt5Xu6U8Yn18/F6Q1uOqU+CbDpCYFudy6LiNaBDb3xObhPsV
tmghBfb37M3EaaNwjjvjEKDMyvckLGDikB0ib1KIvg190R5zAG4KJxofKfP09xwSbf30Ib/x1IPD
oKCi90I5dT2QaxnMEbKZSnIOuk3xze/6Cmasr8TFvxb6pEkg11yjAwWJ3WEJmFUhEiGyTGdPS4m8
E9qpOmScBX/CVHoLFGYS1e6SoW5+v8cJQqjz1KOszszNJjo78kj6AXJs5RBPLH9qYjguS4O4Xkj/
zEEAX5W7vnQnWwLTqqfc2H+w+RvGk8mR5Keo7ZEOo3vAXvypOLetCmAe9AGDbpjcRs3cB41Iv+R8
UgKwHtt/9M5f0QwpBZsxG05594/TRMnpCSenexwMODlyzUkjSk2TtCjmolJyTR4+y4vbqLaA/d1+
jatEIlovbd2da1pG3FRP6KDCo+l9tz37xoBJwjhoQ/gkjUQ2vej7LcTTrYLYMvaW+3zobrrvzkDY
eOSlpbVq8UJ5YtRZ0eXRYfd1Fym7GNTGIEmETjupwGOHiJ4G5HlEhg4Cwul9O9nTsRT7NR2eETDs
+hXvyXtZlztNMmP5iQ0gSjE78rRs+l6CEgdUtxrPt8TB6lISWZtv2aV5DRHh9gDeAgoUQDWfnGND
Qdnbaag5w+kpe1r/ZZ5YCFUMnGHFczR6fIsmhW15Cp4a5zxNhSkfDHpm8cEAGe3vzhkcNCS4QAxy
z0En75XUa0wFpxYdUavQwUhLyBMgUdTRYSn/WnBrIwdtX/YG3Av8JcFJsO7uBXpzlVHEq0eLlKuG
585sUh3jR1zbwNzWcdts9H6EfYV71QbkL7VunM/TZ0l/BuNV75NmI3eIqJLAWrJHuuBRl/uVXOTs
iIryfvpLc762VnDBpXysCeLkhGRNz2dfT15amxpg7YYpzJGp9BFH+zN4PiZv0pwbyUmupX/FfIqv
KhOaM/s233e/2FgwtPIkLEJONGI8JkmMwsNmyo6YCkxtmptCtVrJOHzY0r0dDUa3/XTx7TXxQW6S
5iWNm6wCsCH0qZz8eakIOyBcIE2/EHGq4LzoK/XJr1DhPji9FjFlN2ioYIj9tMDRHfswKCl/xvre
7xRt8SycytnStlFweuG02/EtmVOh5fIbfNAO/SgFARtcIMx4nWEB0e8tTpalD5Zcf/BKaUB7KIFR
A3Gn2f9ar+Go0XDCbj1+c2W0t20H0zVQaATEHt3/f+yC8SbWB1TgENjQ5m/7g9IncDS+CHUnuX0n
5vtBs0vW82vvgXMduGU64AzYPbD1p4fG7FYIf6Xfm043diBvfPwQr17PIsMvNMkTMli2XLzCVb4N
NGBczqs+8N8ZX22Q8Xi3oBJhbSuxeAZBmBWc/2sMrbX6wR2ihj3KhnaEJ375HGSTAHrZr67E2x53
rVou/e4G56MQos3L4weYaevwErnehXskKnJ4nTSGUgT2EhoIhBmxGjjZClcRb6KcU+MZfwdDwcbN
8qXGbL6xCV/pBvR8yJnitAiIaAeDG1+SbmDawOzAjXpJ+8RJGG6+Y+ygGTMWZvXrsJ1FUt37KEUv
Klg7I6TMmJYS4cLTGBRjpzPA80BjMGL1dcj/r1j93vvSIZxnu0+9yEZdH1rKrFzuacfeiRLicAqw
cB41AqCn1AV09xDjuE9I13DJSnlbHYxrfONWStWHLJ6ZZ3Rd1zvA6/Q3ARAin+O/xUh/QAO688qw
cN5UYL+IX3yDa7e+ibVaPd6RV6Q7gVDSdk8Da1CDlYezVae5e9yv9SP8u6GfyOVk2eOhh3ito6bO
hohM5+3zfp/pOJ4HGCUXJhUbtBuXb5mZekyWdIs0AvEcuqVMjzVBvoaEc+4pu9ct/FMqGd/GVRJw
zmm4qDYx5n+YOs+M+wZkgnYo/WAkB2YtsV1MkqoYxTxZpfVV0XeWLrLTgJbnrnPvC4DwNMS/sn99
5p55DRGENcjne3IEqJtdbD+mB99h6xv+h/Eyw9rQO2/8QMqdltLp2+JKRC2OqhWeGCX+iU9Q0Dax
qrN5CHUym0PYVmPe4nNZSoh/vTF7EsjrJyPfFPe9cmHksGu51p2KVttYSmnb4ozbBd+GwShRy/JN
nJqZGKTIxAKqIeI4TyF/zhJmnZJW/JtxfKuMNs0h0MmDUfHnRTCJmZhrbTyto4wblWaR9XRv65sO
LjAMJZJEz6X0m/SQqchDfmMk8atV9La1FLvNn2F9CDc1MkylQRLSAzq5qiCEfxBkA8TkoNprg+dX
ncHnvThgKksMmV1bhA2LvzAILQfwWMzRsiphW/EV7dBVLwR0u5eYpLHBjYn/RJ2RzR0toRBa+jxI
l81f2JW6oW16kN8zq2V5MVdQve8gXuPuANIPRPW5oWhGXFxHiZ7dU8Za6h/g8Pj7AzMKInGnKnyd
k8PP3mkWZUnsqpmDwcFideTMsziwYUcXOJx065r9ojHGQmgozftgwWoCGEbGWDaJ5MuZh9CpzeqF
jXEH/dQL1bzP5UQTf9haU7q30yeiLxgK0q8a/8FZRCeegfcq+zP8SbVZ5mBzIvGf52Q3uZ8dLmj0
xqKwRODWjgbQGF5BgUKfo9q6WetWfE3c1htRI9/EdXCr+iSmAY0Ojh6pkXsyesRnb1ZCUhbXMXu+
YkMGkE6Xou/OxlNDkrPQg1XfIwr4xnHHk4Fk4veP6PIdLXL7fA6nTgiFic8RulrffKcuYYPWyDuH
XT2NMapnYekzQaP5E0N+Ij18EAIqmVZX7qgQ0kSyqHKuRozOIw2EbpkF0lseyDZJvrjOEIfzWx+O
wN+izmXb6MU0w4GGuNVXdOVlpPh2OCCRYan5yHUrRcF9/GHAUR5v3V47pgluDZaMuku8xl3/G6WI
ES2KJHbxbqWYGA5maJ0XD1o0tSuYryd3uRD9Vmk4X9xnRypZYxOPmkofgG+cETvGFii2C+GE2I/k
37wcvPEFbvEdtZCN2wJK8C6qo0BHOTbzNbRy5btUcn9r6fQi39mquAvKTyIDDTguH95HDT/czYyb
FqDjw7DXl2zi2sFwcBz2vNT/OdRxvFaJ2qfeicWQX1lPBLNr16/OSFMt/IKU/ng9mE3TWej5Ke7M
GEZJnXzTi5xrAnSwPrKJTIDDg5vvq7KU8CBqUYM5P2mZWNu60ceoAGm49rFfAN7lKXrgIK1Lf7NG
RuQEFPoogu9ui4ciqyjsIrkH7hKCc0bdmFt7dBILlvBhf/6AmVNR0IMAwlYHYqqCK8MkGmgzNZtK
5gJIOmRgxc2D3i7SjDb/pLHxgTmvVlDXuQc+sWFoRAD/w6XjmZyEgvlTxthLEqkVsLqi2ttIwSbr
F5GHImS2dEz1N9R/CQxLm8V0hiszOnpHh+NSoSoO8LY2b/xvIuYHN2JXyyfvIqOQ3WEeuJMVKZDX
bMNyid3C6vJb8SP8d+M+GRWz0efMPL8S8bHYDH4IJXz6m6HlcgKjP1yf0eACVrYmWLbG/n+Cd6A1
l9h6089Ld+cuBo9TtX/MtNCHt2tdp0nNS4ij3bK+i5MOrSPJcdO2FoIm3/bC3cDqJHWCnV2i3wQR
2MMVoOBYTf+7FHyAw4pBa0IPa53uI8RqNwlmnHoRPgGb42ps9c/q6NdGNT6P6Q4gGpvqvbuCEG6G
nz24YSErLR096IRUG+UuyH0EvXby0gVndWoM2MUma4L+iyex5Um2/xIny43Dw3vCo8feULEpLdu0
GBz2EREVcLT3hGJQB5MWiLwu9hiFgP2RIF8NKePLbOfueXq7uS1bZaSZVEsosGUt+ntkdU+iuSn2
shPE1EsrzDLKWUT9jE8pkQVC4q9siuTXgXs9K5yDJsJeAynftNMLPnt11fi2ubL/sdvo9uwfyaoD
1+G0Z2GEvXytmm3ffElThsRwQMqgcFJ1A44Rt8EeeYa2lmIoSidPzGBzGD3XoaMHa3ONavYGGV0W
qx3zqGc14QZ0AhB375iTuir1xuXXONAr/FmuHf/DoeYa/a6fBJnSYEkaoNOAXwq9ckoGRi+B1CPc
e5lZk/ggP0N0PdXPJMHD6LKnnq4JbM0vifvhMBZM3JYmVz5aIDgjXpyPk26aZC4KIK9HBon80phE
w8O90Oh+0KZhxRgSiOPky6PuUiACF8LKoAOAAAXo/D83YF3yz3/a8NTwuqzDM/MFh5DuSWlbIuCh
rHXya2E0yOu2SsomZs0IHteDjKZ3KGF6WLZlBEXB81JIbVsxNeaE6BXwRkrb1FiZAnUeK07pLN8K
6cWALzYdJ/PZqnzihVn2jI5KP4b3hQIH1IUwG5mjrmR3phdUA+JK2W71G7/LtfscvJVL6BtG0WS3
nLrEIUd/a/ccXDt1OfImwtiB48GFo0qNLh7v60bJGRRrpAsVJ+9BabK6wPh//RYumCnBNG8OmHVo
oBqMg1MYoDyxD8a3E9UAQBivtxFDfnTf1JJjD9ZY7m0GIjX1RCZ5KZWscQOp5WVw6MYqgwR9ONAr
qFwMcP0Uhk+p2ty6hUbQ98C2VTbMSB2CdjV4+ceQuuGEre+wRgtSzpIlCYda6o5QAOJI0iZN4ZB+
SHgKP1lTaNL3aZ50deTnncCbRUHuyJilaeEN25ihu8A8wzZhHAYxyeLSFhGSnbTIP1Cg6mFwY3H1
KR8FW1KaSNZnJrLVBG8O71iZc3fPS4lbFpuS4sm1k0iFKoPYM9R34aNcC6FrJPoZ69q7MA00tGek
ttz8u5EuUnewRgxGQ0c+ZAQVGpxpZTq4yGovpmKCDlPm3sq8FdKTAQ7bOBA+HR9OA3+/EUl7N+PC
lSEj/Tu/PnP4MTU8iRhULGcEdrmz947lIs5okXmF5hz+EkaP0OisfcoR1YJiB+DZmV91AOhPV4ZN
fFJ9Bdp2pE7tWsCQnezwqoz+otMWTY33QJAyk/X8W1YCcZ77JNMKm/D1bsROkDd/9yLoUW1q1VLp
dGm+IVRxbBVwMJ+lXER+48AtaQ9TieUrARAkooSYWyzOlHwdwOkr2nVuy4VeN9KomSCmlo+Xoyl0
JbdLEQf6f4cHJ4Lo0ZAGobPoTysAnCKvcQDr+oEQe8JlNTGTwQrjyD5t0fINXcJaX4aLZ6tIUo2d
znbeSZta7UPIO5efDKbLttf2AyFF0ixLxQH4FzYV5zrqcmmhB/NMgC/TvPDTLzX9Tw4m4x8AlB+S
NsmYrT699jhZ2MpmzaVLdSN73gNek9gqX2mu/aPNl+fKkBh4GgS+M7l04bcz3vPSWW54x1RsPV4L
3KIi8q80/QhljnKw57crFHBy9LhLd/cC0RPbKDrj24FvMFrVGiEXcFNIBhSO1yZmOlY7UQwOx9r9
sOQ6cPeiqAj2G+nJrWZGHiugvKKxMhK+UWHYwswUTClQTFY+2KuUwYkfQh0qxSzwfuGH+OAlf+ND
3rjO41sfX71gd/hbzS3tz2oxBRFVxgjPtNfNdAz89KYdWHzjsPqFLLViHwCPiV/lEzTp/I7peeX6
Vvfn+4EefXT8hoPD0l+bzSuUFRM6f2gG6ZPYFNdjvjrRKWZSZz03LSJ65kB8Q6GFG61PUDVu2Onm
mOzjIjPi6JwTilOCCL27KNwevxVzuSiS1xabLjiL3ZLVD4YFxXGo71W0W7nzNQXV6bq5N8No71va
bB8M5b9Dmvu7JzzPK0eGjT/yCZNNdqc6lq2/vd19sEaQtxBx+5mKBPZ3CBD0YG6l0txfFXneGRC4
M3EQxwJLlDj2f0hXjuraV3X8roFsrxg4LlGPaTUOyDqe+m3EOs18p97/0+D8dmTqtxkuBPmMEvkO
XK46WnumYN8mSyTcUnN/o7Fib68HiQgDqFb+leU24fvX87LlQvwcHgob/18w6pZRZwiAWXOes+l2
08c9uvFv2XCroDcFglV3sBKsnLDM0UMbEvRlvT8czZ/9WHjzTlVH2fnMlk2B3WXeYzgZkdIgm5cp
aS9RshrcJr6LZvGyixcI1nJVOUh+v2zKA7hVhvdA8JHWP1lLPxqI58mSHjhqLaeF4hXXIXsluSQ/
Z8kxvUnns6nA/dpd1gWws7CNGLmMhxT5aJjy4aK/DJcpq7pu+u51eefhrl5zKo00Cj7qT8pIA9YM
kb8ioo2eOmPNNWLpSCYmtMVmELZdxhi5ng2RgdlRQ7qWSDRrGiUF3DutDFigmf30AjoAimm+BubX
LhbXbBCCHzhSrksjtu3pp2v30dvMGUksUtAzmRKl285DsPcUoIfral4H/pn8ZpiB0xpQgnJL7Sve
yDRis9ZCl+JxBSwgXITmrX/bUFPP4VWvT4QLQ6KqKgGa0WSWYdpQauD0tOhHaMDPqQh0P8j0IG4i
6vhsQbe0xHyo4ecgWBDvSf+g6l9NCfAZwMrFZbvj2fhkXh0ibShLMm/7+rB0fuEyvHKxcUupmM0x
Q9N9xnUud28ng0RnSJUwevnrHdub9X+iINhpEQDL0+PU/05p009kq8ADPND7Z8SrLgXpQlNgBpw8
8gxuv0FJiv8KNmD2y8fsrbeVEynQFkmwCaaN7W3QYeVYlnrBCMSG/irYzr3MZqV1/REGDgXPcNIj
djC+7dAHwr67Dg+rmiGiKWibrvMjl+OgNMvnWsJ4CRKLzVLWCtHy0I217PPMZkJS+tKNgTBr1Yjl
/Y7iGS217moN7xnBQBqyR4Nsdw4IFHL3yqWlSyBTGTd12kgRjhI8N/Qqle7q1PnFfLqToB54618P
lkKZxsfPKVQj77OGrqooYo4kwyHDAyeuNmSiieEafmNWKjWvIU6fuGTMdQif+nMOwktV4LoX27hW
9FSNaMp3uHXa6KDSr/jmJQHd7rX5YnOEycqDJgvSyvZsbIEy9dwmLykU1j5tAK3n/EWouhPI2wWH
0Fl40EZWzqj5rNa5HTIplE4XHC5qnOLXScgiIiFOC7WbX4IVz2BOFs1aXfsbJ8Pkhey4CN3ZHeUi
haEpwdPjX/Y6g2ccc/1vNT8JXXVRfFbr07sxX8c3uFRPdQNQQ3Bm3WJWXAJaesZ5sohD11HMAAqr
TNWcgBVy00ZJfP2Rh/QNjFU4ZOwWxz5lEtqCq7S0V6VQerfOBa5mHs9NUcmji7HTbdGt6nYz6Gg6
mIov2QV8YPjRJKJ0aK2Ojcv7gkakchTIiZPsm9NfYF3tO83KKMvXvxK5g2iU0K8TA5TmVDos4YO4
9y7dZRN6Z8tz+KyFVyXPcfAEN1jA5j2WLgcsn7BrPq8XdsfWdSVmNwY27AfKOGhH78PixtzRuJ1V
rec3aElt6j7Eh9kJ4v1l8SxUl6EzYSC630ocixQm1mPK9487R8vbJXXcVudFmOEcxOh0q1OEFnDu
/SSLNcu/YlJlRH4U8JDLOEOMembxua9mJv5HhGizTuQdqbd7AnjDHO18UJUO1h9XJft2fqpUH75K
+fGqwL4TXqA8oYJgju3zMI6UPhS0wP6Gda0CBB7/jWyLFyUHRzAVpGxAjahUr7eWFi0bl3/fxH0m
H7LXCQCR7wTRgBvuS3uBWj3l8B2t7REYnx/1y5gIMDY5ZWAe331ul9SaxNSOGCY8deEwZHowZjc/
sht2mIJYirkibTcKD3eQLjgjvGXM0mHu9ltnSPxb+5DDulHbIJzxOFQthyiN0gVsBACSay8zYjAl
itY0VeCOtRjm+RZ9ZVIYFx3mJJICDkSdRz8jbJCDTAyKenU4Cimh5sfIqASJRq2CQ5wwinSbYmgp
B9Ipmiw+11OdqrQ7F/hDwAFGSBzpCFVfAbtWD1kqu8qL309Sm9ds9n19LhWLMQO1Gp/DZwFWjwe0
jCWi+KZo1KKhO7VKRLerJHuY+dLXnbRAsCbKP6m2JhnUAAG1qWJ3i+DMAwOFtMiNGCM3eW2M+WFk
blf9ORgk/uuPDW28iaBzr0JHD8BwF055ER9sM7PJCC6OmO4+399SKnDdurKG+6tsZoddXBhSo3ah
VQTkEMykX6OfDb8KksGsKTohmqHuIWSXm6IRl8k9dUbyG3ZA866aSnJUwTSxZML0+72gjaSmhx1x
m4SFhRTDY/wMxKL+tN0ll0j/iDa2sf1fkuOzv6VwCgz43cYc1R0yMGpaekG5uXF9NEY+MpvEaJlY
7SBlDZGisChyrCrUBVT4wOMk47TphoMt6Nbn4oK+vDSUyZsRna5PeMU2F+SBD7/88ar64QY/0OfA
WXS8l3c7I8bOki3L7ipWvo0GlJNnVNl/qGxFzMYVZ2ZdjYzGbNHVXXIKzGG0VZP/OnM4nS3aa6DF
LBQr7aY4D6Ehl3Or6POlJD6uoxmgyKh6QuW06S5PFmDFltqEvHNyN6hiH6mpOZEVlVSx/eXANVdZ
Opovvv8BbZpE2+GxjUYjf2GdhNRTCWlgSC3pmQ7B5dTD2nPK6loYEbyBFDTi+ZS8SY/8LpWzYqGB
ydCJyNO0iZ2Y8/fRerStX3JUAwNc0kuqXc+VjqK562Xo9PFCbwmeFDq2qaJnlGFMXszk6UvCbnu6
KXPoF8HDz5XLijSwe4pJzSSfvdFLp8oMyuszBOKHG3SXxSCyF8vcdN9PcUuHJAr2oNvR5fPM36eQ
eGxiPjx5Ceh2Yday5ntDshwre39LYsgi/XiU85TArCueYj69RspCw7NRXnQDgDH1e+Ob+y7pj3bE
vUdbpTKJXp1CMD6Ycd33TSTZYcQIAp5nCterbJuYZbefCTSnpx43gH43DX3z9lUqbt7MAw9CZED8
AYJi5KYXxO+RkYWbg1O2XkXiyaBvfsc2ZqOHGmhOQcZR9ncTwNknEFErzTczViWc1ykHF9pMdunC
2omP6swMCm/fLZ4R96wynSlaBvRv709ZgwEzEiWXyr+Q5hf89J9mEimfIld4qcskExCpdvU/P1CQ
pastxxHH7XNjxrPbw9Rypze5qUOqFQl4PfEr0ryKCATzssXcbt2mAdyR42qoRkCd6LN4piRSdrSE
JjvMD65K7gYbOZkYX+IiPS/Q9vvvhZlEXXF3S17Q27eeyVX+8agUi/5d1y7iH7G4KNqHkjYNHaHF
r/h5jxZWdxrOvAg9KQHF3fuVkBzffdkQ7CCxrKIAsBeFbuQh8B4nsUbLLp/kzcTM4QuGRDNwqBvh
eIe4N7t66CGh3forwb2WxmhS+xA3NUCy+gPvPOyPjJK8izc7GW+VW6R+D8w5PqlCq2X5lN7LwJM6
aDQnt6gZvaRbLRC/9an5qa/Bdcd+YNAZ42hhR+Zb4jVfx7x6EaY5F8votynSxjr2xqve9I8EyF4i
q0reD/eVXG4XoImoxa3fL4AOLz21lNiseBIofo0Y+sUQeIFyEDYVjNvNSNJYkw9zRP/Dx8nsTdQz
CL0dXWgo5zmo31pQXuDiNbS8s7jaRUGvM7AujKyOZnSyPN9qPefjggAph+pmG+6t6eQ8nZp6+Hx+
7G6gVs+Pp1+gDYarShefRfipTbrW0nS7aPTO4YteEGqBkj/B9Ox3QsGB8Mc0ypecwc1vEfRIo3EX
g8jDsyWfBx50elmMi4DOzhHABPTCprrotPhrC5c4Srv7V26VGptdDkK4E6fmQFZHCLy9XjxlCeFQ
ATJI6FZBIAbaCqYc8Lki9dU3K49ChY7jcX/qPCuxqXRV6SYsJbm/PIC9DoA2WuE4ZA4+QyoZpAEk
7WAdzHjG5yGEotmZ6xh4J185hgAD04q7Af5ZP3exM3Kh2+x+9Z9/psz5pA9hs944/cApK/Sxpjmv
BZO4lONhiimolfAM46KMJY9hmt/vK9V3CbklKcJjZUhQo+lOg+W52oZVIgmMdBGWZ71jWPykY1ei
v3IZgNW3oBbXi9jWD2fc1heHTcozQpe6uSxU8dDDoujSoPbd7S76NQWmbOn8C/xDp/KmFGUF/zcf
8Cqph/e29Jv6WLh5gdTCvbyG4KZzkWkX5bv/38+YoDYMqUrfxqMeEUKeEgQxmW1MRMyVVXaJ5HrZ
CpqgdSL7twukv4LNgYVPgWyp+3TOSxh+AfdmMzYgbWWuJfgZ+2JxpC+IZyYQULu9Yv167FAfW9iH
KZps+hKtD6v4rtZxJTPITRFuiuuIq/kiD9HIesY1x2Er7kMT1Ripskd6TLiZwA2nmhhD7ThSppaM
4I7AVRON/1z27yStKhWNS0IElMgMggB4eIggWe9hOvFcnLP9qwvTTWUsUixOpv7fgrGKFnRydVom
ggPLpowEJyP8sDD+aCGXbFCRxOlX6bpToggB07fm8LG1hzhdJmKe5ymC5GZuRNk2406EUxmjiIyZ
6qN0PHvZAVHR1pCyMwSa8/47rPMS4qAFpUi3rK0fQq5XBPrXXsADNFZyO/+jEaAiwzQx2bkaTYRj
0Kohlhg866+mIYCqt4D62ahCxin1wFaqL5pHD1xGLFilLD624KnFYs/ldKdBLzy0aMElUzNbn1/R
UBsXKD235Xg2PtfEolxTk8HHQuRD+VOXE7GA5RHTJkkOnEAqxYj0y32B2jM8/LG3Lrnpt5LVO1Fn
BWxMy33MVe+EE/Zy6IsTEQF0quwujJf5z/fzpXXiz8Bv5kDZ5dzMXohR83HEBdXCAZrJYev7Xgel
AjeyVcGT7xwGqBqPlbXaMF0ArsxcBTih4uhgKX2On1GKl+bKFl+quGgzO8LtXbZJ4eucJJJndgan
0Zhak1dVxcXvoyHWfITTACuvIpU7ooiFGNKS5Er+QjTUd/GeG4u6AQkQCWwnuZguwMi71AjfQ0Gj
t4nDjw5mixlTLC4b9SNw+JSGagqhNoXZtAShKXEUcsTgq/6z1PbrI3nYotDKxaz11UZwF/IcBsqU
Z44h1jOdVpTrq28yDsx9nG+LSFxT6nQWYJUW2MJ6fgs2RQRWcPCta52fyTEe2ZZUKOIpGwsN2teR
ryyBwomVZiRLhtB7TUSdt+rp5qRGRSBkLfoVB3LkMchrl4gs95AK1Hcjqn36t/hgE16eNJ26jDDB
yDPRZ1tfXbzJNDk4ofghTPd1gqakJ0ZnzwymMxCdGP5rg+5JuaospB0/rWDVbKmv7DzhHaNgBu3S
7eTrOspt2NdSF3Gd7JMhSvzKAJxRsqixlG53wvlKEfM1Wl/ewgymEaTikLrXtWCh2tfwdLLraa41
cN9CnzOux96lUJhuxsJIYbmFjTXm4YoC8xprr7MzKrOcszuzBkAkbWpTohw82yeohPBo1WW5ADHQ
UPHdZSZC/Aj+bYPNjiLsD08bpWW9BzzoCD6A/QdGnWLTMlBDA84wIS8U8Ate4Odx6qW1ffEE/JYN
asvXBd+GPVmp8vxpBevWecHFDp/rlCkaiXFY/xCe5AQ0zMAshHEKmFYyKCCxkjb3zn1B+7QxdNHZ
6eK5pSF0cuNSzJB77PUzuo2od3kZBBW5bO4dacL2UQDY2va9nU4TGnk4dWiYMfzucA3BnHX+Iwif
aQV07w6OfSF7OSJVHOQtBv/e1/5SxYN45K9SD0hYS4JLbhV8Ewj9GlgRJEtuZZiOthdxH+fEVWHH
gnCNbfNi5jtIgB65z84MAfAHZgvEScxThtpJ2rIY1kisr92oj9gXj+CcDkA03G6o7so+CW+0KUpM
KCLqL6RG7mJFCZo96XIQTCJqwZP3lIH6K7BaI9Hw56hvpiNZFiSwHYRtnMmA0ezNwpPV/GqE0LRM
NwFYug5VXxztQsIFWhfSBWWzUK4kY5149Vz/zo9LZQm9CWieTqZi8+gYJkfYt1094Mu807CFWEM4
Z5mXvt/y4004abJrP0dFt+Rt9aohmUsbUohTsLHK0K5EwTD37Ati1IKadCxyPIHdrb5S+0Qn1LHI
N5tCHKQufrT4JZTnb1ZcU5NFQ+HTrgCW788e9arNW9G1dmi0cBmkPgvw4Tb2ECSY9Ibv/9FlPT41
/ZeAscplWDWFO9/EQYV3fZFUEvLZ/SR1ur0tWAHNEQ8Xjg/Fs07iwbVKQOKIpjRE38g6wRbYdSkE
EF6+CA2kyzUiQ9AS0JsD7q7hbFzAKc8RWTkQhzbMcxN0VsEQZSNysn5VnJ3ecJi1gNhXw5CDEszD
zX13FzlcLQzQFLqpj+BFnyIcDKWOuZ1ZdXe86oYIJsFg5zY3HFe/TuAWKDkEDDQeYkOnxW/cyLHo
ubXy+lsPA8lBATi9WURcYB9d0PxMfxEkEmAeacCeInUw+vvx7mQWNtG6HAgQIA7V04hKiaooMKP6
2YpWHhVRK4EDhka4CT32PwMs9XXSPyORr07xpebVTIF3djP0FkgQtmURZMEsZExAv+5vKzhuSalV
JWMIS2hfAVtFVGcTMTxjmIhAulGP/j7tg/wlfOXIBFLicR9Xu3CbpUjXHvYknHJeN6MUfdNHNQ3C
4TRTsqYxcEuzlRp1YVe4SyJaagrx5zI5aca3qA1dGM7v80Qcg5S1rRqrlVD8H3yr2o1poIngZOI7
vne6WBncve0ueBRLkPTgiTEX/IWwmAj6B4ha141wWOKBL7DGIVNJzfbXuXudUsvAzelJ5kodU7Ps
x0t9e2m4r6noeoe2qktroPb5BvZ8uAE2cMPydkL6QQsxkWmIXOHRmQtRHuaL2ZumGkVPAWyrxPn8
PcUujmDFAqimHFce6DFXrBaxwCaF8HtUYsNBWleolMpVR3S0vFpmshUP4QibKIa+FFIbZqhSLDSA
xd0dvtdeRv98I+w/SZH2AO+QHclOv27bzrNiqWpHK5f6Le/NtyFcA9axfvn2+vDPljBQmpzv6CLB
92I1VKsJ6alEell1Kn+HGafkw62DBCI6Zj3zHr3hWCgHRYs0rlQybzPRj6XmGPwPvRgfdCnZhkuw
LKsG4u/xOXJXss3LXItmh5W6U6dfrnb0KtKRpWYmG1vACc6p7u9gIADUUMARWlDy2zX6meOdJKrR
7umgIbwtyIS7lunG2kObtWdms4Wrz8UJo6yq2D8YJSMaC2NNZpnY1ykZZVQ7RPswRPpo7rXDwyqA
tFDhzu5uxNITyBN0ukgRsm2suiGhrC4v05QR3BA6eFA2W/WgC6JaVObbtcZkwskhG6UHXXWJ9w3y
gE5I6G9xre1f+6FLgeaJoJLCMtfVphA43GvXnMvzITAzEUvk+U9F4GCbKAuUi59jBKQ/cimYtLUr
1GD6Lfe6IOnhW5IW+OF/xNsgHncmVxnGyItxvi+gtOi1bf4E3BIKOjnhQLn/cw3yD4TMjbZf+rsn
N1rf2T/oGFUnjllMSX2pqAATA+H8v4RV5LDHzhEbdFnVckYKiOe0/LsgIVus0F3vtQTgoayqka/c
g5keqGSOOLEm5FOlgVBFY7fdihYCui47kM+rEsFU2+ppKj8cadamd4M8qqEuF056SaSlZyD5Rzxy
JPJ5PDfuLwDUeb03egcXB7DGLHIugtz4MzRL0izSZ6UKWUU2YP6M0IAMnst+XRXg/tXUnkeoSRtg
fU/4QcNfQXhT9gMQVUOkYdDwTvID8v8j8BoWnWuWVbDxVNEMwUDDMoCECkAZqTTsGD4SGoMTCjSk
gtZ957jipD4hICvLx0A/+MpaeZs6rcdhMsyyQAGDoF1++yjJm+ap/KJAqBz1V/HY616b9vLAoDvB
tDEd4Od1f2I0FXB/pIR6UqcnKFQvm30ryGO8wcuPF8+4Eeb6o5aQdtld51dEjc3tDdREQhT5Thze
LmTvsY0yXq0PKO7dnECaSnUjAKnu3SDib8VKPzXds1T0ReHRW7f4GIJRq1z8e7MxqKxuprwvzRBv
AMOfWx57idkSDwZQXDE529SI8KtTBDAr+nqvUiPylfEorGS/Wi9xjFACLzR3aWWDfsj75ZHffR3i
5+sJwbBVMe6fZ/qP0yorZrNKBOqyuuuYhmNBa1MJvBFAL0hQdArgVamcOzQtPxRcVWSthQwx6vwe
IbRS17f4sLhKKdoK0xokFzA9hFQXTorUcIachKSBSNLFE4zqtl1E91R/ZspxiZBhFOZcT8ooi2Sv
c4BwpY5PLh4cUwodW7XVVWsqbKM16/ddUv1etndVR9fW4x84JxFZfXdyfkQJi/ZnJlwbKG3z2D9w
w8Ag6VQv47tdjZY9gp252FJj5iBvFKyKt5CYglOkuqlCwR9efBpOuOZdExfKINaV+DPlXXm5CzO9
Miv0pbXtt9YCXbNJHt7UjqvH9kwvDyxD6SYuwHfY3oVfZguSusgtjsDLrp8jHClSEBbx59r4/iEq
vJcc3yoVqJwnZErIPp589LqDWhlZseiRoE4EU+7v5Sj9JPWWWHBgIM8n6pmnVh4bUStyVzdVNVB3
lcxpEHPP/n+xJbw0E+dzJyQizMu4y3Ubr5veO1AFEP1rTwuFgMkv8rJVLYpoQAwPLr9kvFREUcjN
Irz+hkzOmpOnXbR9YcNbDbur0hA8TnAfowIkC+jzbgF2qP/7l5aeH+fZslBrPtqdXvbiIptMnh+r
BciCqpy/d4E28+0eg4acVpomComXdYanZQnCpPoXCiHv9qVTfkjy1eH6loQQpi4NinKeWyRSVXy4
VydXzcfSkPZ51UxOD1lqZA9eKf74eyW/GwDtDMGmY5oB7DGimBGtWD9PIeD/2gZwhdEnyjw3MsSc
anwpdok7yFSQBIBuDEwdefGfNwbLOXrqbypsKcBBLVtQQ6vVH6mDK7jfqaSDvSno9jQXvHbnaWM2
9sPCsvy8bGj2uTJ16qUfo1ymNBTNX+5YsbBdpa0kdjY50QeOTNIO84HaMsjUrFpu588Bl/39uEUI
j8Iq5y+zipKVimv7PphqTFDJN6Jw2OxgftmkrLjTpggs0PblpKXjbtytTI1BvQA2SPbg1KuZCev/
RMnLMBDCmmyzsT2jWB/ojefG+HLxtoXCfVyl2UvVukvDq+6qers2KioE5r2+X0WWHYr+vdTrLoFu
EQevDBKt29QXHSlPvRVnAH62FZcWhBSAB+dkDRl2ZtnmwM/0l4v9KZsweZmgjHsZ/ANmgF3BhkQY
+5rq40GQDERoLA204T87zwKbqKu6nE7hHvgyh/mzYegCsMi8eeTGQPIVFp99vNc5ON/9RIPkb+PO
onCwVuanyjpwMxjtkwm6+VoUl4TsbIedS++pfLFnokolhcVrLsYZY4GTOWNC7ZrYW5+am4M89qkg
wDQ8iCuAJ6wuMQmBz/0SilieEIZxKVQKxVbOmqohrxjAu2IgPHReeRppOTWT8K/XvqIbJMfLsWos
p6rrq+Ax1H9bgEOuWQDiUWNNd+BuvIqVtuS95PD7bhtUDYSmMS+76/ITBk5RPGG9zRThvAtTulgI
iNknvqzmkXvc3EAdkW+j+CLhgWDEjReVFNbp6itJh+JSpdh/7vqi3XEjq214umL/F6hc9dV23CPJ
FjsrCkr9A8Ag2jnpFgBOrxjdXKIGKBhsUAis4EnVILf1rUbjt81UdKW2pED+vsxPYNRfH809sNK4
P6qlSaG6anZurWTy94Ud1Lmc6U7ScaJd+i0ao6kgAvQhQakI1Pb8MsXUP/NUayEGGHjnFk8RLbLV
o0fDopMH5+Ki2I59yTpEqXy9/dLonWIyx+fwyU49sAkImK2V3ZwFBBCjszPaV6JNaRFccwr1j4BU
u/3fe6o31elnQ0tOb/u+Qs+SfRqnwMV/0c3AE8SFKqpzsApYw+Yd1NL7A3kWo7m/Z+m211BCkAvc
owOUNPqAnCbMiM3mOt1b2Q0Spf5YgGCPhr3tdKREHLy5uTmpTzBpx02jNTsVoqv2HDKGPxrcToyq
cEHjeAEebludmXX+Im1C5CIFQ8rDTeZ3tPGxYx2ylow2Xz47kPdmrcCC+UoNghFa9Ym83M/Q164y
xqSktbyyewW9CSsaHHuA4+4T9qo9Y87bscUeQxjdjC9Tj6Iey0xSmbwuWXTDjINdl6w4DzrYIXH5
yLitUn1zfYqLyf0gSOG4m6P2boxQSiy+6zJypWNHTLsN0J9I2Z2sgULwgKK4uROv9ur2xJgmx08I
/hcyw3u1VHcB7IuK+WdYwT8Zu6Pgo+gs7BHu7PxQsinUjfqka35wPryU063sfldZ9mzJKEsA7mIp
OPs/vYEuhH4HXTsw2TBWs7rO5u055AMFrqlrnt3RjLNPnLW9oRYhgeRt68C15UJD2lapi6sfSztX
Xjrt90vhtF/sqxfIg53t3a20Y6e5uB2dj0ekZn/OU7pFxjCyD0plvRlNFqO3DoDProclbL0C1u7I
jNduDharmDIHIjN56an5HuU+qhG1YqKmhG2FcwssdwRqsIQm0GPd4yZJU0oyEQWkCzAMHNs2eUaC
kc0Gg6o28QN9PjD79nY0M/+Nrkeq4Oyujtx1LGiFvtqyAEGzADNx/Dfp/tCsA0baPWaIRjPskjv/
NZSYd8sUUmJFOiQ9aRxqAfyxFdLzBAD1JYygsDS5o6+2KiY6dwNa2lnSvqrWfYTtGJRpBczXVlB8
B+ZY/Ibd+PiRA0Rnvf4R9gtPOnvLWtSIfrt8jYW7qI+Mc0BCe9viiRFCSauwxebeDXPEatWjWP9t
SaaW7vxXZIY+jhkZkV1sxlJZiOn0iamGxENbCykvITzrG5IfpUBlPpC52yb/9//tpw1dZ/gj+cvH
+idnIVAs8/nj5Syz/BHdw8croI37BXnJvcr0ey5dyY0IZxfRIzLw5VSi0lEAOGg3RexxTyFzxEkX
/bUkLZ3VMhqSo1cYqV1YT5drHSLtly39sytDQaW1nx19OcDfQK01j9RhdydrGxqhemNAGvu28dy/
JZD9AckosFIuwjYa88MEQrlda9NmWz/fvCL37bnO0hrHQdLxydE82Bg89Iodok/VIah46tb6t3qI
p8w8Z3BIfky1h9icp1T301sTQrC5udn4yY4faiS0nrd5IQnMvlDZEZcQGRpfg4nvxQuZ81i8/Ajp
10D9LvZX5iSLWjQ+fAAEshCIP1t/0e94xtvXpddGLCQ6OBVQsqSu9RKpvaMYBO3xC4RHQ3sRS4YG
q5MhRRMh/3v3ym5As7cEgFfQOrGV6uf2K6Z2A05qN1E9IEhmgbnMWJL0l7OkXz6pbaIzm0KrjjKb
lB81ZPG/Ue3TqtnShs4tBROnOvHbOfvIsG/kUlLLR8Et9adRzJxI/Fc86nh7OyP1Gv+SWpQBUi2q
256y9OI/+f0YFGGXrGdbC6cGzVY/X5EPBx1HFTRebtWvwQdb1QfMm6PV6gQm4eT2Nb/nntEfmIKf
y/3oAYH/rgbM7mTflgzgbUpzkWFXAv1jxHVrPZBFsZlMF/MYn5+4fsXo/icMeCw+D3wjsvV33Uyx
d4487ertO7+AK5769lYHlP3O/VePpubwkcEx5aLGzsZzz9HPQiLZsujBY7OdnZG/ms+lwb0p/3M+
m6ZQ6GplUt7WpextCIymbNhLmOr8owcgnz2oz3jweL10GWQBQm3LqqZOpXbWORMivIweAA5Qqcpq
Eh/ijIgjzaSKOamyUXYjTv6NXe4nvcsFDvOPP9w7WePniRF3PVCdtmM1333V9hjiIjWfSiyTqZW5
5qW/9yHft1RmZAsW7BkntabMjo8cXLOeQdT4iHOFrgrGNZDCNOw85ojmnET34vuWznUd2JskrXkB
P5D3rqoaPfZCZ3TTWkKarVzqpx6W5tgM5hjwLWprUtO3zmnUOHpERCYXCmiYN0IdnEFcVrOxEfXG
iXEDGQPVpTwW0+e/BqAp5UJ/kOexyuZ4Lc+6FuwC8beacv4LjTwzZ8Zugrq4ZKoEExYL17MtSEFF
oNmrbh+LCSXACa/LxPFqQLfYih2zfqQs8RMCFKcJufzrVH9ZBfIarprwjOZewBe7ysI+CmjhnyaL
qkFigzpVlXh9SUklPvLhVoxwPsujF7g8JrjCCX7xvTcQPCVrnV5r+qgBBN0je39/P+JWhVD9xYAR
PbhBV8qFQ7RC5ricrv374yluRIRqDdoeufENPoJ6Wo3Qn6xZCLkLWONwG19riJhG45WX5Qbjuezy
pi6TjDIkmEy8g9T0VJ1/t2tc4d37uSH3HsE7WdP2G2cHv1dsK2wOhQcW5/5qD8pciQFtTkfakkfg
dZjC5pHR7ZVngmFKtwB9iji5CmLomnPg/ShTRUz8h4NU1TJym42VqmL/gbuMq1nIDMG4LLlmjxvb
CgtC8oQiabU1FuASA/pKOvkkPDqeFWBMHZJEJaTc5sVexTCI/e5WMbCiBiyxNkDZatXwHUBXALif
mwpkJu9rMT/8RMNyoxPbt+Y7drA2pgLblRFyPc3pTtj/6+N4aVy7dl9KFvgHzUpan6sBOgwi18sL
mAA6sKHwQyZzGYbmcNjazvPjPzYw1CzfToHqs7wD5SpiOBZcarZCovOHctfVmbBbYXSXUDOCzNRg
2gwi1itdnQypODX3wazjGRfJuL17gIpJQ1oRhrVJi5ek06aKZH/a62nD0ikOK95zydA+WOyBgKWJ
KETqTOJqUo1q3M7RQ2tFYb6GO09W1KE3kwW8O+ZrHOqZfeUqQWeV0Kz3vjDEHMcY4BzkshM7msgH
RPDMuxu5HO1kKVKkL7kMe2rL8J+AoY3FYKxGLElEDrRztVdbAXxVsS8Xq9qZ2EIiqM66czepIQCo
SCkUsJ/nxWwZJg1Znr4WijCEo3ZDRcykZfBnx91xvC5CtlUudPOkxbGt91CMSag2iYgAGM+/Aim0
wuFqszpxefSv5XAvC2T6GSV498z8UE4tDOjGfPk4xmviLuHRZIYw0nj3dVZGcyIem61bQcqk84aL
CV3ujAZFKehAkUSJu0YnYXimYErbUqg2aT49BfH62Sucm8OjZTFIdTTH3wQV/UTM2R7N6XW/ZhN0
Dm9HerK4j+un0RKx0iEGTlNlX8bisvN8qY0XDNsTwOaONloy2jrdsLqHHRG9AxinITKAw9ae6h3w
fpycqa0x0GCy3DN7Ox8BSZKrYg4mGvhkDblmc3EtaSkrphFx8FACwJj5FAeF1YqFntxQuFncx8k3
NRyRoxeoRc6TevRGZoRM9s6V2Ejp0R53B9xJ/0zTVmw/ea0XsOv5NuBUWk+YolxLzPqyXgI5j2Ds
RbFnnansjhu1OZjYUlTTJdjtzNL6VbmeWOvLqGQCq9wfuHQJPnNSeJQq4Zso8qwDXvKngSVoSckR
OxzfVF7gWnqb8BbI+uBdpDGlryIj+3E9kTDOu8jOTyMmowuyKHOVJwQebKQ6YbHyPLoherhGnP+h
rm/GHFzx+S8OpZuAGOr/9lxQpBsxtii91jZ9ScXsdyO6CEzdgKZic/kLskTYUDR36+NUPQcW2TRb
Lv6Q2ZzR4w0B7Ei4U5QG6X24ky4idxavMUCrb+1KMHblohF8d7vj0hazfFNG1IRBtqfm3s3JA/p0
QfpOKk1S8zfe51aiaG59iAoqG2huh+ATKzdyHptzfn3xSIfrhrHGAbSVJueV6TFg+egvTbqzW2j9
KrtpYDTWhGUyBvXsdGJhJ2VuXxstB6xM3RvedvtfwvQNsRvEQRV5BHtADs3Nog3FLWorKh2dsVZQ
LzVH6br0P+xLmYUdDSHJgFNzYbV82yu1h6+MibvYbIFa3JXNyBPpoefsMqUOsVK35/oJjB6UW0a/
FYN5N6l+4O5mOmgU85N8auRhtSTppR/W9tJI/NqfztaybWSnqHNw0nea8puUIJiyfYjSogpM/Y3i
A5EYfr/uJ+9+PwSPpd5Q+PJ6jFyZRgrt4MpW5pKgcl3cvVUj2UNq4yB5tQH4cbtJh1VK9fnNy2RU
ANEsmyp8XdgpTD80flO8OAtI8ea1AqidCluz5IsWO4s5HrlfylzVlMuRF70TVD2DngzQQKdHtBEt
9m26rTgU7i1sFF44kncLedcuIn/KZvHftPqHnRAJILDfsDe0C0lfwLdbH7aSfo4knCC+Pwr29k1T
JDGt24BFRSHW7xo+3/zCedbwRsyxQGPSzMdY1bkLuz5oMzR9q+m/cJ40vx6Ebza9oGk+9JR3/DC1
0fVVtisIn4wfhDA/psMXOMfuC1jdB5S7N8a9DgB6lIeZWSlW30i0FSQHsnNKY2eV1ymxbRE2YVt7
GtN1QFe8svekcMimdmVcIHDAhwlSvzkTgzddp9BntU+5aLtIlGv32ffWW3iWsbBiYnAQOOCtcqfu
ZcbZMI5VLsNSZPBr0880mfTDu6V6PBFj779XqmmUUnDwTFbhhUjUQ0Io8x/Y+cCmJxWee4P5lDqu
v7Falrn9si64QQV7t0M/HeHUwxE0fWCnD46qMaUxUu/yrH7zhwbgoO+qLO2MKR25JQZjGShSc92Q
Jb7YqpH6v+131O6r/0s/QaFnxHA3Rwhv98FtBAHXhJrt/dstH7e3bLNJH5bwRZwSmnFSzl62r8vl
w6kSCACGOx9HfljEviViD5rXbNs4diJchiaocohsdQupKjOv1t3JMaHQuJUzTo/5dV25dF2H02fn
q7Z69Lfjl8vSJzym9t5cyrq7pJA7W/N8/+V4T+gAV6Z9TXKeWViciTwiKyyuOHm53/gpn9EHbaNp
bVldhoX1ZjPpTzrFfiYOUE+saV0W76KOxsieafcpzWehPJvT7OC1mGbhoELRck7oAUfmqi2MyzR2
QjB4LAbvqWuq1rJaWnh8RevtyoXZ7NH2q8AZZDao5f7jKKez2OX/uZ+tJbtbbYvJGqeCN+N45Bvg
Z70a5KK8uq6xR80MTZnIpM20QJUa2PvrEnvvXjD/ixv432IEwdKkT5GoQ9X/pO4C0QmJOb75xHoZ
IF6SiZEfcS9BxQvQurWxGDkjWSNltdCKDxzGRRILviBpQrRUE8YwinKYED5trqM9ZCoplifWO5V4
tYIasBhORdOj/nKF3/vFrbby8jZb6TSKRbMVbRcbPQMmOI0BOvtYKgYkRYv58fEUJZHulx7Ny1/R
s9q/F9fIuhA/pSt8cwkpyFf3MhVoIr7bYb3nzVO9BxkZa9uAai9Mb9D61P8ENW8WmEq1A49iPU9H
N+qwZUJx9pw0stYhRrGQF2z6wOxUofXjzb984uVQkDGZEvE5orN5F0lC7hcmq6JwTUdvH0qh47Y8
TJXo+aMCDxZFUVukdp5bTGZjboTSUO25zJDhN8iA7iWICRDaMKUVXw8/Jh1OgvrEuHMh0VYfI6m9
ZfKx71MIMtdNDnbQ7UyhtNlgmgtPpxHhEhp4I7CHaHd3oPhtuSD9V857xaDF63kCjczuq95oCv4t
FLS3fboshrA3aLyyIwHGIma6npe4ByuPkJxfDFT7gVJUdmGVjrFgmReT953MAqbOgb5z7/AOl77v
+AlH/RalMWMRpe621zI4sYEcoYnvdWBr8RWXwUEOemXqukEckccAeaqsPbdJlADDAVCfN2pCYvN8
vkInPbyhn9iA+kywxQCCe+OFH+31DMlnw3j3EtckKLkIpJabod3kyrY4SLhjzUIGLf6vKLHy30g5
yA3htepYRe6mKXHN/ssAa5c+UBGPa/Lfcqh0o1h0g2hJFi8njWJYVvG+onSc8QdVydymlxwfj9s/
tWlyJVxrGQzvj3gEHcXDmcmYR+R1Wsce+7PYX9t3eNc27BtvdVCiBLnLZhN6B3+4cs8eKaxsDA9g
yaNmeODOYOHIT1CEbw05z+VHgy/cIHhxQU0yeaRZdK0+646zEE4cNS1yq9780p1YrmJ0T1iD72uJ
pFhdOqOKkt/Q984Qa3nGYSDOIVbA71a47lKwiOZcabP+2C0bl06AoYgSYkwe1jzAT8DD6pmK74IG
msaRNeCV6zsh0MxSZ55Q8VgZHFKDoRXDnlDqn1elMl6m/FMMwwHO1s9I/19S5obxpt3hCvjGKpkB
qMAZ3bDpGN/W1ELrFimFLfjcrZYCvc5LQKlLTZUeFJ1c4h7zo9ZnLOHTzXvkyLelUQAA2JInW2zl
Y06ZQv5y5A+TG6xEVKBbFyckxu4sTLWzDlTpbJcOVQ3XETxrvUkvBjPANbK9lgvdzAzmvRV8vBNy
Lc4nUuncjp8RwuNrIgBIaA6/mh+ajsQCkOKMQfnidzV0a3+8DciDXeXPU8N+m/WcmE6KyBjiuRPY
gerd3/yEC9YJcqDRjrWgVVB2NdHeJkPbEkgdeh4dXCTLe5WrqGkTwUfjRPVySsBSrKTFHV6AOGJE
Ttjstbw7q4/FzwGSgnrudNWPSsV7SPPJZIdSRLXX0vHO5p3DWfejogJa7S+WvkPsslVqTMPCdtcE
xkjkpSTsh6fWZCcFGCygaaa8can+bG2Ket4HVA8wqD3RDWwNN6p1TN6RwjC32cYzZ7DjKd7y7Liz
vivL6mFBgGXNaieNm7velCEQc4e/KoE/MbLfKlm1p6nHNLwZKRgON5bNfq7PF4WRPWD7A73VEcEZ
DRh70nbDACaNubth3ttG9w9ZsOwLIICs4M8YoajezMQUSEb2WjIygYjjX09AUUBXRDPFcIYpvh1Z
/FSexHPh7p9kdYSwtrdEOoVbkjd/A0ivBJDRmL1ZR10y885uSlZFshXadany5RtZe8M0PXZ+km6f
KJbiWJQtsA3I4J5ar9rVGEkP0OKN/ykvNaO3VGNm5ID1+d03bM74KBzQ6nuBxfo8ftKT7z1CZ158
2ufzBbpoL0Kml/cDOIjHXHRsc9RzOhKWP3ZmB1+AxbtPTB5TzaMtELgVdg5jgLpCSaWYLg9rFB9s
xYsftxkNYvW1tnF5GhJt29eC/pIU10xjusTEGOJDn1fzyBGrG5IItor2Np5RgrkN71iX1Lsam4oL
vqIT9Nju9Qs0ZVcllO/M9Gr158IxVg4+5hMZ0HqDFN6w4WtammrlzjVqS11BrdiNkCEMfscEYH1Q
+A3CgsZmqAEpyGmEccD8gQnB8dgxqcg2Ar5SL+065MDolgR7zN5+D/izscxb0gFM84qRTqXYW6nU
lYwJa2Fdzebp//hSUVKQ1fyKSguJUS540FgFllatfaRSv30oGuUNqWIFrKJh2uWXbN029LfDvOF/
03OsvWYxRzGZdBgMy4bzxPS5jqKA9WRXaKeFUu3bEIfrFHxEY4lDCbu6bfJ8oa58Wvil8KmEPrc6
JlBGU+0TAfin86oTzm2268Yh2Rf8Y070OCAJ12OY7qAd9PLiKtqMcpSGnoLmiJqkcSMqfJAgaspQ
0941RVfQ+VGtVowxJXwupjKUcbY6Fl53tY1u85FVGZW9ty5iZYcD/jDYyotUnjG0wL612Xai9h0z
9y2B6DUGz4f4f5V2VxoPDeDcBHxOyyDzwYOfWpsQe/CgQWWQmsQPVFv7QTlSjhxK+JdmIhO3bE+Z
DYPXmKTg0Gic8WQM5j27S5OLRe5jNQqlnJbEmoovXrCwm8AWUrAbEoCYWady0SFJGEUJFpV5XTFR
Xli9uVwcARBnWtWwdYXMf9fLoy9um723/J6U8ZS97KLasu+KZ8tZcqMjo6VSQEz42Tc88JWuTJMh
8IhoGYtR1FsZ7YMYaogS2EIq7K8mcUnUsn0GBAmYVeN2QGk3zG7LEFcXAOSdCiyRqHF1LGdLL1YE
juw3a2dnkhCr7lNk/89jqpdW3mH9PUhDl0zbeKn7V8sSFjpirWmhnHG8FrP8uox27qWlF/+lkDlo
jwr4Tv6x05xPDPtaNBmHOqd4ixk0EU1FnXux/PX/mAlRSGXGyhlMEBOihLCiaXGiJcNe7kp/yGzg
vmXf6Lq+WIdzStdWBiS3uMIZl/63WSKDR/T9+2hwCODqrUfmW1MC711bzo10LakLRvixgLGzPNDX
lRgbqmV770hRsFDJro1nXP2LYgTvNpWwUR6jrAoXgO/DDmQ/5Sqgh8xy1acNgZs9KHBaP3so6E46
4mbqbCrVVUrCQ3Xfou/IA3DLT9WapY6645LYOYQL+pgR2qNX+OAoBgZ007mVKV9D70sJwyFCpYSf
SNLI8D9w/sBdU8ZZV0x5uroE8cJvdJHhZ45d81HqopN0AZZffexLgh0FSrTN/J1T5vDM2F57pyjT
kDaDbZNdI9VV5aAhy+ji2bBccHXO80Cho/uxkUgzReovXCadOL1cVDXmj283EH3IydwAvfR2rZpu
B2ycR28zONFQmOc/L3ia635bCgWQ2TOM7mC23tEHzxlXjx0rPSp2elTzExopUwqy4zkxLhF6gyG8
44Tb3rD6zgoLOtAWYv6xUATS4N7b1F0Sluu03wk25hWZTJZ7Y/hFbo02HXo/Jrae74VrgKhsf2M+
4lu9mBbPEVu2mzCPPygMdO7StEp+kp+yoNlhGdH6BaAs4Rdi6UbQxM6EV4wi18IA5UeIK2co2xqU
Wdd2A+EsEF68jUYv9V8S0FUEK6EUMGatxAmdOjjB27K0VfTs16N4zOjNIhascJ0hBIgAX5ISNPry
IJLbK5IT45moc5tUwF3vlGr8rb26u7CCJ0iI4LzBAtf3VzGzkyPbc295hpTft/3BkkNzuMXf/w3a
GlSrO0I/neJ7EUVxEJPRRyEofV743jbOyl5PCEDNsRvq9s12HZDNxTozGTENiT95lYE91Naw4TZJ
SPLIuNVDhVSTBtbcDLiBfJ+1W3h4RHQmkeuJ8qhlG+euj8yZC2V72KwMuiC622GnuPoVhyVmlvBu
v+k7VMwBfm9iR13G3JC60BbKLKTgeqwXdvPNEzLFA0SAdpM4vegx2+qgWR5W2D1Gm67+4twNtsKZ
H5aYS4dq8aUlDUv0pF3mU8bVLhS3+xEgL2YSJz2K2bnI8voM71fNQedIxlNLaUB7PPfmzyax3Cnd
o05ZdxFzFwkgfrMPMhrEUSMl/N5ul53OzoDWD2g0iQRTS0rZuGVvdR/+UReYuHKZ84zaCrZrR6eq
H9EwL5Ono1QGIWQav8nc8/MeWGbvrsHTdsks5iuTachr9/YLQ7Yie50SRUwdno64s/qj308MFmiZ
tCtwsW+0kaYZOHHZhBUnT+draNANAOxKGN34wDqE05xd2HurQAGAGNoTm7yzuuH0jknGKkPfJCOm
OX3DCrYnb95dDHu/oJlmFj7m2pCMxeKXUrQ5s5MKfe0GpvQkIae/3rR13bpqDkVanxpz278hxx/A
9lKmoEQJ2R/b/zLZ4qS4hDC8u0dT7uXy+kKIjcGKoxlpGuL1o0aOoTxFfFUR+ISxbDvmNa5ANbt3
Ly/mvCnlf6BvU1uFcCJIJ25u0pkZXCsdr4HPIThdJVvK/MkejD62aSjBawEuwsYt1lBoEzSf3tFq
B0lQfvjoCepJXCqv1fxC52Q/xkppDX29enbX7OXE0iaJNEO5hGHrhNaToXauKiSjM5tHNUdf7K/u
DjAETdcs30TBTAcchQ5a0DgDAn61uj+XB6R9Qbz8BQOVPWzPwYvnMLRvmm83UIwdkFoc5qsTV8jh
anoh6ehC8zcmJKXSlT6aPuKkwJ2C4elVf1RFvVViZ8bjNXy9XynpBQArihNK9EKIluoUBTEzTpU+
+K4UixBbwzB5ow5NDIR7EPhd5l10t6+6Ozq5B61roy62iJuMI4+9c6tTVHHCxRGKW/tXdX9IZs9n
2zPteQeLKlDYFDjy58pfkGBNX63QVH5TnD6EAhbuUxyFZUyDjDgarK52h9J39yJNSO28iXz26+hf
38or32mgVy2/rqGRkephOlLZAz8VrPexxHGqzZyOX8GuUGspiSMrdnSkCp5GcXnYR+j15SQbQ7ug
ORd6T2XZIJ7LMJHIHAodazZWk856BFMddCldKqEmv7f8fUkQc/nE4lv7m3jiDDeEmhyS14ko1UKB
S0kJat3mCWzILS4g5ZJ9cvPJmJqkEGAeioym05zf0DlkRR3+YDp9Lj/cOVKUL+w00IrVb79RSCBx
FVpM9mUJJpMpaTRHl6EtJ4/PTWJ3aV8juxA8Kf19Aa5KUSksj9sDbACc+qvafQbUyHdeNO5NlHPA
KsM3e71PAJuxLkWvQQ7QdBNEJ/xhqLv1IYWlsqzKYDwZidExwFM9LOL0doxBSXqBsqoMBcctHnoB
4ZIyG8nmTyh59Pp9LWnoEuYAbbcmNX+auUKuk6mvxtSysG/a90X5QPJhfFYhDLokxDIcbTo7u8YV
8XdONP3n+SQoQDw3EBslulO+8OeHCS6fCixNrNOjfcL6sA3cUdXRVGogoUttmMCH2Cy2IasmMswB
D+W94IHlkcc1yHAD6vjOAjUebETPSKKhHj7fsNILyvyLQkozYroTwywAkkFk00IHzxwCl1W9rs7g
LGa28XrI2Xqde2Dg0azE4K7Hm03KjDJ7tOILD+bX1S7tUy39/1Izx81zvWLXPV63RW5Tm2n2Xtsp
5EZXSvVZgRlkiiV/W0SdjiBrJGI/W92ldm7UCiWtqKb5YYsnL03BYP39BJdcsOIy0oP0CvQDacyw
FBDcEi7XlGWt1JQAy4cCaTepXorICL1WyS07eszMPe/I6NyoUYcBxSiWVWQlfrZBIBQ1Rb44XaB1
bbF9iRb+AVLSj+W5JvMXhUw5fRS628LPOMcMjkDZ7Uc7G4S8W/FLJwNJc5u3k4f4tk1BIhY2ZHFF
Cd94TrM6qDgVQTANnL+WLoW0rsIL0bxUFNOhVNHc1kaLlhsUK9MEek4FLUJLVCPql/gPSRevUd10
ldX7hzusgwxDj+7GmlELlrdf9DqberspNjlCIlW11DUO1W9qyaIZJhDhADBzqVRPVfwOtuFnJoCP
B8nHHu377zUGBz5ftzqidDHy35L5wYXdO05HPgQdbBTFtGagkXjQevErA3u3Gy/gwDY2IpDCwXKD
RylN3jI7V3JZ2IWlPGy45L2LZ7Xw2AzXShWBPaLTC/2ZpBqQ26zbuBhYOmt0k5alhGwMEhQjMP/r
jChSwES7MAmlPAGSMunkKH+R6vY48MUNZmAlw1y5InfA2qlMRahqoI63YIhDIWBklwqQRaoSwpI8
ep404+y7rZdfsCxU8xeClE0tQM8Fk4+4vi5ypTRcMXQqCRQM57CapyQpvIyQNbjaSLDIRAB51dmO
9gxMz4rx0d6bB/1vZm8tVHyGS9ifmhPk94yFnKKZZYaqeWvzcH7WpzNT29h5tQhsawuP0NHw6zxo
L3VmfzPxkOYxq5O/UZ4RSCabW38MyQjKsNNJSTicTScnpBSAOCMsXX/EeBItqmbmDimz3HUH0F9E
82uBOphq9JfyLW6fXJtQTxGt85J7Wb+HtNQJIp3KpirkT001193lbss8c04EOUOF/1uH9R0eRDXD
gzQkAzhf6q4UL7ShPN2sjam99y4ZrzTsW/olA+Gqhhjn1ljUqMuUtTlzpksIagDPLS0FoRzGY+cJ
J2oP2Hh3pbDDqBtMIh74mf1AvSj0CcvUkjN5y5FnCEjI6vLA4HgozTgkYakeeTb/oOBiF0db9w4Z
Y+n1UNMonpoIbe/Wgv4suBTNWmjJAQXi2qOc5QTiF+uxD4s/u55ZETug6pe+BQBjeZvLHccFdJ1P
rhR60Xep/cjomGjSAfKZrKqGrrMEhO1NmpQOUNJ21MzDn5ef5/b83RQLIEFXK5GP0vE7aA9sKn2W
LEkxGeFA+txdOtZzoWm0jAe0vJX3PwCQ7DkVKFJFXb0RVW2qnhGqZRMY/mydqz7iLws0GYZo+2Y5
VQ2nKxdn4zbyy9VMRCjAX0n/zEjYKeS9MjCIoqntwwZK/Yyaj7GzGr9g+KXvuHyyfaVjQbOvy5SY
asNkZNpYTmGMZnK5atWIL9tlGysApC5T4dbnh9zbhxTfMheuEa9PmvVrtOGP3nrNIN5ABWlm10uZ
h+vdUWEpO3OXkE4MD+TuHGBOQFvEKSu+Xz/hVj3zmNlnLeT3SRm34dqWe0/G+Vpq6M8fVZQ7O3ju
kaqg6cGabXwiFQgcERT/ba6dWyeWye9n0bdu3OqWAWGLLw+mDSLLlIMDHwXRFKKoLlYh8jbSk/Mu
oqj9xG3ecRR9Wgxs74yxfT/rjIIZsdq5pO47j8oNDVctYlcMiVTsQ9mtr9nEUL7xq4n0L0Xm+nz9
bGPbSSlvvR3V2BAMx43sWm4tT02kJEz0zXTxtCJY0zMXhF2tcWU3XohwUvE6sEalYTVTxZExCAGc
tlSk0wvMx32jLSuGLQJ2fiwJXenQyLcbhCJzuBh7QQU/LKUDFOQ8lfShxR1Cd+ZmvF8PVK02BEGR
7i46dwu/6qBqOpIHWXrJMDj9D+yKmIbKVy9uKB65YXENWnxz8rjX3rDAz7hQYFC7+XMurjcg18S7
MGQcUhSDqfTham5lZXF3FfrPsdcyQkdOEFIEpJqNZBhFSnHNwIOxSGAV3Crsp2g3q7lXhCA4P8jO
XlzjPJzexxr+VXpnFXqK4/25PRRd6X0OrZt81KH/o4lqw8ssIL/NMf17hnpnIDcEYGvVREB/y1zR
W34SO6ZTrpbKl5IyMbJA69XjHsGUN27kWLNuMERZ4SRUaqgZ1cB15vRDOXgJSjUB2hIJKwYGYPA4
rQHgyaLSLjz91gvb6+ncZ4vD0cETvUbU1dGnNSMrfojlhw1J+h/XYdvzHAlt2lLzhiOehjseVryt
m3XGqv0sCNmXvlovB/Vv+1FAeAv75ql1BnjI+tbIIryNmcefoaH/zD13ofkL9RC+yNPIM7f+Wv7T
7Aoi0op49ALL7EsMR3tWhnYNFc79e89S3L1Fx+pbStL1H2gmA1VScGUxY/VVmNHRFFIubtqIhdD9
TcuOxf0wUs+a9jfCniwGjbebH55QTIJq9/02eqhJezHynfvLt1dEdw9uA+fQB1doM/TZ0z1WKOQG
VuQkVQ/sbapCz95gDmGNXiyyDdXOHth5yO4Sm+ZXt5kiJgbOnNi0MgwW+0pvqQloifj5ej1bYd5I
7O8ACKGajQRSHjiyZCX5ESblXj1L4LkRCpiaR8I69bcNXkAoszA69Jw6+Ofl1zzNyeI16CsM2Ju2
FAkdZqOMX55zXaoR8dZ02HFMF44yFNKzgy7YlXCJLw8XXOEl5Ig9VyzdLBBSeAH53Zs7RrvCUq4X
4Wk+tjpADSsqf0l6xZsq3MVrPKbSwC+0X2wOSuQgrUsjVaTtdzXUU0twU2+ym5XgRGa59JYuxKSK
1qBoE7urZpeUyEkJP9bciue/VyZSlQLnnikRdRHNUeCk5GVfmy1XlCxLstfGZsB3/BLRfrdUvqRE
buOPq9kfuNkL1uSNX/0v/Hv5G+EpF+mCFVCmLwjMqMokT6cT7prOH2xBbdDGfAZ4gpdr/ARTcT+x
E4ufJSoQ8lGj5lgvuBC6QEvQkFgD93RvbG9SH9iG8R4qCKHb0m39KgMuewWTjptdabHFI6gh/Uay
uO6Z/th5wofNYWY54nOZggNuou3wtTQsa4yhahNs1GCcXx8bRZfQ84FzVvhCV1R3OjatAJMphBsa
2wvGHVPyUjJDwt81f8U1icB81/3yVAvhmBB2NrB9yL7zJo34kDK4VJRbPh1CYuQnt5PxEwgZZBWZ
Od4E2m/dwLV1A/MClw26wNnmiik6f14KyNHQGGMBu8hPmLDDTMkeZukeeIog3j91b4qx9Qg+dI4v
KVQi9xv5V9Hr3boU97zlwxsAJXhDjS1BbWWzIHmfJmmXK24nwBLxdc94NGmM1Ein9p9AeteiaM3R
4xbiFgQvpO0b8zwTYYGsFCJpZim02ejlQT4qHwRWk8Hj5Fq62oIEIs9nVhdaThG1vLX60kdaB4Mk
z2GXM980fZXWOVSQlf/ELUMJk1ivHyPhv0km2m/nyU1+MV1cUPfgVFkiCAo3L340YPvDwGoe8wDw
Y6F+NRKX5fiO+thj6+DlNTMQbPJaSo2fBXf3kkr4qUHR+4fxWwZJawDP6wdZT5g6rjNdqrde760t
sk8P9rUyZBe27gfEr1usapv/HFAjR/AhPSt42Zm76HHUGA3j6n5CpdlZ6HK+AkR2qakyk4GWK5MU
+jpYt6exQFN3J8IH2lMVDQC9iQcRmXXFjlvAOX8jPk7mggmSWSNfXdABbnXM1FBcAestkYahiNbn
VFJrN4kOCIdVFywXzfbjJNn5uam4qEW+ZoF0im0/9YDjW1JV2De/rFP2bNgZeu6mUehaP5KeIni3
3yHRbA+XWZLeUmlFe50+gZhN5Mcg8CVS72rRs+XRjKROm/J5nTxwWZ1C25c3z5bx42/yTWoDAo7h
14GU4hnk33yLX10tM29pLzvQXDqHyzL7tPAr+8VKfqMF0bHALAHhkAkJRyXLaF9282PExnTgvFKE
A1GkkoBM3r8JuYshHjciVjVTzdtZlboUqter4+5P+od0OxzU1cwtg6rpIjMbntXNjAem24q/aCu6
mNgOH49MGa9sihX7dwHbMGX4C4qXL9FRy/dLdfTL1CWTwoZ0ELxHDZk8gBbfWtscV44LGNfPnvHC
GZxpsjIfXWN6XOhqLUBK4Tg6m5LIYGlLtZvntsVDg0wsTBkp86MpbFsTN6rwQroojQFutZ9QMv5w
zCoKabGcAVsczC6srqXxGl3S5dsZlr2iT6/tXyIHaPUToo1AadeitMg2181irefZ6XQIF0P4FyEp
n/NFrM1nUpBJqVTauNW6M1p5IwOEAQWgMWsLnm00EFHKCaDboo5doH/39cCFWEqSZiWHzOe9ew9R
tojsM6X84Hcxd9/greo9CvrcqObrabEHUE551pDJhAfHu+ZjBjxuBaTCALzaUsf36MZs4ISbevcc
41vnXyNUpAaN6a8CI4FfSCnLJvQghQZJm/broXHEAYfke2MOn52MM38uuNxw139YkjxWYt0IPhhw
pIteCtTfG/o/QzMtNXXIzyt1gIGGp5UfhJq4+lmtru7P6M9tcD6XmoW31SanNi8V8iuchfiLTPRI
mC7+EuSSQ3irhM0JRo5hDe1UUq+pWU7xVAKWVJliC05VUPpa5UxkJ6vS73NYDgFDs5muK2qFJJGG
el6YEyRGoXLe4/fp7uYxYT41e4bWZHK8fkHksHpQ92tE2QdcnD2J7TiPr0zO4mRDReWJ2WUKILIz
DwcmeEpzIXNW/a7LJR4xqUzhSlas5FrCab1iOhuzOllHPOpEI8OGwxt1VsXvXr9T/FR8qooS30kZ
UQxiwHf6pFM16VgrBshQbRjeC/uq2Xt5r33oWTb5ntByecRMS5TsEKFZreBFLYvh3nCU15tvWek9
+qw4yqUOxruHd/9kQ1dJ46FFNwVnJXZsgiK/eg+1y/8mi8/jsBJdQVdAzSiNReBBQI1DcHDzxr8G
DUbAe42sdm73w0GznmQ8J3Gxdc9yVNNQwikuv+w346OKvNf1FXHOKunqecir6TDKtmY4m2F0tXAZ
CxGC7cbSnUKYY47Pz45TP3XhJiKo6LaWQRoNvX12hAQlGhzxSCMHSY0FYoDIQT6sVHEYb0DM6xLP
AtmA3QJ0xPz8sDHtNNMQnj8z36sbJQ5JTczWsKaAKXU7/yEPZ8dp701LnVqSzSv7sRK7LSCmB2xR
nMiHY/vCjXjF/rE1R5Pr3z7k2kZcBS7hAtJiY9xfB/xju85PPTfNNq2mGuDyOmkXaxierwyvtLDn
oO+ssm8zxKBi1utiHYyo5VnCkzHhPXX7OKL6kc6w6i8Z0rP1CYufJBajrMTGvruY2yyTyW/HQGGp
+lEGHM/wznqjSYJUfPCLAF94HnYIUF1H59gZUo/6g1URkdT5kMg9LJREpPExHslKGIoI+vwUqmY9
lPVScfObAlQplj+wI84QXT6u+VfJYW+oawfpp64FWk5a4/tf31sOVynQ/86DRn5ivP9RCIVVRbzj
ka2LpyufJaZ4PZ2jFZm9n0Y956BZ3Zu7SvNbnZVElPt/mhvADjZkh3lHuH7U+P1VifYJaIXb8LDy
uMPGDjvEP4KWllE+D4alpOu5O34ahtMB16swQoYxciW7yPUYfCidNhFv5qLiO920RhaSdcU15Eph
E/mVOwaGfjfjypYA6asVM1ZLRkCFnN06C4TCM3ZPypycBv45c/IvOjzyv2MwKGcuyxM1LnzMCL98
pZ+j7ZlV1tQk83TEewudVdhhh7rZKureOD+9QeHfp+QKXoJ7vcCalKbiFS83xyY7rcP6AGlA9WoF
scYZnFXvG7OpJgEsOAIUV+UL7JVh+Ju1P83HEreTw387apifX+HlWNbDARFEQuQBS7mCOO0Hu/DK
p2vQtB2LyK90+iriUifle3dQDbS/GZjZzcF+ppqXBJsjD11BRvRNoz9tkRpkG8QgXh9OQZexqrlc
S1O3DVrvzBnOVI07/cGRiu7cYQG0OUMs9VoWODex5cw74R/jxhYnwiBIItzv5Bci7f7Tz9mS3MjH
E5m4ayKMM04Yh1p6BhVedvp9AjWVzUlU5LiLW+280jDFlrTai8i2t4XZmAYl3vhM/SjTyTMvaHH8
CdQQfUcTIxpuwocozi+Nn6djCESkTiRjysjMgF9NUPg3rAxgdFieuFtI7dK+GtPBtpqGpexATNQf
8i/oq1ZJ8y+v4fMJ9NzClLlz4CkXTg3NwcprZveJJ94bfC+LwQJpGuyQKZg/wtWVQLJFkAEL4RDz
4upLEzALvbUkIyVVSsmGUMbNVqoFPryjqXM3BEybsk/OWps1hcxtp7Ixm9Jx0AJaXWswDJPC430F
FPwfRTA4XfD4F3YEwHIBeCn3YUE2qf0Fp/RG/H3+Dec9Yqk/E8zF8iNO0kdIxYwwChk3f+ZH1bf+
nd0nhsOK+n9nBZe4F+uGWYesq8flXC+JnEOtcxVx+oHHfzZGzPzse6bQz9TDLcin0R9njUQpbU5S
Z/l8VDJYVQ9RAGGW774UjdSJl50J75sVKdF0Qr5qlHjVA/jLeRYA9SQCiBemU98A1qHL+8kixfNR
SOO4dsBxFoI4ZbCz5WsOJ+KRG4voEqLk2dvBtYrbXckzYarD0LYbJOZ35YzjwUaYIcbGSPXormlT
jhwYmdDS+NCy7iuZDdTIGoqew7rmum8Jone4RTFHeZ0qzhtF/xqRrHxwTOkPYWDlscHBDqxnkkNg
YujB0eX1iNPfZE34P32FzhqTVpCCDsrm1yR1Nv9f3SHotjDoX34BpoVn1+ilgnQx3D17hsEyxiQ2
ieUo5NFbNvPwUneN0ZkOG9ajXqL4/L5llcBJsCLXU3KV6KHOLTULMnO6FYDZc+PeTzqC99uHJpGY
eyTSdctkebWo2NDGZp5Gzn5/DFgNoCJa1BzxRUjmAAylMvH42LAboKV7BTLp04xrZf++zTO0CjE/
Q2w9plOfq7Uk2TZg4Lu2U+TB8bHk4SEitIfXoOsFTwKtCHOcwmgqo0EAM/K2QRxVjhA117oTJVcu
19BUmCLnvtRZOT+rGBO1ycezwJxKtHXzon8TT//APo1EBYNvCPeDXBFh6XvQ/EqbpLmCZ3VirI4r
2cKTs5gw48Qxut3wpmQHA3uSwUzA9XwDKYf65X+9PSZK/s3VNgc3P45FblAy2yDR9oCdiSgeNZP7
0VNonR0elyfxXbKaenOZt/ecb8fAzHgZACt7CDoK46MpvJaHzke7mKFhzd+wgqSHLUkuTK1YSSMq
MLOX4f2aNJKzpV/e9KqQAlvZVyil40feqlVBRdZpZnwKLhchT5fNwpE5Tg6V0up4dSg9y3Oh+L1j
7OvZhJQFRzMRPsMPyZaNX5BIGvNQQ4ANkV2krOWlV+8hV0yXSmigm2gwEW7AMq1x3B1tr8NP9rrn
Q3zKC2f/UzCycq6sCu8UJKY6Va8eCq8Kg0nAxxkXpwDQUdA/ikZyYmM4PU20xBziPgsQxb58w+HA
nViZHkbgvlKqQbYopJtdjUAXkmHfOn2HY03AFrKVBRdTXWdKnVyTJwWBPmN4cN2pM3DiRVhbsgR3
CFhFymr0wcMdMpDo6Ine+aY0IDRZ+RX+2jAox3crk26D6WONuNFJZOHB/TUm2/lMQOG+Qw7UlAuh
B00IDhMSvCzoziQGpncKTEg8mSjDGEi/TqHcijz7hcgAaT9mp3g7DU4C8MGH5K3BtXDNARYJOh/s
lizB8ol2wUQ1V2G4WoBNQwLqlFXSxvTM3gTr9Gl1dbiYTnILBTdgToCQIaAgM2LHhBeYme5hKyPn
g2VS6ZXfnuyjELqQPK1GROIfCPteJM0r9iXx5lQRTmc8uotwmgP7/IeF/pKfyEtlg9IDbhfvIZbW
MD2mk6C3b0Qv5MP0jLaT4dDB17UOK8aJh34PYlCYnYuGVdHf2mH57KQWAO8kZHGAH47pOWeQLgZc
kLlGVx3XjpyVzPFEJgLUO2loIKg7z0JxCLOlwNc9wCHQGFYn42unIpxpauXLnxORQ9FrVFwLakLD
r/yetWF0I53sfTHGPCXIwY5jUB8oXRZEF1ZOl+tzxANL3ecmmJrD5RDFIYjYTm2vBt2gJU4GsGAW
RlvJ4YaDPCuYbc632ADlzDk39Tlwubd8qfhk0FxjkbJ59BIjU5A61z6bjDCJ4OHiILrMtaH3PY/7
6gMmGlMoNqKC2gwW7DJ3J1d8aZFy5gzhNmeiqZQ5cD5k/vfWK9kzUQ6VPSYrl8PL5HAdG2VwMmGE
/UOhjNm8X/ooo04xLN/mQQWwu1UmJvrjGjhm6EWS1RKA0G1LyS99lHMZMiHE2TrIdl9Xhcd35xiO
4k+lERJfFe0kSN0jULw/9+rTiCn50C50QaDLmUFnI0CRHiviJb8nSSygfkWp/fSS5b6FmUuACHRc
QH2wTITmNwR0rhOlaTwTtkWyzgFagcrvDoTWwsTOQC6NeifjaOwlj0niSvlvrHWclpl4nmcKI2fz
YGElmZDKMSf2pej4JraiHpAX0Fxo807C4t59l+74bvl9LjHsvd9SD3Cuk851aA9eXOgSJUxkiZZc
cnsgIOx/vOCRmVWuPoySJ+jzfpdNLpkq1M56C6I8tBmpJAKZkEivrEXIre77nVt6JKMemoZAgvSB
iptbp612U5WlZeJGKR0zVafSLIW7OxOH21zlr89NezGMMRxbWufJWe2DRrHXwD5ewRuozcwGnK+I
0Es59j/1GKtSwwzwtBqMd1bSngLbsW7dIYX83dxmG6ct/klTe5x8+TUyNpxpCbTDU7g9O5IhPW5f
OEHilp/tqk89YWHRt8rFuDaQpZn6uIE9pkON1P3nEN8Kz+fGdRfDsmmWlY1JGnRd/Y6qnEYmMHTU
4nIq31Xe1v6ha4NV2teQVNds1MJCiCDmHmRHp60YnOlo7Ar/TGv9DpI3XxN4KZgF5poLkUBSaOV3
u4EZHE2ER3b85TZNxiPtkhHVCIVcG7U1iuuNUL2QOhdavEzEnMV//0yrFGaRTddslvooi7Kbl3mx
amIf0MD+oKMWfweSLGEyKdxPNvRD6Y9p0RrmOnOURAD1KTVzwiJvec0y0JEBU+H26CAy1XaMmN2Y
lUQuitd4oevOMsZJgLCCH9jOjK7xM9ZDH4cGsk8LG3RnNPtUp48v8kClr3XfPFeQmHXyE8ZEDScD
g312aP2b7AvMpcHAw4y7Sw3jTxPQBECs8gCJKl5rdVojroeXPtO49jzoZ5Mh9kIZPB+9bw2w1wP7
DT+uWB9MHiY1rP0SOsXJrGU0VM1JlRpC9NY4zDohl+eTHUS4Q0cEYJnMyB2il5Sw4X5T8jDzmGnK
Y/s97uEipEA3UCgkTh5rFaP1aQeNQyZsxEOwbLPk3qSvj9j/Nofb5jUb6OeZ+RNm6TDBDzXuVQ/5
CT1yMcyRfTw7RDnhGrEOY68juu0Vr9DSozDLz3qvgTgRHWBaWD/eMoOTrg18Sy1SN4KmFYlhoRol
M0i5vmm94pQvMW2QYCICk9JG3diop2xlTLNotlIJb+P7a+V/il6BqZ487CuC/hDAYl9pKIdMLxnh
Du2kwLPxF268T85kLw1fHRdO83VEsYFYHmok4QQZZoDylq5+vhPXTjQoA2svdBAU4V3LHJ6xgGY9
8RR76SxvbnVHCMTVTcvq9Kt5Uuo0F8w3gyybCHesVMp0Yq3tYAuWw0ct1JUpSwdYVoPCbpx0o2ue
BobRjfgPrxixV7xTN4ndP/P96ZItwZGTuVkqIO5Ikua6u8ZRh7UabPEZHy6s4a/d5+Yrn7xAvbEj
6k7YWzClYIGXLKjD21GO3EQhho/iqyQUXbwPHIgTfFb66uK1eVfrG4pbNoQHLn6Qk5/FR6bvs+U5
XmVJlvbRu52LJU93WR0O5ckY3ZW9G0JPnlZor5s/NyA2bkS/cXaMDNiX+pmUHQbd5HFE1+CLsfm3
YUiXi08A+QrYQm2gWhGAb4j0tgetnbSXseTVNy5lfFd49w0+Xupmt8B3olj3to7FcbGKacXF6VBO
s9YZiR5AVf8MgO61bRn4BHHRkBcLa7+iLT4SQ4EG3MWUf6/9sJq2nOUhX8oOhIZSIfi/Bvki6ruc
FaR4/C5RcEOcB53zTwCmV+uF7tIS5zL8PZD+lDl7CUOem4ua+dklNE0t0XZN4UGrCvnymuRVT+RL
IP2sTeOLOBd1mrFD/QhsCbrP2D/Rui4uBJpbu4Y6lBZuY5Cu1W6ij8z+9FHs16AfApP6f6yAMwlH
79qq3tb+DzbdmmWDHkk7ty1GHKJZToGPGUscH+a/gPI+l+paAUAhAkVNq5stw77ZfTErRGG6OSgF
75YUsjHUfwwe97p4TPeS6xLxBOm/eAwgkg29pWI6Kvzc/tkO8SVZMIUCpfP7WAoZxYrR6tnIlpO3
czPiddhhyE3bLggbWAOEBevGHG1ehAHcrBYC0Vm1+IeaJSK4cvZcbdP9QsaocckFlUOQ4nxwbQNi
dKp4TgF/MkeqWR3uTvtvp94V1GAoa18WuW8aAgPUUtI4XQsGSQJP8n/qox6bJ39QtuqB887l9ZtJ
h9iaYoY/xv2mNNT5gs4RaBQO72DSGBcaD0P7em8y8xQ8Hl+pGQX0Or6NO6vFM4rySj18QSLuS4TG
5Tii1oRN6FPk6oiqRqZk7uJMhrfBPbVoaV5kujhl8bK7DhQsCqQt79QPk6qRo8E7Q+qPAoObhaX+
kaYoPnDM4eOyrPtqmpA1FFOVjkIB6j7wOxyTS8jitY7NibHxtma2IJePFqeQc1m3piNUlAm2E8J1
E98VXNdUN/SJzikWZO7EYubA5KbAbsG9ToNf5P31NEhM0XPm9VzT8u/8kCNEp5wwjua6p3eI2g3v
O7J0O14bBTekwWsFHef4uGUjeOtdReTze/nfqZ4q3kuBRq2J/n+v7IQbxZS1S+xcIjDyoNgjuP3G
uPCsYgaYFsNZF5w2OrR/hRbRS9imsQZ+PeapEMwhCuZjA/0isFHzkc36QLahSbZg8Kjj1uY+Jgib
kUaldBEKhySHx50+GsEqJ/KrhqgQeTL7/YAw+JR7vkRRQj9GsKs7yRzX1AP+WJSaNsOJE8M4IlWt
rmKWfbChYbnvXdREd6+UOgX2HmwViCUdEuHPGBriFWotZ/2sujzuRs0KuWqmQDvLza9USI+lmlFX
I8RrqJCLf5QF/LO3wSPMyQ+PzT5kGNUJC1DzPIyeQpEH+2TrayIDcSAOjQ1m/EpaSyKoZZTp3ARJ
/oZ4xeFTHa0fYYkPnzJ402AJ1VjqVIWtvvqsk6KSCENgWRAx3w3LPMvFKYcMVcFAKghuPOfpJDKu
FzQ+UoVvqGKL/AC91mAbC34OQwiL1ZqpwyiIHBL+zqehzd46zU7KdK/XpGNbbEEJRh0d8+WdrGs9
2jYAp1K6ZfYOY29Ey2nKEvUrBCZfc4N30zUN7qHa533+4hB50ZfoNpNJ1qhHXyO5meGXErTe6SUJ
ERsN4FUiJw09FBfgbq4OumleYO2Hpuweg4aVXokpGKeOsOZP7GozCqbEXoVusebnfacvzehAUqK+
7j1FNlC8JSBg5srHD5m6AyC7gIKckNcDLl0uAbnZQxcVa7Amy4G6hdpMvAHV8Ilislouboiviccp
4Y73ApqxLvVYUAlX945jRt1VUBIQbsjIutw7PFE8bP2QY7iiHuFcGhf0ozdKRexz/EHMMDPGtfH3
K7r6Aey0oVo5AhhIY4pYCekzf6Zva2R4aOQFWZgV4OVlLIyvKl3Xg59atnskqguosKYnImutZFNd
4Ys6KZU33+wcyuY8DihjzH7vUDAbh55Z0r5ZHIq737Bx9+bdgD0k1UiwCDrW1A7tD+kEq6zYjf6Y
bA9FlEleFCxTLXhl4Tar+17Gdq2jqiUWA402tmGeTUS3QpLQRyEStKWuAKGlKZ2b0tuI7zHfLODz
jO4npK1nCpv/W1CtQIT7sR0i78MtUUiaYQ/glFRz9XoXgEBxn+avvAwpCpNXnTsFx4+HLFabLT7B
Cs1qIVsoN9LNoNFTbucqSvPqaTmYjXKl8kgPHDe7Yec5dtEHfdDtsOx537VkVEpDh57Lj5rvP7l5
93EuRj6V59lV3etM40ve3cSRfckbu/HFu3k7O3CQik0UZ16S78e2ShInq0aPHvnlRMxYIC3PlbYQ
u+benXP5B99drSezpWtAA4yTZR849Td9RiMENivsQozBd8VD6IBuzo+pJxdKmSNKJUvPDRc+JZnG
yX/zqCguyd72SaBV+5cWFCR4iqFqTmKuOUswy8BEHJyU5uyfjdMpaZIIma/KPIC9G4uNfMYKhrnd
EcmbCX3DmU9K1RawXhLurVDJ0CqZyAuAsVB/EL2FDRzugW8dnwfcWaaxOmZDd+Z3Bc/ymLFcM7Yd
5DIPltAN59ALUD8/frMcTAL1yQVfHc/spA1ucaNzV9yIAoDQ+OGVQKlICZUNInW9MjwfXliefIgJ
pRgUcFcsMBN2cQSeY2bWY5nIObvXbJ3xTuf7eWZzjdz4AIuiwrU+irksIbZdOQUV8X1LnZQWASmE
42FdgXadKd9aN6E9yd4NVL2Y6fDKZHXfSLaSYZ9Mtq5EPIVyxYJ2SFwk9XG/VuvDP3EwrPIQ/yxQ
HCUp1xDp+8c8NkTRDEUSQzH0XmzxtNP/RcDNt0BHhG86T6AzYWoUzip7LDHx9yozo01CT3KYwPkV
mPHsf0M0Yjlx8+REERgSev+s2vfpfvd7oNofw+GENEQCQGDc1h/VZAO8e6Ks7QORPuTWTgabk5Fe
dpRoUT7kEvMDNo3ilSaF9zbcNFDrhTYtTjaZtKEL4GVD9Q4alqlHM5w+n8fq2W07pJCUvWdMfB83
Ru5/etfgQ4qKcB0c58lTy+jxYqsCLOMb8eJPMymHLMBx3DfBReX57CuunCtfJSJgXpt8Xo9YXxiR
xu6OcGIbi2vP3B8i11W1l/XOR2ebhxibkpxungfDFiyBhoCr8zyttuuarKiFq2OmABV4YJzdSDmV
+RGpr3mFiMrRbNhWpjcriUKQBHkNlQqXbNMyj7E11NCZHVi0gJ/YBEQ12ORnXKlyjkhQBKK7RtM1
IWtaPZ0mzf5tb9AJfSSBSUgK0uLmKbSrS+7G9fA/qwAW4K6O5VR/BEJXqpAOo49DcGQTlLmUcZ/7
2OHR6jPJOeVhnvOUzod38jYQivskibf5SsaBXFZBU9RhLtF6ctHU4l6dH2H2fWDVNpkuOwYlyUbq
Yj9HmparmzyuXJJNLvIbVO3DZcKeWcNuIiCzunqGtz5awL4Ndq/k7P8PAh0KkwnYY64+tee7quTN
2w/TrW56wiEyBtR/HaSDThH/iCoK6V/3YBBRKBKfCtLIJQy8BTKL8xz6moiTYeecGL50bYAEOYnO
ULONO+len619CV7jsXOcBWQo16ZOdioxpO/0iJY488ZIXAI+vWSZzziryjjY7/XgJ0vQ1by8p/6X
366ETF95sj8YOiRpTUPp1hfgORbdIg8MIb0a5QLNse5XKVcoLTFteVnB2SZIjT8VIovF5QfSJrIU
sT1TJ8R3RCpBvRGLp02gp0Mpd5fh73bA7Wbq+hHl2kl/mw6CrJM+pwjdMPt5ZuuSHpxNtekPbt22
cqLtloWgXFDvo8006o3DLPUYaV2LVrSva6z+VCOhaaz801Q7upvHa1ISF9eZqN6Zvco1J+V2FU83
q7n5FMRPP2Ky2VSGQiXM1ZCkzcrxgC3xRO7vYNjmlZrAb/L9a7ZH7p2Ko2dYgLNJweAYZHzC+g06
LEQS43+bzMei2a4Eby8x1ALGT6RTji9Epgz0UWUNjQ4YTDfQj9kG5OZcwfJSoDgGaU8RUB/ivck1
eSTm5EfKVn7qZ+2RjIeTpQITyAn46Klg4FTYPKAJieeaqGoQQaeUhnsyUh+O1qEiLmaQbXnwS7ty
ehP3iJ00w9VSnYJN9Gs/EE2aAHHgsY3/7xY/pSUcfL9+5hsXY26xazZ1oEIBvl8jDS4LPMBnKv49
WEyciGrtKHFs4iNFEzYc+RXY1YGTqGvBBJCCVpJH13nzkxbZKfnUUcxB+cLVNW10KdqYtu6t9BXK
0LHxDdGgX72F4DDHXNVpzjFkgO4b1VsWhHdjMaNYD3xUyYVLpFJbtomqXlLcUcDzGgsOJOWYoLvw
R/zwmrdl0ZLDgxzLoNCrHLDk2wUTf0i2kysL9afCJzqbO/vEeNlEZuyhREQnq9C39JDtbLqXuy7q
8Ei35OQ1a/wuXrjLOa7txV+I2evzApwwKbUZMetj9XCCJ10m+oUFpxFmtC88AW9Y05v8vvPNhXNY
HWK2Gvj049V30ZQGm9h+ngcgVK2ew6DQ4Rx38JtdKGQ6+Z9VKVeuN3kcNIPDZhsIKIEO/xF+V1pC
KG58spx2Ouy9KXqFlvONcdvDYAzjeu92CjTIAvePFb2aQMXG9AS8TdZD8OpUdQX+7jZmanDyYyUE
znAIHJFiCmWER6iUt+hgJPRA1nhjLFKRbd/vntObLCsmDNFLhAVfvYYIfGWc5JTV8LRjgVulKZd9
UfVAfVcNONxXc+HTeJSYSN6uaevck/2AV+3oGLPyt+qlO8XZCU/4KA1sL83NyHy3EW55hHCtmWep
I8G2Cc20gDGz6t+9pOreHAbow85d1iXLXtMYtkVmrt2/hD5duNhGq2QdyH5mzcu/BX52yPL9UpvU
1ZMytAZBFWqtQ5TyZ/jde3BD2g18Xu+hrm/xCmDT5rckXoPXT8HKEYXjujgowHqLlfGwduCVFNDH
H21Z1P94mSmGBUx4L0B8pgahLxY1Ji520dMSgNF+w9u8I3C7wbqBegTXLwqL8pH4iBADbRZgFX7K
jBT9EEiypoLxEi8D0crFRiZw5TJr38+iNHTBfC9B83KGo4lU9MpKdzo4Zop17aHIfnUzMkHdgFGw
ZaLTT13xBWTDAUmIFfVi39JB44s0BntiPaqas4dPQh9f2U2zy6oa10fU5n0jqSA1Aje9S1GfgIkK
Qkl1YZP/6hwB/K8LCaTz89TNApKLtSl3m/Samg6xLcwpBwv4hk8r64KCza5RMFIoBVnQmHtAwjKl
KMe150fliBfeMAgwqXn256QgJ0hxgOwxy88WtX2td4T5eJWpo3d+25iZcth17gAkkIx2Zx8q+Q80
ehdg0KAXKDLLTOa4hLN5u4Ob+XnhbiHWZ9kVsQ93Zpk0FezWlPq+XAphkpQ2xIXzHzSylVSqkPsI
CPxlXCKxqmIw9khG/9E/ylH+s4EGOBlureS54dNDxmzLmumXn4HsxzwrfPMPyM45g7b9onMZ6eEG
orNfRYVePtGga+bYIVX6GEyjOc0CFrEkfCvnTq36dom9zah7nqufDnA/64/8BNmQ3WZdaYmfJmmd
KfogZ4Yk/hUABtfFw+YDmQRscu8vxOWlQEVFPTihVM9vriC/48gs4WA6jTXHQ+Abl2T4di5UVNOW
N9UgojMq97Sqrp+woDPGUFgBRAuPG6gA8+KuXLNeYSQyswREvgZJ4DebMhnnotz5UDYx6yinYggb
bzFRh8w7FvRKXDgXA8NnNJHMF+GhVwZ2UFdgIzvFdgV8HIQkj0WCGz6H9DiHY/8TPVambsj4hDrj
xe+R8NsHg24ZDlZ/MJvz+zHdSXAUHTUllVCdWbDVDJFm/tPuuzN5xCAurD92i68kIyVrRBTemzmX
UJT8logzZ0ajLCFERZA4jIQgG0bdGOFm/DBJG3F/FNR9KqWEZ58L0D+kvJiKtn89NmFwqCUHlZNI
zhyTYnG5HH/oxO3zKSeH59NDdy0NtRxMlC29lQX46xLEJZ2AgV8i+haXSIj5QoHXIMyWUCQVy8wE
bSGBCX1ObW3oWnKDHizTHwzL2KCQCnHjwVQdJ2CCuQRTpn/tVFsKyDaDmPVilaEDyS+DnvF614OM
gYKm5MjbCr8EltA2ahAVhO6wM6XG3hnDGYc2PNyJtOZHxIjwjU83Z2T3AFNrrlOz7dT8ur4DOTus
OT984K/6Gi1HmIbH9czCfCj77koPAJfmiJOn2Jq8j0BkZ5ios0cJ3cUY0+16AgNrEnrC2/VRziV3
CmL0Wu9EYdkuomyWG2EXjFVNS8KelQ5HAysrDq1HaWUuvP8m28I5vPQjUfGJV9A4RX/RtbVvcr9n
aozHcz1zTeBIgecuCmqQuUW1nJu8Jcs8Lgq3ykCeNCh0rQvWLBqAeTI/dxYjk2vuDR0ry0gJxG6U
FXuYvoLIsPZbze2Cm2LFWySWylCjQFOO/VkKOHfTR+rYWsTouMiDZrHg6JOmMeezDp2GEwvfOZrP
Nb19uQDh29ldUr/MlrlKkBqjLKgb1d/ODniaw4bYGpGdypjpgc0DSScU6u8PqoUQqsHXD2HDgqUa
rW1K7oCsi24w6v0YpmSPBSc2Jduwnr56Lplc1yNSLlXjuLtuwcFQaHnNQeTycvNrSerc4ZtMUWsL
SjGUG6Eif6qTw1LDQhtz+wGQ9ahcGZGDC1ebKffiJhH23y15eVy0Fm966WhwVmDxhwsN18qnpP+m
uL8YjEc0RD+nFST/OavFVqWAnuwZYl6KZXK0GOp59rXsBIq4iZZUJ9zbw066YUi7cg79yOpqcbkz
f7hOvMEF62Ro3WLe2e9jUFoV7HD6dsvdikOeBw5HX2Ul62qDIFg9xfBnWIktsNQCcEfnpS/R9VQK
Cy8YWEzVaHf5qVtmdEZ13rJtY/1mPzyiuL+ighymrG0CX+tYwaimzx4oNuNUeYeRh2J9jSiWrCNC
95Qs1h7pE/eIRvSdZnUDQyVksv/KWr86Ncpkgth4JJKgeVFAwOUEoV+jRvESlKMsPH4J+M47rgPQ
2d/1jQtLiuMS2PDNjvGqmfF10TqCH4cPSpVCMEv1wtf1jIT2UEO0sx0coZh5xui7eP7pU4Y9PkSI
ad1Z+i3m3nUf9TLWuTH4yF5fR559Kemu275vRj002bdcQCKPSp3VUp84fT9T30aost/4aNEB3qb/
hKeSal1c6w4a0mbPjMTeN6SwciHJhNFDv1zS7ZBcBmagvBUNy3hjxmJZhp+BGnUw2LTkAD/J0nBN
SSyv89lUe+FmGrXuDNgFr5VElGb4a5V/XczYjRTst5C+BpDS5kXnTgcdA3+AcdlIpxkR6gWADxYG
nvsKiRn4KkGLQkd34zqOsI6UJu+ApGIBAvZcnG6E9knkhhFcceqr6LPguvOSSfxjozdGCYeCHwyN
er5IV679uM9hN6OZ0qXxtUIv/+kdfvx11BAw5t3g7IE8GcIceC8Evl4RjieXnEVojbhKQD9CTfXf
9q3i6jeRkMP258k7HpGOLi1l60gBHYpuRa3amqu0k62tlJH0wQ8khJTqfVYWaA5LMtzv2ewbYS/h
t1SVdfmXoFVOaq3cQczawBhj/NJa8YJx4hxh4FCIRRX4M5ip2UPGNX5cF/n9NE5bgRhRoAqwEzBh
ktpx4hW/dX8Dytzc8s3hinRVDNF1nWHO9XOCqCBj5GGXo7R7T954VVf54zG6QHU3o9mHyaMoq6dd
DQtQ5vaMUps/G3lILDusztOgApejiDuGyDKEfog0HcUgQPqOxmr5hHJjN4yQr1AkD/GWvqgW6N5b
jupRxUgGSildjNAHfgt0OpuWKZNpP8KpLLx8TWGZzXzlIASQYtSxsEo2FZ9+Gc+yP1c8PVrq0ELz
xObK8R+bkoEjmD9WjzVvYelLykivRT5/qvsz8n1zkECFTxcwF6u+s02NwiJLvhdyY6e0XfVSJDSm
WnkQXGf1mTOH4GVDdFVgZDmh86bKxNlecazC1Ynbrmu1fM/eS+diKBwHSZGSfDfeDChzvtYV0spp
vIois4IXs0zhHaq8xmGvoh62aL/CG53i/7b5zBmUVfm3UvKDDvqOY95QNGd1tudFfQh0Me7dQbLu
tUqY+0Xntz4SV04NkAJLKa4vCJCULwyYHufhBIIEkJRtoYoiJLcIU1tCD8VqgPnhylSLyX99P2LY
sXEziggdrddjKtPoyuX98r4ReEmGhPbfjEy3+4zdxtkoKWxQdkB7Twryh8VdmSLBrs3oJH4EYTmi
ZbR97KgubOyRiAlbcJkHe6+YHg6OmlZVlLX3TupnsEJ/HtGAAUinmajGwOkr8gayBPZA3dIqlwaO
C4Xl17Vwuio3xWzPpFEW/bV/cT/mrYjUinGD4tnI7UrzqF9v5De90Pw4E0yQwM5ODbdANUH6gvWN
rifhhutCJ+7epK3iGVoYpmm3LbScIZ+7UK+kpeCVkU9zneAnrQgcWhloBGriN+8b4eXUsjqdec8E
ueKTwyGR0oO4ug8vdVz6ZLCrBJNyM6c+yMyk9IPW21KTBm6ukBmpwUQ6c9tAex1+XgV2S7ly2tai
n4Y7KvKP94FMR7f0grO/+1eSARNUiANsGC0JNy8Htpyq7mnt+xTiKedheCHT1caN/n+MCs/znhU1
eSdqN2YRb6SLaDU6CiCm1MB7B4Rn28kmp4DNUDIbxD2S3WeaoBooosSyzxXz/6mpGpLOVyhVWMOD
YyGW8MSKg9Tdqx66NbepXJbpxUHC0OpCgk778U7DncH7FAzG/MJqVt48iyuZC8eTHUA8Y6VYc+kw
KgAQaHrarHJ3RwUZpIhqIu4yiEIoe89ek1/uDJXTvT9Vral9aIxzrWubdRPMkndlgvf1x4eRe/Ka
EINwo19b9u/eUJoa9QbXphyvIubdGZFgzoLuQ4iT4xKvdSTBoDilDEdlZVgj2Lx/2QzIwhmu3dIa
P8JAy80ccInVPHgF0gcA8uh9AINmg9ZDfvr8CGdKxnGoBJt0r5tv3YzxiY0aq6T+NIWJKEYS5Hul
A6Kq7Vyc9Tss6kASUx+Ea38byAIhVdDB0bUyfpvDf8ROru6Z+w+ZykFlLAj9TevKx/W03DHWDji+
VfwAMk0LYjSx/K4r1rnBVzhV/8Qdb6ZS45HSK9C/H4/8yzG/shojW1yjhj6Yq6PdilKw6EJWEYXh
WBnTgA4TL3t6GGgizLKHnw5JBBoAOv6cmF5SVEUcGN5/79DKhcrPtFcFxOxvtY8yofVq1m6heckd
mRGH6Ya1XsW/dD1CnBbkmvk2HgyyYHxpieoRP4L3NgJ1uoTzh4GKISo/5l+1xTXlJu/HSyjrbONd
ph6ZGG4GH9gaqs8J5OHk+reZ3kX0u2LWWi3FjWxWAdJ6ATCM8wUBrrQMX69IKae8ez0AfQp8HY+k
NzyW/vSJLU0+031gisKcoiuHkROhGcPt+mKNWqe5jnK4hK9mhVETWOcAdC1mZR7cun33lopAicHl
YHSbTt/HwRYduoDDZKKT7N1HbhTsT21EQF37nJUjROewLpWB25qzZ82W9qVWv+DiuEZxrPPdlMwu
yMcCfPRhe9tb3nWivmNUgPONP2hQkBWIzLvKaJFVve8GDqCDqaiL1GGmPWmR3mO3jOIoXS6JaJIv
EVeCbVRcT/PVnwsj9POwiZa4nLLyrivxPIYXn6C7RAanjV+l9LEmGO4XnuJJC3v16jDQkPOWuWtC
dIDa7ovTNgHUhO84zjznI2xAmCZisFkqv+t3DtMfjnWCFBjOkbKBcb0KduUSCvALGpzUVBZq7rA0
X992VhjBox/nja02eOfiJaRMFB94dRdh2Yguddu55eJV6R8DNaEpFc3FoEEI4VjZdrOwC/D2JJFr
f0UQvH4ZcsLk0a9OeZjd9MahYAO5BJsrTMwTWNrKICGbg6K59/8kyDftRaSLm05le4KN3J/YUWXw
bVo86moUPcNr5DlVya9kLGi1uzyU0Kf9pBeSGDVwWvd+hylxqKd0ItJBK9KSPO94hfiODxOh55Wv
D8tLkWLGw2Esh3xtvMHTq4bZO+rM9bStXYiw8u+0SJ2xNVt++/vqA7XsHHI9Jq9gc/k4of4sgLrS
U2b1sxmpaxO/bpXn8i7quf5hl8oFmMiCL2ZYdwjucqjxoBjyx290phVKQOj6K9k0h9tPYn/ZWpv4
SYZKDHTkcboC12TI/NClwnJmBrGTRkUqb7hE87ZIXHnEOqTIkjNawxy7bRxzv/3f809EhH0sZpGq
lXSOwAGIb+z3Cn71XP6CW66sQUKCz3c4wpRIlZvsiNa76PuAE4TpgtgAF3ANz5fxLObW6MHtkV4Y
Ym1dof4nTOmQNWJB9RixLgpZ4YlIpqaQ4ZR6djGCxwWrOUAP/q4kn3BJPfEvdSWutkZLjgNgstNV
hoVSelfCWreYDyrZNjoSI07LNbM3eFOjXLEaDFJDxAWSQpqvvsJ4oNyvVkiPebEof/Jjhk2PeJJV
eZVj5vshajhCEAZ+ba5IxCLvZ6WoitiHQ3AzrjllnIRoRFcn0zGHrDgSGhjS7QEqLOepDVAfj2cp
kM6cZNCADXC9ao5JVjzxZe3tq/KcRMOAI6aCOPLSzIY2SMDy4P+gJ9OVMiYkRdcgDrmZdAMItbJQ
E5/mHI9JNLM9PT0S9+CEHy0Q/T4sf+4Z6p2oRryQR4rwiQ66pGIioBOb7eKK/iW/BDhA3eTZqxYH
xbkfi8uiQ83y8RHDsvBakppF/0/DC2hHcV0Oyb5e4N5juPqM6MIaGsWQM8hCLEd0InzOAbIzZMo9
ugQ2ZxRReaKfG5PtowzRRlRjAp63C9Cguehl53i9698MGzO8NKNI1Lq7IiN0a+BfPTQTaaRz+sFL
4j2ovuZRnpV0W4E3JoVVO2aKnfSOG4FEhhlsdUd1/etM+XSs71Fwx4FOIV6rxUSCqk7+n+dd7uNk
yhyxGrBM4O/PWSLJpkdK6zvSbfMdYKtpAy0hlptBoZjzqT/KNVn46cqa7gsfcmnxxpJwUaGXYNfR
582Wzckf58IJVJXhg8O8ajzaW5I8H1THFsdnclinDboV6FU6u9eLFUv5JpuILCd3R/NxMm6LkdyE
o0MMI3dQrIe0WfGdU+jHtFNbtGy/oToYZ9IzM979W8xfy4Q3HtOBszewe2G107ZT2HDIuekMRbV6
3mYqGxXPKucITW6sBr7wEy556SgRTAxr++/kfhQMehGAvnSwbS9xQ8esezsL1lZLvORjrQ1BKs+4
lfuwpkFvkszqX6O5+uu9leHp19DLT0ZZRMo//Jk+JnT1OHo8rxez3dFKWOPy7uxWW3B7npDgfWWG
Ro1tAGbdAJn7nD4pCx3ISWEojWVjKncMokrWtOAqUSexo1gTq2VKsC4XPx/6yZrjLsv2yEp4MzkW
duPVuCkROlh+nDW1BV8jBBntb8Ayk1XdQvPrAyPWGvkCmKh26lDtjYZ+v5Lz/qDQU7kc+tbvDrtH
Q9kaG6YBsVgFOZ0I1mxvaXampsersHfDlY8+T+Cmib/SN2dan5v7hZUiwijoeSh4rCfglisr1dZo
34BkfHx75WmOnixnBORs+9Ux/4sTph+rSUPOHVVIkjoNv9v7Zul26+y0kWudfkodojHvZxaTPnP5
O1UldbxBP/rfcIXa+4Jt2EXJJKB1cKM/xoZmzUhkRJFlUKz7b7p5mpxlKrtXF64GUFmRYj4wAoqT
7Xx1K9Y8yY9pG4Bb5+/1VcHSTce6LRDwogXX6qquw0+2YifIr7rtgAxsJcZYwiH8Xr8fDEgpWgUD
TTj6Zoe+cmkHzseqNJH0wxyKob0TsYxwuj+l6ZqjoI+AQdhIUp6eFsefyvu6j3txiQsLzXpXeRKg
KaBA3hFyqJbA9rug5Wm62uha4QLW2nSFu07MndGrbfhAHNnBAB9I1yY7vU9cyMD3/vn+P1UVGd7D
KmhK3mEjCzyMYgMpPCcOFVQWubSjwC1AzQJoS/ElT2d3OJsZ/8pQVX8c96/naOVZzJaPsPWbkV8k
3cFo+Wi+TmkxLFxuGDwM7LwUO8yNnCbMGQq4SwmC6aLIIJWhGA9qxgX4dYqp7VmG2g01ZBBRbAPu
eqmwwEtD5GU+JPV70QZ98THYfdplnYm4fy542fClsdY2bMz+MKK40nb9H+6Jf9XR5wA1ngakfg/9
F0qXKM7QqZMJx2u6bkah0O2SIQvn/5NQRujw+EYN89RS/cDQWdGvZyJDz8D/OWzTroIAnIcVkmBP
tu9Zpf+GI2lzZnhpbl1lqjcXTNFZQ8gsPPRP+OtoTz7GeE9fRpx74DRINd1yyTh8akOD7OTLHvSB
WG3OoJ9qoDbGh5488xwpYKDs6zAEMTihJpr1EKzB56EpTpO8avLLAglxcgbzXrBZUGv29Ni6MsdP
HTNFHZZjl1IrFQLjli+3Zi+HiuQnkT1rZ8B2yOz9tYh5gES4e8aUI6JajtnA45X7MEs94HxJIxTu
BmiIviaTnoN63TMVcQrw5pJ0WQDWUtNmRBYiUnD0NZXLZbzTdTfgYMvZtvLpw6s5nEM851rIHStT
fBhLRrvjSFIrhkPVYBKFdcZhTuGwNiA9bOT+6bJ8hnLXKYgLxX+l9DZsMYGkhaCh6VsX6SC4SWdm
apEU5jU8YiwZbeZxcS9fS+3rcbn2yG7CVucbKIxHIjBNMDRMmb99outPAVsW/Dz85n+nGdVrMIKu
PruP6egX4VdxccKmhTtEEDd94pze/KZxQ4anmytb9Zu6sXTbU3xx0k/heiw7xXG+OURkwe3rydOK
rcPjn8hip9BMznoKDc6mfOkt+sW6W5mfNnck7N6ZtvSVj91V2iqyJA5PiosDAlgkSszhnwfwnbkq
5Y1WMMVZ17jC7I8v/NO8VCytSNLVx6pqOaGwnuoivcakGWCwM53i72Ur5RnRe915kaS4AoPLxZqi
jxKX3duOVAJP/E7x91toJm9XsxIhOJ1rfl7WOrHCI6dIMR16u9x8fOtdSwoM8QPywWzodcij5qZ5
bLljUDEc+cSXEpERsm/7Yrg11tZT7e0YO2H/98ymLzS+q0EhjWC+Cc0Q315OJUl4zPV2fc/SVf+H
nKoYiTH1GcxvBXxNB9JlHhBWEeODkxTCWtIDfqPdtjWvGJjbIpcO2yGwtpFOxu4p8BDtUEZPqgxb
prqVY6nI/qgzO+sPASuQdvbr/1x2QA3JxfWkABrZTXuaXdZ1n/gG4FCbIiEviW0Eoz571ED3Uafz
r0hX61tx2ccRm6ScBIZ8vkB3YpHBoWm9tb5k8nzDYkC2whItLdhY98PTlC8Oid20N06c2ltJuIJU
dLK2jNhqBf/fyTALraAAM+uZm8jM22q1fXsaq+n/cJAYkdNWyHuknygUDj+gVAIT2maxT38ScLTW
5LAO3fgC1xu/MjtkVGRvMBLuaKKQQb/6EMpXCAe1IRrDMB/EmVX58gjViSdfnUvrsFTqk0kWPA+5
FAJ+2naFjQUruMT22Bd/ws6ZSGMdf6ai8K+7bWFAzfpYAzFEovGMA1bccgmSSGQ9m1AyYJ5D/1Ab
o3AXrCV8KHJOmSFQ4xu91crFGVD/ctcjVtfK+0vzofSH2vcUvE6zE/tWtVUFbNA8Xd5F3bRCUIwD
T+9fiFUQGhh2j2vSwgyBFLgd9nODACozMoQkGAbTJ2IUUB6IzG0qHp0KHevL963Mlrx89eKFSu0F
K7G6QjO1bwl+9pgTMfPqB7Py2iCpClO2VM72WgEPv8QoDWcGaV+1gv5haPi1PxBdT4RNXJxymkxo
56SQ1zR3RfvBxYMOzK+QoOD7W+nWm2YqPxknSqHZ8Rhv8ERqgkchhRtRO+vmHVy3Cp5Sd4phimVK
6NxlphSTATxzCAxNKXBe1M0p04iiORRgwRZMLrR+cPUf/pGh+/RbgRETG4jepsWDQzvNgbQVZJL/
vOXN6jHerAYBAoVS9AiaUcQUcIor5ficCl7pdm8aHMrSNcGUJ5QcUKsS8RSxNCMN6szIiaypDl6j
fmegl7HkFR4N5sP7NCnN+2zMkt38Mp0fXcAj4SbI/Q+2YVnyqj/6WgRd8LhhR2QeeOu9xzM+1PNI
UlxWcORF1cS8+XLJvGeKy3k1Ee5FeWpo2LkQWtIFCTODRZN3IWuzfFlQ4ej0EibH5V19xY5hMxVQ
y7nNUplKcPPOhKhfIGNJcmWgxAC/mLRdRN7HpcJYR79yShx4fXygLysi+/S0MEuXpKBT5Bdi8O6v
oeZ/yKojb0jEBNkNtcevInOCfjc4NwKrIB2R8nneoltSm16xo9kGvSQu1AdgSaIe4IcdDuqqKTEJ
hb572kE0uSbKOzF8W6b1edMsf2kb2xfWNJ3lWJayLzmYn9nW6qCYxDu9UaDOQKLPO/Txoq1ilUoL
47bQKFL/bDrxpaRbk7L1jToX9rBOGgMsL5I5lri7hNrzaS7Xhy12qInutI4Es+/0JpmwDNjns9CU
IuGylccEGe3QcwfSsbhuMoNLdeIFxBL3DCLipK9/IhukuABf66QPqvMJ+CbPeM8l/SiwMjmJ+FkS
XpxCCX3m8diQKgi8zu0RWMIEy/tCDLEoiSzSypOj9Aup84AP6FYp5qf+RoM6/sHg+n1xavHhp+dw
TmDRATt5vCe3lU+AJqOV4/mLq7gKvS657SJ034vRk1YCtqWkqJJ4q3FSSt/OeUtZQZbsamQBlD/f
We6vzT6on7p0Wi5p197D45kYtZG8l0XpT6AvXG5/+aZ5lpQoJ56/5ICu7iRlPlKJ6fsmc3AtVjE4
cileAx0oMzxubFtKYKnhXgkxVVhwUGkHhFN2OIzW9vU+O6feTefWsj8ICX3ra8z1vkFKMwiNAqJ3
8XP6bTpe5RexECnVk6EiNcFv9v5a5hAEZ4c5RbPKSEE0ePqrIbbn6mUwS7Q4cQ+HZX/RuMjFPDwg
NgmOioEJjC8D8yR7zamuQgsBJtLgtZnZlcR/WH0qQ50pXGe/cXGCGnX+XaJZlw7bCjbw9AMIRiBf
d3EQJAPrD33OlYZxMo944u2VDw+xj0R+5DgM7g5sYFxtbcSxvuYQ0xaQeJUBPfAjOEt+Ur7zq5jb
cer5Dlu5VL3IQyI9niM8PXDo7t+r+xf6tWbzFBYL5geJMqY8Y8DDmWAqpe1xqwegZWUxJP9OZ6u9
Gu7g6C9q3OsWb4Fm3+AymzaAdO8AexOa3elNZ9negp2XmxhBbaL8+K90yXbcDFXkAxYs507sIqrY
vKfqw1nCxjodml3sDlY9h+Qb3mBfXRcT+Z47yrImgqMQ8P5Rg9DGsO/HIPAua0fmdyn2xOC6V7uP
Jpy0TIJ4w9EFfzHQjDoU5pmmXki76HNqcbe1G23AP841pVEcD0l8dy6ldH3//x/y8Q0VpvgI2/gA
RVGwfq5jEyh51dfEndOuTQy2gioaVHvdclnnVIXY6o7CmQeFp1FPsb1EHJUsjjyNrkfLv2iaZaq7
7sHPmtCRfDj6g2JVt75UmU1qeOJ/GP3nL86lRW1Hc1zZ6p7oLybOaKHV9YCKKpT12tJOIXefAs0v
oVQVDwSposv9768lkO/svIBptCIAgBEGm5Xvw8cyNKI0NTpfObUhvE/Az5OIW8ZmW80sbrJnruE1
tnU9uM8VNsDSKU4lNE+63ICJqS9nsL4vfosuyzNrTijeZv5wWo9Mcu9wYkpU+atA+CqrQvIOl8DK
H1RoWcECe0vcqAbjEl13WYhEpR7C2DNkdlmuLk09CSuR3FSHfvyLv9QpB2TSk5quyYKiUyuG4ViP
5xIOkTVhNB3u9xd+zzbrElIdQESTr9sk4RSjj0szRSABDon22Wnt4USgz0/E8uFjWoEyGA7gd0Zo
GAa/7w2IxtjhSDvPaGFYr6AfMreoSJoJ5yEKdFm3pr+hl9ln2GstuAU4uvaL6JfPaF9nJQGa8PK6
SrtdOsR11KnFjY+r0JqBF4Xm07IE0ivB1/LuE8OftG6MDJCiBeqXYs6eR4+tdH3Fz9xcP/khMWKH
uBeveQ0fnp4U2WZeoDVcGGmhMWXtUvnNl4fsYcoqWimaLpyUz3GuKV1yxbdkm26UNe9KuzJ9n4lA
tQZb+U82G3ilAqgEoApHhV/RtlcKiGxepIADlj3lsYoIsFW2Ffoi/m4bW4PExi9vWbMDbKN9a3DN
jDXvTiklE338rT44sHVBJqi/e7C0lDJ+RTW5aYjC/cSd7yfGZov6wEdJs5hSak1Rsxa30WNbmG0A
23g20thbwdF7Ae70g/fAjYIJzg38emsGq50Y4rPFkaHT+kUjreHCiRS2JDqoMul0XQAaz7CUhME4
mn0Vv6am3FvqAieZRVV8g9Ucew3uQLelwIr9dTFCNzXDTPa7Vu/Bd2K6SKmYx5qGjpQGQwZc5unZ
upIWV0nnYgNUJg98MQsNY9TMOReHFxSjWkm0+z7LrVTLIigcAZ3IeSZ+4K2GpcKqjYq/kKo4jLw0
OiViZjj+b6zYyb36inmHVB6Nz1Cf8XxetNkHPaA/MYkckY6d2yc/RZ5b3yeHhti6cS+75TNqdST5
ihS31GtyDelrRX2gE2o/dX+5L9IsTHNV0ibiWQrh+R31bkG/fBrj48E+SFlX7hB3W8rJiQvZOB02
9iE86eG6NzdK3CxMhDL2+d7n/bEWg4zcZjgLlCJm3/aGNjCRp1yXSW9uKU8S2e9C05eP235U5gFv
JYqxq+sFPZkcr2TBXLbINeYFefaxgX6ISShUct0ZU+xMvMmAP9PPjieNCuOVfQTze403u8k4da+X
Pa+w+IIys+NORWbOfkxEXDFiiKgnoW9mmoMT7UZQ79b3EAoHoNdfc4RgIXibsmcfstw4Dwrnv6kH
Qeadw2UfcqOZN21W0w6I+KU4y/tgFIemkdkwuTYLwimLBKer438aC7Mu27TSU5rptiC/i9iGQcLA
zUsd5oawiR0kpSTeqg+5OtuLNhy5vqC8TYzfU9Cknyg1EAbMYH2oAfpjgffmnQBsHsJP9BLPbsgb
V8NXqz8FKtGxo+4Aw6j2gcghW37tvN+ri1TzbZtlrrBoSEMycpT2sT/6RCW731yUq6Q+JhiPahYU
iEohKCW+IAcXWGPaQxFZthv1jp+4jiaR1U2K29y/tbru+vRwUJY6gjs3MG3rrQBzkzgiFQJaP83W
ja8LWfyHdX17zvs6Bom8zfsZbMcTCtEFcQG3vm1aNaujOl2ja/wfbJfY9kglYXfEjDhguPFpZT/S
FABx4jpfu8bzYOBXgNX3E9gRi8gZYZMhcf09LIbfgpNX/lU7m0m3YFV/mhyC/sPVuXubKuIFMhxx
7nU5wSSWpRHe0R5CCxwMeiGeWGp4cZocWQLbJj32meGgb9Ahxf3VVNjYQtjZKsw6d+azKdUnzxHX
Rz4fLz3yzVQwjtvtxG7orBjfKgW+vcGUYIWw9MW5tv+hKrCZQQWa2GXalCpacCrfkjnhp+zcyHlA
mcvHwZOGVhLZDAPB//o5Umg2ubDO4aWhzN5c4Lw6ibbm3RF8U5hHfF9zggQ0bVjm5n7wzmppMiHQ
WGUVGzh1TDxcN9h1F10rH9tZ9Yz9+hO03yDBmKPOu8YjxElvEAumX6iB+mEu6bGgTdBKUeJVN3kQ
xKJ1nY0auvoL9TBZLgRQUlslh8nNfUdng/BYCnH8XuIh8c9nbrvXJqCYBQ2CTjJkdYK7ve6ifhqV
LBr3B3r6iXl5dX/4wizvhEszwnHjceYKKzGMomxa9p8B/fk23mjfgn56y/gHr4FJIkvIb9+e15OZ
uX2UrEgFF1KxpJpPF19Eltgisn398gvg2istlwzIKPeEWWWgZuXVOEqyP1ERgy9Itg2/KevRsJcg
GisoDUtkaTxg/CMnrN/+ksNhY/V8+xfQUytDzBD+xaroxvCrLjSDh6Kr0MqUHpsZQ3eSZlihY1W+
DYqpcvyl2eJNPio3d4NXgxF8INE/EDA4vgD7vqgMFhMFlZAl92bKK09N3rEppT8GeIg0MdfLLumb
a2xU9krF07dpwl5/JhUQSzdmNyxlBSD+K2RKE52G4pQe8zM+NSVH+lEZhvfq2N4K5eM7YucezDRI
ejnuD0Wyi4shwWLtDSW+cWSb+qzO2J6owwPKsckYnbhz1ScgSp8RRQdwGl/21pEJeCk/Fwfy/f5g
lHcGiDPeQdWNbgJIHRvOHKM1PG+fpbta0ujIxnBLLhB5q5OFJgzWfYDSyxshdxH2okgNCNyAS4so
ps2nuMVEtIrKHdPGy0TE9w/F43I6oHy0nJKHOSu5ApRnGyNWR7IYSw1cluk3Sry4luzv3aOcvs7S
dXWqs/BI4YO8aT8hH+ub6MJC+pGd6oqSlgNp/tPQ8e91FulsOBn6Y16Xo2vv020kJIa0S/2zNUZ9
RTcXPDVUt2zI4gQ5e5eyf599mwiFRU2KNliRiJuYX7ZUpuWqsjMJ+mmDxKykkQ5ces2OWsgYo0UM
ff1/7hdPc5S5wdjxYIDxuWVSjjx+UtAkqUdxjZEbO1ud507OszWD7bKEKbe4oQLy5oQS2S5otmN2
+AzojmgiTJKAvsRp17V6oPVLWjLsI9ioZHNf5UqI9QM8zuiPNP08vFCW3A0SmiciTLwiX73FieNE
tA5G+FAeCYaen/kEMV4UCrBykwJYsW/ldnMKgjEafyldN2EabXqnf1+wbGhyNThsvqb5/aqc8Sel
3ARevCJie4pSHZFiBrYScFLB+BuqDGCzGiArvBTRIHwdR3Q8aVuSFw+pz3nAhswDU4PXw5wr1BC8
Hi1Sqgi9kHYLSLWIzMIDTQ6+q42c5SQJENIuOTIWVyMsg5X3+CVmrq/yivTVVXj2pm5EuM0pVUWH
bn4ZlcMQA9921jwSqHmGJEi88fDguH1WfWm59MuZOR0CbLzXpYzMrNJ7CFUAU5Hvnf6N4HKNfcO9
TBOtyChcH0LMkLTrh+sIFzQ/oK9RUWoDlxjGdE2q/F+UN4NFgRs7hHoruE1TRPXCEn56pjGz1Zhn
uNAD61A0FIM6e+RW8TVSjAjOhioNS/hoCIGFIx53jINbfUy8QdMxzMMRzyDKWyCzq0GScLzlTZ2+
K60pa9kF/V71r67lMZ+kaVYc3Mmf/ImobNZSyaXCFgimBXfL9w5cGBAicAeMYuO582sH0qYxBwwv
YdDcAZ/lLe8FG3IYD6oGLfMF7Oh73DwSXPfZuHjQQehjgRbfMvu0bpHz3ExL07Iu8fsMNxyM3saX
oYV1FDr0iZB1tmcqw2BiuKFDmQNmWT9A+QQyBZnSG9ptrqkbL8qUDyuFLL7kap58R5MHa73jY/Bb
rWQNMcY5U09fYMucxpvUtG801MLoGTXuahq1ZHuM6Fm2mkTzYpghnJrSvVRdYh+0AaOThid5dVsL
tCvIog9VzUN2ncNtqhJMJJzAHYeho8HSN0i68zrIqYcBuSna+Vepitxhg7vSNMfu5D+Q6HHcjCSZ
MH0f+yVK+Zr2IQjL0gpIyfhYDtB4GqO/dBuF6I03xqoh+eSIYWiI5pCeCNvWuDMLmral4NsgNis5
EOmu+di9LUM4mQaN8b9MXPdi+noBGllA8vHLG1k0ruOUXCmoAiLUvZC9q8D/kNiAtJciTWvYnyub
oOP7Oa1ujAhwGouokCLWa273LfniWNmFzkA7bV6rJD9aQwvmkY4SWWBDlPE5XJgHJAnBPgZDh145
2fdwwo3Qnhjdcrtn2le72VamLz6JgRFHJE2ogU+vBU3VBF5zIpLp0SxDVGHUrGOCRwhwyEZ0Y6WD
/CE1CPXgpZNMEpzjKYPoIpXPju+DGv3BdS65PlZdrXzHt2tp3g0lUhJY/tKD0ZJNwc85czabNu8R
MbEt0GHteG9ax8oPLp8N4FGeXGiCnPWKklbsqs8yzfQDTDd+shOylMDiiv70m1ifmYyQvwbLf+C9
fNcqq2S2Dte6MmxFLE42czI0aKvignZQRn0JHdoAs81UohELK65glJMPOCh5mxtMdbe3CqQG7elv
2dbvfsXKFuvA7aLp5E0NilXi8BdmmqwWBkKLD2Rc+GIB/+ZueV+UKqRDXJC4gOUylBQ/MZW/ABX9
QC/2o9lWOCE0JEvG5/cFnF9yx+npxvCuhV2d/fSl7e3BT2hNmyCUb6blzGgbHzdeaUaoFPfZGGdb
nmyxrHNpNSytLuFSJA4LUVdme7Am4VfRnio3GY/G1LiKyE2byATWuCST0euhED7cBDcESc2M56vG
jzZn1rZGS90k3H2MEbYn84mEgUxoSVk5DuGo9nkmGpKqkv2c9wCgmNCQdv5kgCJrFmsx5rBsxL1o
7yUA7Bew2px5eJAPf1BJmZhfANNGinpveyIPjbwOncxzZfF9nOIWURdo0pQpY/PpNSmc9sNsZQwS
QdTgRfyCiFarwVO94VEgmUTXRSgcryIsT6+tH0pFRug1ACg9N2J+K/pMln2hbsqaL9i47rY68I8r
MuLwIdIX0MHLASnxOUKSmiDMSyKHVBp6i8S0FZCjtN/cyaEIptIFLAP51fcmnoNSb3TjynINEzvI
riisgbi7xeq2QdXPp2bjkp6GkMW0em1wDOOuuMVNu9KKRx88DW1LIIC4tAZpB012q25H7LmfUKli
fq2RreKRhrkSpU23V4ILms/BJx6OK3b4aUoWVWFA9w4kX3z/5G3D5v699Fnwbs9LTeHK4k+nOCKw
2jJyZ0PL6AvrzS0LbprtIhwZIAUk+A5V34uoOtV6d9zO0BQ4vFy+go8gyWcTivgrj795A6r0kOQn
Hk4tfnoz2Cnuv+wsidDh9FigA4EU06rDsql4wXxvTMFG1bXVhjN1D2rfCEQ0MiJk1kf9xkxvHrOx
+yPn+k0hV6sJugCuc0XiRsJ5NmRzL/pcfX6hF5sK1XwC5pmlkWauYj+GQQnT+Ne2FzA2FI60sqd/
goUVaZcV8IL0Xv0Pj5xx2JygW2h9P7mYnHGDg1+ZwzUiANz/xjYZbdCHWNkUXq1kp83SLj6HLCNl
/EkaM0tkmOFxVXpFVzpF4I0qheIS0Vf1naRW+8eeasA4z94GUJLZ/oe3uA5dF+dNm+UxUkYee4zH
Pi0MEuBob4TExwWDgFbOMsEl1ti1RemIXbliCf+/x8RP17gu8iJqYHicqidIIgAifYsfs2nq/Gon
SJZoLw5vdLepGQuzzHQviKmA6PIdbVHQqRtXjOHz03+FCg9bOiZrQoEEXwVgT+PaADy+vtPUfVGp
l/KUI7MCyHMnPVCRZ3i1AehRbdYs28pWuP81hpnXGx9ykoFk4A58+vuKpgpdb5pF8/Rp6ihubWPI
p6ZxULaKSTf4wnKA+tybWgRsbAUUWbb9qdyhitRVDB0PAlPku3CxOQS0m1zUBc6LeGPJqShST2Lv
PhnRztyBWbIWwLQkvhBFyJ0H7bd0lRu8SSeD7qxZdJGMhst9dMNFCJmFz8+zhVlOYY3g0m11qD9T
L8H1YMVgNRvWBvwcNLVF26QOYl/ceCXJCt36Hy8BeI6FYQYXb3b/p2YGONu2bO+ngPv4/EyLq1Ev
PHQ0PNGQAyvuE4yS/Dgn1xWIV0MHLaKMGiMcgerO8RvV62oFA1qsJ0xYRWECSJMpoanhUjE5eC1n
aizeNulGGSwMSXqnhpFBrfsOvDO0iWAKsL8rPXgg5+coJ0PmDHBn1ldkBB72+Nvmyrt5NN6uw0pp
yg2LMcdkNdGAJHAvdZkNiu4S5eTmhacJDEtQfFhULA57rHg3/JY7oSPLwGDxiuvDUzjt6UZEIW1f
SQlO39M8HtYwd9/DMKPDwRqcJkwN49JdntA0jtOjGk+yg1OcqzJX0xryx/wZQ3RA5nOWlvd8IC9n
+/Ug56gr+R/zXMRIgyTRlEUZKztKQCDBiadc371F8SHkfFL2l1IPnbR4G6C2LIOzFi9Lgbodk/9H
e67myzj1tuSNt1RQYNVOGGoHuRVUQ/v0vIN55EkA0OjyTDSFdlLjslQWqmT03ioTvuI+GKAVtmvZ
C+k1SBX/kEeqt+cQZuYjYicPaJt0CzWwqJko3t59jHuWEn7g5enPVnoXylGUYXdXuKF44iDOmA6F
otqNm5yyJ5PQ9lkknRBrEZSM57oUlkGrymE9m+d1WfkMQY/tAZe2moeOvoMwHvAPtb/mnNl182zb
4N9J2qZd2pzND9KVPCjHOeDSSSNwckFhWRNRtv/UpYwsgv6qlb9XJ87lbcWuos0dVS8fZ9T8o0nV
O1bUmTxRO4LTIJ77ug/a9UKv5iI4ck85ah7bcPL2DfB2e/7faO4dSKaY55b9y5DtvNd6mCr0bOqM
9MUHVdbzP/XqF/brvYZ0tTesqtd913cMx2zyu+dJzpCQKBzzvMiO6P6rqd/Rdj/43XVOJkKH5G14
gc2NKZ3Z/sH+m8MlQKy/ieJx7WXbicVAQONNQCmPMo5PCHJHutk4EAwAkop6oojK3CJSaFcO1fSc
A8QWTTv/UOekaXseLgQa/uThC8gUbZnw4bcTustQcO6LwlIwJPmn2MTMjtzC8xCnGFtXgWjq1OE8
SOuGUiK0ouVJgquy0e0UVqBi8CicdCgLRDaoVkWiCd85qnJTbhzwHHNVQt96/qHadQDbDkbi5QaZ
fdznGMHyNWF+zOGdm5wqkCBn6c/37pwrGLasPHnQyc4LzwVKWP+XBvlP7xgZiLKmgsG2B/UgufLR
DCXe1ji8fqu3L2lKaeTPy3OuXThjBXB7HYbGxQEkZaDVNswuo05wO9wc8OwTtWeHhMsR77tO4x3T
aibUU89DmLsObxZ47Ma9ZO04H4pM5itVcS6aBV9lqEpFG1hKWcDVivp9OmukOz7tnBvuyrgB4sDW
JnKv4d185FfBFtL2yzzBwAh/Ez1v4sOpOE8fMjDASGjL5Q9f+5oBnv6EbSgi1sItZtgItmcVLiie
dOABKt81xHnsV82DnFKh/Eoy8YickbKepA2GYREPBLLDldqdLqINLUf4kDsOxtgOn10dbe7nfH+/
A1jkCJ9oqAHYB82R5oV3SZyzphR0wrXIXwHE/UFWVPzEjrWbgtL60jZa5ZZfY+MI0bpjLpQwT8zE
o5vMhDIBIcDTZdb3hdOYb5bOx5LjIcBSjmmcZKCz6Z5pZxUU11W5MA/qOIE3o5FSJNEUcde/DJ2m
6God/tFdu6vi4rBe32Z799QH9NSf/RO85Kwk+oWymvlljvoOZOFHNnQK/jH5aCB7YwboS9DjG0bG
SomdsD6NSotcM7bthSJM7C2c9ZHmo05nZT+9VMOuxxK9nAX0gGveTeHUdh3s/dZTrWYIFHY4ajhN
dsH3QrpIZqqUaaID1y84VXJ+cClqc1PPzr9b4wfB6Q0D7lHYCVOsyokk0QglR06rlKgClsiJWQo/
HS+DwpvshQMmlcCesxqnJIw3qX6lxzGR9BL+uxIojXXfbdZgIrMt7s0ZD/dMLm/RObEf9/VPBJFh
bCvbx6ptkpbQR42rLzMFLZAVilX0KFhk9PgH6Lw0bzzgF8trDEb57McOBSy9nUWdPE1CLEZeVlRk
mh8R/PHs1VH6MHJnEoYaa4VOwk1lHofKvlLmwD3od5AEhgZs5pSXlIt9E5Ma5Tu0PLps9MJqx8Tq
gu5Heqc4NYLkqCretpnql60EgU/Ndrr+SaCBiDNV7bPzdcUt8cUFkOMRNdSg8NOsED1c55pYfe1/
Kt8tdg/8Rd8jqqPJCFxyPsR27d6Bagwc/C/+Xg4CedA0j/pt+fqnc7AlQKfZ8+zKthqbP8dLH3na
HIv9uSUt0HrmZOOzHyK+h6GRirw4m5t1HTeJinnKtvHuZ2Hjqm90Nrau5LFxli7yzy7DWTG6GG6h
rV8rQ8ogyzrrpXFfqINwn7hSlIv9v9tlAhLTR4KmvvzZzxQHvd1qHMlQ27dUhIF6H8QVhnmrpfuF
LrPT0qdPnOgBZCoE2A+ecJmJuqVPqcpM0lV1pIsT3hBgHc6ybFQcaJAX/N5HWWADHfPHskIMF33z
jTYnLy6S7w2ITbIiCGCudNCPMDP7nn4wA97/F/PtRTrsRlEzqiKCEBTrtksMuPylNHyrq3XUdAHB
levApSbMn3N4jP5HzhV8N/QL7bxyu9oWmIpbexRcRO//rXqwmY9JbjcrgXFTx7FIIejNtlGcfR4O
lRqUYb4/DPbtpKnJmhEy9AKad+i4wWnOjGHIq3W8lBbIRoE+wBtui0zEK7gwnepP0dqm6Nb7BGTQ
R1als9xYsZO6EyD0IHg63Ty+DuNxir3pmRCPNT4tCQ4+29qEG20Oq2/t7DULiCwFpv1lk9hXv60d
PsFPmptOl8pNcJ0cfQ1MeGslgB2lZM2pJWtqIumzQr2BkwbpqVUXaaiS1Qm52QXyGkB6zlSORaZl
gqjSjxDkUOq5kPTrYZFgWN5e7zT3mNmtZSQDsK6HXDWGc29omGxUBdjfQPJnwRuXmIAZZbgUwzJ4
tHFJDXNNk7Jqz+gOgJzxLYMjV7GRkLfP3E5Y4fhLqlV/spoeNgfjK//g9Oy1d78WygVfUL9T0Jbu
ezPU+6POAv5CLba6HuZWBYMpPRvzJCkviW0yh4gbLYGKltzhNbwbRq9CFWC/qXL/TxVm1gA5kXMd
aQ9rZXk2Qz17tq5PBTzZpzSojD9Z6vrYdTkWqV8hmCf72WMlq3D/7SowHqUarvCBqBPmRPThK/J/
yNYxuHmXzzuKVLUIkGKbfIK3HgXucauesWL4tDIkoQogs0R7lJAu5GG6vKE6haUJhILCMDUH9WD5
FK7LG1exDuxg+l7NpDcI6zFeFYrRAbcXQ0ORcSrHdE5BYJFGqAvSVbL0TJr6dpdZmPIwsi5SERns
im9WCe5OjVT56Fw8Vy877XZm0bRQwG6VpWpvTkcN3wczwlr7NKNPNoxRxFo31NDtFZuWOv3/GIew
YAPymePm7MWp+hl70foDQQPpr4HdEzmsNHL8/eTF6VCWdNef2+PwrT3bz13sCzF5iIsfwqj8xB0L
lhl7e9goeE/etYTXLZVrgUw7a5eNnEUvPyNBoGbV0YZSGs2SK5HbqKLbOEiJFYDrjVmfrBZj4iFZ
hLHytEx3nnyKRhCOx50nbKN6PETCgbKxnAAs4WOE21lx1VBYyCgasBqhbbsBh0qUdV/GpnOjaCRe
3z/BT4ocdKmJK+jN96OF7PxLbtZXs7xbXWuGBdXGZtLI7W9gY1zU5pe8IGRHRepMWMu5v7SC2yNf
PoWFDbXYr1WA8gcF5U2VcNIKbtaXTp4v6HBl+Q6HYkvMePCioODQ5FbbRtUP/vyfTtYefiZZEH56
PhhIxHK86sTRIxjRdU6KvYIOuEKdQ0BTBXo0qLgVQPNRSwcjtaUK6dHehen87cM3nXAxFJm66f2F
KrBjmMRjRBtRuKO1iJtdFp4GTXivWxDfME5TuZorkrzoFG9Q0dpPAx3Ku6Li2rsP4qTY//5Fu5yR
6meeG2TjeSFdiddYV41w3/Wbu++31NuAaws/S9232UOzsSx5YDbcf1W5i+VD8uSTc0jOZGwSnRor
GsBaTC0UsAE6ggR4d5AI5LiXkMcc79NM0Zw4dDbHx+3H5le+SihfU7HB2WJh9tp/EbZJp3+AxKeS
dgeMeZC94fwb2TCDx3V4fz+APrT0uK0iOtWbOCpIdRk28MkdNEDPe8v7naxxvD1ZuhXfBLQB0M2K
Shm0I2l0yg+/JLsFkdMA1UDQ4mnF77IgK7AU1ajTqiNUe+JiNH9eJQ+25sK208eFutgHp6qWE1MM
BmCUIN3KWsqJxCc5MIjjP2zSu+OutyudHgeWoWxwPTfCwXHqk70/o9AaGrUX9CUSx06LQX+Ac58t
H03DQY77TyEYS0xSDCpfJkuKFD0Y2p8v2ma2ffyeuqtxea6hlXC2JzwDn1YOWd78ZGHfIRBg9Rvx
n8xEwykOdczMFoHwSywYT+BxkuMmE83BLWvsvlbLEo5N7D/5JAwt1M9W0t2kglavGuVFNM9qmRr0
QfZTUwm+Umgn6OhSJqCqyRL5JB9pbNbPdElMP4HFOHsOPtJAq3w1Nldtj7RwLIHwOMXjYKl9WzIB
9jH4IyxbY2ZaiQoWCjEGdN2A0btldEta/Tlim0L3IqUUlpVRkYwtP+pjIvX9Z7ISAqGmPDOVRJD8
zGdjLNDTFt9DRFh/J4Vrh79+Fe8qGWo44gvCUqesklsWd4pRV7z3VBjt3XbhkFw/pDv6ccTzoOwI
Umfjj8cD/WS8ZqdTPfy62y+i6x26CnHCYfyjtGzO8xitmSJ1niZPiQgdXI/IbR1YmiMl3LGijvNS
dh/GJde8EhIom57assjONnLEyIf2OU1RfAO3ANpAHH1cGrSSrVQ8wKGfFe/W43GMLiG6QXC2hIW0
jhgYqE+MTXAC9HhDvPODiNtdL4HSpnBrRKWl/GXVbp7Nma69FwEsPyZRdsCOxrQ7l4BurJJoUpUR
b+UNfXf2oruu3c39wyN1nrRx9RpNarvVmh8il0N6Zi4CrfkdbL3K7SSETztPliGmo12sSlRUlX5U
52FW0v6EUUmpBsOefqaIKlJdsCOWTqBbqFov+1W9J1oLo3MXIhNsjlGOLTfESaJMGvGSt2uRlJCL
M1pYggDH8TtAGaEfc2+8kNYNtHUc9Emdxq6t1GGqtnyS1kqFOO0WDoLM1+mmj0U9VEI4x5XeB3XN
r7Q+UPUAQnaenytdwdWOjqZHbqUICLmFbkLkyxWA8ZyxJzhmJtb5RHx7VQIeAAPt2uxLxGljHnov
ZX3vqQHhh9fPtN2f690yCANAjGzSqcHlrGi3VpKb7+HFwHEm3hwgIU5QuMvqjDLZKunOmkeMTG1P
uhdXGO8aVAp0O3zb/TmbyZY1RXDnalzK1xSwU/vOnBI6npCFJ5uSb7O+aWp/1P9CLZevO4MidZfD
kdYTw6j2sfIncpN5k0lji4vMn4KrXNAPXa3/48cg1s5kdAlCVrQqH/hks/IlvX+167BlANArWQ1U
BjgJLtujVtbc8p8X5WukT1V/vG3EHc/eCA+qcQGIADAx+pALUa9ueF0sAfu7NJGLUOK4f1Gu8XGy
3xsyol7tW8kdi9cih9m4H3DfHN0koPgMv3VomgNnecuZMTdbpiZP3/JwJxZRozOavNHD4QVpy6XU
ZClHAysYKFiaEvEhAaYfaFoiECS4QyFNDjNbaoIN1/1pdaX3yntIaba+eH++Z9qcF6fIHrSJKjdS
RrpbIOVkl3S4Lk4JK7G6gcQLygAKZwkVqWsz374lJ5rJ0QzjmNFOeUBPWND0ydDURu0jhU4Z4i7O
/ib0rWozlBZGhvAvJTJbABZx/KO49AvrNrz8l2S2Ktm6HR5C9dJjVwACoLd0IoeLZq94sb6MdYCY
9EHdzxWfS4R3n71QYj+Nw16NLTBvC/CNOOsGLQ3XwevIAJacf3LhIcu6/y3Auke8+bEgtfY7c5NK
fBfOzjt5I9EiVpXNpYyupoWEYOV5QqU+vPbc4QwXAGoSo3pTQh44tgoN/hsKo9VKxi7vA6o5aKwj
/X8fHlfqS976k5efJJvesvehX9a9cSbfyADj6GSp9x1xb1S3pmSDDOtibep9VdtlGf2ckP4LsWgk
fvlB4hVEEoMthGKnvooBhArfyY9Vaw1tQz9bDv9GRQ8ICzj3jMD8rG29sC6HyyWXpn6oeKDnkXuy
xsvf7Fx6ODNY7NGwN4vN0c5RyNtnGV1Jub/0u/yKJDnB/93Csi0ELrVS/3X3QTNnpEFXERoqBnps
+OQQf+x0upC1YgSwrUCZqgFF5+cjGhwgt7xbU0uETUhGrEZUL1NHAvRL6MgBvDjIRzY9cE1+MLFu
x/5Z7rdtdeq9li9zxlmRQLUPio2SDvftRmvup60XFM7K4gvP4KjiJSRwCNfc3gpMz241xFkkWYdM
Rh3aeZeaYCUSPQfwGfldS/Dg/7yrfaZ1GKvLidpEGKgrFwqOSv0vgsMBZwQ9rLqC1AKnnsKt4C3K
d63+gpgLephDNoWrfs0eVJRzMy9j+1B61dBIrccMlv5SFX/2UbpzApDkOvEm9ETte1LwqLiULbRM
5Ugk5mCvS3X7ul0B87lsgLW/e64As95Or8TV72whUaLURgBHAk8aHFeO0hotCIlctUTUJfTN86lS
WJHzGqS05r9BDzXNErNJJT4yyRMMWxbOqBT2O4Lt42Wzz10gnrkeJokMpAOmtT6ZMj4gerfRddHn
jgefIDymUYttlIiopr95meIF31zJXpaCqR/8oL+KKuvEmYVY6GFdlTfxXX1a9zkpFAiesF1cbaO5
Tb85BbA5NrFenKJ/xwV7igLaeYyBWwkBDqBL9H+00WU53Th59qxv85K2A47hxlc65stevvzeNJ7V
xJwJ2IrKAdZ/2iG5toutNL+Rc2RHbj6NFlwdv/fqwMToIn/YTyvTXtIw41PDYrn7mgvcRqkqp72E
tisNN9yb+oSyDdnZTjjCtyPy7LmdhhGwtURyXZjyqnSXCUj+/S4Ngp95Fk1Xt5/6em5LQVCb7SkD
XG6NtXgKJj++KuHx9xnW/jkSqlKxlDI8hwnxEffbe8XTE8hsMCon27WLYG08FDuIVfoI2RDSpjSy
6epNLz3N9YSIEi8htWhPTI6Ecw6WMRRrvsUoemStFvbjtIFpQ7CBFo2igfAgx85p+/NJ+5xKUmJw
3A161i5MA2TCY+K36uKthjaZ5Jxobh9xriK290rwfogMzY6GBfLYw3jbXMLoCB5Uo3NuCUltCRr9
VQVFDs8DE5sQ+e2U74iNT2S3D44zkg8qtB8fK5DlSAAntJoEkPP66zJmNxO70FQP03rxaKohv8zJ
XCZqn/BMDFNOuSOep31eBW3dHKhw+aGjUTT+F7ILvAI4X4X1x5hp8JFS8zBcYl3tB8QD+J7vbTNG
KdEEcdQLglrfwOsk83SeHttjPSdJJJHqJA7EJU9oTZ5O8fwgA8TO4dDF/eY0tPhsGa6YIYkDnAK9
vj+ogzzPjkGOC65yJsor6ihwmQjrTam//r4IdHKZIzRp1CLj+a/fU8Fl1UnLoCbnqg+/aL06eL3N
Siv5uIuprLlJjCh3GTfig0cGLHa2Z5PZvO3QphyItuP944V3xvkNi5CeOdXrQ1F7YpqI0UtiQ1GV
Rcjmm6YhO2aVTpvq0S7eDc1tw59zdnaT5i/VE47/C/3Uel2GqaVR+5GeUNm6jSbMsIE2En9l3doF
0SmXaCfyK2NWMNGqAFQOFy4d5GfVIg5aXE8BVyiDqdifoFpztr0viFCLNf8r1YK0eNUh8fYoFz8k
lARzfiid4PCppezycD5TusNIYsx99lhLlTibvu59dcuGvDI2XJrPFXjNSK+P0p9zBrquFejfq8gg
haOZ8qjZgmpU2ZepGq5iWKW2Ink4SNsn62Ndr8b8u2EUAOluytsB+q6jSz3LJB/kAGsmAaIqG4eJ
dKm5SqljrAIdI9MazPDPMVBt8tzn+m4UpFXcd4pfLBh5unmoiyuA0qyie8eZo52e80qp6bPW3N32
RN04JD74n7Cz/KgkPwfAjr0xLTYNhDQcvv/KaLf1LAiyiR40xPauVfzqtUx2oHWU4PmLh0VrNvao
4o9fL79onIN576jdP7snsg9vNgTp0nR/KIRqHatc2kSA4B/pmxS1Yry64gU30ayPCuGNaRVb4IQH
66qG0ATEw7xWYHY1l7EikuVI9kVZki9QD9Squ/2Leb2b8iGyamCGj5m0lhH1Qf9nduOWyS/NXJ1m
6bz/aeXTaHWAdpN+mPgdE1UQzorzZ787+1djtwj5UXY1D6npR+CcpDOcaue2TowWkvyl5mL46EN4
6m9KVq6VqlbRrxNIbszOjt2m1AycQ1fEENWTGlOvljyXLZ9CI81NQx+0yi1IjxcfH9pSQ+bWyDFt
KSEudN4H3cLeNCH8x1KBR9iczuNJGauDLq094C8v2WR3KUTaWlDndG3uKq9GnjRUQSnSyfDfZGKk
eZ3T8deaVCW0XCU9ld3Xfa8OE6Abu7JXyx308Mak0RDGVz+jpiEZN+xS3XfgJHjnEyLq8E9ivx6y
Bv6F/uimPjKEq2gpoZ2mPplax38cAgTm/2DXQ+bVykWEbcwknQgS7+G1aLbbHg10b13x/sS3L0Jd
SdR8/lPNT3Nu4dyxDwcNo+bITchIPxTMqVM3j1BoilryJ/YGWj/9o74vBX164ctAO24pEFsTCzwQ
0SaJXyEOV5xW9C5FYOMbaFAf0YPGnnnbk6MMGrgHj4oH/MNunkamkURNqvfC2hY0UzDE13ouK4AW
Bkr5q6AyX0nk8DUQ5wirWjgsGx9/fFU7joK7P9LZl4spedCzNBnz5WkIyajslU6LzXPIT6V7ezxt
8FDfC//VBumDA3CDlddrVCZiKJvmtRRPvI83aW1nD9JoY8CoipLh1W2m8C3Z9TTkjikYlogpPzev
DpyfBGFlHuW0/wohN8mDQZgUWsPHaL5Z7H7fRX3LD4HxC93zXCyI+zBqUJwopk5F7sPW+cefDIeF
Gk0eSEhvPGkH4tYMlDCrQFCT/jcnH4MZWZiH3YcZT+1nDOqZSyBLg14GTZQRpAUABp46qx0agPLl
w6hEa6u8nDhQHwWjG3LhVeCRrlINRsrx9BJFPqLNfxWGsjm5URQMxzW3S7DtJvnVdlic+5BjGg3e
E3mVQ9j+jxO8gesIilvZ1XJ4UekzIuES0etEAnm0svHGbmv9yLrpkBVjbVvRJbpzSmEvTTgLSRFq
m63IixUF0tkcrchCTsX5WGLH75ltinyY+hmwHfuuPPn+I9YRd5/8F2uEZm0WYlfb7zW+qTW+vTjU
FJmSoy4joQtOWLJYc3+k36XTyaSvvNPZQjvaDpbXW3LiRB2EmDfhH/3o+AuQIj+/8U5kPVLBDUK/
/XXYWsKrT8DikiaOI7jubwvS7CnK0CtlqotrOSXW4h5NZN+1Hob2w9DzcKk4PQtKqe8eaFOEibit
bsG1+blVO12Zzq4GLz+QHvRGYATVTQZRnOdUlfkMSi79cgWqh7Z8BDzRlSW5g9absjWVlCcBEN3g
Hiz84t0TN4nBtErEmMgBWmRyblqlvzEFVEyOTP/UF6A6qG2GmJLmxjMRslC9nnPaxLZFl5pLiyb6
c6LtgOFGfsAVkym4FWmoX53JmsZRoNGUuTsyjYHvPHufc1MuuY3EFvsjkhBgg5So4W+PwbN9R9Zy
RWZ39113GuqqCu03XWwFJE6LB7rN6QuoOVDWKTlV/DVDESwKhRMRyP6yr5LhRs9DUCWToOq8h2pZ
pKfEU9HCj+Ax/j3ZZaE7SD9ElnOZWfMOwy9u8LQwMZ5AFxbs79zAk38chTdMp9Lo/YyYrHbHgjpR
zDkS+fMk8PSwuPaxIHW4uUcXppxlkxI4A5XyH4RoBDCKbdZxvcujBVH34jz+RHA84phJOffAbuES
ky+2DK8fcJ3H0xWwxP4aAplsseLW43eAx/3QFlm1cYcPzbkuqAeV3s+R+dGyFh4CrYeZQ96F0XLx
NYfjEAB5n9/c1XtIUEjj+2GtJbYkHXqjbHzH0SUSqm6Kw0tEgz/i3lu5I59TZa8NwlvJtiKtaMr6
wN/IO4tETfVoFWMJ92cMasQHyjvunauPNIy6rtpv7nmUmHXSYI6cAdHWlXqlm3CxpTMX16rfD/EB
KrCoJ3q4LK6SSkC1I0Mlg6CCazooVVeelpILwY6PHDZm1I4ozdLiGLQ+yKKdyJBbDH+WogARUF07
bqpc6ucYcCQC7aSSCh18kJffwn8pSsrlJaftCCwcDrVA0rHRieKG/2z+EPg3cMibroiDeKHLOiLv
UlvcoTaPmQpwt01LlUnHNBVyXs4Jncv3J+zyjhRRp/n4b2M+xYoC/9kJs7wWQeiaEWiFFnB8ZQkA
pDImiMAcWXOR2gt5ggDg+HR9vQF0vNyROA4xJJyJpRQZmvT80tkxvet2gWjkHJ9M+yr36d9p0imf
rAE5vaHnMbIo+kFcrnuc0YL7LF1rnpNQ3oUJR4P8MQW9q8dzLj88mlSQaoMtRVLoCVTtnCzE1jIM
AyUxEC4vmEYeyqRlrmYkPxkcnxjPJARGCEBU0SnGU3WcVLiBXkN5sD3jXHzF8IPBdiOa1lsa2Xma
d/GJbtliaImvcqmkOKIPu4B2T/MClwwT2r7bthUzeLAojSJLW4kLZJ64IP7ztP3wOfTEVEOYKSOA
kRVlsYjHtTR8D6IXNZVXDYH3DKynzMlHvWH052qDtDBdfGZ2ijE05SodRmAkqzhwZp936OHOjNaJ
GBRYUFEhtwy7SNHXIufZE1J4zkC0nTBJ2ROzYPcHA4XGegQTKo3jfciAd0qE7iDjETzKDnpN9w1E
TSrcFl4n05QLhqDNjZDPrI67V/zY1n5H46L0DjKeicgb0aih851G2GleoSYVU3STArQIeOIKHO8L
aNG5XBwbDAlTWn1ajsUDfy6JoB8CQO9ue1D6p7T/X/Jjr4FMn5YR2sTOLq5o3ivH5yOhjgMZx5lw
bc9hR32fLkqUgGYwAWGBgztsRv5fJZyIO09kel9JRSfbCEs3jZGkuulOpU0Gb4CJ5AK7yuxfKSit
aNdh/QCpnkk6nqO+CKWe25KTTt/a/vwSIkWG8NqRNADzgTnW7T+SRpGnPz0mhZd/Mbc5F4iu9CID
HSP+Wz842PjDGPNQsrKXIxEQiGbmhzSxyZaL6ZsjUpyHXeM2b/Kk3cyB6T5JEx14peIZOH+kbuSg
DZEOGlYkQuxiZYIjvrCTS0XgURI3stv6E0NThtock2lIPOZVY5CUM/Xqmp0uNRYs0oL4wVxFhIwi
nsOF5gQNBOfExflSXByCbE0R/q4TXDWuE44MijAGigs2zzOYbxxImkPTFiC+G/7AFbVy4jmrcRSV
iVXa2uZyqj8u/5k5+rwsXI6oIDIq6HH5zKWyLCgej3vlzzQCuwYmsRwPqRi9PtVp7FTJyloigNIM
tmZ3SXRm91i6n+7CnfFDwsM2cHg7gwtYyXMVC+oO5tF7sk3+T8PxTnkPgZonPV2Q6exQK4qq07Fb
sPQNGtLLY3RVx0HEbwNkgaVrOQFbT3SC5UKGPbdZFzxTjr7oH57x1O4b4snetm2Bzx47OldhJqB2
6ojzCsRWqiqUibZmemv8rfqScMsn0h6h31pTShswAwSxqE+UxD9ZeiylH/DTWACdBSZBYqSx19DX
0QVAKlKAU5sXdoHPi7mddzh8SJV+wwvkuwidb/18podXMoZKDXDrS1Me+cXq7qQUypgM3SwffuBK
6K+cgcF2Pnfs72l6RQPI/4u4j60P6swIp4mxIUQ77ctbgUh0//nuLN7FRNjNjm9uDq5qvL5XDS6s
RlDYiwlXTdrrBEOGsFJq7Ji57osiP/EJ4jT/pal9z1Qjz+kP9H3BXES1VtKhBQ9/O5wQNSLmUmHL
M/pPzMSi0ztpU74W4HTXGyqID5jvyjkKPQKhWHuuZ7ZSdMG9iNx7FC0K5h1gJQVvR9FXdI6hE0sH
7fFaxnpe0q5uDHNoyBP8eEaGpa0GiDrQ5rrS8FKs3Dw3PoLdMsnc0OLOKa+qdrREWqxpsQt1iXXf
199PtnN+iwKNpC086hfDGXHKBaslY8jXKXCqCt72Hs1jHpzEUQrEBzl310ORzls44k1rP/bl1S8d
YeLaKAs3SmpUi/F8F9c7koF6dmRQdcBYtishkJcnbjyVjwz7MzoDCQELgGMUfF4aISyCpUyVfBp0
KgjZaKk+aXg9No5KtTQnEp27dsph/QAmDraoZTDbk3cMnO/F2ogL4o6sB3c1nvSPDR9JHeRHsHXR
PeYTO3uwxIvlcGLT7IJ6pD/XvWklNeapXyRlNylO9/VoUUBjM7e9FvUhAheC4TnLnWrsLRjBcENn
1z9H8Ms7JRKAzBvtxfQ2ZvUXlaLNb2oJLwmkJW4M13UoMCi5UeJxGx78akeRxYM4XYCX2uxqbRZd
ZQRpPwRD3BmjL4Gsha0PLai2W3CX87qVm7ko0mi4psIp4xTmvo+Ndq3HlJlc+dXkdA6nkcJ9/AgA
/0txOpfXKOU1mbGnLoFaRHAuWWneg4PHWfzc7ORi5Gb5U6LBZmc2s9/ZGz3veGs3nGLf840dj7UQ
bbYU1STC6CSV0i/eo3Z2z1ad3JZusNnZs7PoyPI8FGdWeJH1P+CIJ4yu4rizUx+rgvq4CK60+bVL
LbWhMKiaEVzvNKVhPhKE/rcZOTM+jw9NQb7zJclDANOOUYiQ9R9yX0lj0kMp2Uudv7038JsSwo2B
H39ctCwh9Mf3cpNnuiyQRapkT0v6fOj4ySe4hyT5GT2LwcNWC9MMXYOFIxfNOPOV7P36mY8/f3Fe
wO3eXJ87oEobHOrW885W2/vN03/LAbxdcG7bF2WxbeHOfAWdqD75UqCqln7Ta2xX5xPDf4ZIhp3M
eRVs2Xn1EgIUlOz0Kmmwpq+2BKIIRcCRuhFfridvrl9XHAnNzMYIZcdvLUFPrEuwOB+nqQrU2ldf
rDlG80+LyCXjTToGZdw8ys2Y5h1KdJTFqu30L7Lh9Q8hEfV7qulg/rKUEkf5X0ZJxtLOtrqflcfL
DuWbf163ugulVfZdRk5WmPlg4goZveY6G6DR1u+oHhJ7aiJmpyR+UzKeGmAFoVgmhdRggPyesFHV
cFWmLI3/aKOtCLizxpV4NvAIMjn3VRT3eFSSIrJUrRalqX0ui+ddP4fy/Y91bBtTQ2o2vtLDme4v
stj8RWP6D5lGI2+70wj9D9LQRu3dwSiif8FqQCcz+/EGUX1qfCZ30RRY2iKaJtv5sMSmRtG7Cjg7
ydva62TGo12l5vCe4BpI/nvOunihtjcEWq3ynTKV5plNmNcOFwDHeCdtF43k3hsT/naSgAlISmq2
RKJ4kUq4/Xp4cz/EXDOXL/S6kJeE0VpYeyG1BlrqF0zD38aQ1pSNV9nZefemhfwglYUx5OOxV6kB
15Ccpo3XmwE0kFuj9vFIhKfmQ+ytyzNBHTVO0C5LyaLKsJIRDhVYbZahpqlFGHy5uY8kBK5l/gQ0
Bexx4RiUpd5C6+n47HBzH4tEurnv28HNIW4udyO9ERIFpQRANXrB7ozJAJbdfkqdeMPpX4XeOjEA
D3wv8xDFwb0mNXBodcU3dcOSsOB8vah+wdlNcPbApqzfr7HCdmwTzIntHud8O0rMNthdyco3qAsU
8zwqLJJeGfApkZu9/FgGg137XOC4R1DWsD5rT35l20GL8v9hWWMYuGUvJO+BhXomGdkdei43+KF/
yVm/hDh7IfHGjA2h9hI8//p5WZlw7ZUMt06PAwBSUZQDNi/4kKT2odgGAHKSwratHRk4ywUWrbo5
XiHI3WFbPa7Y2emdeZDoSAOOPdzW3IqCKqQoe/yXY1jwdwII6aqmmR4qo4o33Xb4FmrfcXdbY2mC
BGQ6hH3mnHQAkXf/mh0GeOFNV+uu6+jr5NzCF2TRnPLSFww/ThvQJTixET0x2KmiRpdhz+e/WJYg
Wb28g9sD9PhjKTU0bSiXowrOWISFrxxMIVPrAdJc0jYK2VRsRlbUyUL58+cqLB+g7p+kaAttfGgp
jyybKii9YXjhhdQh9q979LuNYw7lXxJVvgrnnlaLhWc7MnHR4deAmSOrKdFZQB13BdHmRgjJZxL6
sdpOs62WQw5f5oGwh+EVQ0MqDo0Tv9h9hmxb7rG3dS56gOWxwPIvJDWgBOo7yxbNS9l4OTffLWil
F5/g2Zr8ouiuipBli3u/6DIixFboX4my9Udm5b0u3WQpWgO0I+S1g7PcbdDoRzcGdADxrzAjICG4
7O9E+4tA/QDY7/MgIVYKV0LE6P5+RL4PnuRYjWw068bgrkyecyZMiVbOAYRFHgzHH8Xz38OKe7eo
Wcbw0crcPs0oCRacA/SyqW19Dy1Lr0XGC5jgrYTyTqd8xynQkS+s682U+MaYdQgkrGeWRmV8vUxx
Ufo05mystdS8SreoCK830Pm032eDuFTAUO56QOm+V3PEx91cFBCMbJcmqp5W0zYWT+ZfhPlPVhwi
JvG3PVXf7FdOLqPXhXl/mpjjxwt44lLI3MbhMSBPW3TJmw1QASDD0hwslek6W6Hip3NGTqna3pcd
xuUVirwcGMf2CF5uYOahj5vv/zT3jcRK2RD542/Np85LFJkRSZX7kY2gcEyDzpErgl5uz/7DbbDA
fpNZxdE3PCod4tWmld8PmVPKL69/XQSNC9wvM/W23XyJeAH+vzZ6lQiS1zc0S7qsweQYtzBwdT6W
VX/H/WKG0GAPKB7FrjuzKp+3TwoACpAE0GfK7mzjy5FECVFaXMkOThVTOKLWehRJ5Kxy1mbJxqwj
byvIhZSZYjkOdim66F6DzK4QkGnu65DVhMEzUQEY9bX3GLFlNacqbFcPAVIsZjDbvFWXBvuazFt4
cpKMuhDuAGkd0c+Tkl8Urg0h4O6K8Y1Wa78vGtDhs8nMo6JwJJ6OJkLwUEJXXEZCrU2ZgTUdwiFX
x9sO2B3DBq3yrAjg1VGVrH+Ed+PlWHh4z/NzwktyEz1+ZS4zRwzgQ4mtiOuRDlbwjCl4qFF3aCOz
ADfwHRGxDcUSuMMTAIEneYZi3LuQRVW+2/5BK/oEdR1AnD9k7RALNJwMU9XT5xb3MNNwtro3TNKd
w9X/uYR+0ignVftWqj5K51yqiQTapTtZR0pzyOcqCG79QTXWGMbCG4WEqpuP2mviPboETjndxdPu
RiGzJStE9DlwR71swWy+qXTHbZdXaghi+AlSroc58nFiEXBxw4pfm8JYPJ8fhcNlasZ5HwD3yrid
QRfVAzXYO97sXD5Wj2Gb+DjLZvohGsD+tOQ8uCN4oLlQDOEpFwMmDFlrAGzjSHuuJ+8kDhN2lYhd
edcc1xgHdpPdXCM1uxeoDMwHlb8FsMDkYg0wPwFW2iWlyLyQi3YMt4hSFEF9otGRhKNsiv4H5x8x
bZyvBNJ3q+bIuoD+kr61kbXiUGe710PPFydI1WavIhkS7oQSAj/jnw8pOd79UKEIDnONkX9GcsKh
8VtBPml67BS8Ul87b1zvAyZiW866hy3oXzuLoNLprVWqGp/JI7STHIVFiEQIq2S6z8T8GM7MsIOB
gjcnovXWT0cACu/7CfkuxOeNoWa0msBUr5eA5Y7q+TkgFqVNrWuSHI/sTL7K836zyQEGKg3qt4IJ
2ywrKP2XrJzzAvJtfebvFqKr42VQGJhUfgPD6hFI27AnPI+UFApry5VnxXwmpfKuSwyXTb3EvyQu
9ORB1oj5QfDx3UJAAYlR7lKrw4PQAW49KUiL/RxM6LS1aOy+Tp4PDV0ZbOSsI6pW7X9L3deK0g6O
XOMAyvpIjpTWlxW9hxJP/GsNXntgaqEk3JQpzoT8+8ebgBXi1XnH5N+kS4nuMcR+QngdahrR0KrY
QHj8wNsHAKnSx29Wtxdhd4CbMuxdUb9QWKgWxfiSvh33vyhKRmPbYfhEShtKxy7RMbUIr1NCb0AQ
95Vt/PAQu/Jqml1ClCJcqexWniG1Aurbf1aA3EjSGxPpYPo9+iF6vm6k9kyLlfBZbfE++gZ+a0by
DQzSOy+c1KGqXTwWV2WqcKhuVt16msgMiO7Gmvkf6YbBPanpwLGfHLRBzm/gtTgXHU2Be42iB+bv
RKRm+yGPJNJwjR1KyBtgsGEvGiTbQOMFMgfi1ZUVdmLNSIODPCFfTFxcrZEeXEHY2vv0BJ67PdbT
C991/LPrwKdBGNhdAd01iEpXNrFffjI52BE0cLR1aYFFaOZ7gm030EomCePhk336jbU4hSlCwttz
ZLD1yFp5ur95Mg+A66UC6r8Zw+caQsMITdhz/z4wqUsI5kNlliyJxUCvq3ydDl79c+py8ST+39qb
CPKlh1E1r5O1Rl7yY+Sm2guj8di3Ate5Oa1odGe6uBQZdCxIQukUBrrMX6j5KiQJKD+k7huykkwN
zokNAZGFDwsj5z/beay3YGu9snvrvxuAks9T55QAeWNp/nrzeSeRqXPTHMI61n6aVbuntE6JD1KV
rLBSjqA0ogmZRXNWxQDHbOtNnBzVuL2CJ4zT2jWDL+pfPPefo9wKi1VMJVG73KVDOXb2WO/F8v9X
A+l1JP29PSqTqMWxWmwBuvOA1l4/oy6WuBtvhmqZMzYwz0IolwfkuM5aUj9ck5syveVaOurMc7WC
JavU3JeMMh5kz2Iw8Nznq0NK9OYZMYsYipNulyMk3ItffOko1yFn2iIZ/F6Vs/jhjGSyypWt33ig
4vsqi7/d5u3V+ZWCgHJqORu1FfoBnFXhxGvKhV1PKaL9GEbKKYH3VsA8xbcW7YmEpQnnWcqzpNkJ
FdMDZ3WhBHFXOjQe/VMKfuc9ZCziYuv/eWqCn1FTv6CgPi4pm90DJl7udeh8rs6KVO5y/q4eiYaT
pKCy0ktU1GtyV2h7Zb2OhLSXkUCivZFJc4+egSzk/1HtATrpJ7CMEv5s3NscrUj+nQfaJQSYHfPE
pRm4iXnU7wUWsjZTMs8O/E13crmtKWzx5DmMMx2MJDR7wU8mqiPHx0e14hgP/f83IqnWFgWJI0/Q
f/8SKqJgh0ry8HvqEE/WEaMeZQjvbU4p+ZKUQ20kkoBA6iUKz0kbrBspURzLuMdEOL+sVY6QS6Gm
7OxYTaKYjxiL693ekwlmsuuvGTMghodA5GFAl5SsZOV+0flWddLtz3V0FOHzCdW/9vGTU4W51J4z
yltXyXkQJTfmXCkxOyDSBxFhebutQqTsKB7QSmiTkhz0+1CXJKkuaETrkzSGt/CCuhYZ2s+Uetjh
9xc3nihUteFl1bQYLbCOoudswh5gLHQBkXRvksd9uAmylwO7ZXtnQESM7bhglyzUsYx1R04Rs+T3
Mqghf/6soyMngQl8WduL7Tfqf0c8Xggg17shwDmrB5S9nYi7pcXkuFJpyg5nB2xIaDXgLY3A3gtT
WmYMWrcXF39jHmcC3UAVbPrAlnSEUsH5QliG8DNk3o1brWG0OuHQw4QHbpM3HY3S+Chj6mO2QalP
oRLOQAkgIMbwdPQ6JjK4djD4uiGqYxb8ug+N5TaGA13CKL6CmS52AUsGTNj54mfBbxEDIxF7xmUs
2BhwD+tN0dzhMwZ51PDiYfGLalZ4FOQIk3aKqOfy3XVyedZrLtMGpqZfIbF/2qyaqUE4L7lpC4Ux
4wSsKvWUpt1j9DP+e4Z4GrWxXDJ+h4N6ndPLYPtx7KzoP6pAcl81uYBisTyiNgQBtWhbm/4+1BSB
aIehCe20WHIxvZu0KbCmm9qFeJDLHaW0s/AAhE0/y1ewYJMD+rAskS+bt+06wNHFEfXFWEr4JnZY
BCXDXv6kBeJbmrq09NJDw0T9hpffEaJIOFr9RzeCTLUPsJYWJ7JLCnVn2n2I6HlS2E34XTc4XpAJ
7aBzOz6PXRAE5hs5yb59SrWTwfusf9Nr2iEvPkRtu53WONCDvNRSJMrENhr33iknxTj6HoBzBdqN
ecNd2BPvmNAzzBRoV3RZyMnNDB15b9J1SmHzGcF0KlZSKQlvd2QhxDCk8ZZvD+ZOwDsVa3knaooM
Rjsbxc7x9TLDC1mNsxmb/FxARboemWhBUZO4fDp2rNzBmkMkVkOHQPglLO0tTxlur5IaptVw17wH
KUGH4igv+d0/GyGnYaIp07bBKTef1ER5aj8pvu/gVMMPnR0ZfdYJZS047S+RGiRvyg5U1sQYHnyN
jWZ0IayO9vba3FnShKNPN5ilUZg5/I1zp/74uunYrSJn2bvM08YQx00HNy5tnrmHcWg2ww9nVC/y
+2PKIBO8QTEOhdyqbjqFt5isgopt8tx7YNUp5GxxkpF4TX6WW/IYnj3Iw6N5t9WN4JOQl1u0M3z2
jQx1hHQkhu0g3UFne1oOovaamOxVs3oBoBF/FDkyAvpPzEbApuV66LQj2eHpPh85DNxHfcONpzWn
psJHpGcS6OBm96MBoo0DbrR1QbAYHCMerPq9ciMd2NyUchDZGSQgMmXuQSabQkW6Z4Zc27VRjMvW
xL8tWsNDCsNgtMz1Rn7Dr4l5okuVxyn6q1LahCM82sbgxnuw8aSypJv3jqEHJna2ONdvdicC61+I
ELabXNE/VqsvYUVj07dO3YmTRIEJOop7sxxcXCKuaHCHwLHEVsMjJNqm84mBNZ6usxScXIxqSqpw
Re7zGHy/rxmlMccIwHehUKvGWtMpROom3mESU7OKfxETKvLAKHpvFCnG2wCBlOaiKcOv907l3oHL
2TVgh0Jc2ReOhX+U2B/2COoxtT8um9nVMZt6ehX4vNA94tjx0V1YnMefDn1Tn9T+SxPUOmIAGlHH
N27qtTNA0vys4piH1Up5WA+Nd2SYLWkhD8bCUaVS7RubxzWmm5Ee032P1GgNySUINczZBDCBACg2
/97KXrjvwd5Lq/csrgyxtVnPGHXfAaiPhyWcZdPnz35A7tQa/mo1iNWoYystcplI3rK7FMV7Pqb0
h3hiGvdjOh6PcTDwBOO6Eevo/4rCf5ygN0DRKH6xxYmTWAw9hxKbo3dczxZENw+WJlBj82MB2jJH
A2ZazsJp9I3HNK48ryQhhubxcPDuW09hd7dLzT6L3X5z4luoCpJ+HGzqZ1t9/7EeCMUiI/0/q4Wl
UApxiiR0tBOop867ljubQNzwLvJ8aXJ+KWJSfU0gS+sh0Ns2WfiX+CiR/NPo7HTpCcwWOYzNmmg/
Hiqwy8eYSK/WuwuVUbq1/mVCZbPp/JdcKJCV+r+vArQEmU4p31Pv1IKR+ZmjN2Jo2tmwagmSCUwO
hLdNc+Oww0qRc8iLuq8hbYSo1AILrG5f6vyn42AdDQEo4vnJ3aODlRbV1nQ+bkCft7e5wAFCM/bP
nbaO2xDR+m/oksoq0Wr7+tn1zMnrIKUnO9cYVkzkovfZsDacMntvdEvpy3o6QKBsLcNQPd+D7YGD
0Y3T5+LXhDS/n5bWFtJs6W8b8TYBDa2qGoOiF8wSRBf/sEE4fE5eW/Nwptvo9lMqkfZAe2zV4Lm6
KiH4UE/c7/DI3DXdmy9hjYl4USGtwE/xNa3OHKUiZ/mVmgpuQ2WXM3n8xXn4giG/KSfqYM6wCtcb
fEREOOK+Qhp8XQ3y/g79MICUTg9zU0Fbg6D8dWH9UDtT7/FFf6PQUb6TyGHjdEdE2MmT8pZLnQ0h
QsCS/h9SJg3lS4GtdJ1MHjzYS0JgdlNp1A6azBb4+k9vrN0VcqzK1GnJICZqAX3+b56grJGWAkiX
036/bA1jzZn5pMpEkflA4rzpLmnx3JNaVN2+ydY6ATrkSMtMQhtrVCPb9HCXBubFZIQ0dA8RTGDI
rRqZBhYH1LlP6yBlSuJVXCT6gml6SVINSawikkxWUhXA9dvu2qweVKEPjLmhmfdwBC7MvOde3iaY
eDPF9f3OC6+iZZb62SycAdtNk5qfQW2waZ8kq/OSf/g7LazVYa0uFjYOIkGY+osZ+QOk0gFSc238
jogbyUcSk+efSyhWKp+NTpsqQZ1l4uo4LPUR99avpxsuoR9yGxlJPyZM6pXdPdQlw/k2ZVTLBaRG
m1hHIr6/d0nKINQuqLTXioi1q/wQaGBNwFzZGb29kAEcxdMvLWFeHWQsLkxJECxR+KWO+Xdh56hv
5807LIfcLrQXAsB+njxMfb3r6hk59EzoDwKLYen9evc+iSOtWPwOqgsrDtorN6RlX64dRGWRbkmw
OmL0lfWAQt+2gyrIcig+Z7zTylf+Tji3uNYBYjivspHFQJyIcLMa5c2Ic+CKPSKNl+7iBuN48Ocy
cAGXYEn3KodPdmqPomMj1kzZALKQhvAPsJskvBoV5/5zRyUcio8bF4UaDQTAoU1bxKqrR5ViDQMe
4cPV8f5J2iaZPniqYaDFL9TnqkLnOwuOOaTsM1hdV55CdFtYNwdLqQKhPuUO4RfFdqZyI8hJczeW
vcWmGRUGSBdTmfGuDL62PbxDfmeEzKqa+auDFpmH6vpW+SB2RHj2tNf0STqrrsxOXkh0FbgydepB
3HJTzUbbj2LZY7dOQyRmK8jtbrF5a0Itxrj6S5IF+aSk+/MC1CEb3K/Jl2enoDXFpiyJAA/lpT2f
z6QB9GE0IHVv0j+4OK0RAlLwf0DD5W3R4sY+EA78K5fE6Vn6j7Hmd2+QxAQwQ4ach9472//XC0K+
W+KyF6wsIJfCzN2ny3ya6Mo1oIbq0kI1x584keWK7oeAMC+aDa/5tyMcN8viNXP1Ko2SrQgLZ5vJ
sLwBxXaLeocxl9pguHWhDaMe6R/XcM0uRWFJ7BM6FGzVSO6ybnvTFeb3tT92sk/xGl/9Ni4ZoHj6
tBIJ2iriTeRe3v3bn8t4cw695nG2RTf17Mlllwyysx5NKeh/+rgWRwOcYtmCv9P3DeRqjAUElPIm
po1kFYGQizgcdzKIP+E64b6RCE4RwvIJdsjZSGOe6Ai7uT9nJemLNmm7Uk2xT+ubSURXbMByYaQi
oWz4rNexMjkSiYs8gMz9axPdiCZsiUV4fY6fQNN7Kk98PBn83s4eH6okLJmP9G0d6A3brWcOkHDd
c0DDbyUTjV+/i2HSMp6XMsBaeP8fE2PNyTkFq5Scd5Aw4icm6aYvQ1MM/tpXeyPu8LZr8CiO9JEn
BEZTSvnRIxKyEV5FAW1acOgnpaX5jrd+Q4tfZ+c2OdJhWFAJjNBzh2ecSMqqfwMHiXrsLfdPbqMb
OqhJBS351mtPZZeOZfuj5FLuJS6yVnMoAf/iVHAPMh3p2A3+Fwqdutv/7cWm5BFu3to3NvkeVzqf
STDguCxBhYHFRwHzJS+6vFmQ30U4vg7Q+EEMqtRfacA1O7jw7OZNrBSM0Sl/4o5GAucDz4xu7P13
4zm/bOqXk5u3yBm9N+poPWJTijkx4F9LRAE1XuUZMJYGPHCWq70fgU81PCBoouXbMXZfjkcItBqP
msAjruLS9csV9TXVVUIGNeWKpCA3bKwIquFqeBE4bqBbN7hvuSpn99FpMWRUwW4NCHKRzjzJfDse
ma4ut1o30jG6b/36UsnNdp6Nlk4kCEhC4p4nzrKC3gzlaDPTozXr/m7AIyy4pyYNY0iQ97u2kbMm
Ki+4Bj2ZVW69DWco32e2RJh5WkO2+701T+w+7xdWP0drDi7AUoFXThn6E5U5oEfZ2ZRZ0kBG1OhZ
Zg/v2bPj9IVxQYrOTHsTMA9GJ+6Q8H8s7gadpBt8snp0ir+fgJ1ZiWVDXa+jkWtpgMZ3glKuThOW
4L9YtqLjN6gm7ycJOVOFW5IK5iqHoWVE4NpXMuQdC1s7tWBho8n6PPwvwhvY3eCd1Nr1TBNlX0zv
WIyzpmwlXiZAmpyY3wwPRaR1fxXNnZCP3nmjobObZgRoBIVgdlNXV3CVgrK4AbG8UAWaoyev+1Hm
d7lJhnrTMbXjz4HInm31L5LJBMwylLR3vEZWaIGuHN/Zk+TdDd15utqsvQil/adtXzWoPSZMYD6+
iGzzf1RI69l+WxmvShY4LnDMRVzD+Sh2QMSILeKFytAzIjUkeNqSUsPP1MVrZukOZw5iPgsF7UxB
DTocS3qRvDky0LVgWuAnF2m5CX8x2pVBiwbT2njAFktgGmz/jJ29Cf1DaN0giyw3OomvKz8W2PO3
S0UAVkeDTSC3TfWPY4KZQ5jw9rHXbYjYlZ0LzWSzYy9WH3zKwUo9CrCpsnRZXgjoLS8mjdMUlyxE
o+wM2ORyRA52ppF3hLBTGmgtZ++6rL8xlxnXXiwVk9rtDonw//IeDXIzWkpoTHWiM3bF8EAP4eju
7Rn1MVU0dWWaJtuqW79gVAaAdAnu+ffkRwCJ9GquVclF9tiz59zkSfmhHUHW9WtOLBBy1FGxX8ya
B8plRRIGaCA+u2aakdgBBHcRJQ5Izr5uaAcyb0LZhFGzDbSWdhqO5iubtTfNI/pceTVM/r5lCB4B
dyzRm9aTNNkjIeZ01SjSsA6Aao6cf8TwmzNcgOl5UMA1bFMkpntl9aNfVJNdNm2gveSjMJVf/a3c
swVaUPTMZsw6BjWvCwdnoh5gMUsWvZ996emRDNc7KJoX1IZjETZdzJVg1LUc9Wd8YFsw9ObM551m
V4b3W19JTZ1G82Kr0/lmVsI5nNdmtPRl5e/mBMqMhtyokqeCq1FVjChSZsjq/yFkCusU73On/LbI
jH6LVGffquqa2vaCky683NAKXvmVUZP8Xi17pItQYUhxaftAG6j1Zj1/sjbUs04gy+mHgLa8c1cQ
Wm6V6+wraNQ9bIzed0RWrWpRrWrcf9c3Qo5eEw5GWQSrr/jDY/xiNl2OTqpZd+46J/0Ts+Lp5Zfl
I3X9FEAOnLRPIuJOxZM4XF9mqp3Pbg3Ky+H9wk6B8yBpHPKRw9R62BQLZV4JakDgt0MC1T2RFumu
vj/+SCWmEnncWdg5ozJYPI4QjHYR5es+aojGS9N9QOZ+2sNkqPIT74+V4LpUj8JXD75VbLOy9Ffw
GevnxgCAQ9YaT/bnGbE4NL6xjERK2UpcjUQz0TcU53GVMthMeyu/mHZFLpLakfV3y5Bbl5XTOyh3
o7pBx0SN2ovafsLcqxrxfoEB/frJEyLXMwj9HDgAodLEHI/vzJd3kPJg34bfcqq2AYNcEzSoXtG2
L6W0yhnF2Ib+VDTOtJXqnWhfozrba+tMNctj2QDI/KdIeBGbFvQL1pnkatan7/BORLZDoUeFbSdE
onsbmTimX8wCBCpxpyGS/3AeZZTtEtZM0B8DKxhq8dk8QVKIoA35OxC65p+SjSyz33Sp9KK2w6cF
aDggixriy0EoBNZWqpPDuol9lgRN8X7BFPhFff4WxV0iGCKm6zOdVfTmAv/iU5v13VYfF0ArFuk1
oYTc7FGHlUZdVCEvgiZLjlDcepcqYdIUhEQ3SHmM6w4V0TfEs99r9YefiAMME+XyZVQXMNL628lM
1tI3STp035L3vQ7vA2Pe2mWVMcdif9eTwVKsG0thUsSfvZn3zo5LPKAhnLw9FzKiIV9DEkG0G55L
3GWfiKAVikXaq1mpd7VpQafl98tRdfRriNFqrzxTu0FsiHT5X6frXVA4KO3lK33VVAJBEOXs58mi
8fBko18BnlABTwMBrohzraD4Xx1MUSF1usRYb55dvfoAagzTd1T2XPOfi7l8rqErBgrzjjtMAoIH
3Xh68Sk71fuNIHUjbmTNGImZ15rt7wMJtWMk8YcuF70qL93XJC4aIwFB4VD5CFNajmLhnP4kM3g6
pQ48x+2KbuVniCJP+PENQWWGnNDQo2STrogv1EuGOLjdZbEqBuVPkomhsup9IpdffjNK9WsIogZr
Scn+qydN2HmhJzkcGVH9Q1k/qsl5yCG3zZjv57EoC7LwPBgBBFGqMuI2Tln9RFnVS7kyOzeG2gu6
IYXPDYzStJE9Kd5XVbBsf6oYdI/smNdW+e7ovcFxhWDungZm/sLm/0aWrwVTniQ0T87/ttKb/wDp
mENkKs8HE3JATEgDMVYcrjpUNEwEYGhUMIvvlu2791bQHykwdhXjqBSHXBbEdBXv8PtVaPVqyvEQ
ALsFl5gcxgfP/tG+1a6PdDVWLYSX//5w1iS0fASXSFRA62QiT7vPdNFyGtSWRJWpE1U49RstYB13
6KpxGSt+LsTd+30PkvRgxWd71n/XBzL6o9oGNGow5mGKP93G61WecBfgLPYmptbqmbuq5/GZCDwI
Ri4TICH2FGgVRYkzdgkVZz1WvagB6uvoIe+lTgXFvuWvjPo9wPn06NKG/ifA+sXX6E68BiBEqKt/
pGHo/9+J/QamxlNsLFxPZZBoP47X/qj1IxSC7Pneuczk5nFnRlZVP0EuUwV1e3K+l6rYVPw0q3vU
P61tAJ6rLTKh+VK8EQLVPhis/zXB5ZLuxrMkbiDHij40Xch97oFAoLo5TzLtT3143HAZMoICJxRH
nLrPq+5FeoIK9XbQFeRcg4gL5iIejPOsfa9oXgRxaLJxk2Bccew3vODGbZ7cJCPLAaZ0/muT20Z6
Qvob2RF1OzDS7ZfGaFWBALaxoROi3YMTkn5DDgoAc1LiR9gNGeoYHHBDss3D//ABMqaZ9N5TQUw5
tjmF2M7WIjhA5dShDB0i/IB+pum/q8i5jthB1ME9m0I10vrIC7YJFxnEkRSzZQwzz2WUvgynpJUD
Ym4/ZkmnKnSVK8XFkKz2o2+13bmuDKDyS2UpgW9w0uS/uaDyBC6Hv5KoCeoedfr+QgS+ppGHpKLE
CtGy3y1J8JRUH/1CQOmKp4kJpjN7o9tWi2ufVroG9UzwOQagvCJRlzf8VnnDKkk+OEXPmPs83k49
RS5K2omcdnhC4ISD4a18u5/ADFyEEynKqcfG9oZ8N66qgNXEd0+TjjEwwwMLF6kJPD/YzvJNNJR6
iRClu052d/khV52cVxJJF2k03QcQAGngL/i80ALKR52/pb4oCf9wpNvClRqm8wsM73iU0AZ04EJW
AK81vQguEIRFIxmXbM3Bvg2ICkKHWF9rhv8O2yyLR+ymDbgBqBf4DGtlPR+ydjjwyIIqrmpUyVCq
aaBH5gQBVNLLkfn51c5hRo9nNdDDmO1U+ZCKoAMOCbeg4Eot+ZrHERjoIkgohWiAZROkWOxAISPn
iTHTxFXV0eb8cqO+eRjmQIU6D706FyWjIplqwj+GOZ8jSLRhweDgIG3KYoX/0eZYpd5wt5LV8YXX
m17XBi+ClxprePozI8vireZYPLqoWRcxxtqHdJ56lCw+FynZzu8C7APrclnSxwG47ntSnFHnY/oo
5ZFDOhwFE3Hd79rnCefaYb8V+iZ3jspoBdS7dbD0Nx/mzU68+CXOz20ZweMFTgxHWV+DSxm+U7Y9
UtZyONpb0DEm7ElPgxcAKMcFCWsAMDwCrXnE6Jx/hQ7Zb3Wa8evPB1+PYi/nuX476w6fligfG3e+
ezBByBYAUh/4rcyXvsixZMt+0dyZVLMAOljjl8jtb+udk8BeXVvGIYbA9DM+SGqaZ0YeAEDlGKFi
mcUcNHrMpUa18scqGbDH5BpnMHtl16sMv+rc+jkRdHa3ogb3ldM72b93Klff9ocfYQ2tRQ6Uh3lP
IvMYh+op7WOPFjpHq8z/ya9Tkx/VMnsbEsUMDBePYovcoMCCVJNqgqIvUxOo0DB0JEpI5KOHmByY
UEvQWvdOOzZPRCmksp2PZ1tB4WbKTxSMVlxkHYHV/Rr7Rw0o3EzY8k6PW6T8i5984f8OsP7rkWgb
eR+e0FkjaPWUrklN+T6kcMXExq8ITbL3Zx665PLDXWFtKaa53PRRj+Hgb24QtxE64q5vfmIhvVnI
UOgadvwSAxpmLwmNMrkPI/zLt2xsm2UYfY8GCgDPf3Z7NFnFolrxpHeJsIYYX5NQSNrFh6RIfpnU
MZeNe7xRZeMz9ykuYWgl3RJG/vViPa8T8LcbSibetMKqZrCyaKTh2Ms/9p5IbrVSz4dvcfGT5WCY
dvBwByiVDiElhFUlT17z1Niqu/R/UNK29fHl3QWuKwb7t0GvPvKvxVpRy+4ZjAJF8jyqGji/ZHCy
bdXrjp7gIfHhGsAYaI/MbTJZ9J1W77HQ2qIsU2nk9ifhqvA3l/LP1VH6ieGaNVXPGOLkIrj1g5Iv
z3RWwtnJWdFT3Tu0LFKf43qq/VlsyG/1z6ymvUbeVbC3cKP39WxcFOe5PGeF8YiNpd3FJUPpnfiY
iRCBvV38IGl0zONfKyR+ISftES/CQIonssiaiBfPRToSfmIs+nKdHvaKjMvhIMuwjdgJStQYdvC9
vKjUcFHVOxqE/4PtcszP9UYIhHKDH5tIfarBOsnL3v4cLvUwg6l5ErBbCuyudglRAIfH+w73ceG6
kSR4utvXttkn6qkBuZsCOE8Z+V4JtJ9dh0RzltMRQMdDhNz/XY3X2EGnAV+uOPibXevKVKSlMbS0
FRWdFaDX6rKwvsUx+Zl4wSTQlK8s7c/iUd5RRI0eyHc9O8iGcVQs66dh7qPLqmHNSgEqzzp+xDTO
S9bb6QJGSeuvwhStAtinSa4er51Ryry5R/I8ARWZhwYrO+9DYdj3zUA7Xkt9zjIwvSX/f8jJHzjD
5GS/XzugTDTpulWG2joxbbZ3I1tvM32aLZlhHBTEyREoW8qgg0rSy6yvy+DZEYb0P9r1UGwMJ8EC
cB5UmgjmlkwaE3V//HQ+Nl2DnIVMGzbxpGH+M1RHM3TbZYFjuWwKvKFJcxpO4+mqn+frBGHgbvxF
/Nyx5U0+EWHn3piqtq0F4c0Us9QpIzF8n2HBmmZk+8gxVeNlXhnxoP59OJ92nL3ni9SLO9lLSp00
QLkaigkJIIvbdLsr3OuL8vj+VsTWt4y/dfkL0+bMPOM1wwBIzXq5UB9TO1mNvFnDlnrdaaLtBeoY
DUZanap5r0LaEeY12ki79u5apn54YPLrs7w4wAQZvBGcOG6WGJG4VJwhSyw7v98bajSIXk167uxM
k/gYeMqoVOHiMc6sGCRZEjvwZneIzhQvSv9vF4XCj1OuML5Y6wR8nPpbJ3R9EeRRFOL0cBjj5ri6
EefRKiWYm7xUtw36+C0lj9nBrsQyh8jbZVc66IBZlkHRoFFUD9N2k5WmALqMpH68IY1CWveFrsxs
RfMj+U3H4NZPl/N6fXbAClElr3lddV9/SFl/EBuCm+8TgVe/se3YaSRPszsGpGRCtjB4hHIOZFmW
RuLpEyARo0TC50CKASK+BhBKpBxPj+NU1YAOAdPkNHb2cHpIMRhZcH6IsXAb8ZPyVdxBTvQdHqL8
BJKFDGoX1d37X0mL7L9AnEHXvuGkDeYHW7qFsB1nq8GShjslvIBZ9s3JqjjCPLxwwMdQWLEJ2aRr
osw1Jaye5hbOU2RiVnWaUqUpD2yKxROj4IkvItoKjRJ7E85GxcNzkAqVlO1erJGp/SjPaLhNgxxI
gRL+b2nnKTsTaVXewXjMOFT+N70KL4GA6c5orAy8qCbVzQJ9xzbf4EdH6FG4WxLgPdFuqMZAdjdE
rU9t8v0jE2DxkrAQG2chr3+NZv8Z5bKg2z4rzEvMEq5XrY37TMRbdWypoae7qDgBqlgQ78/4y2SM
V384uY39UaNAbve3ui/6qnvuijI0KWWLa8qpatE4HNUtoCE9Cswei3eqo5odXGPEY85vk5wX0Y49
EcyQGZI63x01/nm8A3VRDmO4VyVt+pPXsfnWfbkrdyjLWkMK5XXj2GYGtAqJEUq1LzlY2HLeNrWh
BChGJZDn1p9VL5W09dbG+TX5b2HJ/yTWlp4B0s+roPACnPuKi8pubIsYYhLmR0eugJQIC+MXc9C8
Ytfy4UqoKWqWzQ2j26EFvtdcQrNDUJCuUN5q+EQlfdD1AyhI2avYvqivi06QrlKHdN7j7Cli+sJB
aFfPntiFT9anhnfQASGBEFuR+B61R7mZvlAiyTSgMHywNsx28QPVg5aghy8jbqqATkV1xwT/wmJv
I2Z4jlIdD+qhv8YZDqpd9Nrt5ZtcpnYtyDLYChTTgfmlNTzWidW9xb76WZjPbnExX9TP8p6znLAb
vSKT0tTs0zivbXD8Yupo5yVOl2ecCnjGeqpsIOXPUZMUQbaLsV2Oz9jJbEN+4EzdKBvY8pZe3VQG
gal8l9HwNVms8jSqBq+rhUKkXl6df4xKwoZ8TJgJjFS/gUAIXQhvbTpDMJ0Ur/ND0NArtllx0FGa
/A8sm1ABmfO1uj79n/Fn4m7bV5dRBOPDuLGUuAAtJg24AKD+VtxgdOpxFr3iGAhKwKzv8q8fCkxf
OS2xj3qTuINgD8aMAqZ33JAfjXC6hFUWMDvadezTVgT62xpuh+TYmxgmVp3qf4SRN6yYcDjjqehs
Rc28mEYGbX1VJEUocP28T2P/i2bq4hWkMAQ7bz9h+6BRQdqpgc+L0mmP97s9rYJtZXGPh9SncApG
6KxZtNJBIX+FdnyAJVY3g+Vt0TPxscy9qtSfkmIgaOTMBMwcaa+ZB3eoELP2PjC1kA+o66P1pAhu
1lUJhhZ6LBPGiiQD+rYNt5XzsEb+zTqm1nc53Z4haT9cKTCtQeJDkiR/WIcAzNcXzjfP8L5sNK4m
uyPS76JFsNapEB1hD3Kos12Tloby6w4lvlScnEqKyDcX5cslOv5d3Iwul7qJpS4edkYqIiafSUBT
sJbHJRarGAQpvMgWtvotYwY9d9g1nhvXz8UKLVIE5JS5vQuCXtXqIk8EqGYmH9uC2WZ8Vaqotu15
bodj+lLkgDH+oAbGaqSgy+KS0s5OlC/schTVXHrf7g4kxMNJjU6G4IzRo/AAidP1GQlT9UEwXMG6
5pMcUC5dxMCNeHfSXPAdGkzozzJbPlBBMNF2soCUYh1g1bnI6fpoYxwOw+1eNlHLL5seW6fGc9b2
S2Cmsr/pPrH1lETsWDX1x65zVkFok5oXfG98iJWjaTeb+BnU77Q9Kq+ss9DWe4Weou7sqYZPLrPb
FjQ/feZW6SyZ6bE3manuoQ8DBYtFfTJZi8+FwodKHQ8/Lmjg+nk+02z1Bftc0wEGTT+kLbDZtLXl
hbHMA0ag6RBbZu0RAtcgeA1KQfdElOrVotCaUMPla/7vg27j0T2zi0Kxt2ADgXorAz+NUVcOj/uo
tlPrywC9Ai7PHEVGaveoIZan+xxgQ5CEkSPEqa7KVe8tl43QA+vLrwlsxBfro8hF6LTC4EXKeKv4
r+4m6lZXt2CrBp4jW7JS0Bs7+18jCMzRUS2Dxv/O8Axp+oxJA++MtEDdQXa0IIRQ15Z9AX7yHn+o
lC5G4jRDMEGlnGEJiQjfmky5T9bcciNmH6vAgaT7wIUvR3emln6lPEb+q157zftPF+5m/bN9MHau
KsIPOL8MTh/2t3KOS1IfYumpsabtl4Sthv0veVFW6z3R65xS7A2ZVbyfagxlBHJiSDK0+LCGODl1
JEQZNP6aj/8nO5Q/vdjHZzX1iE+nsqoQaqJPnuG3JOjU9Yy3ogaRut6T+bPeHqjsBzfm+Xv7pBBC
awPVvjKLiN2MfqqGsujM7jLBJP3Y59GyA93+PEfrxxJ/Bl1TWR/PuuOtcZtFUmOFVBrEF8cD9x6F
1s2+r+4Sulxv/wCjRvj84D9QlJDrraOly2Tsuhn9MUp2xMuQ8AnVtE15HTIT9i+VkOS09/Wwnn8j
m14BLZRB5n4rRl4EF5+W31RWlsVnXrBMChCfqpFRqVrW4QsJ1ziGsV6ASMlzQdsSuR97w1auiUmS
DgKjZ9k50eaqSDV08iaSRIRMYGCr1n9SSO9MDlxI/AKvo1fE9+V74eNIF/mbXRLiSqqtdyMXcA+q
CoIIbe4AsfBwm7jOGYSgRPyq1+CcW/Blgkp/GdZ7aK6Hz2dQXDnudX2FVrJHmmlpGaP7aW9aVbhF
6cpSUmC9UZo8DsOVue02HaiVZeF7FcKuZa6mmVSp4QdDzkIK7nCPTtTUcFWjIL3Md9EbBKRooyEC
2dwVkVH3M6Cxic4BB7B8uDmE9Yi5CUG42KQ89YaigmMPdwptScDTH3dS184Wgv8Fd8PI0H0QTmQW
Df4iZGmnYvmsiRavAnQEIk4byhMherSwl14hJWiiNdaVo68gMmMT+PdQDSpJlhSEfW44Ej85ISqW
A/5TzCEi/ydGejn8aQdnbEZXPW9Nlcnubv/7he97jnw6PsmhU5KuSpnjjMw3FRrRQCFspcJ2OT+0
2nBpWCiN3GDQ4LvKOm0sYVPY4b9o/QgoEmIoKyjqhFG5GlitB38Pw97jbtQ4L3vmKei1tb+33adg
hGGB5u/KIVhcQP2zW23jnjpYGLTMxfU9WqQM+f9nLgf7WaG5AWYA6lHYWpudsDaddf7Jcb5lQGqU
CFT7DN2X8sFvLa0q5bOsoINo/NDWc/muNruzSpLfqWts4QRbelygQhEf0l3UD5S2lsEucD+XlwrU
Lr8BOJ4zfgJ8vU4873vdybOA3sSmn2Cu4Qiu7ux7Q8LgtvK33YyUk9xUOpr2FBcZpc36Iuz2oDLo
GE2gS8Wy/5lz6PsSBDyrqlWYFLfioy7Rk/Y2XddNPb8XZwqSrsmCXfY555SSJRANpZyVUa2u1wtQ
PP2CGF55Ze5oFkLmRVlcufZwM7FYccAWFRj6BbXVgKJHbAAP/gduxR0zuLkfHeefD+VPiOTyBpM9
Li4tV1ch/sj8a5KKfIlX7b9OBA8IeV+SS39OHEZSagn5Zhm8VZGu+bviqlCOMuFAGnOo/h5DavaG
mSZGFuTDdsnA009NoqmY+60wi4AWei7IMUUr+Fr9JfSOSDBI42tztzFZOCOugoUnqqg78qYjCedv
w6rNaUYD/6D5O1sXXLGw2wEyZ3WQDXtGJCrY16NONOgR4UN/pV/ZY/OrYVIgLWf+v25AnlMDoLmd
kr1nzYze1Dm/djNy/wWBnOhaLArFapmevp6PEifstpGCa9JT6sC3TFm3QDqUJNrhbMaS+EYJDbNt
m2M+zPH29JGajkUE9GOwsJPMnXp59zvHSgsfJ9+xr/wpXdKyA1iTfIXnvQOTmOCkV1kvI8wKo7X8
UhrfRWI1tMbbRG/XDJWejiICkbPM/9Zpd7HFt/i6tI+P8Tk4DTznzrsISHobusCEVVI4R8DWNm6Y
57Knv83Cq6205KjHFtbZgdHgzFne9pRaVJa4hZU7HEmiMLjg2KUCZ1i68pLr0A/5uVIFpLEHEnlx
idV9rLhCQkH8xHWGsY4llkWL0+GUGT926TkEtiQIiVzRFIRkrK5jlOEy6/22JrhsM994aRzsq8gH
giGVNhIuv0AGKlqWNcLVYgc+nRs2Y+LFfcgTQxsCMwyX2md9tjMOLkp/Ux40vvfN3qAJcK7Z0/L7
PWngiujlcq7n4FN86T/GnMkTCiIxrBK537viZmW/2eSpnqACXPBjDXxrk/dqaz4FUJpyHQ7PCDFC
5GHocx9GiVlnovLOGAkbUIkoQXbzqZVSXfvHpp7NNeDXh1sWXUeWYnm48uV2EBuxZI39g5zvEe6A
sEGNUvXHJ/Xqs7djM3OEy/HsDkEenqz0DfmCF+WA+9vY7O5ySyezJs7fg0oD+W09d/TQ2ngSjnT3
TT5SDFnqlYgQhgnTj+PsIfYqmRDX7AD7QJzy2Q69ltuCk3XfHQo1NwDj3mMRpbEieeC4kxpmQWBF
sa33ao04FBRfPTcNS5qx/OvCKNNJzi3a/+UysnvNy/+ad3a5WMXqZPBMX+bbjy7UBJE2V3c5PJbs
aZl8ZhhoPkCRBpOg+hjIjVvJtXnw8H5i9AGrVhk7DF6faE9R58DyeWcLGW3gTklABOPY6IzGqlrC
t24iHbVmYUbIo5SzziKzUJg92NY1R6QClC87Avg9/DR2JAfP3+VQob4wB601S/g9HaugBxw4CAio
wHpr+QWn4BCD8EeIhZc20fqQ2wWjzAuh1ACSzCrKv3Vs3xUWQTOQ47dkSk+E0kJ3OEtJypDbDZiv
gbN3yffs++3rksYgKLtQ/ujz6x59txtfWumPSzd2dW4zyqgllIv6U7/GKG6PxfQfdJlRwy24QRQo
PvciRAA6MVef25ijm+1+nTbUpjuZ4KLejK8njuc1Z8P9eocLDPoHKYl9OrAVRJT32cWH07Svfewk
fiG5grWEd/asquMQsAcK6yENYlGzV96IJUBJVEc/2ETMJtv/t2lq95nm1HbmCPnsnZSxwB7fZQj7
pucUCbfxcSjvYlaoa5JLPgSTMJi+UDhuudPK+XcggGOuqnSXdiYpX+NGEXpFyXheWsQco6GDhpPm
dIOHjrZrjSepcPRKT5vYQ21nfqmGGRXdBHTF8r1JsElCoAhTj7114grk11qdq0ASi6HuLHLShiiy
mbe8LEqjSTGm5T7sOx8UmuHAMYfvO/ijl/3H2ycSvnT42xqfyQsHTqsc9EZO2l0a0wOU56wfpnY+
fiB++rguY63frpzdZcnMABNI0YJJPc59PMrdUDWYQggXnm/PHGLHcOk6FY3O0g6IcZWwXoko61B8
ksvH+ztIY0pGQObJ3d+fx4F7UqU+/o5HwG1rnGC5dYFxT7iby7+4fXSz1HtuGw48J3G5ChNKtabq
okY6/6fqQOnP4lGvc9aQMqGXdsHmMGBkzaNQQqd1uJKRfzmdMQc2Re1+f+SXoHEw7LoWfVmW754S
8yeKWjIIkpFcoxV/0o6DVCD7yUYW1ul6fTNp4QIV78j/yTrclcinTj5b+9Wl07YQbHzJc9JLCj8E
u3w0v1vk/xRP2GHhrbVOtbJNTYxVd/PNngPByB1vjHhdm2Kaqm6W3xqS+wLhS2MhAppEgatPp30h
6oHkt+ZO+H1ngemlpr+edQ+y8N5jycnSRQhmYL5xQkLPeoKuMawx3+OyLcXoDvRBK6jzro1Jk4O4
e9ICd8R0gxB0e7ZngpZlcILZ1rEqE4iZI0WnK/EHLkmDqW0gt9YKJyrtHKShJHPhu1XEhhAILfX+
q9lBNg+U3PfupVHcyFVJNGxOUGBQmIptawNxkXKgslNr7SCGUNu+ryOJLSE1QCLOoxD30j3gzgFY
eRzrcMiVp6k1jkHxjLBAsEbGQjKzHjcuj0HGX1LKhHGlNwOJCB/M+3LcZu5KBSBG54aHXuf6O0N7
S+e52bQ0C7Y2Y35fxY1SWsUN4RYqr5Z+bt6q3rISYyIGdezVlbV1QuersS7YOpsagBBQ8spxIG4E
KS3he+zCWZaT/e+sWwOcwC3xNdS8sgd0xH3Jdsq/x3Oxym3VJtZEEiryTUVFpDnsF8kjvAQZhHD4
GOIzFP5E0w1M3SDg1gf0XwbH4DgzDVL+MTqu+CtOYfNpX+zKssgeSTQxUnJYMfBdDSeyS/55iF23
z6m2NmKj3mSLkSHzb4u8B/cqZtp/enXWwu1WazO2jaycMPR1ypJ2yqb0Q4/Bxs0pLxXEmlIEQGbU
9phEVmfMKyN+/cfYamlfgxQSNhcxqbxyiGmpcvuyJXrg3jdfUzASep34gEPE8YVXUQ2yW29gjIHw
VWjk+k+jD1iWl0XZsgij+iSYJqVTCTyWdXhWqGP15MHxzAAnUHjbWnsXVhnlmDR1gz1GSg8lrNcp
mC6SG9xXf1z5Ejn1Axt/6fRdALl/bcCZbpijkDhnc123or6R6DDKu4qiA+4jH1A8ykN6ENK/Mbb6
6VDSxXsRV7KKpXiJUHHR1C1CBQFRMPGMW3FZMuRYVE8Wdl3IEyl+VhxPzGAnV62Y2j9V+K0alKH0
OYhBEHs+TjMVewMF2PGe5T0XoVbkufUWrpNDzoEcu2qJXzyz/XMK/mEyRNe5/SWZphP5nDQaaOSO
myWET7/dawxkwC7oIiKzTbBoQo3pMqFrHQ/DVY8HajXX97ew6gFu9STy5RPdJVTsQKX5wCiAgeFB
K+2482Lr9kAwn++MH4vziocJVIU/uTbNBX0FBbJEE0aHLjAJagqMtyHd3FtThDckl42D4TyqMEka
orVtm45EFAlIV5PyvpOXjsOs3EHHtgHvbCPCdVuFkgV3//PHvDYDOkLD5EnO1qxbynMLvGOysKMp
neNgApBie64UEJi/fXKI+AUwG4H9dZF2wrqIbv63ObkMAj+3nhZhSmWWpwDgswYqAjarj4iwVTWe
WE7VkzBvLyLnHeU3ruZs+kj5/OeP/hBjyvRxlfjuveR4I3yV1GDA79wsiw+nXK4eofYu5RXNNEmY
MbPkUh1AvPOkiHE7uajcUWMJEqn/AngrX90SghBG42A2Sb/e6AwdByxCvVTlBqcC1jnqR0mzIsmh
U680hJivH97RnqrAM4n8GT8jY8rvpFKM41xnjNAkdpfWSH+pTo5Uo8v7c7e6P/QISHNJKdT46fNr
GOZh8xroC1HEsS142A7DX0IGNjyJbd7T3mYDZzHB7i8LcHz1e+FNtNoXhTwET1ijdv/09NfqWyd0
tkTp8jesGcIw5cqUIva7d/Bfo2jhqJ/hnu7BVU64gyLq7cVgibe4ouIUw4mjhmDFblXnAuMXy3YB
y8+Zuh/54AHbDqQRQo6w3EQEXz+2cQhF9X8VvxUEQtOEkc9z6tjDEiwMpQG4PNJEk6+7h44/8oYO
pjHEtZiJyHEJ6iePZy1JYnQCIXaLMgMdO3K90oLYIztlwKvV12x8X7jWKHeCJbWOrAt87dqLecJO
Kc1tKeFdrAcdjRS6V+Z6yTdHJCZBY/GKQ5imuJttPVbsssbR6hH7dkHP8IWNvyLPtoNlg5eHCNhP
duQtf/zKYtoC53PZF2eI7+inHbiAvUfo8KGe5usQk3v6ThsAItCHvcfyGUgDbdxSFwRv5rW4zIff
Bcek0rU+FbfQFjcJwlWd2R+qAzqG5035LeIeiY1i7/0OLd3lJAr7CcSdzO1o8dNZdRTmJN0bBhgS
pkgTog1eSzYqrTzfXfl7pPaagWbj0oK3zcCCoEQhtS1a2xUfkrD6h9ADqSiBDaUPHsLdEniRdKZo
pc8arQ5lDQcqpepMWrJcv+oUQRT2e7y/eT8EyrDSH8YagH4kgrBk8R5zZpnCO2NNWyVavpc2I/7M
KyIEwSRGfSrPv5oYfKwueysf8TzmqbVd0j8BfLIEZAQbr0Lw1INv7EwJbKLp9PTFoaqPAyD9cBn4
jV0E2yhzabHrBze5nI2mv2YMFQoo8CwmtCMW2XqUxQ3ReV4m7MgW+11S2DPv5zb2VCeKheZvuDKC
DJygMmc42CYhvYqepoboATH64Fq6aEMIxfTuPqqfuDIThqFsIaYstWAz99y+b/V8o3e4byHuLJ9T
uQg71Zcgqm4Xyg22AXWQyuy1/fMUk0y8HY00ufU5PX63opmmwldOAA4cRYv3f4pZI1m0hWcFoerC
pfIencHOQE/6r7uTX6dUBEpYCJdm+Xv4iPrkmdlZfeGferrXP8BjFfztodeP72vAM59KdO9p9kB9
p7Ct42B4VHcxbwHgXp3mbt8RoYJeyuD1Tgsx2PWKxIOwud4JD4p46yDMw+guEHJGtkl+xONT5imo
tOoeM0T3KhuJq8UMeu0GrvKqHvfU1HlEkOxBL/bt8us8meRUt+on9mbcEll3ulz5udUj5JgdIKHW
Ve2L5k5UTwxN5g8obyURyeX7XXzGk6pHRNJ3ZghIjBT7tujqMGsV0GbdX810F/FmBhxEc3Cg4Zoj
1+HEHbXiqPBBD70sCdBVdDkP23qfchtlwwmuJKgKfkOZTP+QZ69XK1D7atj6CggFERPR+crxYFWL
CHtV68ZdrnQkld1Lvz2CEEKqCHJ0hcFUxoSrr0X022eQLqudLbmaWN14rTLFuLo326HShHEoGff3
R8FxAytYDqHEwHCDVimzo0U3sw/fDh/48IUoUsBgsvVD1P/odjkPqNVxwQzm+mlt7GqZsH2F7FUB
aWiwybdwIyr0VG+g3RpVE4KnUfv07QTbbW9932TfBwBjv6O7lfryiBAjbKrplivloRBT951kukEe
sWmlcwgLYgwSM920PxF3UyVm9lSr+m98MbxijlTofDP9gpYPm/j5SMsyuzoFzl9Ft3w3OkJEFsAY
nqoZCgun+JULXfCPJ4To0yvWaiQrpA18JjYyN5bMx5y5jO/+zcXKFDR9zSd0WTnJ6l4ACm2t8Y1y
ECs3Ss12BNAz+08iGgkfJA4N4NDLQxTF5W0ibgjjC+9Dw9UFT02ubzjGoJn6dd/VKXp7HZ948ruX
v8YGZaD0xRAyYFyR+rMaYd7q77FBs3cXUzzN9QJxNvn3zW45nPdQJb2Muu/Yc6x1SfpARMHBvs9E
RNpzI4mQ69/atwyN4bzw3W+AqrejHPwxqcXtprFgt478o0h+qh+aGF+Imqh8z+K/+DwqQ8D29dfG
AAu4aU7i9Lmpjju9PTLugc6qFbV4F0FzsOw1O+9XUmVE/+toxn7zXz9w2cMQN+ayWMz05rwUvN/i
2e+bactKuCp3yLETSmKjemoPjnxE5ahCI/0eZCi6kEjLpj64HMYEKDPLKTrpo8Ba5N5VLsXTy7Kf
K1FKcexUcHmwv0RaiNBfmC6NsUiC5Gl02rAi+004vyYY0mKToTp8d4HXzmGjGt7k5GtFDPBJFmE+
nbjIjNJLTxw9H61qFIJzxTVpYLxeoJ0WYmsZM7CK7dmG6HxJh7QA4eiqK76Ku92G3b/xjyIzbZpA
qD82RnI+HRk6uVVkYUUcy+JzS2n+aPz/AIw5R2DHwTerGzRriCmq2qRtw58todX1tzBajV1PkhYh
kEFjiW+AnbotjjGhr0KmiA74EpngfJYoi7juJv9ztelCc37k3heqA9F175rAgbw6kZf4N5eyf2oJ
lY51Vari1a+JmunNyPI0Gu7SQxM0ECBw/zGcwcXN9BZv9KyL25LoRW0JABwgTcSiY2lPf1YD39Xj
OZmjoLlGLJ4Ec37OXJR6to81UBC49cZEocrm9Cm6i4Jxsy4pQ9XeSen0Z09vHbIcuS6JIoFalWL+
Zq6UU4W+FNbp0WoqBfahQN1WXK5RfbBgV+nwv97tvwXYB+bwoy2/1pBVpbaYzkihBB61DJt4veOJ
8GFxnJWJ3shugcmGqjv130p/uZin5ypSs2qrtJyQq1WYtUlIU7EDdburmoKT2O9+reNZ1oyPl9xA
RkcYFwQpMtNUyFYTSZP92akBNnC6ZZwga86vCzlSpep9jsDSKSSiinbZ1pcah8JlwiPal6LPRpfj
CM7sotKof0HB9/K9EN22vRl1MX+pJRVAq3Edq9b7jzAcSOWcbJUck/7loGZi72ngok8aT0YfZ7d9
41YH/2AtZ7CdyYEC0MpIcTCEnAxtUdLqLEBCHLDmyFtOCg5TPmm53hYmUhYGYtbzgNyo5QBTAtzC
4qNB82E6sVxcuW5kQ9/KX3Dl9gUrNv1kiOWeUQwHY2mPil4hsT1e5By22iER0dTpMt5/2CID0Who
qB0OoIYzsxC5GrEQTkvLJRxUpEd0AMeAbEiHJO/Of46XrJKZU70nkOxbBHXAWUhoNnHbI/9pQupT
sMLxXYQxeDJ+wPDKFZblrPQ+8gYY+1raBs/tPUeLepEoFUt6hKz3IrVcJ5hpUaxzLT1N9o3aPfoG
JTcs98wy7rWAzygBUJj9mpGo+WCkHuIK9hf1VafX6xAqqiMOutPZwMl2tM+rwkx+OwLUBrLIlB+2
TnnxME69LmWJAT35ccl3d51dtiOeU/012RVON1tKPHxgndoV37lzm6HDHO0qhl9xhQm09RWZ65Dt
JZrfZ11XzJ625a+WjVdSH2WYhFK9Qn+bGPi5XpZulbHuh4oC+0Ys1KN2Ckb8/VZ7nKJ1II54bTir
t7pnf7JTgBI+WRzyu/2mzECDzTBOraggZf7LGfR++c2cZIvewBVGl7jtqTEktWQS/s6HDhmrbih0
TlboNOAZng21s7GSCX4idmTFENwZ977eG+8Fl5DwAtAzx64VVO1+WUBSCeT4iSJkYLDUrX5VlGC0
ovnolPbjz1WtK+qC15nRp7gCb9GgLJNMdPORKTpLt3JovSQeljoIBtVWT4ZW7CUp7nHw+1NXUjNh
Jtbg9Dp2Er53kTTLeq9U0Br3bGDEy17qYW1SFqFBz04CfKyPmcRV/sxzU8OsdG+b7DVCw+tN/AaA
DjOpeiGwJGWcUWjAbS/RWbXZnWMAFEP5h535p3jtLpRluIDArpiYPF/5iWugp9eBlH8Qj5Eibdip
jVnyUgyiqCDcHY2CebVwxYCPks46rpLhOxWL0+Mo1D5QW4eT4i6Yzth6J2l7xVxQtrAx5n5yhXEk
M5gjOR/2n/OqonCCw2aFQecvfAjgCkw2w2iNVpzaKFEvIuL08Zm54IDuCorzqUI4iW8CPg/fTnrv
QH+3foLDHxxM87wPP6iM6/sCw0MKMqiGjl7QCLziL4O8xEVX52CceQJ9rrFpmrznSC3UdNdHfAzU
bdzvjpi5HxQc1DGZA/996rocsfrpWpIyRgTnEzAX87y+rPiQBjpq+UT0Mm8YbdUjP2cp2HWeQ86e
gq/pDfPANCG7C8Ieus93n+W350MpTIMxDR/ZCxT+KcUs8GXdJMaqpgGt0hTyFxZ/Gv3VXbpWco8l
aKPUGtihtv8Fya3sBi69bNGNhJ2pWNFCEb/RsXA0Yylk1TBdLVdA9zqMiBKDvFBfF6++bW10gNY7
Z9gXLiW+YfK856r/hA7Hi3NQA8D1xLWEyAkM3Bn5zEuIHZv13OA3HbsYIaiOuLMaUZnbxHGWt1kH
6sI62d3gG90JkX+jYfrNMF1UZCkhguCxHbzyijdC3QiYUpYUAowXwskwGgoc09JrDDv9GCh15vt9
DHXUxIUbDUOfuflFzHJ8ysgueYPpaCkG8TZPyBhU8Vmucg2LhWitRkR4Rr95ejClFEXlXT7V2T9o
T4EXOpubm+WcoqZ75z+mPWVcO1w8V6WA54+NlFAjsrXZBtGueSb1z+DrR9XHnDaaPv8bEImmaML8
H8B6hBpkjW4pAWfL9d3/F6qSO9mT7OH6mwOYJkihxcabiPiRDdrhYCxK8k7VVAMvr6L4vn15b4LX
lEX1ZeO576fcCAM/EBKytXrm8UDhAvQ7ZRMT8JTHVAih+oYhu6JM13kH9tvS5Q2SfmYU992iHvwS
C8chMeRQzLPkPwtt7tGyWDiOXWeWEfskKUV1z3/olUpW4rr+Nf/rVPJzPpCUBztkQ3iBt+7WzpwZ
g5/bCNimK3fXHaQvKY+BJdUdkmJtKv0SQLFBWr6wtooStYqiwBII/LIPPDBdOUrmiP6NHWu1SWjQ
zdGekJzTSZltVI9gkhdh1cE8BegLPxlyLwYi1Y8FGVc3ygCpVO7ZacfZcft6QZ45S8uLYwZ5XtGH
cUKQ0rz+N34+f2q2JQFzBD6nZJdKJBWKitm7Zq5T+Z0RnJiNya+4FrWH79FEWDeYhQP6mGhPcUGL
APt8uzJLciygRBeb4YNlfVaPO5+eU8dIjzu4rMII+Od/wy62OIL4qdf5khF0iD2WgfEOAVS7b3+s
2uY1ezaSYjc/BFlBCfvw9yDCtQqMcoO5XE3b7bhAIpIDFQySLf2hphw0kHQq4YuAJMcjsEfOecDZ
+oc8xIP4ntXw03wTo85bKP0Wxdwk8ZlfS/4nGyNiOu8dJOLsGrv+C0XFX/xyp7h7cbMbTLAejhZx
UhI82CUiz0Fghoqq28CuHcsddtPDfEFxqWQHzup3/xRmuYqaF3Abzy3Urd0eD0JLpt6FL7JjtEVF
e2JGd4CovVidO+2eDbPuaDevZpwXraAflSbC0FyfoIz/n2AhYD0G9ErGfqmI8RLchuQJTCwP31wK
f1xrAbW2Sx1/RgRy5e4rDY/FST/s1zN9r7vZYXwv35KgoKMn8C/ld+tsXK39SPzETEcnte1xzgz/
fr8I7bV9rDcaI4SBGblkV4wKrCg5puM5tanl0NvNBEKoLI9fNAIXqQ+FBS5mkFaTIEb0huFiqONM
eCGu8UQnUBxENwnC2OeWQQWE4Wla8d74MFyPyNcL0yMM3RfMHWdyvCJ4P4i8Xoy7AtTMHDjQWuOg
RYmcFp8VSEDCYphXHUDwVvkXFVzUtTTbIMqXKnVq4sNXA1/+/SKeUbj3EKKFY/4VvceBwmwImXkF
CT4hEsfEziWyFKFlPlJlzykTdkfBcKg7nunBfFMTj/+nLOFbQZuTLuWC7/GPeZM9pt0V7kP9B+Qz
jAEe/0xCfEN8oU9DzWZ+bouNgVdCojaWktjMwjYNeaxgObEVi2PZ8mOK+ZB9HDT7JxClgMktFxVK
yX6yZG7jrc+N56gYJaKciCCe67GikukSKTxFQDLpy4O9m58F8Pw4b1U9XYxNuuPSPOeYodoO31+p
SbFrtUlEaRCgha+Q/VUywu/1iihInPS1bEvKdO6XzHV968Stin4G6sxMp4s2sXtWHTgakE/qxPRj
E9Vew+kEJymIYkovKXFntGdLz9HUFUFdRb3+dLAYclew8L3KCbqy9FPbiTpSqtKz13ozAAI5Jalm
HVcUFvhaDD/8MBRO0x93Fwr5DPEG//MmYSvImhh2rIWg8AWXzhYNd0vxKcEVV0GWxAXVZ2ykViNZ
Li04OO0cGbxr7QdbJEhUtBKlGEYp8PzcQFg30bJrPbMeG1+wma7biThY6z73VO2eNSO3DpWHvIEg
1/oKN+bgLqaT6c0qNuIuazuEYf5XwmyBRcX+tweWyvVMGiChsptjp0EKqjgNQTGyEHeI4hcVG/bu
5ji6B45AsUsaspSOtkR5Juv3VBmiFLJDxXIofj/E/t4h6OTYynimEZaqv1pOpTGIPWA0lNXqFqen
t+3pbamTaEQR1d4gYuKr5lTROONbwPTtTp3fbYyD/YOqBS9pzQ3R6wtu0zJDJnW7utFrBsDFSjTW
sRp7zTUGZkU2AFanzqDxiz3DEprOoHNT0kG2ztvhWn2Q4eZgvK6IIq5PKZWDFW0QzmOqikQRLI2M
8gqceMsO7dJef87pATyTPFANOhMMcXCTKSwyoeMMVClPCnJufUL9C4NLkCmSqDmfkdOfvTqltulR
DvvJ42ZHNuzJUaplgmJigs8Z/A4SyXJVJ3fuDPWFXnPrGm4aqWrPUHkInZh8sIO4O/eBanq+YHC4
7NI5Kxtd8gn29/8L0vwPC1pPiLFW0JNPddE8UE//H7CLpghZslvmz54W+xYgxuSJ27fS/wGA52fO
w6rHh103ZAt21rc9rVcbqhGjNwU24xkX0rkucG8CAmOSVTXYy7hnF+OuOG/U3YlcV5Cku9v6f47/
jvM+zfBZHc0Mbuol576SQvt2GseVXp/1Bu1pNtaJ7Ut7b+5ewbgHgkrgQXHDMqmZfAbpYS9GaAN5
Tpz+xQt4VPMysfwjI/H0ln9CnAbBK9JKQ4VDGdSs9tHhqumMbxzj5PEM9rgP+rfMXvshtL26hptR
4NDkbUeErclY3dyDpD2hb3ivbwuIA1evuF5vUVKjSdnlNzzTlG52Abz6fZeVuHdSC3BaEslOt//T
KEeDyotfNP9Qzvh+caJF0rfdauyHnlF8lOBF80J7SFbzV7lGtCLr2IQn/QPtmpCjlNXZADIonk/N
zIDbmv0bOQEYw7z+eEKeI2xhFEcqecdtXgvbrah5vvwvwtAcvQ+tfoJUdgmZL6+XvZYfJDJUOVwe
/XE3fWip5DfZBEJ1P4cstfoMxG1js9wsV9tQpXXMN2Dfs+6B2pIaXLVr09Xid8Qs3S2gC307RZrr
JfIuFxPGQHQFSneeStNgA2aTo5fN6fc9rPw7y/5cOtkq5hOjIaGNRO1f/yBin5ro1rI13pBEXE5m
65rXbf7cZWoDM9Iu2r2lmHxo5crc5ytpfIYMEeAFGzmemcQ4ozqXISS8J0ZAo6n9O1ZSECxQIJtn
aEXiVsWf54klAFH5O0RIznUPI6rqC1uImnVd9lH6tgPrcE2S+EPjlvHA1eBLOoh+eYIGpvTnGxb5
37KdLd6+PDjXfnNTPVEUPh0p9MxSRLzgZs0LZpWvN9Rjka6FjOfM467jdSDvJxIHR52I5gGOfaWw
bKu4xen8riRynCvaDRyBzZNEGh8lVhNszAwnwpEbIps9VS3ao1c8+ppGAnqJSuOlyq538fOD/Pgf
nudphF9Ph5jaQEeSqn19JSunoEoXAv3hnYL+fK1aEFdffxd6sPOqOu+gjJ6nc4Pxj6U23YamDpy5
+0x/+CdrPsx9PiJXHLt+7gvPVB9P3GQ3Vp/Qjv3P8WFab+tHCbEw6LWhPTWBlzcHM+wEstEnZdcm
JlvDBnYqmoM3cbvOMOu7TIDXeULMmAy/yN3NQwD7fBfRZZfSOzf9gg/v9wOpdOSFbyqHuI696Cno
VIVwTspfSOc2qde3LJWsUGkP+HwCLdt2+K6i5u7SUKM6CwejzPVh/zTaO6AhzPLmK+i0Yux8/ysT
06B/msACFq9KhC/8gDu7IygtcritOn+kHoc4Eg66VX0N+gyMeAU1p88baGw/B8/xw3U5rox7vywV
YvI9M5xc2b1E1JREKFpfo2m4NsXPiMFtlGRPpOVOWYBYWid2sQ+/D0XAnYjY1y6FliCaiVlAXMm2
hOF2T/lVIKvSVTosnvDifE9FgMvPLIPCg+JjXu6EWLgFTbKS7YdCkhEs1LzIRhE7t7F+r8pt9VUN
xIo2n+u/tkBLasrCO+twlyHCM4DIkh+M2jO0Lk5BMf9Wlf+qwTMi0jpZWs23imTYQiomZC6yAYka
PjX/s59avrvsy/wMffOq9miuOMTQBFUUceuL5PgB8Q2+AN79kbCIKGynHp8XDIA0VUwOkrUScbvY
NlklWVhXy6BuQ0XkXhL+D4frHAj7fhOatDGpzHIdco1j2qzSkrN25+zAnHvtTwJow/EXesKiLm1Z
rUJumeEmFUgOfKgfrrAAT6TX1Ws72OKx7H4Vo+fC2zFJVABS2dfHg7vba+YCjjaS+FO0+6n/zkKH
zLoPRzy4ZZUZr6o4C9innvI8WskvYG/W63NHCJ+0gVaGr2TiDLC7zht7u+qXITRnvKNpEdVancSK
/2dkselspnEFkr97AWE8guwrmH5TcVGoMmlerd1/sUvEBUdQ8hcaLiuq/I95rTQHyvXY8jQjKbAN
Z3WaGxzRXBHtPAzpfEvTDGhHr9Yg6aCX4J7YI1HduqByvHpTvOwbuzZ9Bzxv9AlTY5Oa8Bquuf/i
ondLOkSUelygrRZe8WOH+Mw1MRioZh2itG04nSvyuhrDwJUofzvjvh4qbmdlsWiz50cMrv6lCopa
U3Ejrvf6tZ4Kxo7wIjlZHzEG/x+7Ake2wimRT4iVSn1axfVE6fdriF4cn1vtLT+2iJILVuKtAm79
mM+7lXLeXoiimVxHlr9mGAamCNBR53hqhSQ1FHdywwxE+hIRfdii4EELCW2vhK2+YK1pEtbE4xaF
QWvq8BkGSl650WfILE9lU6wpQH+wOIijm89qoz2eE/qfjqrWroqQPCG5uPVpuMLuD58o82dPmY3c
mgacQUeabtlhX1G9Mt/z76O5xwEvjBQ7hpjxo25/Q+Qw3e0YUfMJY5oZle5+ga1EX6aWuZl9zhu4
+R1OkGpk0EE8+3JAzJ42g1dI0ohru+PnZUROqwzFWSOyKsqJojRYkK4sndapgflqQLTA2iYoWpl3
5o0TrZGKvpB2vt+r1DfP1qbIEgUC8PXPm0UAMUOJ9rCSlfgDVDI8UKuimKqO10fVJigWpiqBWkdy
IBJZfNGUEJ/DLAcYQRGtOVP93iA2BQNiIR6V+5c54YZSgCIWvdET2g57WrRdrixOPNB9hPGf38TE
4qeufVirXTZPMjxjyHl2I9sCTAzmb/4Yi9dr6XLTBMD+4ZgDRuckR5Ktz1lujDg6ex7SKMmqofuJ
R29ggi0hwLRcFwpNgZdC3GusKa/L82hM9ziCTCZLvj0+oneqIXAPCgbHDNVLqc/YGI1wZ9uDN2fc
Xn1wTa9lk62uB8uYTc0lPRYcp7qZRaJYED0UtXXRSP4sBkm8903/6QPdlV4rEq892hnF5LRkBb3z
UzUWqqtrhwC/5pqfMf+pNq2zxbfsfd8sc6Kzsj80w3BlY/6yJvPVlM38lA/MYim3rg6YCIQ1GIfr
K9Gi9+QnWTC4lBfZhuWhNPLouvprW+APT/UyLp6cZNhjBvkGjEv1FqoYBkPmKFu8CsMrKZfe3kQy
rMJozhc+ixCqvPq5ZxI0CdAH4W9Yf66e6itESgol/6kMwYgPMhJFft2oVUsxVLRvD3efXbSo7Tyl
ZjixauZSUNmHuqy0ikCUHdNNkmw0AfHSwYoM5C4TPTtYQXzDVpu2ri70vHyPkoj61wx6NPJvxP4G
ot/BFJMThXvoxEM4He6cYly+8LN/uUJNHgpYp4Zp3h92DRAbgRF3wqExNGh2Enhki+m/vj2WGCOo
LOjpKXJ99UKeMz9ZUOJD1YlvANdDkdBlzN2A7Bo1SEsUuWVOFxVeLTyIYMIdNdudaoG5nJgGAm+W
BOei3SPCatuNEyq24x7obymI4+gTwjH4T4UuQG9kRF62OAUG2oYSgtmD/PS3sowVFFi0A0v5pU4L
BfQbRcE8crf8R0A7c+bG4yQP0KYSPr074wmopRxInrXIfwKaA6lXn2Y8mkP2gh5PelY9f3GjGU+U
Z2syD2U/XLf5ieIxSyyNzcLtNZZwv7s5gpsVGHx9xJtlcTVXNIUL5uXXo65dQhfGsrp/fAWbgUru
IjAbVPhyepbGbl1VTEmVwxWTDlqFkGFvZdaneHQHYjv4PptPmknS3nwC1ZcPWtqdua3B0X1XdTxU
W/GmpQYOIiO3duBgzfHrylCWGzuU116/wjKmHHwL9BfZnuec2+Lsh9da3m2aijDc6oeRzSwgPu8V
U31ENxvaYWTLbtQSz/m8kyU8E+HzLJ/kgySIkkF3vA7jA0PNcnqYMPUV1DZxKlAZV2idDqdBgoXx
iUuYC8csCi5AE3B6HCY9BWmpQ+XwmEXr6wVNdRxIvVBTCxHyCyu0ktMIanlPtLY9frglNurh4zTU
0Mzqn10jDLMcnvVoA56BnD8y91picY0FpTRMu1R4ggVee0ZNjvxetDBfsCUneZ4wkmgY0FgUKND0
DjZaVXD8dyFpDqHAxAWZeMb3LjHwzjoUNfsi0u3T1xpxxUdl7l1FGfJEFVCq2M06cgYOsuQem32+
3eI1zo3GGLyNQ53nyBvEV4LB0cks9K8ZvtuADXwdvkNMET3gR/D20BP0k/qhq0k0hjd3d41rhNqI
yojy9+TJcaTIfY8K072dvhIQ0QYjxjdj6+884Cysu9EBm8Z/c0ypVkmyb146huOFKU8LVGQQVLSX
T/mcckWaFllfRQ0NrxR9xTUhAvbM4bMIF+KDmNWOzVj9+UKh3BvyrjoMTHcNTw43Ky5IXSgUB0tu
cyF8ZqvudsHAJHWBhqnne/8pT9rJcYJp7NfFqlUVy+RbZQYjo4VCaMdGpsolN9mx+zrf632abHni
PBbMRNkGhPPcgw4b9IK2C9QxQRsBDRGX4pYb6WapPOqxU65+50W5auJ5aLIg5mql+W3H1/BXf2S9
JIyJKC2Kwubj7YIwUHAXf50iHr0rbweRRU2jMOd1I7WB++AfZfglWijBNotfHmZmOevcK4oUocZb
Efk+GmdtRggAQm76c0hfHfzzdqAQI7BwhFjMfYYigxc52CbjxnM7Qeb4kBH4tBOmfkJ++055Nir4
sYO8myo6Xpg3Yu8QfxETFYhdt/4NbzaELdBNRlvdoNFXz6ITZIhTiES5yO5xH7scOpSUFAKY+MQD
0xzzlaB19ufpX6/rPy3Ry21BPOXRBpL5zNO168P1qPQBYBEOCjYdX5jp/yNx2UCvfQykj1Stoh79
/cFT6A76g+xGqzjwItqmaY+H34PWCO0Rr3ePqH6XIBflfBltRMYtxkYMfGvdO77LrJghcSOFxJNO
d/K8DcOFJ2y6X0kTZvgyJyv26vST3L/+IHKCvY8aNJPOYg5IDkRe70459S49ibiC4HfiNuTC55jh
1x23WfOCkGVD9BF+wycPcD/TVqTWeZKuixz7e3WldzmXyZNwREK700BfIIoypFUQ8c5hYTKt/heE
08kEUED7WbtU5xrStOwRMWpA45Y5qal18+Ewahf9Yyk6uvh6FVu3IFVNVVPxQVBMQQIn9CVDvmYj
+8U36vYL/gYU8OXE+lA9W/RpLLbdp/x/G2yGrIIxPhxU2ujqc7CkJUU9OhGALB1wQXSO4+FII1xW
3+t+asiRqJFBfc612zAqoDDQIr0yRvr1tHrmeripl9TSkVdZFIIsNeye5M5RB+yQB79di56eDnK0
4J8mBkNPRv2pNESo2h9gJ1CatkYZFSqp9B5kQyqeNDJUCEvk0ZpI884TQpy99pVyBpv5NWr9NYS8
91VNvNIMtAiFZmI4nEGZLqWTxKGrplDv36NsGZjFvDIjSqLkCFhJxbhRPIeyqra/I1S6Iszt2w3t
61aiQFLuu9TK9/Mp3KkcZfvKXnLHer5L1vBHEXQrbc/TyAC4rXJN1M6MxabGhJGsWs5u1q0MYAB5
XjeuSoiyDq1m02t+ouL5i0B36FMm/oRovRSPQvp+vQxHqNYeIvwKcO4jZaH9MxALvX5lib/f1sso
aX78gBgJeQysV1eZDR3XegnEg+HAezOTF42WjZu9/qc+WMuBxiuVy0WcME42u3pXuUU7j6zH93oV
1qv8dU2QjEqhFNLC8+b9Dh3Vq3QxnxhgRp7MWmHCsczAX3o06z6GBRJ8gXNOXXbO9X544B6uuT9Q
GCmXilJornBtz0k6A/6NaE1SA3wqUhK9Tx3vJFL0Pppj3jrxtUTP5jooCTlmwwr4LSFaB9bi38Zy
grFednVc+eBOdXn4cz+Kx/84n0n8jLlOOaudsAs+PuJKkeaRiHklPi7k4t1u6zefNEEz/pygN2hL
3xKOHnzFi/GUMuPZLwomafSGz7jssNkiou7tiMraYVjCTq+OKpTBBUpgSOdNikVAX8gC0GAe/lft
7+9HJz1pCk90fyx+wqv21QP05gfSiz52xCJP43kcFadr1Ji3nx9QMpgz92w3OdE3m0sM9+1TUFOK
Cw/1QIh2mbBG7BcW7GD/ofZLc4t/eRTYBSQPy/19dg5wtAXDIDRPsV5mC8o7iWoQ1m7skgxThoxc
bDZFanGJDZY1CxavRsrwspAHrbIZrcR3glx03ribgCnrRi0/wG1eItOzesvruyxF9egNYr7duemR
M5KfmInm3BrNgjwIp+ZWfIX2XsbDASrrnmKUZfF4N1Wu74RKE+wgRL3eO+/Xj72HUlC0Pqn5/eyX
hD2FrlK5122xYa6+xXxT3wwzgiYxnI/UE9oGo9IcPyt7z5f0SuW+z9JGaoXVzutACLPAeflpPpz5
hDHWHfkin6xiL0oLlYIKxX8zRyANxq4NlU3An9CXX1npJ98FvmRjDKGf7uY8KcZiotB7hXhlPZdn
HxlwjgTzxKmR+lofSaCBCERyM/RcLCMXgZdHWSp1fwSjribP7Wi/U19vkrylKHMsCPrCtzCfeOOc
xZ4huQMV3uRpjef2ZYRQ1DxYUZvCBSPJxew5ZMsBCqiiWhxVloaj+CefebmWrlPUSoDUkr97zEUB
bwXOPONSsHkxr7+EmIfwfgUxmGLNEjfuGJ9/6jmc/FuLbpNp2OUMLdEj4wdYuYKgC/IUxQ/A65IM
rIxZCEhstRvm7HdpxocBohnFasDVdob54I+CdeRI8RSoi6sAaMa6Zdhhwt8YVlu9L9lqCCuZWHDp
mPkcahxwqtJZTzSz9LN7r7Bwe3eJyttBGmg1iDvq8rtddENkxGIGpuMGQX7E9hHTZ6bkmAm86G3Q
fsVi9iFKCYLDR276K2HA8Uqxd1IiKpBuYUZRs3C2zLGEvhBRzN+IshMEod9ZU9JI2Ato6AyAQm9v
vDnuxgAPCe1rl2wIGxhPps4y4G3tlXaQZuiwm07hidDQtztEpxT5WVDiPiECvJAZO/YCKCiC1RVX
pR2dxqNUQ1WL2yNb2WYU7Azx+o3T5Q+winXENKqOXR15xAME0KVPjnOkxQjSAkQdQz0M1faHrBXN
eWM1TuIOHbPuPjz1qne6FUVgpmyLVMYXS/LXrVyO3ME60uvQA+BlS8YMrmyKRPw917xE6UTfoSZJ
tQeH4/YcDAOvFqK7JJvB4ZvxO6/iDFEJ2DJyEGRW77xyFbPqfYPMc2/xGCN4WshUOFVs2/k0BCBT
urfpXx0oDYTJqYo67W4JPfHq65EgmhrTrdpqEfdam44giYCMitLBAMpB908kYndWyExh//S3CAre
S1a3Ac9psvZufJgxsup5u/m2382azfQVE/i1/jy/q66UpQVsCOTAusVTOXG91hfbSy6bcM5vCd3X
My3/vyx0q8cFLce6HseP9rP0zDExr/DCFwDJkc5jxwmZGwUB1qifisampndaFIwj0jTBRYsTP8Ix
dUKQz8HQPxA+FXMbrITdic6QCuomeg8aZAAzg64KZtisg+iDJwfdj8Ar16b0fi90HMJ0nXp/0Spt
+ZDcwuyux0P1MZur2FErtWuHeenMgik/SqA6ppBGecfDvEcXzg3i1Z51hlJiU8YpjMxednOtyftF
AKkCltqVU/mdCjryVHHCbNLR9uJtz+943JBA04hZ1MSMH5R7/Wf17NKhQrjXPoPG1DtPeXpX9Hj4
SAGjU5YmQjSWIh2acY8iEdfzJmIEiETFhUZ30XUiezGSSMzrf/BqDhnTIMzj1oqGiioyGk7ahUvK
RCoUB0FI40Dbewnv5+Nvx0drMTqUFcooOp2OEH7cw+of1cwzJ0nsKvG77cYyO+dNmWeWa1ZBj4t8
RZPSIRe8B3yGJaaIITz1E/ezc/9AxMEPHfz+ppJa/u34KU5Lp4Lsh0JUrjW+OgLc9cAF48iaYhqJ
pGsHdmXrJEJc9XWOI+DsVE0R0J6cNLuYlKtEtbJbU0wqYYWz7DVAHUeU7NOpXe2e6MD1+ESZmaRe
QniOJOIIuBeebxt0dXDay1auJNdQfX+eDUcYK4zIPXyZQCcE1muj52+/ANTbq/zlAqmiSWXvkU2k
1IW2yQfxrWB0xxCYEuPCIqRM6EWAHcH58x5NcALMHUuyly34RBq8L1Ynd/QZSvomJewz9ge3PLGJ
SwoY0dXfALeEjcn8nitLBQ82dOkbjxw5D6TCGayQrMDzQ3ijcv0smOjS+eiIr/LxHHHYkujx2BJO
vQLHUXO2Qjm7NeF3PgU9YfTavbGhAVScn6PK03R5HpZ9pNhGoL1fIKEd+2oCoaZLFtS5O3J0tXLl
dgqPwxw4bTiwdGzrP5+Z5aI01dttF9WkRm+N18daVFBgvSAdkVAyoC8ZmP/qmBdZsms4YoRCzAOy
YzTm0kMnGsBOSNfGKufyaivgqJMMAvz8L/MV9VFGR0lGxroKWA5mMytgA7CDM70yjFZ9/Q92eBTH
a4nqJDXyURbJgH74enh1othGLrdMYj4FlqRSJVUcZ65X+h9vNyMqyg2rcP6ixgl41ZH0+186WYxr
DYnP7Dr+ds/fBl4PmKbS96s8dA/acGDowJNon7c/cRP1KIwHs/paLm4xoVjSnNHy0s0QQBmTlOhw
IUiZDGIXEfBzQyEgmkuiuJQmKNDTIRXqJessi8yLRLt9bNTeruhwug0ThfycfzAQxhLbSODikqWX
qNy77Dl9yaO8ZSJZxrdGnPeS4/RVhos4zpFErliI8LL+3wFNtDPybWOi6S6lIQf3VlY7B/kQTls2
SngzB+JpCD2l47ciLUsi3/9G23SWNkVIucU61zdmNQflPdQi6FfjMRcxyCBXamzyp8UsQRFrRPJV
eyFTri8nXyi+kbDwluUWXZG6OJ+KPDv8h6TKxL480OZNddZiPepAFujJAxAyF2QH/dUz2gFvJkyf
sjtdgWsMgMkBt9AHV0XpQkKJahESFIAzOXXPg/sW1cKYG6xObR/DdCLay9NgCuSJJoLZFxgW6lc/
xMz3lBhM8JTLLN9FCsAD6FQlvcnEaPgm0gXk1AUyhZpnLJbfzMTx2dHIlLlp7zraIXLB7L0Svb3D
TpZlSoG9+esNVf0fkt0lp2W6reCzd0jlIHZk9XMYLvM3S3Xy8JGxDEb+N8ZrgojiHTQTr6yMC+hk
4WTMQ/x8rkj6dYb/OSQ9/YCscJjZoZo+BxOgVy+ralivGkpU2Am6gsRFN+lIMjysWsoE7GTNyFl8
/jyZS/gVACfG9U7oERaSczLmvpWHLXNBhqXtpORlfxlQvdV3x4cT6o3YJHPvVAhLvMLbhZBMtPZR
1hBtorF423RdH2d9YGIancS6sfx9ckv6Np+VHK1ANIzZ/9br0GnuvsZ2abzS3VisRu27x9T8PC7R
UxOqyEB+rOx6CLktq1uCUBKeyf4fenX0hgbOgHZ0VzlLISdOV8VdvbqZJCuCjMONRBUiFedEQKbB
CzITFbIh8VPQM8RniRrTKvs33xsvqrnHWWDPIvfkvfcAF7qQC9xL+EPuFPyP8GU5q3HNxQMHL2PI
vZotkJDtVqfjVGO+8mo9kSO/G/JTlGn3DMrWsDCflLUFLt8ZqSwA+XdBeFvWQHYNnmH57Q9A6GWX
hOI5DZOwqNixgaCay1hZNz2wnDeb7LtVSITfz6z2z9wKcgc+q3EQyU+JjyqFp6qfcJDgxDybaN/+
f0BMCvM8oKBzjW/gmP88K1J166EZVzh3lDvhuzBm03vuLZcPYJ+VhicV4etKTfflyYHH0PaZVCvh
zPHR4wXiA/gMGCqHt/twigyjpbyvzhVc3Gjw9IOhx9sKRyDV3Ydhb8q/xAiZ9ORAxy6dWJdUI7CH
VXIqnPSZXZJpX4Tf4Oc4+VVlIj4ZNvESlgZu0bDFR+/mPXtL92PH3t/v9UVzTl+ldbaPJ5BWTQ7n
2oZEYQkXhqn1pxT4yw9wOogVRLWXGViAwz7as4IhbrivEJiraVVGsFq6seDwUW94DgEV5buhJkBk
RPZTdfxMjqpTOVannxaxMrAhZspFriOI4c1A47sOpZO2rFs4+1ed3aVl1GTtrOIiJfESyDdOpcTN
NzL016W7OT9LXqLNkfd0QEE0Fy2cfp6Da720iaKc/RXxQn1NEyv0ye3O1kZDU+oeLnen9JcEwNoM
me6ewzVlf+JD0LfiFOEjGOQPoBMMCZJvkJ8NYl0Arj96bAx81J0GdUFBAvvr7ZXhL8RSbNpnv/my
sGAv6qWNrszw/nMIupnagR/kHbix7Wj3a7TjN/SqB9hr7NJUaiFc0I4gjeCl32dJMjVntbLUm5XT
ZtT8F4+ZdHOZPdPgAl40keTRMSW2ngdYwfEs5GlbDaYvBKeDU3KwnGH9ujT3iJ0moEekLCQMk+E2
u+g3hOOlaCft2FpmsWqTer+wQg31QODqRenvepl68x2ejwABce+3KTvBCF4uKJk4mZX+i6umMXaB
IVgXelKp4iyC+xFEImj5RpGzWZ7JdKl975PAH/JgzSEy7Okl7FhAhdsB19FGYmG7Z74Zr0llbJPy
VHyCJG0IL4UoBY4hrHpRYq241tJy7iy6+gn/Zm2tOlSJacTDmFTQJ2+furnM9NCX9K9BifEbMuVO
bacfa3F8e+5Bpulu1O/B4KjZH4J9qKJOEnpE1IGVdo9Da5CHOf152zmuzXMR45HdAQppsofPJwnb
f/pMxxRCQ5A0lNclbMzjqAcanuW1JlMxTRxllk5oOmW9q4llEg4eJCW69SkvXMIYQUjJMb/TnpOi
uceJ8Du70g93L4qggzoDcjGN3h70AQKQaXVOU7VAhhvqkvtpR8vJ2mqzP7cbUlSyUl2TNcd4fR+x
67anYe1lYEdwA3Dw+43vpBHQkznUwwvpNov2d6fUWEgQYN281E1x89R3zMWbJ3EPkMNYqyeG75HZ
mBZfsdYHaFxs0FTc/HwoFFRpWqHsqqjEcimyMhWlnQrkAOzFlK9eEi4MjlfMa/mM3LjBY63tfzHm
wATf451SQnqNkrlrQbdS/1HuNBGHkBFL1nh0U7jH2SjNBKXYh9JHzeyibhtzmAbCsfslRWsS3UmN
rNJ8YHPxGykMxkY9lYyA7/7FidZquychLFU6aLHIzDUH4zXJWJpVVIUn4qQZcT8ob9ELHwMM69U2
bs8VkouE/GgdW//s9bztuEs5uDUv/clA5ZCI/y59lYtzK0fIChnOyTZw/4U4VynaQgj7PtMtxe9O
5e0X+OoNlCSdZHjdOcZ31Z7j32umigt69LaCeSOkdvyZzbrWsNpNrXz4veAvpR0UuzeGbgWkihyj
xE7LvhD+x0PzR8IdnlYsaquzcYFA0xxQPM8QPp0Tkk1G/fwxcCwSXkUBvWjCxRMQVS/KP0dErNyL
yvLNliJ+39qiHGzG+V6xRnCQgMvUGel9b0UcmVQ3fsYXwH1Yk6qVWS90FUuDS+7+LajkMONafwFg
20DaXkKKLorIW2SVB9icrIS5iz28fSgHc2eoeA4cmWMN+Dz8SDTKq7CTOIWHz+4OSkTWIy2CFZOs
JGBq50cJCs1ltNYwpluC0+qnpHfNN4e5OGN9P0LmQiIoT6lfQPi08RDDTmh4rKlj0vS6BnrGR0Ud
TIF8ueNivEaZ8PHonQ7u4nzpVumUDuRoARtJcwOA2GXWmTQCo7MVA8B5KRzmccpXud6pMjaMIo7K
NadIkbuEQQCHw6hock2xA7Eo/ogPSu7Z3Hj0PRBk/URx2aeHiw6UGChHnjZo306q9PmGaEquEo2h
ZFGANyrXGXSkdGHw9p1RzxXsXSsHrUXrZZ1N6U5MfC1JsD3VIkjmOF/kh1S+ITIYCKHrcg2F22gA
XJ76BhT7OpDymvnLQ2JE6j8zPe/80hMaLLt0/E9YNl1i8YXIoimwE9w5iLuE3jZ6o0Of44jdIt4L
x87dcXj9nv/8r4dboUjzTXOoLYTTupYMEjmXanhA7Bf/aXJZHlEDfjRr4Y3UxFBm2MKzoTFovd85
/v9fKwXJtRi5FvyqB/Zox2Bk31BRXB9JHWelB+nDgC5IWvUTXeBPoWRqGuIcq3kKsJNOQcRI0Q26
HiCYsaNDNnipv5V8COF/EsGGfBXNDIKA5Nqqttr0d5se54NeCV28NFxjmbxboreJ31QnFb3TilDk
DsEAkZ68rPC1zi0jIZnGULRhj9yOIf9SMgI0C+xLLalfDA4820MI4S+VrTyTsw6hNxArFtI2jBmu
Kud0RSOUmyFBUGG3msTU19ClwjE2hhP5EjeY6WVIb+wdklfeQh82C+L3cqPmuJd++D7aZ5oQC6xl
G0TTTBWlyMrLRmhD7+2DpPaSuVEEtniYxMYzVh8VaNSepQTDNXBaYkR8LAACL8seFaRy4PguqagG
DL6GvwYaIKz3+RXo0yxZKOcvBoZwt5WguzoI+ofDn6FT9Gv7LY1mDnZoI7nqqOMMK3RYLhSBuSNZ
K3CiaeXt4YsB08875L7rIa4P5oYD1VMiXqIYijGgzzaLB9l0tQXM9N29/l5/W5bEfeqU8EntuYwM
YLtR3VXz9w2KOiLJVg+H2rmqMb/u/c/qleKvsMHuLrn1VSufh6jmDQ0gY+VCNW/bT98s0vcESURU
wyYy2Yv3ridVIa/Kk7DR3EFwqBHxvHcQgIilGjxb3A/km61jTIZ4zHmQCsvmQwzu2y9MfilBSsN9
SwKihN6ip0D52xzGnjqCbEgF7FSJ7x7yAyXh6Gh7fsvXL2KnLcSh4TlOEJuKkkdyH6qaDGFawIR2
+6JQqyE1MtIVPbhPYoKnuAAc+MZsiS/6DTL9OqDkn745RbhcYKpc2qAbzXyxyUbhObAETlHz0TsY
D40MpYl6asSPAPJ9CYFOoNYUvxBPzG8sQp5ww9nbe9EFq6Muuj9bi+i+WqUK/TijBAXB/Pq37J1Y
AfcFATt4oELbi/AyKcbg+LTYLhkJzZ4fEVAFd8Oq8XUBZCtxJBdmDkcpDTlbeVO7MQGDdvl5ixuE
McyUjR4rWsXMgavRe+r3b1X9rbMUD/dzwqPZN1prWmNLL4LDeOEdumezeC+LzyTBRT8CUsR7Lx3e
ImPECO0YkPHs8N3tGWTO5tDoMn3QFNzHYa2yjs4HePn8LPl/VPWr5Qtf3WeNwCTTv8yEoQcZ8g/o
eyf3BSshpWUo6rvMuweRp2Hm98stvkc9JyiKP0UMhAvdOwly4KSBzccmB+snoF0P4XjSJtwMRrVA
JupyWXqbRmqyQsh8bx+0DMQJCQwaRiANzCkXE0PBGRzGZYMWq2VTsHnQQPcin13W3nL+a6rV9q9s
OWbuROrZBqTJedRIaXwwjU9c68aDS5xGjdbH75qozSAQhS3RA/GI7RDv+oUj0YtUpC9a4/YukE2Z
ii4ZBzK102kACdjd2gejc/DWgXLmvSaMH0Flx0AmF6CvxfhK0PbW6FoWm8/4zkfOmtleb+OExV7J
sO7DvdlAN3UeLBo13C4Jr+EaSx7jpw38yluSIevXu137FXEUtgco7mPgB1OWDSzgnqg2PLnUaESv
ES/FOVPBsvUN9Y9QaXMQjhZsZ+UuE7Ean6oAaqT7yEIbVvl6Oq5dPuUHEsqeaprwQxeFMOmnZPTt
WVVStolvTEPu/u4JOOaW05rJAsaS+iSxwp1pQTR+6w8pUmXSu0cSOzOVm/XAnAkMOsRioI9GJmWf
H3+nJHmCfUsX3ESfeZyOiExYgcFx8SRxIFfl5Jg910PtLioPEoVvtJhPtOHoksbfOQc7s8o0XFMm
XhQchZcOdwbMvzEvZBULHYlhxCzlzNIWXb4oURA3XtiusDLgvjrKv7zLl7tuoFrucFgZsViVr9Rh
up3SnuqIEHTQh9vbTcjT0nvZkasL4x+DReaGBBRrqE8e0gVJ+e5Sm2sTlDIAGcSayqXgpLW0W043
yyG9+ruDSjQ0lpD6XyekQJSunKVGTC5UZidNdLHFmrsiEsPlvXzyyAzfF8k6KK19V5L+eG8EKIdW
7pQhjaBtK3uzMrHXE8b/2Kuw0wknQOtR71bDTkAamA9QvA6uWB3uibFnmWRGe2UKNsfGi1JEN42r
pVcdh49rigV5XZl5WqNnKB+NHcdaFY/HFLuxkzobulRS8SYoGV18zXTyNBRvd+Qo+WANaUtvq+iC
iTqD4EeXKnGvNgnD1diFCbqmnA3OtJbt59GpgklTeyimXgyrjUhMliQv9f2EllH/q25e3uR1nvoE
ljyCpeNyWLNZoNCDOtqNs8c8y0hM3k0TEJxkbGGuoKdPjblxrKyBPqQ2nRBS6ZzWjc596RtlIhPl
6V6oYWOnf9tLXJOWthzI6K9YnZhRv6eAHINdNsGCf9TyG4Bv533wLhZr2DcWLyRVV40MDec0EzCs
CDcpIgyKRP8iIqJ9moJzPbsMnI5/jSvAbLMw0t2+p0H8hqxV30q+Zv/lKvyyQa1qF8gq/A82fXMK
E6yMk/axiWDjKyeuhBCBmlSb8usg+vVwA5R6SwqeLcDnqFiXlqzmah4XLQeRnZi7+mIsiXOaYDVv
vrWwTh5iqNchIbp+Mrb7xSmUU+qUYqJjdp+xYMJMp2cR00ZoWBmj2b2SUUryRx4DfNq2IDk2uUfV
6nQAG1DD3KUIhj1g8zSK8q+FssdboQIhaW/37oC6I3lbQDGTrfM8OFIXjBbhaNQGtACBpGK3ldWd
RQHsIe9y/iljAPzobOWIDp6IDJISGO6poOfsXMnU5VntVPVdcrPe/THQWYs6hR1FerM9ZVz7R4px
medc3BNJ4uCzM2bfU5gmXMswFH2pgUC2pLQWSNvJI91n+XUqDJlI27EBz1rBRyZpL3M/RhWEalJM
Nz39TOWN1g0Uqxxft3EILnxdbP/BD0IP7aPwMY1uI7Jo5bgvj+NYVjNRN0v5KztyJ88iezr54rNS
dHjXUvwWURFg8gilmGMXBjwUKPyZq8DFdXrdJbBkDJ8q72L6vV5Wgilv28reNAbSIWJedm5Et+U9
VJsk9e/pEIgn5FP9ixC1lEa1yHa+uiLq/XJ8dU+aiynAKL7N/02wZ5SAXoa28WJlm5nuRxxcVLXC
S3GRx+8boYVhBNJD1ovoZYOyCuSrXjNpjtxg2ue4JTKjbubeKKCSZodhAnoipFET5cvYqzf27TkA
PZqwEZA5+zPuMsQ5RHVC4jskZNfeLD2sSZj1OTL0dOv/5cIaFOUSnVfULVb+BGnvcdrXvBIEULrl
xhTRuaKyFAUzhgOXPVLnFDCuZZWTvKPH7Wg69GRI6RgsuxuMsPpedZZDbkAzu3ATsv0IhlrlORiC
EQFoGB88mEniwRERvZ95xK0xsLj0qeds5jkPSqReWFTOna5uU/JHJPx43zsKKsu7btMZXPdNkot/
gvfvuWXSOnip1bar4JZmOls5JREHDg8Vsud17oG7QZgvdEkDwe6c49uYjQcSW20tvT0VKNE8EQtI
acJBHPHVOzMG+/Qb8IM+k6o8RSJ4Ml1kJSoN+LO1QQmmDjs0e8PTuDhtzJV2XlueR4DSpGp6xDuG
FXLxk6kIRWQjZRAf6wJQuziKRJLKsglGssvo8I0KgTOv8pC6GhyJfX9mQUt6kcwsehneT7L7FiFd
g9Un3k9oAxS2p2BeWsDEl+0w1BMQCnd3oiwGMQev4CrjTly1sCqwwx0tredH+H2Bqgzd6z29PBu/
hE+PBLnQBm3DvV/e0m5U7o7kSacTcSyPVce7311H4X4DANGMzrwMJF7MDaYzd3eagd8FBc2F8jCg
98nu/GEy7dquksd2z47DqxRDHWx8YwmXM2gBLMjfCTNOUFbgFzmIT1fgip/r568ytdPZ2MxDHwM3
2xrWO+cQtAL8VgwNiiN0ooFIxj4EQQs9dDNFnzoFjEo19E7s/uH2SPMfHKHXxij4AwTLPgouV6uR
kc8Teg785uJPRmaU5etmbpYn07KNIIUqSAW8LYEeYwRMmuaF7bBi8LfPZ2bmWnP0p452Y44RDZGn
Cj3K44JzfmeeAwMsqKN/6OtluE39SbdlTIohjUwC/JAzY2FbAiNVv3kCxGfE1bUFBc5BdDpXyj7i
9lF8eJtH2X5Gv52lxleIZ5HhKIGLLRMN59Qqx0r+xoIc3HvzvALaq2TateIaKTP4euI+zNXO3Gt3
JwI2GoNSjHIe95hJFh3OqEL2+Ldr9fQpZTGDH6TaTIfTRRvlQKH91N3vbL1jNvb2vKsCi7oRyxR0
ElvAdYrhpker/Z1La8UqKe6D95orZ6XbkTlalX7IBLBng7RdNLTWkORJ8qqA0sbhERE6XxwvXTZ1
NClP8yFFLlRNZqtSeeOS/2VvzMIClfjtkw0+Qt6o/GtRHhAVNPwQA0ZpOJwuk8OF20wFM6PRMBpp
sFzSYNLpKjE1uYgq42t/9Vhrwkv2RG0TcwQOgVGZAqa6JbHyPoqWsBJ8QcyqI1u6OoB+sQEY0jK2
JNS/sPNx1AwxFyxX8gcJsU4yDjsnb66AqtpOeejpg3itvvn0bZB9QnXVKGUgZ5Fs26JFnpT/I5pe
QwKsXZxTuTwmsD0XAjEcyHFW6I0LFBCDc4STsNSGTdrPh7ix5pWgXggUVdnDdOaCMM47gQKRrvjb
8Tb1//Z7a8whktAuScho7xG+BsL55LQSrY5wUPoftGl/DdXJHrfQ/2w4W+t6XpgpM1QvYVhmabCG
ObMmiyxwhPncor3/rd8GmZFacemDRyDS90jqxT4FGtHEl5cB20x1xdrz4v/ZFdYM8+vB1gxRpjW6
qfidUa7mRXVSN7sTexPjz3Y6f0VGnFTnQEMKnMZv9euRKdmb6AI+gDFl/QY6Ob/pjzy3ZtoCNHK2
9pa1WUdm5VoOBYhRED0leFvuDhcl62WFNTkmKrV9f9ihv+TvsQ/zQeETV/jrxkSPDDqENlFHxCVL
sOkEgSpcwSQoZFXfqrOePtCbvIJMMg2IfPeEL2ksUDjiWijZxFrG1/TVV9xpGq8s9pLZ/p6VMzii
2evzZyJ9N5ROlbbz8W0xfIeBpUKVuEMZ58TgKxxXjgyjZMIicfPFudV6fIr57G7+8bccxKz5hRc/
EUuAvxt3rX1gj+GHaz+GssyekAYFE/s3ihZ6s1RfN0stDCvAKFUz+p6VtZTAEwTTfaGn9/EmniTo
HYmxAemw2KlvFuaRj2sHzkDW61f6RCt/KwRsaDLV352olJvlSpbl+a9Z5nSUilyxPc3J00qodNJU
CiEg4NnaUbV/IYUHP5+vCFMFjo+lFmmP0X3yfVzuXb0j9AQ1dk0WKYr8wPRqhcKyXLq8XEDQRnmg
R4ewFONOdE9Dux+vmVAFlzUZ1jMiUAUSa7/MCep5bjXGm2CgsxQ4OL6K+2JPEkBsu8W+/sg9AfTg
jcJhfkAIXSt9JPXaQkIcPS0i/4eAl86zn/2oerwWYmy4Xink+UqrKGFwXxW/QYPOS1zcV0tmMdvp
auDgqor4NkZamwf6Fo3M+y17qEeoUOTdynQDciJDrwm4AkFDpXrqUxYpbLY6Skd8ZL+jfctLt6yi
OCjQZZXyi+XidideYoqzvzZLrIZXqn6p5BwuLE3vCNOmfsleAcQoUHj9S9FVsVf9wp2cKHlf2Qh1
IyxFjgcmt1bsJ8ScJAF+l28BHeQOmgd/DHf+U1RP8grCGAyr45T/qIEJFampAYKz9tYhGNYWqXUY
+uDpSSMHeEpEeTR513DU4gejKKyvkwftljfgHerjC7FGylJ03ggQfHBuTVqpSV9QOqEoxDqEBjJD
eZgGqtQhFLtMnyaMf45GRBi+9A9mG1Pg8PsADqJAB/h40R6wDizwefRGL/EBZe9NGffFAKzqnv+3
H6h46cDko4ZxObbDrsotA2KzoJhcjCW3ff0Yn2k+HimJJ4LyklpXUIqV+g/2BMlQuEuczYtKWs0M
HD1WeS9autvmizyAyrPo+JMhl6Wa9XGew7nZ3I1CsLpxXBj89KtKPECytbg/SQZyEOZQTEYSl1cq
gGMni58cXIBSmsQJACEZEhohngKB0XGzNX+dxaHEYiJmHP98LgKPJe3sluuayWp38z0OQEoLDObV
49N7IGI1/vGU2h79YcIdlcB5QmFejwYVydmdjqp8ZsXFG6vEGnlwgVKOj32jJFiVarB2R/HZGBH4
pamaiPS31fo9Lp5Ii8wGNrXjEXwNIHuMZZ5z5cofDQPUXsPFuQPppsI7AG652SdMlnvqVqVILoqh
hxcfzH02+tp99VxGbcVgkTEG+x1N0LnvvEmpHdS7G8Kt4aY/80WM815ow0XzlF87L3HmGd7u90jh
c0VRtp2585bI694OSKQyG/XiH/XvWOn05MHMap4AtqS146y3vne3gxDyFkefPTIZT5gcrhAqd0mo
cD3VXT1KPO2H5EzeM/FFz+Y+CfB349CJknsTuc3Mktrkl/v53rC5v0NmLnktYlIvkAS8lIx6YN1m
n1ci1z2wf+LB0BE65vjQ8BTrXy+1Ml7BSi+jbQR7D1OozWTHg2dDpyAJ8BAjBhOkhYb3PimvPnTz
ViwfYDkJmpQUR/PqQzSzA2uwXWVnVSY+EUfbWiWFWVj3JUwjW6m3GRb3rJ9boW6D9nKtTO0ofGXP
0PZo+rNnm2JAyJKs2KHMPYNzFSPph8ej1+tLirkIsfCbGhEBjLlS8g+zUMHQr5H+kfNV0FtXLptJ
Fr4xsllXtwhyvZ/njuQFrgsTpP0m7nETdbTvF6fXMAT+JhudJxGNg+ypBb7K9+b6XxImV6htYmAv
tejlcbmIgn2OKtRo2QWyg/ZqzHPqtVijfUj1bB6e6oA7vsjm6l2dN47ZgJAbK5jTp1qY9g4NgCO5
72B0SGLdP2fNFuy7GsggoiNpbALDUVCGh+vzQi/DWV/2OGbaYbWP3mdEK9xoNuqE78byxdvsmXyx
t9hQt1Ok5tM7oFyWN4Iy/bRMch6EIiisNe3P/k/95ix/9jnPAuIgvn828gbi2MBKfdAXckB4+Psq
omiW9CUdFTl+PtTWAqJ08SWZZUtbXtZQDvyNOtcFKDSYm98vkmqaCe+sKIqLOF6tlZTpX5LbUhPJ
OtQGCnp8MehyT6jVriFiFwlAZUwUg8WaEtcLHpz81OjMSTQiWfXM0Z/TX6kG11G0Z23cg1+EN9FK
MBqQNOCWtC2fo8m6rgPQGbHV9zBpjX0eQJ2sDma0MG6lzFr28KMicV5PaQDU5EM++73aQlJWIOpX
MkInuJq199kR9ReXbmfXHL0G1VBf7mqj8CJ2yapV41dj1oFxTWjWvs7/8cDzfbzI6GOmk8JZq7vF
sUOdMEdC0grTnPAio1c5x15M4GboNMAR3qXUJ1unWQ75bdLHwFHLWX3mOrgMl4aBnmcB2mdquMt3
2QMclrYbPkMbHTJENzD4qNJAoHTaYp19Oi7J5uo1ca3bYGnET9Zd9zGq260iJYzbREe4tPowEkCl
WDUU9wtXDGH98lqPOFgzHp/7UoMkKh1ZhooN8j6gqXdNGGj3w6/+NylA6CPst1zrpv9tyToQOk3y
1K3Nyvij/ujOI6kRXy+74uJHTk9IbhZp0rn4ZBzqnyNz5h2Gn1oAU50QnyOcuhdNzQLxErCyIyq4
zpuzeKrsO/vxckgMliImTA6NuzPR0grUeqKUCq4cHYZXOvUj50ctJ0RW7etDpVYABco0iX6Z1w6M
aVkZ4pqm0kbfUKKjZWLCqxTBNa9/M4mbTv8Bs8JS8FqLQlIB4OR0ArM1f2IdP+2+UjkePScSPgmY
aYwUis+YtGt+8o9ypyRehMYCgaOwK+t26jutXgqtRqc7PDa+c37ephg2DOW7zXfZ1oNR6VjmnquN
GI/6umfpMuL/OpT+5Pz/nU/k36f334Y4ROrL3F04sj+xhCcGqIsuAccaPW2NBz26QVh5UK1O5hE5
amNDj0+rNTUE3n8C1kFuna+nsAxGiYa8euK8K5aKPUIseeh8t1rosQbkDbkDhUdiTmbRAtE6Jg6M
Iu8olExqG6d+ichaCfyCbDlIU4efPVuszcD8N2tVrPt42PEwZtYfr4nsoDov6cvwO+5smUg7yLiZ
FiXk0ul3Eydl69uoWtgmmyx7G1k81tD0a9P99RI4JcH6yMInUcZ+3b3K5DCfDru7dAjPGS+HhSv9
Xldj4zvMJ9s9p1hFv6Az8a2xN79uTFGJeaeXIne4n1pxyKwv9g7ygkLXOgJEuX0tLdYDwPMRZV5M
M835npjm2/mE6psMETbDUmDOLZ+AKvK9dcDeuZd18RgUulzhGNAfyISK9H+HV056MsDrN4wmRrSN
12x5Ute7PGawJbvaqhddcW+qUAuChJ/vu8HbDIS2jY7VZB78XH7aO9Ly9Bh+e3E4nxRXJbIv1psn
zaLS+g+3zmSXMQFhF19RpciAvFJS1FBINpT95eqUOFHwNtftf8TB7UKq/g/0WcBa5xJIRfD8Sw5F
jSHTY+fYTYcEMvywlR9GfQioQSIbWWlx5ZHYZoJ7l4gvgdGBkfYXTxEf2zVVinHY3ZZqtBmoYAuy
WOBWvb2RJcB9eMNDy8ULi54AsI1/AS1HDzRjt2qjI2+nswoefrpA2UfeKcCPoyrbIXLIHAzB1L4L
k0j2rQUTlJC/nz3SxDOnPUYOVY8kBrPpQhEcvOH5dxhaiyAhZZymOuHGvvEuO5RjLZpT8fr1kE3B
IU7BF9DA+kn+AyaVBMFa8OX2xVQk/oVvK+rqDeprRDU8cIckf/QxNgWRxuhGAycGSIkijB7kutIr
U4s7yHK2DmpQ+lvMmfd2eqxidyPCJ4nUZXJ+/ZMkKpLqx0RCwMw7/zP71c63P+a3lRYxAZ8ysDpQ
N1m/Zz1BD3/j/8zGMPFSzC6cJwQLGqS+OQP72K0H64ISuChtY70UA+uxmY9A71a71YFpe50VIXEs
Ye4cSG4fNCf0BEMwy4ZLsB1djBokdu7hd9GnNmku+1fzjBvMyA0fX62Q2mdlSY8DS79uPh+vTh11
hHm8p1dMgavPF1x3/KbXzHFXP5SBBuY5Vxr1VFVgkV5r6rPGLLGUH0xgReHY35JIyoh9fdHk0PBP
VIGvqhKlf2LzNpBcO2SmzuYhCCDRQ2AXvQIChsb8NkplTY5JYffTNUEHuMc1sXNpX/tiyrWGBhRk
fhnv5kCAGEL3r6dPFwN66oE9fRZDeGB1p0kyiXdWUIcski+PLjWzkbfC9SCewNmLdYjfA9v0SR2i
cXp4vRnIgUGVTxXKs3LsCS8J0SNQc+XaRV7k+lwRVbpZ0lKrf8n1UxJabyDFW0WrWwyQDTtR6U/U
f/NoFZtUO/4Uw8UudsbCq4YRk8m67OJUEaggbtvsmBmodgkx+HMukSug6r626tEfGNYuJnp0LOoy
nnXWBrws9ATSGjc4Azt1fKsDOoq1GTYnkva98VY9YqIFUUtcOela90ACyCAUvnfHsGUC6AoU/npT
lxi1qLbUDR3g9Sh7sIeOeuY8HmfbGnYFIz+PrzyJJHjZUzArkKvJLVNMFZmTV369VGxofgoWfRJ6
waQdasSpVwa+za9uGAZZMcpMYsbYpf9OPJbY5a/uT0LNvEgJFU1j9be0F8ggVLp9vvKOCLssRhIr
uWnkFWBMhwq+vHJHEUL9RKoytcVcdiy78m8HifXkaqqNx8UOgNiVsUwpWuksLhQblwojuBUqZrj4
csbDl9FDEJdEkfdgpnCbXrzcUNXz0il+FpfSLlrDYqO9YIiUavkUamhm76Ma2tyOeeo9EXRfZeUd
q0G+iA7khEImoZUtYY/hY2Z8DDl7nsGlZEaJmz3teWxuxL25Ef8WWtrRBpS3z46mynS4aKXHVxyG
NQi3CV3brAcrBkF1/gMlTffgGAUNCZF/9nUVKqDmYPTULlWkqV3HojFODqtxpzN+JkKuJmNrJG5i
6xZRQzxPWpMxVnFsLr1mnlODOztyv/xXoothb22iI0TzmlEaoSBGbrM/qp9ye6tfo0iawavOOVrE
uKIeeFrzFoe7kIhL3huvoNb+L3Yg7XTdr7yUfF9/pvYBjwzBK0WhxsH+8c+F6tPbivJI2CEbYddQ
JY/fW25DFZ0H7ukYNI5JdBX6mozAKwZWHT0XVxaCwRcdHfyrftdzzKaTHGsq6riK5gquvaRuvvpk
3gOEvpcjKFfxvvd/+Z+7h4x/sTESZfNhC/y0yjacyg5Fl84a0q26ClD3N21++5s+MVhRFRfS8+Ml
nuQsIxyAF805nEtpmPtPkLZVTvMcZNX5o9OfbGOvAhFSDOdk8RG3zBloQC9lWYPblogR/bMcd8ug
EhI9hywQY0gXkoKVnnAh4DzYnKvKatVjeDit0P599/Zg+l8fOcX2thW7a+fjZspxjT2vdKWbjx7B
WEyEKViP76yIyUIiIqsKkGcbt5ZuA0dg5dMgiXZFpxUNZqiQbvDuMCSWw/GjeEeSeqwD6sX781ck
3afoFSrSPMdgX619x9DZdo3nSF6J6CDbiriZWGU8MaNyzm6tZ1IKrHSbcECP9XEhu8ieUv/kYCxc
cHVGyHRrWUc7hF9XI4ZQt6RT+1PeozYgOKSJd1GRyh8xE+genFNx50dA0aVs8fD85T7PAwOMNiht
dqgvGHGv2rZANjfpoYw26xE6FiDGXt1so+IFY3yeZyrf8QF0AdUVyfrRFnQDCS79+ksY3g4yvqT9
QjcgvctfUMGsmc7RvaIv4aVAn5dzsETGM0gURf3YOPvFYmVsB8IxHMrxTVCa4vH9DC5rcPuXKTgA
fdgoYDjyo4jE2FlgFLsTY1mNssodJIRCaNiblDcQ26JpdhCYDlgkwGfAtRtyT2a55VCIs7QKNZKo
mwaGdXH/s60lbWN/6H+5aspCR5T3PWFFMP3qTZfCqg5t0C2r5yhz7gxDOr70BhbDsXkN3uTxJL1Y
hP1G1k8ZIeQ+xklSdv5J171ytxu2xS/iqdqGhPEhel+sIb587XEEaWtMKzQtqBkrTzGdp9PLyKOr
POz0zVRBckRdMLN0qjPMeTkU67zn1oYnfX4HHxix6jNWk2O64Jy6tsGCHAOW0NPVIZAkYvcrZ4lK
Y9RBg2QcBgZCJ+T9Pr+9RHE2gd/g+hYh7sxks8fq2TCdp+2sttOnVoMrdUXhVPRIcwfWsFGiZrJc
i2zmupY9ScHvKVA+nDS84RE7HrqSoCoOtTPgXz4+z/J0hb4Erfhoo7niAZ/GJ3wsGOw1xdA9LLjy
RHaKao2xjEyhZr6KxYyorPzaX3pDC3Y4Rz0UGSyTxbCYXPUzAHHylpS+niLfQ1qeqlUm28A3/lA0
XvOSwdEzefMb3Y8vTZ+Niduc9O9ZbCDzAlOTWRxvIqohfKQJt1z/sR9eOZdsqX6dZDVUZGqhO3Uf
P/kZKu1hWWBEqI9n2G70lpLKmScSdoPKSmZw8lGcOhs4sKYqMmT3HqvKYRX63Sqi0tKQM7pYSreO
9DqsESG4wgxrZyyrHOT9/Sfrh2YuEsEE80K8qXqo1azpUAgJXAyL0r05xFZq/Z6oW+rJ1hWoh3II
qPrOZsEsNI/50bqpxd75R5dm+UgzegG0++JhhA5+OHHghDmQeASIEI3iSwOmrByxB8VXGLsqhhWN
4+2a/WUyMQg1+4XN62UAXTMFR0257turvcXhfc+3MAeeWgJ9g+VjwgC430fxod8k+zYJxiwbHX+O
bvFn6vAbW7zbBtpOR2RMiLu2CFe9bWZrxFoecPALvs1DsL+U7XGF7DZMu+IKW2VvT5n8KVGTnQZv
guKo+/V3luH+Aqj5K97P1ElEdNNyBmIe6R+tHZjj/gu5HXd07szH796+xrFtO8exqu+C4xWCeAiV
/i//0ibzKKCRhUKmbVTIVTq2hfP657UQtnQuGmFhkoQbLzIuHZ/9p5nOgybZVlmUMWiLbPD3C03h
cUrfqZBsGkpUX0TrhXKZZ90t6z3B2Vo7rCCtRtBl/xDImyfLs9sUFxvo0pU0Jt1wfQIA4hjQu81a
Ga6APXTngK/rFM0AnD7zR196wF2okUde8eUnaI+Q+t9dCO0rLXSz+YzefW7RtwKOV7PSca7mjMdE
5xlMbKkcPQLBUiOxGjbilsC7GKIWwDUJ/Raxjc6B1dsGJpJh4RZm8BswX3MF58K/ZZCQE/mqPkLO
W+ZP+cn1Nt4mAHfN/gtawa28e5U+z7yKsvyvf1366DAStApB7SSwSm72ICDg93b/pl7VcngosqAj
PSFrL3DuHwI+Z4EG7LqlmX33jRDJFAxs4mI3sE032gmyK3JpMFVA/eNNsjx5LbR0MCawsJOCh1ji
8NuBUPcJiS+qxuVwpMOe8ZQl1Ff6KdRWjmkUjpt9PQoLWtXgC9eUmJYt/NaRIg1ptN7mw4otjbwG
BZXCceplPSUPmzv0t6EW6ghYomNwxZLfY4dCf4cwonNkWObydXgUV3Buna3ybMIi5BIrJHLRxBKU
hAIisgXrPnvD25zgB0VnWagssMJqC24CtR8LehTAhChKgIL4oNlP9wOtFbESVMNaphTKf8ESQGxA
GxinYjtWXNraZ5ICD3bCAu3nWqCrTJIpWSUUhDOo4JOoHkHHS+mfMfp5zcyIy2UIMskUSgwOUWEE
vFqnriqm1GttXar+ZrFNerCaGtQd2kwxqUKn3gVmo/yYbzsmUe9qS8EPCClG4qriygC/rc9wMaE5
NwSppVr4NqRQzC4Sp+Dktpj/RPJNT5mBrWUzQVZ2/SjxJVwir5s/z/+6RS9m1/2PrYK//wr9L6BT
8AT8+zCUvg9m6FOjwUhb/wH0tqndUKlcVqNRZvcJ1jJGpfbtW2r2zXENHoh7wP1B/d6GowX+OFU4
NRr9+tGMdRbTy1kcOBHGgw7riY/BjRk8Re/3c/RHsouH4HciovPHkqDlIJIe+r0DfgpwNW7VpDk5
LM3ptwIyL4jz6LtCz3hVGDzKuqAtkgVU2E9vqRgcL/xU4LfsDIp9m6MAvihLF/XtEQvg8VP5BSS2
4q97Qen4SsaL21TcZoZOrc1HHvhu7o5+tSgJpnr8Na5pQYOkIm3yuFBtMKwjY6SCFxcBA1+z3TpQ
NKWJsmjMTqpH4P9O6KF53yzt4mnSq+ZmPUKWXJQokHNUEwdi4Nhqv9ktXTNymSvQDtmIiAHpTEyE
eNut6SY+xfaBCwN67fiW7qo2/NB/0Wnf2JeMAzyzBwkj7kiOlc6DwZnn/F5IJp0lqgyhv0wKMrwF
BgutqkB7y7x1tdg6OBVNA1CZWCAQkk97bfkl3B09bKAm6swnB3vlwnGqQj5bzx6tVmrxi5y1P3IX
iKXHfbN0LeI15UmcjlVYosq55TwW1UBgNO+akXV3ejNE7jpPAJGaCkCLN3OjSnVS6u7buKOq7QMg
fKRC0IAwK+GfMp3k9+gfqznEg9Yovym7AgJT72Ll4VDPYpCJtlzs/rCdW60ZVQIbDivccJnBDAP8
AQCBLhkyJOocVmueI7R6nAJfBTjBXwe31vKtMgniRVM/5g8DKGHu1sU2/mhDSVCdBNaFtziWS8Jn
urk0WoGdYTMogCfS7kXi3kOJEC5YxcTwWL5LqmxB4PXnkfZN1YUDQRt4R8ZBLaBL9g+AVSPHWmh9
WtfIknlIPzmMoVaB/QtW7uLaICGte0AIOVFHpJC+0djQEay9zWPoTGMDs9F2IeccUyd4+/LmBduZ
1Ik9e9df3XaPX1JjQsndeKCRtrRWpmVkCLtMIwQVpHP4ZyiytwkeoVHmZBeIldBE3xZNB74tvpJd
JScIUdY2bN5C5EAvVgTeGEHlHMPpFrafJfu9vZoRroe81Sy2myyyaiGb7TxXZHBG5ibPqpxxV1j8
shtpMmsB+4DdJcefgt7liasz7fzVlBYSoaapgssi7aMCF2DANR5YLKjdwqsKg2CZ96ZIb5x9+RY6
5uV7uZ5Qd7HFkcvuH1SoEvj5dM/c8Y6bUFSlV9lTnJCYk+dnSzXqEjaJcPSEC+BAJAADANowWzjx
AIU4USqZqfgFlt7B+1LznBHYjMQBHlFfFnf/Qcx4iZNU5JwSFOwOxNfA83DSNmpAdcSrY7J4YX7J
j73ImNb5gXwaVOg/sX42gjdGP8APL5EOs7RwS5AYf+ATTNFWUKSydx+OTATrSTvi4IzsWMn9DcdS
3YuSRjXvDg7X6NPStIn/hLivIUfgRBpVaMHNgHvGeHh/nL8NumICwIirMFYutWBb1+tFmX7NH7Kz
2hGlx9oeeWViN21UGpFstVV45+/5v43A2QDG2MIEByxgAMqcexiwsOJI8vnYhVv809b1tHtlIZ9F
l+lUmYmYwMUnodb5EZFSgtFA0IRkrRwQ1RbSN3QCfcxxWr08gSIaSkP5BxeOhOe6ocuWQBiY9x3z
xEXM38IfYYyvjXWDMOk5qCBrjxmB/Njsjm56xdk6DGj82LVPxcTZDQw+MhB9CX+sQ/FqVXQSPlp3
00wLRZzxaTWgThcDVRRckpIabp7JDDDMgv0vdauh4VlvUcWagOF9ljG3+upLQiYxSVKlXn+bCklo
IXvlnZZmjbBVIZTAk9jQkfaibAgwJxsnX7GMqyfJXAMTYDRfE3A6nHL4od/0q5/d0q263OjYLyPR
9eqyu1x9EPci2B/5YEguWN+e1Cl94v2cPhSJgcP3g9YwLXOiQuBn35FVYpGbdMCBGKYCwqBDIGu9
LpO8iItcAb+duPr0IZsIdlI3wk8o5IfpqqY9RWf9qReqR3ysUHRmc1rtv8E3eSWiEdl/z/h9siDX
D11yNIyGmr/UglFrnfDbEYIFxCLEXytrlx8iQOq0aZ+SnkFFvH3PdknBzjrTQzEXSA6/YZUcbHDi
gC7anuR/03hQvkWjuwx1LahVNvWBwnIRqTF7S99qtPX0pKxvx14+QymWnGZjXGlTs9GVEfN7G6r+
aSxcQhhab4sCr4lqbMFGhTJiDRpx7wE9O3ToEzTZQqRq9clsw5rlmdW0um1ci4/F20+xpiz/X0VB
ggzZVJgekKGljBngBKB+t3VqAeDEnovznIVoBqf8BqrQDPl8qrQEMkuBhcCDIi00qwuOIE+ZcGls
CJ6kvRcCKOYhTxsRLikSMx5hPPGQkOuDXA4JUQ7wKzA7ODu6HuDd7rICfFb57wdBFrqDFVaR/gK5
1vqtipgG+KOafyj7ko38zn1UiAYqpXBlGv9guPaEJfW3oAP7YQCEAho6OdcFldorAJmi7MvqEkZj
KjpCNAvzX55mWiYdMJMgHre89Cs8G09y47ISI5BGy3VDLscw6oaIDcptoSBulx/GEP7gzNTtpBpy
T+vXs+zqiq28Z9NKQ4jD/l7p46KTTepqvQTqFjFElet9Za/XhHpa4Qs08XUleeF4O0utMMZAuFPF
Md5X5EtN2Jb9tav/jYkzfz0X6yBV9Csev7gmNfJjiQjWHiX9P536FijW5EBmpTCeASW98KSfrpYy
GMOIOXgU/DNaQPLkoOBcFfZBng21I5AuJ9HU+230EL8+LgEg5pxlSXvKRXlpFK6tJ+AbVt7aMccy
6B+lACusorumqgvjByeGIieG1yPQqfwv4qqnUXtrR9aIut6upFSC4C+d+jOML05QkRVMu2f8WVJK
zKS7Ciz99zJOIwG/NFEDEJvhKb44N+g4fpFxKrtML2utxoCQ+9dGEs3tBXj1IPJluQbq/jqZviwd
Bd+sqVEp+5WQEfXuywGvfamGMIsrwjC5WTcV/WT9hv5cYmbk7t+TtJFBAmt3n0O58LTf5Z7Zv5h+
iWaa1eU1FjNNa+h00sggXWuAurL8E63MnV6fpcfDIthQJWm9Os6ynrQPxT7/gfx9RiDOqCXR2xFj
0Nd3cvOwx19R7MJ7VLpVFBUT7WpW7PdLsCTT30EqRh67jLZ4rDdoqzhiPhfuLfsZssxdZbwB9T/p
5XlKkvBir7vrv/xn0/IY2+80x4utaSQ/k5pomU4p1TwG4bQArb0OVGlqNrRpzxhlH0i0tAJzHKoH
EXE/Bg0ZIPN4g0IdExZD+3QrSrflQbuLlEVQYeBaGZjsw6BTVAgjNvB6kkS7avayZYLIJUdZ3RJk
8SXL4yoQZt4snxYWaWRjfweScU7wvfnjwwrOMvw/MvJXOgRpLdG3XAeoF8/dY6KjWmHHVxlJ6SZE
3l5Cx4VoLQEStJU+m0Z20YXZS+M7pRnbB5iUdNrYXD/YQpfIv149yThZm939HLMiMVEXQUauGwFl
W9T3SVVE/1gP0fDcqOaLc+Q2U4R/Kbpl5d2sFC9zryff2ixSVPlQmqoO1WhpadyNErDWW/swmIlp
Y5MgJGn6RUkd7J46jnzxDLH2uOf1PwIDucEUhM4ewZT9GzeQvZZOcXY5bDy9C8AcLtfEL+IRFSgj
0PNWubcm27Nr6fBF5AVyKBNy2yrV9eUkdcmlPvwBIJXN/8cK7wzpk2dHoJ1i1BUhZaGggdNRnRAP
SG1joUMOcuv2j/M+BApr8w1G3d5DZo7VraNUxtBcziJWivsbwQQrvSpsVoI//qZAZHbtCpZUTWOh
U86sTXl4Nn15wN5A7sEL+tXp0QorbnRX81xv4k64q3RmMKNcOG/C8DAs0l0KkoP9J3nPCV4JOLzV
Dhq0hWfjssM3xgt+OZtS9Y4YGOjZklzG8CbVm58c3yvTS4bI77njobOC6GtKfYVlOiL78iEpb3I9
RB0sO03QfCSJqG44sQR8JK3FPYWd9oUKpYsM4g8VHrns9VI3qOxMnk7cobVE1P/+9wTTi21sE1j/
2tSoR0YWTgFk/cZDotCIZ7RxH+6PKTYGGJuCh6oioGt81ZE1JYEkQEM+75seLX8VTHDS7m1qeUEv
rRUYHEvNOtlu6hIDViJKzqSZRoIiLWDtzbj+9uGBmZ5hxnz+YbBLMhp63h+8WH0ACw39i7bRAfGh
22Dv4NGvUfmGUqy74db7XACXFtU8WTvCJbs1m506xQvJBzIyXxuvSeILMTefYnjPc768ABbLZfYr
LJJPuTmgJZ59ku9W80GNCsQjKyUp4RegW/J6mrgiccEbr3z01gm8UX49WPr/g3fUofzK2Mei3DkX
PGf4czEK6o8571yAvozwYnKtqpjGcWNoNXpPJ0PRgMyoFXmeVHMsYc/+z5G2nqdn1gYJ0bseADEA
OrIyQsdxhkgGbUoy17M95rjPxzU/7/wyC84/pQ10buY5q3pAGc1ZTLgWbMqN1b9nubIE6qV5PRWW
h66nVN6G4TpaqsEl2Zm3qQ92W9Md/Y8SsvD2hPiLLQuNyYazpwAvI4W2qDuKWQwnqtNqRHbbxrfd
CEWtb44Voagpa6epkudyrBEklcU0AUtd8pgMvsKS2hiU1obcRUTwA9TWEQ4ofLaUuF0Y0vHF/Ah2
eRyEZbT0Fzu9eJHYLcG7DtOu4F2aaXec3QI2AsZ/BBHPIzQDYzZ+mKsyrVhOaasEsAEi5n41uhnO
UWd7Q2k8H2LnmLhkosO0hw7bXDsgknbQI3lkbugSuskjPYJdMJZvdGwdIHITwfjXoD5aMhnbn8Zn
pwCZ3cFhAI1EDt7beBJk5F/VWKEsbnO42rc2qRF8ifDJUBS/UFrQSXnpXsRE5kSmjBrYMY1reTZS
NN0Y6Uz9+Z5r9usOGY54Dnxjv+PaxiNL7MbQXn6wOAGYBerNugnIBXfmznb4+ENf1VFgzQgWTrgi
+T8yGUSfDe5r4gz2bPRP9G9ZWjr34YCRibGVhl9ZPrTq0Nx9mOSYNhBAQfVFqso6TI0q5O7Bb4v4
rK5pQ0A/yNzIgcuZa5UBx78+EkkXYf8OamHmtToYOicCei17iDxjGwkabt0u+TIjbPnvoiY3N3us
6PIlE8VZca9mgYcNuNf9rK+FeOFTTcX7mOLRgol/jqDB/ktLHsr/sRB662BEUIH7fvIHqUX8f5Kr
744aK7xmr4dj3BLTHI9xBBbQRm1c0Sre7vn8VLB9fu0FIIlcH3r0CTJiIGMxjGABbIESLz1Oq3Kc
NHYTEnTWdf3D1AMkuw+6MRuCOOU8pJiCcJ2WEdD/lWnhaOy3/i8h99yG9i3PYoUmNzqDn3qIJ7FC
7NxNvhB18TBZfXIdn3ONasl0LF3j1hGIQ07yNH0Z1+geF6ceSzA5xFgQBGpauSdQbYfb0sV780X2
W2oHQOyajrfNI6mbkTxNXXk+M+MGeqb3L7nSx36BFEId+EaWDrq3nh8t1DjZnhtsDj1NcWCPKbJb
G/DSqJVvSAg1JqPNhVFk+qyYL0cb14XFK68WsBuN1K/oBxXyz/enCdq2Ru+15A/9qVlMyRlGdo0R
oT/W0ELFQp47m0cItkUp6wOHKq9hQW0/nbNL8UAczLNOeh0J2URXmuYIsCPrwAh8cpMk+z7kqzd0
rxFLT5z34aN88eUeTrMzTBu7FNzlSatr4IxOypXrf5GEt7L7P+IQdPFrpcD8CThgDTY99HLzU6uy
cHH1d/JDUXLqohll/Av1mv3JY5Lmekr1tvSztSE34HAtSmFYOdT7wSu10f6agPGtfTJ4UzLr2CjK
bCBj3x4252OyTBoXNQNhVeqiE28e3v6xBVJKhfKYZjfICeJNrSz1zf2k7nxW7L8B0FuTnxk3lq4i
txSB+yro5nuy4sk7Gb/2uZRO34emZZm7/shN6yz/j3ppqEbl3pJ3Nes+7UuDeT6xBAJ46zVpFt0L
ZDPIt6eh3cv7ENkKQpFSVznNDp6d/37673+G9xtap+Si0RimmqFjjMbMaSoDSXPceXMw7Oxnd8zj
1Cd8H9baE+tNoB+F5+8bYN15RDvX/QuYn7aCb6m5hnYqTryl1GV0ur+M/6i88GOy9c9aKS4pqCJx
NyHgClvxBb3wn5gDimqd826lbYThHTSiccaPo0xO/ZceVKMP1pZp1gw62DQ3+YZJNh/Ksvm1BLXh
ltbwQ/m/RvfjvKR1IZueJgqOUzYO4ZhRnF42w31ioA2ofRpn0OCcE3AlJTZTpodvdPaFn9XLf0i7
NMBOZoWAfvDc2Akdx6rAdqnybyWuv0CjVieAhh0w9PEKSIo2H/Cw51JWq1WEl4UFcMz6yfAEaEgp
aQoMXkIbvr8j8wrkhe/FmFYQkpIiScvX71jikvxEbNsvMNs/AFyIZMcINWJO0561uU5k3vHFWD1N
NhgvkGxyXDYTskxhZkeY400YGoYxeWGbk+zmAUao73cq2aG7UcI5oEO0n1mHmmhazhvP0Iq3qQYT
DzpTseFF28PqgUfQuDjFHDPoMeVtjE5QKfvYU81+QXdvd0htTVmYFj1cpu9pSUad46CrSd5En/Ok
2yGR++5SuUmDqHKkg7SHXGrqS3PfgA0ejbyPPW3vzSy53qxc3Z9fkAZh4It6Wk//vC/pzhbySPBQ
8Q/z15QMMdQJ9AIkf7OOIDyaOp+bsOPzPIxaz+6f6LktUvs7ol7XEqtTOEGDMYNtmwNNsCAJ+g8z
xp1oBfyyARkZT0fAmi64N7YCxYPgaZEByzZOYX9o9HQeaXQddSq3dLC2a2IxOcl37hJsmH91j+p9
V7eA8h+woG0bz7fouG/JtMCWfEl5NAIcq+Ge1+S458avNRABzadng5MMHwzhUyPkHKc76XqfrgXg
6n7R0KP1cLGJOPsCIcCDOVI7Gp3OSWM/hwfHLUmR7Zv5iDaO8J6CWeA6FhkpVzv4Kg77AILa43Vx
JNgeaus/fjqIJVcjz3aXX/suTKGS9hPsmsQR9nFyphEVtoauRoV1JdVHC9R0UiCfFGMgDdhifP3d
2zqNXab9mQETw6O9jvveBwbphfGuJXd3OUJ/xyOjujCPsffyy01xCGwfuMtdY4jcHyZ43ejQqIn/
WMfd8m0U/WgR0PotQgpKTdzW/ibh3Na7VgI5vAN5l92UVCveKe+/3kYhWv+gQHD9fP7KOXjFxnyI
y7QBsN/pqQc6SYZB/uE0rXfKiFL+jGOtZqfQkrkjzyDP8NqxSppdQAPheD7fOjx7m0JDUo0riC9q
2NeBOWIBOwmCcWIreMZj3t7caTSkBE8hJJlFRiOuNKY7C5BBKl1/qow4bTjfjoV2gbsx+R8ieCOp
alDkHxwrK32M2XpMn4wNxT0yAhJBF+WeKbFVo2kn3srYwWbBR1M4R3T5e7KZbdu3wKYWCIxjIK1V
J6XK1oTzLkaF3eDXl6i961QcARJIzAnq/1z9waK1SPGYXTKVv8+ic9HkFgDSLwzt4qh/Dc2g8w/m
48b7buYM0HHFDlvnzTEg2hsgdwHYrFVLu0rlFt3eUmKjppDTKrxK55CRNlgoCQXjaJP7U4jTz6Yu
CMG3NY//lFV91jf6133+X3rJdER5ieW045mFG+iesiVRdju/k6P2fiBYbRxe8znDYpaqCNadEvTw
1wos//mloQot5aMZA4/DZTFPUpNeq8Q0SGbSJZCzRcx0vte5On3gHY7u53gPHKFIgp3RFKIT1204
jLUfrbiPBpjXnnwlpr5Xwk9FdR7S+/AciKas1sI4eruvdTp6jfd8mZ2GRhjevpF4mZV3ExyqMFS7
2v1GvZ2kUUErrQcQUcVP8ntaAn1LfSFQBTRLjkUk6qb63k+ECoFlF0BP+b0HdfNK/45oisY7DJAt
aakZkymaYn8f0fzpr6fOwjEtgnSpODok5MpYfXcJI7qj8UEcScF9sTJLwyePR6P0I3LzX3hMYVNG
AR+sIXNGqAZRVKAydYZCkbm8lUUKWeQxGldzVQ6nBxI3u5I0R8SCCNdqTgwtz3e7LkuTiDUcNMXq
eut0TfhIWIpCx+7g8apsx5iQxfFtsLiwO6kCCbjOWSG106mXAVjfqbplDwcTSHEAA/CWKujJHPNJ
8AKiY3GFha1DOtiu/vEYq0rpAtwLXWEYGNgQtEo66hP4Qm369iIRrm73VsnEKfVcctaHjcz6o36o
i/3QnZeqhokIeR/o6MgcjrzM6ft1MBGjVCulWOv/uLbb2W19tiaIHqwyBkDDYeLr9ipUEM0pCaGu
DBH2hc3A7FK1LYfQtke2m0qQ88GFhVHrzt7F7qug3ANryOkScccN6mNk3jUXQdD08AEnp11k6IGt
eWTfBwC+J4q7+cqwZdur24pKD28pT9aGyibGubH37Vg7O/hyDk57anvJcY125zH5oZPsx90SbsAl
vTZMG5xWZMaC2f+5gzDcpD3IEUMzVTodUKdOIdmVJ+dMbysWXqpBOT2FOlsyd97i25aOmbdvvL/w
IGnppLnw/PfYKT4/kN8SVThk918lAI2xI9kv2KfYi+czCqkSJEiAmJ2brBLUa7sU8JZzlWy4fEQ/
UWBvNJO//bKMoseiESqQ651B5rwVcBIXZhEPlBDv4wWao9PmfkRkFKmvMNqlGeYAwVY3v9bkGwzC
h8xHYCFZVPsEQwob+oZcyfUJcG3r695aBNN2eAiNiHBAkYoZbWumaFkn4EZ+EA7y1+GKp2RG5yVt
2YQv5eUof0vEmdzj8YdqdOSpsReBkZCfOKMa0xxzIRMvrCRpQ8CkCoEINODdtcxfgmoFxeqeDKoh
MXgSPMw54Zto19WQIBGOR3YxPDEJgq0aP5GEg/z2KMFh1fjGJ4lZtlZYI9qCsrqna/FulvnnN8Xx
X9DjKoesuzU0UE+g6k3Cd82Yy6ijwtMV0WyP+yDLbbqg2ufCxFNa2Ik/3hsoige/v7OYunkJ+uP3
stsj+1U/0PSShFhaunsI8dSPVG6CNTc7Sjb1cUEUeZ6o+L56OHPUM9X2oczWj2JdaptmOxybSWj3
bb2wDgqac6eznM4zJTy6PSDtSPAQmB3SsYC/tS+xT5mYcCLd8NcqGsiaQQR5eEnxurkDMJFC3LGo
YWo0SGY3q71AXqdzb6C3kFdJejViY9ydew1hIMxG6pI6dkDFwj0GXt+B98GFyVlx3D3MOxiT/2l1
cYSpoteGPAanaDyUpwNCCSkDoXrMLAHcCtiqxZFOtP9PDp1iW9Z4NK26Cgbk/nxjOs1VIduPw9m+
0awbMgX0ee2d5NtmRwqV2RfdB+5CEprs+r856vt7v2Kd8romslMORaZidaIYjKjeKUZAfxgdQeZD
6QOnQX9kLrEzZy/CJm2WTLocLPwtxc3vI/tdgpFNH07jj1W1zX8T8e0VxNY1MbBwuy7L8Z/C8FKk
AYvZO0XsQYp2MishQq7/ftfPJahQw70p0azY1aFKML0RzuNJUEmERdKWN8pGJKJezrLOaHQ+xe4O
qz6PR5TvObuiLLVGse0C6Q3TN8MYBPtX6QeISzQQqTF6jSNvb/s1J2GLt7iGrnIQ83iPjDrSHZme
iaAH6myJnAkzYL92I9Xcmhs5cKeOtHJGjvC/7EOybmJ4Pue10FTaXI3qZWhxjG1wGOpnCMg2MB12
EYTarrxS/y7m/IgnEfPUKfuHiGeAaysI43gAeCx8o488kisdc89ZUtORvShdQV4wpZAt0jXL9c3n
ljCnI0W2Cm1NiJpkmZSx/sgiFoFQoD5ltHu0Qhyn4eY2k+jCMx+9lPrAMrhX9l/BNEY1fj6IM1N5
S//Y0tWNevIBWfvqA0HBQ8W40/mgTpIj0urFRFFPkbL7w2s4lYH5XYLP1KxMSFh2fVUIxO+vZLHy
OdLUXnKRc7edQmr9vJF/WLj56zN82VmbGPuTNT3LQAIzHh2utvJknGut1u9O+ZdrCG2SFGqWXfYv
wa+FGyC+18JYbCXnNSmCziB34WhGu4bNmKGVhm3dagU1o7TUcZ4ylFWg933+9fe8gAONrHbsFIvI
L96hf4u1MWJ5hy6HurWf+m5QQh23vcAoMD6a+/IoqHN1oS7Tmzy/vQcBsZKAmCIcaBY+jGc5QyVF
/zmj22CPzuTXIPCQikIqr4Ana8cT/QPiVKdM3pbHZjHcjSlY5SRpNsyuPuEbED/Bk4ujyUIi9H7N
7nw7JI+rbAPcT58llT0rZjJ9F5oI8t2G4EZm4xr1uhm2BWsnBWT+0UHRJ/OkO/23SkDiNH79aAYC
MS9zfhL4V3i2o/OB/5uVJhwjj1Kl7/vlOLr+MwKdEnoPc8YV4unXIyIc+vIINPZLLol/dbhJINA0
wZ6vAh9VMoaJVTTloMlyTpOrk2mwQBCiQvSWoHE7jo5iXK//3/5C/4c9zRGHUn8DczlidSUOPUnT
jUFXAYQpDys6JuWEvp16zt8Hj/QBbJ3X6TmqHDsiHQ4QASiEUZ5lXj2oZ1ilWAL0Q5VNXh/Pxe5N
lIoDsvx4DfnZgPRLXpcHWzWOhPfzyQsbCkKtkW4EqxSUwRraXOkNSzORgPKS6BtmxKi+7gKy73Tt
IEZxAq6/w3Yj1PPUB85D8KNQKgh4Phe4Gvhelz/2IMLYNasbjGVfBB04LaPMCxQxBZBYqnwX217T
2HLKcmUj33vjU1qRT7MZY3TVn/pxycS1dldyDdb6bEzpqgiyH8eu6UzYwV18IvM4AIo/pj+iR8XA
HmcFoBAgcISKBxqn2ZuFfnJc41IdPKP2k0AN/HAjkFocQYkvd+YqcjJYuuHdN4OMQlqLQ6Gsn4tC
k8jG7+ad4RjZWMRphL982tk1g3Qnp3fErnF2mS6tOqIxrpbhfaJJpcHicSDRGQQxSH7G+paYOIeg
8aLfJhEQ/vW7BopGV4vVufUz+L2yvimGcwEa66fMyBw97iLYMvgJU2BNiMcOwf3CpILq657EaFtW
BeMKvdtaupbKnlCdCbOWk430aPZkWh7oi3+1bp14WFpet/QvlML3AR1Sb1onyKnu32buv0pOwnkZ
plo7qkTai1mEDWnOl/+OUYljM9+mZVxCdnB+2pRzf9y8SAFKDHGtzpbjQVXSgAVTIG/zZ6x2rs8i
H4M/yzNgdcEB+kYbcmm/PWChTKxm1p4EHXyB+FkIJUzO0410cNSRCJml2VNkJ6cm0C5PElBOfCdY
2cSuShMWOETMeSwIdZmmfCQk1WfEVROwMS1SzGOd8Ygb6hDyVP8VP8IFgp2u499elHwsRiNg0J4Z
xiRVj00+tzIaMUPdgow7cUlKt9YvhTtBu0T2QofeINXGxEer5/HiJojxuUMMmhHcl0HapmVzO0fN
m5LlFqhhuusbLGcbeBEBs1cH9duzaa5C6D/vT4MTjS35zFSgEldVaJ6izWGH4uMYWBJQM0HWzNMW
ouoKKcsy33B9US2Eb2f9AklS34rjW61vAYufHhkjCTWQuzYDF09rrpbevM7VNslJMPwhbaMWsCs4
moqRv5QKCbECMwIOzVEBkJSE4ADO2jRxJ4CDfPK6s55hdOD6fqHWBPsYGtH1hHKWVSg2lP7Z464p
8rOs7cL8srWFhDrcWwbztt62T2PrQ9Ojavo8yE5qDpNCnw1qsdnV6noWGUYb4bJjxSE5Q656P2bK
kYvlhlPLfVTwwATVv36wGxA72jKZvMzZxpiDduw1jHpmb+FgCJOWMRz8TTL9u8T9kiPuxTFgiC+m
ENXIwpZEVmE0Yfp6UH9AYbJpZvEsbn6hLCK5y36MuOo/TV92r6+RqPaGbKUzIbjRHm+S4w4gUqVZ
BuEl9mkl9r/20n0a1B4rls202Jagp7tkA+UAoo7blp73rqJsgiz3LosXgEp4/XHkoRH6NLmGwJAZ
1d905JIECws4fsLegwJDnYd7g+TXBQdiLS3v3immQ0bcPoGrHDIugRjxndOMGeBPh523YoBAsAH8
7yRjOqgKGBL/EcV78pSaxODnO92erTPFrW+JFj5P3CvyGooNY6h0RE0S/mISGy1MTrznOLrXkVIB
nKgDznlkCAVlkLP05x+hfHeumntddhX+7htUJ9L61Y9OMoM6i55fQHsIUDO3VXGfQ+fnlHNF1zwV
OnC7FTjtNHW/wyfzZg0JkofQwR4GbaCKYvTr4lhai0HGHSl+tXZPdM+dNdO70Ws2rt85djOmVGi3
sbJO/sB17Tc8pA91sxPawVT7Ra+GToBq0JaCfbO1g4vNSGpp39DxNNwuZ4lsqlZ9zVXma7A8RDPI
FT+GFROFSEHQr5fA+tOdDBi+DZc7TQ/zgOnBesTVwl8ckYzA2frQ29zqoYCxReg4h+GZltrfDaP4
1LAZj/77FZiBgMlrvH5dOPY39Q1SDxshmY3EEf8GjsjsZvic9zZxCFVAeqV8KbZV53scCe+4ymgP
MKWv5M/Wp66K+objwLGtLerqxm7nDcz/psINNnaKMMZS4QIGhBdz9YGgvDoffqItuaGUUyOhq+So
2pxYJukVJPmqEpTP9ilUSmIE+bJah76i1LWXq9MfpGWVIHtwQWvVg3/rKZ1Q1p6DgBkNQmE5y0Dh
xhyFivE7sC3wUBAxiYKtSYszZHO7KaJSljadkabcwQ1J6LvBzGY1HMiLXhbgRA6JFSq01vzLlnQr
cUlymSkbuekHa7rwgZNBzNu/6T/AIbzxoxnnT51PPzf9PhsjNM5gY6XbQYPEZj5d9Mw0jUr+D8Vb
4/OoufnJfMMJLXDWnM5g26wOIZpPETe/NwAB5mzZWKVfcesMk8tbA7e+UpoEGDCeVqxYXoHdOEhH
Yx7lxEflsCRai8cCZR/smFh1i2nZj//GX6Hg1qcdP/mNvQUzEV8RT6AsIfRjm01odaF29hC17wHv
Ht0nVbrp7PFbpXYhHLIR5KjtjG+yDRpNG7tfo47q9YJb33YfBbSWFWCXNB8C4XXsrw2sKN5S5oUP
M8wYNLlcwItp1T8koskBz6BqLXRrsSHhrFY3eNZZWZlWB1vmKYLhUuO2cJzahM/XPcZMRz86q+sz
y08qptacWZ8Ai88oORjkWot0NOSFFXFBj1f1P8RTxz6gh3fAT22jrQ6kLejOqszPDZsEQ4QJCAW8
0RowSUn5PNB2Jz4Z12Q5HvXc4UpBtUmbl7dxEru5eIJO/1bJcqhAHdNJByxLdzC4SKOs5JlCBtXG
6O6NHbBpKMv73LMGF+HLB9ZmpenY5Uok1umDjvdOwubxwSn6cIwLVAywp72X7EaO1qDMClU9DiwU
nh5r1BqL74rIzNiA75N03yP/6f1q4YItfGx3pWRv0LbB00y8+AE+v/WUR+gSRYDiBUbFSFB8YiGF
aU8MEM3bdRjMeHCV7nmlfsa+HILmhZfeTvItvYTQ37k/Y8Y92Dpr4c6oHUqETiJWn4aCzP/jenBf
F+61eF/I1rutN1v62xwm5MWFfDiV8CIUVVzNFOYggTibgg66FCLDJI49/24LO38w/OMzCMbfzA93
MgkwO4LOYYiTgnyHwoCDe9IIQbKUYqsDL2jgxxfhKH5OJw24L1uzPYiz830A6QDHZO3H2cL9wBki
wSEvPvPtfhCFvJbsoN6anLeqEz9uULrUGKPWojyn2jK2AMed6WjwtGbHZ0WmBG1iu0fdBzi8n+zN
ES/oNLwG+FkfkdogF7zu7t0K1NHBhr/+Q1pFsFusbswkzzpFeUJ0WBFcpi7ENAiBzNd2lTcHik21
HbFRbKKSajVf9gr8/po9sDO+oMWIY3IKwVdSut8q1D89RcTmLZN8Q/wS0nq54aMDskzOupiEaQz2
c9DTjHvMduG6uveW+s7clEePgtDq64WTT7qMsGU0skFPocivoXxppW5uVrHo8pQF6vq5NcTw4rEy
i34mIsTHFWD78tCRfw5KnpyJ9J7lfe36Grf07WU/GGaOzQurhApqD3cP+gC9yMmw2yJTdWCWVDl9
i7rDNnVmqWAuEphiYqTs78UOWzoLDn3i3hHgz85HGwV933I+GkMITlwZNcvE1EwrDZdKrx2Whnv2
d84BXpcF3yNfT202THouRVsAHbCV5UJ1nFs62SRFz4nKXbT+HOk3Vt7Lssh2XfLRRTE8WaorixFl
m3uOEQ0R+ZiSSK1jm+oI9b9B0hkyGcfTFwr2xa5IO1+Bt9urlB3eE7gMNAkF7xdWv20VENZaUCsL
LncHcS7Q8gRDlF/jAJjelSPhGB+lWoZSWfpKa2dGtmNuw9iTw4dt+wSEXxU01iYGNU831jmCbgXx
fZtSB23QSM9z2CTb8OCr8jQq/pJAbnYZLVfRF+jd4kjqV0UbbLcCpsfhyyWD8PGR4McZzo0kfpHQ
I5+CeAO/5yBchknuNFBEwnLK66xWmMhgYJpbtAOrpmOz4GTnYolkHA9qMLX1QNXnk1f0t7yjsmrt
hBdtmfXmxbtgd2j3mrlUaDzhJhX5nins7gUqhrFGjnK2VYSVpThzdrgzsvxiqelH838u9gvUyhvW
CNh+fUP4E3cKsdbTD6+LNNzUyQL8ZA20UVBb5AKgurn0IV0lkJT8hn82Dyr/BCFYGDWamXDoJo5u
HttfvNC30TBhJUQvrnFZU5XPIm4+nR4cwJiJTJJX2wOas3UtlyKMEXuzBzq9GYE3CHqi1BBjWXir
rNTkf86eUOclWQbiy0lHE8G7l+zZ8GJnIVZ7U5TbgEDpsJKG54WT3/E95235ZLcXIQwQsvoG6AQt
DuMYRme12mnJEP+MkvaC7LRZgpmgDnbvG76Ugc8TZbZW12859dOiCCTqEWd0sDHCHO4QfmEhBpmK
4sc4VQD0YGefUUWj1thTHxFB53BU1IQWFdWPSuHXViQjBvPhne+TEOqs+LS1415UVJBksNsogHQT
ItuJx4yJ1OpdBq+xaio95iCVvn4uS50zE2Wf11lPKzk0nziNeQGYqHzq5xsyWO9k2h9Gr9L679PS
QiMyU/jbqLDMxZ7bZgwW7xVcjb4+z36w6yhxbSBcpVSDsLrYSurXsY1JGhNL9jolEYbuHycghJVg
+Jn/4DHkEmq5ZewuXvZNHbb72nW+AvEkRDL0fxGWDJQFtpUYkhnSyjILY3fhVjm3wLI8USihLbog
fZLgdI6ZKjH//d27w06J7MLL/A5HrcVFfU/Ob2bMGuGmXWD3RpriMvfGw+BWW5PQN88iOwwtPT6w
2n8vsj1wQFuQO+fHco0UfQWRfL/n18OtpbFaDPa08QwH8AsGK/tAs/dstY5yICqjfcszz/N6xU+5
YEGIjD2CmcLmeDTlZ3vYPkPdbYTsGt0o7zls/4cdi6yCWXGxHJwJ81KcVQfV+y9Q1Ak/qo6avIP4
fujnFFs5v1pkRZHBdBQmfaV1zFyxv7nkbSIpRJYmKoBcOyiDPZv269BZE21ECZadnUg5qF8x1KlO
ibHRuYqjTd1WQ19+HzzZpKhqEeMZRFQ/3Kk7wq+bcuGQ+OO9GYsKwoyBSRg+bNXRtKpOWQNp+RP+
4vjxzkiWc12bPQmKos292Q74tYekxIYz3rfYuI2O+CwLz8MjDhpqTx5Gav649Kr2tKGjZ6F5uVJS
GeASyzRSBiDdr53O0cZhUxXnPxzurlTxyGI86N24MEqZLjNdVPm0FwkgZwZDTYCiL6W/x3xGVoRH
odv4J1VWXJ7C2zPF6O30qIdYQZvlPi35n75pBCAi2Lqj5WFD5tyRNtaSiLVc5nPcbMwFOCXI9KBZ
x+wqXfqpCiPo80DYukJzp0HvqebAMk8FV3CUgdMKT25h++8+P07xgYoUCG2Ied6QRTp3Zku+ZAKe
cUPtKIh257Sn7RkHIWWmgeNFql3RTBvt2s7IWQ67u+iyluv3HeDQXRinZ3i2Y4LD00APc+KEfaZn
S0tM4d1hSNYf2WaW8/BaTGE1XssyT/rLcJxQLPuhXUJlgX7RNUumF73Qj24VJnP6s+OHGnIRAsR3
wRSrz7ZkfdZ/uWpohqhQn78uku7XBKXiZeQz9Ya8JdbsEy88aohjEXoo2PEuG1W1Tq471ixr5rSI
2Ww07h/zIhoAPM/InHVqAwffvJxGbq40ecV19eKfRr78DEF8Rwo6Zkdmydin7jN+HU1JIz8nngMd
J7pwMTBxP8FYVvNPauqVBQMIP0UDiu9idzbM5AI37/fNQVvqhTnt9I+Vu9+G2YoPVRWnVeRxkz7N
Lym37jSTMJf7pn0aNsFgR3qJIfvjBWnoIP3/AxK0QUR1H9dqPwMAYWyyLWa8zWe1S7Jx5ZKX09PO
CMnQfk2fOvkF6XHUSqWjovu6nBKLaK64c+UaJKcQn9wgOtVG8dWbtgA7ZYAJKx66Czf9uddnr0SJ
y+DRUOxTRPVtIydXT+gPx17J+SJ+z2vzJj6ZZJi82gJOBioYQxnaZDBey6ML9e4KcNurKnBXOAlb
YfdNhLgBCK4udaBUKCDiVGLXiL7p85lMpxo3ITW+FGPN0/nKamaUufk9YSLjrFVacojPMH44xYa8
F+ZLlqe5PIYS/M7auEw16BaZnw3vKZ/gy7kVH/JoKo1lBwan9jCJXNBrEPFUdoramGO5JJdt+xlX
r+g9vRLczWukULSftqAH1tMFLhXe7t7ckAIT2XHn6jn2OZCBYVc5XNn9NLook9owwkjqo4Q9lKej
ND+21JoJhWDnoJa+BUAD8x6zs2IBRfK/YazvhHkBunK/dUF9pTMd8FyeFFCcbV241tKvOK86q2vy
AH6roAJN91TY/kQb3CRZfrQvpcYnCtYbTJLMHOPFs9LihWLEnwK0MxxXGkCBeELLwu0rql+LEKEM
b/Ciw6go1YGISocW2umYBnH0N1axRONr6u3C5LGl/+01/ZG5OV1kQ65VNUJ9D75j+4P/iGZeO7QF
7xkVsVA41LUkxqZVf92TfH4VPe0O6qWFI98u0qAtD2RncMbN/83O5Aqy+sE6mU8KEv+Di3KGQKbP
1p72mNR63gIoXK5tNl0OdM+Ij6GMBJxbSFRPc9+i5SS04NAOl/SnBdAmER8NqjEESntq2MS8CM+G
fbgH9hHu9yg83re2C+EfYVfdA/GMBse+DyGB1GEJeob5zxdvH+QtHHo0oyBazgzY4b7zfG8irOGZ
VsNOi86vQAwUyLdjYD/cmCic13hlHHdhgzKjJq5rNc/0fiWpMYknQQDvKI4NXlrBHFbT67OLiFfA
EECX8j5TUghsSyRe15rsgGLOKR0VVRgXN+VTRh3yNY9dYjoU70f90OQHgAlWEjAMiqCKVZ3fDwTP
gGlqTrlwyzedORQjiWqfkJjItItHjdkclUUnqKXq+tlMD4gDANF08EAbcd8cSHchv7L13Rs+3lTo
S8QBdZnoDutSnsyvWsm2CYqcqyWO5vYU4wvBzSlJBSgm8en3pru8vhMc+KUwc093kYI/CL1+i0Vl
OqsmCPzROdPG2gszkS/j1hVjjOxzuk873tYq/JjLeR+JOZzuybhInfdOlQzhr9KCAuo3jI5l/tsc
xgD2Q5+cWB+uu9SfKWAWs6FDNxKhJn8774TKxZwUZ7bry742ACGgSeu3p3PSdSdPhZMmaPqUIoG1
L+hGGpE/FKXsQQJ4y0dI+3n873M9lAV1q/84y17St3ApPDDesBgBZQg82q1J948Z1bVOYMQen8FD
T/h9xQ+LXQo/AwWfeeMld9qkMOza/ziuu37EvMRWYQd4t660uUUN0BqEgWBsXjBrBydljSOEcGrL
SPMdaoCN7I1XJePKgj4hBOV8BgQfSPlumjIHHzO9Ozf+xcKxlDSws9/TtRzjmO/ePNA8MY5UwIjM
p1Z0CyfLkXktY7xZ+mZt745SZWp0VrzsAU3XnRtSx9N0uyr+JwZNa8bONY+/QszXbzFZyimeyKjz
WYP2h+n29bxd4yxqiUEHsPWZdkRdTaIqtlkxH+iESsdB7XzGavqJdkmZqPcCpuoRXbrwksA64MOG
Cv2aT9z3SpPCCOtn6ULh6WGjeCg7BoSwiBwNyU+jsdBsOMKdWTH/zOwGDrN/gpcZloiobr1BPK53
PbbMhJzgnQTdDD4trrezjLgb8BLjW+JnbPsXlbsw5G0Zo89Q+4+T2tNlHzDc7iLwhr36gS56EvTF
JzlTTpaC+1KyjOxjuZbXzh7KaiTtJZmyJcJdFzwamq8hqqOLTeVuMNFgrPyjpQmTSJMATdFXCOnU
Y58zqgEosrFOfaIxs9S1SvV0LVBkORTdTDx8/E0brhabgpxqeS3uqXjqgjRAn6tOZRXuj4NXCbG7
K1OPnMINo5/9/doPuHNnTep/73EJmrrCh4gDBuRDrTLl7I705usAN2qKZuQ7ttn+EGyA8X6Mp566
PdT7D3Fbhf8vZcv1ZBEhdT6LeQIeL2I+vCU8IPsGgqDPZOgzn9uZO7EKlT9u1+iQImu9gK9j2GpS
CmXOudW4BrMH6xjhT4f6tEIEDEm9dFFrViMEMQ9PYYJ3GkogZuDb5Fg1sjsJ1UgXkDKSAKMcW+Px
XWZvmDQLdCHhhcBf8Gjp+wXIF3caxPUzNDr/WBkRS/eaRtY6NqzyWEWVLO4vhIeW3sRuVpopP+bo
H/ilA0P9AB1a8eaTocMgjsXUlweH7fgMDCQLZiw6RdjdZbGxIYck+YA4xJWeAPltaEca2TJEegqA
ZMtzL2DKdwZIIVaGBUueRMv/9FeUJRJhXV/6x6j/I0gbVb2xzlGkNVfsR4XJwP29xZvdyQ3+xMC5
WDls6Ei9TrbSzgKay+TY2PA158j9VwZ2rFcVoEtX5pKcRh1djBI+Vx3pV3RArjQdYv8VgIiEYn1c
bvsgsFAcJIYxGSN0IYFNUnuQ04FHFnwzCXr3d++bwBlZtiDAWdQGNzLLfF2mfnuuEBNqhCa+glA4
jxMr8et71rZsWQBrr6BaxIwPLZw2cTgmYs4i17IJPx9byBQ2IxWvV4FHoFE505gbOUlUovGOPp31
Tk0NSDnfvcFoIuCKyk9WHRJJmKn3T8x+328lsBPruMVmg25ZDjTduwT+QQ6xvkm4xt6vYPOnsFbt
Fqg4VciBt8lnIu0OAbZnmU/onBXs6PbPNCCv+AOIoVpzbh0aUPSOLp+o98oP2nNou3oX1ETXqydL
EeUaQy7qfKzYWO601BTBk8cruywHN9Livj0i2gh3optSFt16SOexnH2rSRGaRQOWUNkVSk+EyRrz
z2gdgzuAjI7MtZjcwYTrNB0bmg45rzrthFIxkPa49XGDuvhzzofRkvudnWD7DiptWmOM/fXhWO7R
p90JMSPrKdGwlMherrQRDzApURrA6YaZH5uEh68Ds09tiY0OVzBuQ5GaR8u2y0qrJz1Sdk6MIpAf
9exYRsiPeu1OAhNYUsAof2Oj4hqSEtHE1y1JWg3jxgmeJ2crGdoQIYH2yNKGLJGanXdchQIOq8g7
XOBwXUYi0nSP7jJxhKeDAZMPYsoojKfk8RqshMLsz4gOY3YYp6g23vB3YY+NuTkRT90i4n4WiXSc
4Zd+RJT072ouFTSKYwumlhcuLVjh59bBnVcG8tzmaxbsNdhZhK7Azx8HZyCTvhr2ZzW3HW6g6JCZ
3eE0HgozboGLwvrwgm/VttSA/P53c07BltiSOVN7fk1ysIOVB942S/SmXz5SlPxt/LidVDkaVQXt
Xn7bAJrp/FhRZioaZ7MLA3NcBuVhJsWxCFQutccwiTU9Pk2+kyBKTQ2sOl+eH46ZvtprV6h4WUBE
b+S1cfCma8NFBZuW+oagXavnVRK4PIF6Rk3iting7m9VSFmnr2hp5tW+Cyux/gd7A+dJsyLVr1dq
SM4H8KcEHm3U+6RkwRE8beE1QHLdvWyE2je4Pj1Y4Y/QN5WQCGso9F7VfHJcSdK2FUwTODW8tlD+
8qNyNwFQI9HyyKxPbtRtrkiNdwr7Xl02QIzaf40RGIsvD3WWl5Ayabgw893vCe4/2mi9+lpeYfVn
X4iZshTRaXxZGrMH8ZnwHe2uXQCVUCh+m/PNT+tQ5jn3cuz6qMUe8MZ5bIlPXgPX0nUMMFs/JUqG
QWr3a83xOFOlO+aMKuCWfedVj/8mHCUxCRl+ny/9Kn1GUMqen5zWqntymAsEEeHcpI4BNBoGv3Mv
MuAUPtNoomt2NFIU8TDIwQy0fhND2L7iAWYFQOWcW8L7MYSiT/REyJzHteizr7LOpdltB3hW5H6Z
D06BNEu0Ft1NrcWDYPzy9a5MP+mPgH4MvN2m/WomdaKbl94+E84Qbr+ZY5jkz9dGMfGAZ0dIzPD5
2W3UG54ySMxwT5LnKdFzxyFhUBdb2pVFe8oPAAvF+mCsE+zFjHVue12KfIXn32wt7KccjTffJ631
mCEl5Poj1Yrb+cJoQobEJpXxr1PWzgnxoP19UKn7AXkwBginetmpqqMm2yeLV1PBIWjAcjEv3riY
kRIA4AQmm/W0/D3Db6LvsLWrFes5MHE7V4t8ACJ9l29Yr97s4hWl2qtR83vMfmSFy7ZBtCjy8ejV
zpfOA/t7zLKY0NTPZbb1RdwrU0dmuQfFUjzSktCsb094asAZaLt+itD00tVRTSRfPmlsZ+PyWEcU
FJaR/4tx/BF4dENchgUrSINqSpsskpwJfFjeWszfWKiGAqP+WUa9hSC6ODjFiUOFxBB5jHoLgg6c
Ge43yH3iH5x/uNJI9dVZ1OYnVJkkiSwk8FG8Mtudzu6Dwmolbeezg1W9z6IF93RHzXKkQ9w0atPj
sxHD0nEizImYWtSCvaL1SC7d8tLeDPrPzKjJbsRJDBxamTBJtLu6cjp8ORiPanpqqwHlK8R5NUUd
pwJ4jqMvYRahz0qzUzhsDjVkwL1dNMLGQzXWtiTuTCR5bAEQbQ/VHh4snN+T8t3ztNbOd7sn+a+m
manyYod2y6aEujkJF+H6yp9usLobeRQDcSVA+alDYzYiwnIKgoWfk8wFUXxIAfpiqOsKERAG3qKL
a6BULeEtLa5cyG7KSSStPJkx+WGJ1qv876dbbPEYaR16TbVOO5xdCJvwfKvrcKizuXi2+KbBnof/
mZVZAgMUgp3lWs84rA1dKTBTh+Vg6kSMmd2Ef/+gRZuR0IzARH42BkTR+8yW/HPrR9my3gA5p3pG
kr+q3qkOD+U2548VieyxHGX9yU8ZGhueVS3/UIVFWxvuzUtFrR8BG7/XMJMcVWpOIWGW/LkFKoPn
dyCB5UsdPjrExAMm8xo65tqkhXfntSGzyB2b8hPTE4utg/JYqWVCQmH+bH5FF9ASvVaRk8U8Z2R9
8yH+K5n7nNfwxJN+7yOW0zJAgc9swNzVPN7AZmNsDnsRldlG5uNlXaM4PZN5Ag394RJt9AvsreSx
oOyklXSNejj+ReKPSfvl8JILYbh30hXZne3uvCruyak/S/6UJczk3PClR9l+uqxXzCfrBI3ZFTH1
9lmlRwX1E9/Ff99qHCnX2hGaiHvATqYkcQx2N2izuO7TgBoBgl5+Jbe7U0VCpIv4zeRQRL3liBYB
iJC7KGFNSuB3ZivT9Bx4xQDyJJG16r8NxzChdWwmONEBIZQ9A0HEWbJ01RKchhRiHamv60bpGHSm
ZSUB9oJU3GOAgoedaRux1eKfaGD5Rxbk1UIGkfhfGWklwJ+aZVIdYhfv0DSDvhgtVsPfC/en50XB
U4VO9ZdsuECmlVfLsaH7wGygIrCVCclKiUIHwqaQKyX+SsaTeY87jmG0agckNyguepwBX+gKcQLA
Zvn8x4ieK21QFhDj0MuRr7o5Xfs8jQqxnqAR55tv686PMwR51uzHUTw9Knj7nA73fng/4FXPqD/p
scWMfqhdyoWV/gBNEaMbcwxTgPBC+4RL0qOBdCWfaHoMTEpYUdM/8hV5vY/P5gAA8o9sQp/MUina
AuwiKnznkNTqV6mchEi6iGLVlqLeYDR16QLngCtAg2UHLNMQfvpUZxc06gPJZzMGB5Wf7Wju+H7N
OE/s6hZZlKE1NytjD1iXveY31hIoXysVJ70XnveRbwt4Qn9p85JsP0QrSgbfGpkfcj+BQD8fqwpq
jQ063ajdDFU3khXJU5x/ZPuwdWREG4DrBkBad2eGE1gRA37v+o8KXV+E2Qte4kEp3ySDdRgMNi0N
Z8liMHNCPErNBnspXUdkvPC0qfdbPWaXfZFa3MvaF74PQUUMfZSAR32rtP747m7uRylWHr4FnZKe
yil10v+5EYFCkzT9WpqL58yNSR3V5XOp+iNULxe5mlRU8IulJuTkcGbXMxChfoAArz68f/uL4Lek
2J50R1xZmE67SJk49wEh3FUFn9d+aqSrgiDOPnXgadGNDgMq1F+oC8cGOhWHpLvXOTQ9/1eI93x5
hDtDY1RN+Ghjys7rQGVCeeeEVDL9fB18sDwB4FB9a3VFIz3866yqvCn7I/vG01RRokZ33nFxDNS/
btOkzRgQizSfxXDMMyaKL2CjLxi8QL753T0rxZtOZpconVtm5nCsXjzySdmgK3tvRt2NQaZvzZFY
JIJNTxJ36IxGkRDeaF7Tf5/iEajYJVYcdWKbOWaG5doKfLkKpXfDndF288Teu5IwGclXrRC9lthK
GBb/bblPFZLt4r5IocDuEN3UkW/bzsM+OGeww0X/MNnp6XWubJuIsDQdnC99335JXM4Kzkc4mvc3
Bv95rgul+WUiOMiCFlt0WrZ1xHppP6pcpnabWyvGcT1CtVdfY8pQgAS8H5pYZ3GQaqE4+01HdiTT
oEugV8lHQLthE4t0yQ2FV6RIiQZRw1suSC1EhLRNNvlfkozF7wU4WuS2ZQl1rENfdcSqCk1lrzpw
J62L3oWluhf1IPCwAVcv8PyD13+zXN98+Oloa6OIAu6gm1wtrYsyoZpkthjNQwin2ZAGT0lwPXZN
zewN9G/9s3RBK8NvgltEExm3dWU17PMnpBUetNDjNfOzM/ilPYempDBA7pI4pson8jpBiwWMUYzh
Aaj0TDMAGdl+RNC6OZPKrlZidG0S44b77is63VHQU059S8eaNUhEaMbqyL4S/3s4v7iH6RwfdT89
bhhCGu24z7Q7/+8H07IUVk9g2mPf3LztJeR+6BwyncKQ3hAFaTySZRIfGvab5bfW5d/kqgAYNG+f
4pqtG7eR8r4t2KEgoKH0pwKXxgNpwyCQ1xC7gUJN5d7xubdONmxM5HCkaXHJ2c7JaTCiW8lm0YVd
W6r60go+42NhMM411oDoukqKRKXsR1E5XS2XhGJ5TUmjh8PTM1aAX9w73TDV/6kGja4EdJi/eMhJ
ztdjpNRtQDt6cCHNjtzh8MJNdw36OBe1oA/3wGhMqYFwkIbnJf/htOY64wvPFIQuhSX+PCZscSzn
EjCiRHFindqke25DDzuCEGKbKMrt8MLTyDhLizNg8y8Y+AYZKVuKm2aBalrHLA7clyHuCbj5cwe4
2NZDCfF9cj29t2K6VivqGHJiC/OF5sj+ZduPkWdMmhVRexWKawht2+/YY+nTR7GU1tkXKHN2b9s7
Xlftk47AE2Ry0ZYNvCtgK/I5vpYF7Hcbs+54ks8CN0r2kZwwMSevuHUyb8YEOdaFNxP10PKsdtOM
6ybV3tdHOfhEDzPtWhH6hFiveamB4ipbG6ZfXxeJqJC+AmLXCgbeR/JMJsvIGt8riFNtIDwhMr19
ORs0aFZOgczbY9jBSe/MaZZXwL7JDiOL9GCGF2lzqmewdsZu/DGTAAfRdj8pRHtqAaWrqdFT9Mmh
N0cBKTyjRaxhocoBuvkNiE4G4h2GdjK4uHzIiE7RWRWYcMABBbynNrxpYS2VDfkaON/aOKG+kiLD
j5jeMG5DHg8D0xfFXCiK21PWXXftyLM6x7vUgywSsHJTwSyeQ6NqoyaIsc3JIrqq0JvcOjo5ETez
Q+wHin3VMbb4tFudELV7onYv3D12bbN9tzYHZzx5sjF1qVFj2bU1G9CdGGevqd/3JsFoWWJoMoSq
Bx9y20lzzW4vAlR4l/CU8FrbymmHtRq7K5YFezChDiHkFrcB2aodtgyybDM/GXFcy4bzkVj5934B
dJ+b9EOoMISibHC5qjoy9OLnyqAnu9qtLSNl3sMKW7AC20ptYtSi8Mj+5wgtMaNwWZyVI+kmG8do
47NZHUQnRJCyOWsoa/R3Z1RupAmzYHQY4sWX8yfdo/a4/wr3DnniCWV4XPkR0Ef6waUVia0mAh8A
jeL1hCZRt1WzD4dy9YvZlW60ZofLJYmj8ZusHXMeox/shgoIOHAP/DMsw7cCNB13mgqrApHK1IFo
LxBNUBvS9Qm6N5KslIy3z7KSu4tXCNawpeKWmjDdxV+wYKWDcIplxXfA6CYqZwXSSaA5IPvUXNc2
dRxQmAM5C1mOihJrK13w8gLu7h8kVegQrHKRSZHu0e44buDkPF/SIqpStwyXF2cJLljaH6nU3RUa
aAlfkMIiu+nyaU5K0DEdT6RAx3YAzVH2EQ1qXw8+2c1h5VR7db5yhOOyi6+Gtu98XqZVUofEW7Cd
cCB49MHT2/PoOY9LkypRdmh4+yDaZ3U1p8YD4qGurKDRmt18ZxdUbQFQkzYwU7Ynws1Mt6qc6YdQ
DSEJwIFMWMpHYcsapJLoGUfaOMiQgqUJlIHpVL92pOTKhF5Np/HKn68/TpDEAw32HkFeLm+ZstjE
kvrKz2ulresHVx2ClMKDi5e4t5MJIVu7xc+mf0LWRKE7cUDxmbZOn1bNiW7o7wKcg6sQ740jQ9QB
nJs7C/VpPTYWv9/QOp2NFz/cSqd5xzGmnf3oyxh9F0JAc883DIb7GXrhgy//vMlli1kes6rQADdW
unFCqlmmMAfPnoxDXwsk3Hm0OjA1Ug6aWpfxFWckgciI43ZukIfswIAusPfWcSqPvoqaRqy5cgUr
4y2xUx33D9jMNShV0yGa0NWrRnfeX8MwCwHJ37xuGdha+yXWbcIrPiQGyMEz+fh9yfwO/ppdDrob
v6nrfIuIUfRVL04AHDt0zbpcps4n9I+RDuRsLZ2guqzab0AhKq8Ky0bdcCTWFKCIoZEqWahUwQoL
PvXjwRUAN/0XjYbIv+jmIboRgajjRgnsx3+tJA4wNYDS6EUujXbKigC2b/LvHRykhJp5D3FZ0J8v
pS25ltVgmBUqdctcbrCuw5HvCml5Ofo9Gd4u7HCJnoU+hm5vq5svU3J031+sqzb17T1OMTwCoHCa
dzC42uuDS7j6yDuVGy8XoDcdaX6V2mXzCzUC7dpSDQnl1J305jqbr6LAkHy25npjhEVDYZmYsTWU
WAPlrJNs+zeYEF3ZM1TRs6W0VM/obHx60EmgS/4VXHvVnf4C/H6Paz96kBgrWnJodLQq6hlss5LW
B/8IijRtyCxTtXzJ4FExG1VO//fJUY1thJIhwM7IqSRiu9HKCM3uAfQXs4zKMBxZW1wfTo6jPvRU
9D5tlqmgiOA4uyUrA2MDey4edo9Q/HgXIA94n9xHtLs22nY5Audx57LJwfjyGwRRFEmzK+EKR/uS
F9wjJN1VeH2JWVMf//v9uZiyxwt+QBgtQ+0s7tE+gL0JFGm66UnNtyohG/fINFoWkL/C2F88fEPE
XACzv+CfIlopDEAde5elnftInuSlR7EFauUE/iLabG1jyvFYUGGScuKm/cGTAJrUGi0t2l/cILUx
/KWGqlSOR9njJHJZA7oSsQTvLSmBB9PHC5DDpE26Dn1EdLplFLJfJe6WMUbugi20M0DsTzQLvpMO
a+Is/5g+2ooisM/AhiSyojKVJ95mv09J1UYDTRCLnytezT6nHgvcrI6i/eUeh8UuzfXVJDk/Rq1h
RFNT9YMqx3PQq0DnjdHZbBmD1znet1hnNheN71CTyVN+enIwz9v3bTKVzKYUHl+2ZPPlpHQEqGk6
JE2rMYFZ+w8gxb+E1tC4s+Uf/YJBr1jM+5tNlYznhtdNd+g0LdIjFdj/rRpHCwem8G3gioM4Lnbk
1vQTGiCCVoFgKi8d5xi6FNPuADabEjbGcMICoVxYF+MvqVF0nf3u/TdWmoq0K6BgifezSlGWyGaj
1HhqYg3SgSWWQaRb3IMVS7uxq18czChOx/dAE7zQ5bs9SvS0S31Yl/AQtOcuSYxklFLZ6YLcqBQu
tUxU6vJGyATYP1VgDh8LB6mGhGjhGYpUIjtjOAOElkFmAlpPhe2+HBc/1GgOoF/SMXLn9dSdHbod
Ui0BTmouvli0O+FJdXl9bEhY1R7HDUxp9QclB8B/fx8/P6bkfMfeSRor5aDd62OImatpLQm+gGl1
Mjv0zviCVt+7XszLQ4EMuAzIsJkwHz7y5nStpRgh4NU7bLOrc2BIRsGnxdGa1THcvwBuUVpYqFCF
OabS3jSI/y6TNRZE9qrS6b+Ijv2LhEOxheGSHn3r4vASkimvyIop1M1Cw0Qg9O7kpMsC/OMbPrsQ
J5Kuc869kf+CO0poNO/jKDx7pfoa56BdjxlMp3gND6emvCLIL+C4xyZhWKJNEmT3oz2iPifU0Bph
i2PeIY2u69662+Ug/aE+QzUDm0hKXZJ5C9IAcm6ysJoLtImpwnhiTIsNYJLx5XBp+3DOBqvNiTOw
0iudlZ542mLscbEzfbHBRJxSC+jedZyMyCxfZDLp0cHUnWXlQfMTVzGWBW+Wsbh9ZSbq702BqFqv
DYAyxXevmN8t/5iCcwm1wSOU8AQ+HSpk+2KZ3F4V7zrQ3mRutcB0Ud0qfCqGUyethJX63W8Ku9Mk
Tt9e9BdDn03mB45K/hyFIQjx3Nz+BLZKqQ4I2f6D5n5917uZpmls15l/xIGHS8pCcVDehJwk6VW6
g16aalmC1TBIcQrv5N0vSd+54NmNgLoE3fyiUBjniRhWpCh76Al440ChCaal6F1Gw5GxoLsqHCdJ
Q75KSIKceZ/rIchT1HlNV9Q5q6Hh1yg4f750R9j88mJSwqMQKOTXGVOT2GFvCUkRIviziVEPiOZt
hEa47oQDBDPGmc4Ud4r9ncZkZP4z1TDJ6PGyngZzX5zf1x6T7IlRtjypI/7mAwry9tViiRJNIS9v
26XBbU9yNYmUUkELT7e2IlvrIjkiRnR/2v7rqvXbBTZpuQ2rJ80OsEgpPJJKoB9QX8BJ5wR5w9ts
bh1pMnGz5Fd4H36CE3aFXaJ75gjrHKIa953SSpTvoOIMeQqiH3HO5MHNEqyXpDKb/iPyE925ZFo9
BMUl8pCFMEebHFon9fNnwjx+YGz44XbVIjN8FwcJo2WkCg+PbIKTFkat4L3IS7j+7weVrEtqG3XO
E6cdsO8aPyANxlucsLGPYAnH5vqVaXc12G7xTHTtQypWr36NksprXjL4vaGIqr5xpZPbwTkqEIgC
Ql3G3mwNGb0vLKfND0NQr3VuQVGnOvoYXvEgoWjkeBgKiVop3n+9/XlVpEyC5RB79Aqn/JgJ7ju4
1JRZ8H488zurk/tITCnJ791McfnJT2GZDVw1ruhHMyc4m0lcCxJSS/LxgiTMa7tL/qEW8Mmda4z8
/X2P67CgvBGHFpL72Y71LAUh3wV7W6k/N8nHhI77YNHBC6CS3GsiyIkpaTyH9C4vrMGWrqSVYzu0
lH0yyok6apjcUkmfpd66IgRamNVd87xtorNR8kg8nMEwp1JrzYHWRvx1PPHBvLCy/wS/9tFxXPY6
ic2rf4BdpumSPicPcXJeXUaYY/sRZkrHCVHI+foDDBkHph89LqaFWz9Jimphvn8lG+juYd9h7LeO
2YRcnXSII4maEdvH/kSXG5h9+4MvU5xlYTeynEc+cCEjN3klguEOaEFiLvztkuJfm6O5wKFyXNZT
7Err8KePgXE5dxu7nqlUSHVTmTd81rbO17gb1XxLRqGUJSPiRGgfXBYkuyEFeIKJEFwjgO3pPq1e
C0XHfPkM54e6UloXjPrzZMzt6ilNRtrB1OaFJiCcKJk6wQ5ePj0pTrYv9j2fMbZvqCO5mW2Rfr9k
kOMOnbk9OqbU9tGTsNTIYoAM9T1wzOWAQegbI6DSVeZ84tp38dEwtxNB66uNo1/mMxdnnc0VImVS
v/D2Y+7ShEfl0JyP7CldDptVCDbg6zcdNjhDSBUfK33vpqO31/yGINzJvArQZF/1OEi9RKMxnirV
DSa++fC08gQ5usWCvQowGb8YLzKadB2MnSJNCP4sxCeRk/Np9I/Am1jfs2nOIM5WEdTz4o89kwOZ
9avIrCmeEGeovm6kewWQQxwoW2jflLF6264sWMRZkjRPCkRHr5P63PhhmFC+VaxrhYwcfL06PVHo
AWj4n7nre7ZHohg/0fNpa/22zoCbawugjt3OaAFNyWk6nuRkD9xQR4GBQ9VJa1dth08l5eg5cHn8
5eHS6YPTCbUyjKc9D5nnE9jMFzT9zVrfh/9GaGcluwyjzVes/e3Xqmjk/j87O0EwHRHGg67tCrcj
2NVYqhfBX5YO3S36Tdd6j3YCkeryDBsyZkF92QT/FYqY+9LJa+7VJ+Qd+BFvddkb6xcVr4X8fAe0
CMU3yo/MfMNQfj6GlYB7ehoYGmlpY9zaqDMjaRQPTxx/3IZglRwE7vPB76jl5QkCbNLtVZwKUq1v
kqbqRUgSRb4oHV5MIsQbla10Pt5shEtjTXwsOtw9+05X+qvcgZMCtTfeDsL/WqQPkdqWV6ryMN7N
SDgmXsvJV2lYtN3WBIgedf+xoutLivfSDib7XbkKwgHCikgUxgvPS8OJ/vyV3I4sq2T5P+l0/J4Y
AtzmxxFfZONHAcTxjlYe/SZTR51uQ870ydWJvTwZKczUIxgRsLJg/C5Zv6F1BrVE88SCTIcH4j0D
Eslz7odZOwHtG5A8fGDTAnKD/FGaV9AJhe9MVGLtt8L+JCfBHFj7EC+WxIW0sM1B4JZ76R44uegx
lG5OdAb5HUhxb/uzs/KlWT+iW/3yUUVGDAadviFdyxrDSw15m3RnHmDotRNwKkIO3QTSJIsivsgO
E13bogoZEjSC4Np7ZRwL6/3Tb9b/bE116sdV5hg73grIx9kIRebigAlNiQLkvCMen/KP5NC1na1A
4YyU+jf/w56sMVLgyuVO+NV84P1susymd42LDyQdUyIwaMxQyhWq4kXdXYia78+f7OGnggzT+vP3
H1s40HkPLaJju70bjNuonJX78OKTiKDf6Y12xJ7KU+nvQL7PTmkXVyy3DuwSg65C+gsWU6xhz+OI
uIorhtD8rFzuvIUS8MK7oIlyYa2fHgvvV1Dev/4uCqeeOkf2jWEV1V/ft9wyYzxlpKU37xdehLYa
uE5FXpm0uQLEIIjquZ3EiOl34Psj131rRr2u0xmuGyn2AivmLze0iUN5auzI5XC+bX3U0YF4+hdx
JZTMUYdyU8RMzhm8zjo1yfBccQFuD7txEaL7cStbbGHNDyPnz+sDGtG0q8pWUUK0Iuns46tMsUB2
nXlH6jruAiS+FpC0sxkWfWKV4g5US6pbunGfa7qLS7MBfr4JlyIUGLvstktohqvDrp8hoKr8jXTk
y0rAMDOhuUUyIJOeQr0CliLsAcSTyxsY32coor8GlJ84SVsb4ojhEqGvd7YBOloDJ7+WIGbFhIxB
WB5h5+ImhEdaHGXGNn2MHadC/OInKdIjRol4uNZWAq4Ckx55FAnQ/JridPGlJKYgrb0laWGxSRkG
etoo3pF9Opx4mtEwpkL/kKPxUF9dnhLpuLk9q5XsexD0vErfDIZ4DIF1W2faHGlttg55BWvEej02
x3+0dEK7uCC4NJW0ZxbIxHwo3noNPBOhzvbF2OmuUT2SI+GkL/rcYgqY+DxZRYQRNt0LOF0r8jcp
07Q7ZEbTNGVAJNj1d6NeVY5JYyf1++ThIiXHtD1O1kOWqTQPpgA1LXY8epklZTeuhyaxhjvTrXrx
HBAgPTYkffeiQd3YdaPFErM8UnRT5ctHU53jYvJvkVUN9NboMzm8DdjbARmT5LMQu2xOaaGYiGef
bOI0nT69bsT5mhex5WiKKuftoNA6U45Gg8XU+SGv7iedN/p+SmeFFGDVYlSZwZRn2ZDj+WYUHt8H
1kR9XZNRxatZ0WOwsbjwuMfe2tDeudTOFuwviQOKb+AGCgs+en7BdQIuzbsJmgCyLJ1qsQBtmrUa
g4ET9LNH9KyuXFKCvT4EUL3PWfqscp/3X0nWV6mK7vinfjIcOJh4W2YazBLA8EldiYt6s1meQsY4
zI3AN9At7q69G8bIxXox3wguZ/aG0lms0k++gIaeZbUY75BPppYxwGNFNafSih6SqLkBuzh5Txkd
dUfBJP1kJxa5NTUSs4nsiT2wBscGNn09kbas2O7s0axV4kAE88cVPVtn5+5hb2Wya6d5IXtSToGW
+WmYYln7OGKumpfHnYdaaDKZZV9FDpRkVyUyS3DfRn/BWenLHOLOYhvAIdMLS8X5aiKtt78XkJR8
ZGO4PJhU1E89RbwD1qIx8kXs9YJ0jCaQUV/7TCt2TKahzUMwvzRL7j9iE39225oQRzfrzIezyQQL
pQSNuB53MkYKFNf3lHjy6SNWckQtCq4nbYvf289qWmLF35WbQJ5xk0sBXe2ZAjf98jJddmSFRiZz
avr4nrn7timEJv20huG6OU3BbitS4zzElHOKVIAx9RXNmq93IumbHD6jz++2Qn0Wh7McL2Xl8mgl
a2XM8YwSK26SW/ibBjXp4s5pGIK0RLnr4ILLgOtVzoRhgM5WCtsGHjCvpwX8mITNha6gz6jNY9Jj
FptBVWVVx9O67Id9ZRSdvN/2eVHxxWn+6mRu2+EcCKT6c3ouQL9WJtgpJD1YLtKip+M0li/48DE/
1frAq1QQ6ZWnmm5OjVrYmCrUdMeDgGyy+7FVbb/YPtGP+0Vwk+i6Y5wHoU51cXcx7VWLdVmwGKQr
mBbWlcikPMfvloblSiofV/H8d3mK5RbxTD3zWWu2+Q35LAO9Gt+tdKYqzaheivTsAXUWX5n3OVsA
Mi1q6DlOuKHIV6W6Ps15gZhG4DRwgH6ILgH/3rqlmubDGVpBEoNgS4tNcAzmD4JZUzz3vWYdLz+u
ca95Y5gfu1Kk0Ix0EaVTMqZSMtaqaAhz/u4+2JwZW1AEvouQACjaVcf7++9vArh+4IhLsda3qBN8
mlcv/lMX/gdFkIldR91JQ5FAqDsJXs37CWaAg/jokzmyRYXVEaNvSNzgVYK/9Um58mhima57lz/H
VsaCxrLhBD6oZNEN22m9ZfzHBej/rVBQP4N2LHPQAC3OxcqM7MGG+vWVrNvMvAe0een8cmLdvlaq
hQKACQX13E9YGWAwYu/nOV8bXqUf/zylsuZSNNICnKkr/e1ZarlO8I0XnnEm2G1FPc70qLShhW9p
2Ji3oM5+zbeHIIvA46A2pDJtoft7+bXsclZIL0KJEeqLyiFCvBOTFbed8o7SsA3GMt6j6XhmSiVc
k5BP5cfwhmSGVUDvJWlW/Sk1KhKGIdEs8Gx0QsMEff01qHcOQUPEF+N/0A8+GRFaANUvwVb4OpAO
asPBTeploYa0MUT6feJJrQDagCsdReUHs/5yWgfAdFr5o6/llqZza3TYnYucLtzpoNIHL5+qrAVe
dr2CEUsD3SwdFXM6M7onANLy0PnC0Eb7RfTtzhrJypg6RseFxmGJ0h5mV3e5lRMOMbuUZnSF34U+
qU5Wy8M+QmHuy07wKYG+YJQrGMBbObYL+V8JQGh2w7xFrizD/o0KsCOJkEfTO/A5NzJxU/AALOEu
qDSUwG5AI0ZcDnq8A7gdh5eBeEemOI4HGjge+r4vDhYWo5WmWCkDMDnS250jC1D5G2oVgTwwaPMp
UcH3eAE8ov3f8vmHbKt7/mwMJmx07Rc7QHhnq8kQje+jSZnwKTKhNB4EPd2LGazneH5lzrBI46T8
VS1pXwq89YZiI3C9H9UzCEGvQ9RYed0E7tL8dSyDslXG3yuhU2cB1MWdkpRKL5CEyamN3ypIc8gn
IZZZCHvtjABW2IrAKh6C8pKxiP0PlKDQm+Ev3V/PWkV5utOtYddFB3s0E5ybD0BmukZHR+X+sL4Q
loZrtEe+z0pAaJmskl2WnK+flGKoLy6/XSzsOjap3CANuNFgm80YohXZ05fGOL8iQs/m+fYq5ZnR
BV0dAc6cKckCQ1PIyVYk+squ3rLH2zGb6j6B7j6oMV/5Yy7BinnUoMSlY05HNj8HqJ8DQ55J77zC
fL5dOasld6EQTyNktNafgaHZaiWLVPN1jSKBHxSnBaY8A6BsAxXiZFP++Xm8CgukOO9GiRDP5fq1
jxojB+Wxtd0n8VJT2ZVdqmKl+UfKOQkINbg3CBC3LFH46z0dfPJL/UDE23OGKRo+8qUhWFJhiGea
sk2EZHeIJA7MbXN1wLLkv1T3Ah+p0nVhC6VQ9RKd8QxgIRh4j6BqVMFAw66L5hRA629OpIIz5mSJ
ceJo5QPBVFk6nl5yGbqIb0XErkGjSU/NOaWog7AOZN1mNmNqNw38pnI9dQhIzfttkS5VS7gQO/ds
8mcRHtFSj0vPUSdws5u7t5+Wl6yZl4HuSeJfdd9l+zWYAEnRK33x/6hHw7Fh5OfOz+Kn3bT+xAy7
DPYV6VwRYjulRnzWxy/XnAmrTAhMV0Ps0JdW5qkGl+RN9k+7B1Dc4vhdTgsWU8jaA6Px3BEch4Sa
abbj8KgsyGiESuInzxTJVnt3+pm//AUrMfuhICWqzxl1eCiDdDAzia85X6Gqs49Tp1xE5WtEisLC
tww2xBkVZbq7/GLLIowRFzjvd/Fhzc6xqzrhn1d2SZO8hMkjLSae5GstilukLnaxQJk+s3aldV0+
j6RJP3P2Y8nZx4j2BfVXISCntGuDp65sC9ati6e/GuxoZZjh51Zb4iaoMNomvv93UBZPbF8k1gfc
gt5DvbikjkvouvCWrxqc4bJ1E+uYqc5QjuM1uE+RzX7oqSz2mvck6Y1AbiEtiCJ15u0GSAkHYY1D
OSEpylwy7wBgfqbks8hyt0hQ95saFg5ZrSyeCLhjpml4ZpMok83jBimNfIi+qjuIyZBueOSyeoR0
A3ARB1RcoGdjchbLRgXRdhf+9CwYb6Lt0wc9bNovGJfxu6GteLfG2JtNcWoj2NGnuDKAb0PxAH9X
1pW/M7TszzXcRm8gC3ExXIK8OIXXcAj7CwLlSh0MSyeLIPfwyncVNL73bhA3xDGK5qc0gmhmlwM1
M11GqKTxepDQuzLNxHX9UlOHWuhJ3+62GlmlNArA3Wd0Y5kLf7yHHuJNraJJePjkJB22a7EXwB7v
3x7tQqhLrA7KlDMoPTG6/mEWlq3/YE56X30nXUi601UFVZzquIdWmedR48Hxg+r6hOMdAZ5TiBSs
NJynNQdKBoeeRKKMbGLSS8v42D0WCtwx1F6MayuBMAOYZK45PhHf5W/nWeVTFpSOMGV95eqsfLO8
PxvEptCxOjS27UkvUw9guHC2YMjdzhslJ51CGWAffY6II0dxI/hobhGGXgLnhBMAdAwj/PTodvX3
CDPH0sXe6QYJSmWqArviOY7k5UV9c+WmirKypMGwjgbvWhuCP5+Rk5Gh64/kgHDVo9i2jcdoAulF
aIjioVgPt8fz6yBOVSlwn3kTMtpE8ewQMEhWWiiLRdpxpRnbFWYxC2XUP8oRSyYn0Rvg6MHmmnr4
1flu+09M0qPd3rewjUc9jQoIB95tDhfQWYeUG5Fhfc78/RQj0YER2Z4NTpccNGpfN0dxMHCl26Ca
l/pJfUYYDQkfteTc732d3tXqXHUSG8rIsSpo9e+WoSicCCcemXPpX8OUUuu1DMzKAt/TeI5uV8dy
lZhYNOGDS17kKdNkYvvMvUpnzS3hjTvo/a3j5fA/Na9a+aMcggKe4YCF+UEA2FqYljkcZsa+dMUs
dEBI+T3hvzYAaeVdFL+FlzhQTq9k6+JVQaTki6wMEIKddhWb0OpgIG7MU2tcUxKAm8SyNwY5CiRd
Lx8r4gz5ZBiw1q0czyjiwlJp6l6MjXVlCtsd9Lq2c09cC4DsIbzR2lWzQZXXLku4GY8X7uDJmeED
i+DQ1tyrEQESeH/a5fbE75acwob5uKtA5ouCvis9lh/sXhk80FNpGg0MixnkWwg8algjO8C7tVf1
hl9dTClFvg59rooigH8mpjPrCfLa3PuyO4u1EHj4TIgTvgtloUTfMzhgtlDY4X6H6/RnHUy1HqWM
dnzNZxVnOVL69J4iYFHF2fYTD+UlT0+l9mQvJY6lS/0KFKNGuXEPJrhSh1v21piewa079nrd2L9S
aseU2wZdxlAlaLa6K14k6N6VrJGOla6QaGCZgYd3ggoNnL39x9+2s/JrGiguyq99XyUiz6d0mNIM
eCf17a9KA8J9EzSrIAcS4o0t4tgkE95A7AGfEmwd6H4hLJezCbcMrieoBypM8w9XSWUuw02Pv1hT
k4t0989O5Z+KV6+iuOqXGFRxUZxBVISA4SGAl3BqvjxP5L9ypJ/jcK6p8RUUZ3PrHMBJ4bkkEbh0
JRhVWjs9ENTmvduJ2invEAXC3C35ciUkMaGAXbh5+eKTKEBV8doNGFnfAjw/JjlICU8tqEfA+nh5
wUcocmoMbzf85rEB9+WM57JTXBQGqFzlFXNI1bhxbsxtH3fJqtz3oKllMj9Mpv9Ma7wz244g1kDK
x+8TD2JNpwieiCKC7vKg+MzXA6z+5Z6cgj7gZcKUmJZRIzPr/wzg4hoZeblNnRER3qb0xRZeFN5l
CXDs0JE6GIyBWxZpOnIODi/c+YZv+3MXsNVvV8tVe/9w7uXRqpPUgbnpjDlM9YjP3QGciJZfc2ht
WiNemWPCkvUoVHYzSiTwl/zQVfE2SQLDPGZMaykMxCl3Vz2X+ZN8h7iVWNtV3rKP8xvktoZKmvB9
cE8Pr6rYo4Qv8qLlNyPKZJsSJEFjy7OW83Xf5XucEfsE49t98GN0zCCSEnxfXyzX121tXRyGSret
pA7l/88y/ctmY9bEjSQGWM+laP8cj7YK3WFYwyMjm56sVtjaJBWA9JTxsXI61DEeQFfJySKzbMqU
Ri77tAFpT4Gvyt7qLTgtDrDYSBSbv76ibkmkfuDWCeQDNENntKHqZ8s1l468e/XkCiA4ex5+AkBI
Ng6jrGbNowu7kBgItgnuatvV8I9QR/XlMrHCYlp5ufvypZRIGPx/ZdUWIwAYaxoKi/bBPldPf7ws
1dC1gepXHgDfLDXj0NfYTCeeMpzs3wVNE9+6zz7o0ftEOtmFSmCvQ/6wa3OY/DNygtghiaPvu0ei
k61bMlcDuEhOUqMJOW9SAiyq2F+kFefAIHVtK6SRnp/1F8V/ImOAmy/4X+RzninwK521NUxqrtiO
R0ygEOnkwZGAnflr/bzPWoxMvt6iJYVLXcvsC3RSX4977kHTHwK2bKEGBC4iB4yy92TjeNIqlEin
Qvm9TtKiSQy0dsEH47SJM2MojfSl77yFhi6DKRH4OMOGOrtcfyIMh9zBXh9+fSajNX+OTrHxs//q
F7vfE40610oTsb5gBgObcMoiX5QxeH9f7CAVLDo72GSiAUZ9fBVRaNyx8mDFkDs7TiVW1lDgcVtq
IJLfJFYfWQt7/6VeV6yA7yo3Y9Rp7kW9zADjptHnjZHMJg8yPyYJuueZCjPnHSo8Jf2jDHdDvut2
OGEtxUfN4Ypvo5p8Fl+GGXRp7t32RccsFJECnchqlAfr/f6QnfY+zT5/brWNAgz0mZo0OaeYZDzI
UhI8juXKrVkc2/b3QfuVzLr5w5C4sidECHEDiqECw8XIiDX+f1ryKLd9QUcCutb02XeIvuIlBffJ
z/aaKqp6oGMk6M9KMhx8HOEXMW0ivWulQvhR30V4jNIPchU77NnyZkIWtROIiy4B+aQ2BArzadks
MvOAtrfgoY8KZmgm/11aEhOWv0M++J4OCFpffiXbARMg/FRTatt6eejWbpPfALxcJqdx0yRxXF0o
ww08AOAyHKZfR6WW6YWSRZFix4LqJRKTREBwQTE2C3etOxgHsVmZJsXe/obW3AGRc942Ba1At+OX
v7CMON9JgvGtRIZMNExw1682EVdbqSpp5Rt5xgM7nxYr8n1v8uYmYr9Ozf0bR8/SxLwG6F/Jc4qD
qXN0u/ASQA+eiyThTwGjujitJsieb1nYynjmI2iPr7AV+1VgHr5uSzNJcSi7qJ+zkBLx7BJAjJCj
i0RpvWIw1o5RmgwaztxchVow2FBw/+JhBnEt2scGaTaZ/JUCAF5HwG9e6lhbj9klOBHWZLcvauQG
HmHL+QwyHojWM5h6U6QfDBLws9bVyr4fKPAl4tScIqWLhpAoLdWvJutqvr2Djktn9IWbD6wYSy49
o9X34N4CaFtM0Q0K8MlQam86AIWRjv96+2cML/jxmFs3ywMjDjX4v010ExsfmBcBZXXyUN/b6OTO
FavumJO1g4u0UXBPheYhMtC79ftKGxN6ZGRpCp4WHv7728Ty/9Mul43n4TxW/6zXMKoHi19v9g76
EYFFtL6JdtzUOIxkEfQfVJUSruMaTZ/xAi5gXduO8WT9if4uP+eBcNg96RhzcFTZQbOF0rbiwrVp
PUJ3jjXQilkjOhRUQQIc+XQUwomJ4+w7tNtMMuoInvtqnr9wuPZNAGvRf4fCwd8cfEQb6sbips4y
3QYU9NsssyLPsMPYeO1C+LXrhewN6jD31J80mqpfrqJCAmmgFaM23ZSRuCAbbFOwefBjZSCdBwIj
/8A1kZMmhzrKyzoo8eqEkHAljlQ9kEVEFtpwYBFEIvhxwxIUGVFDuGoL7KAsBGels0uvNz/9g/p5
UIkQt5AAH/djcGk5J+SuPYk4Lc4kn5CiU10YZ1Kx48d0raP8Yrzgk3+QxVgNJn5mdGoxu1gCkoux
izntUiuhf0ni3pZ1BNc5L5Jiy/0+++ar/dDF0fz6OVi4xQY2NGD/YL0xHeGPj6ymC//V2WCGewrK
Q55Wql1IIGA+nLBDVQ5hfXJ1Y4JqnINbBOUk1MEpVFQIBPcV2wc9aipquQUnmapJ3JB+FpDyR58D
Z+T9Xbgzb3jLTPmpzrNLSBenOpBY0B/4xnAhwhl4MmeMKuch1O0gnZnthqiIABCacytA7jlJCgT0
tr9gfJDlWZNvhvnhdQDd2UO2WQC8e2rkbmB+JEyOetQHxi8/omImLrbXkBqMI2Ari83L+Nfjx9KK
60by8XB7d7GDxdkhW52+wVaP+lRXV1YlXuoI41olAqCeYhV5qREVH1prLRgrTaDKmNbrLi4IDHeB
ibrt3mdtBACQNIVTnO5Ec5XrtqthVUwXdNUl9RvXp7w4+cfm9G44T6ce0XstxaIE6o3onJf9Tlu+
MRwY2z7uwi2yk/XyehYsA1y7wdb5DxlaU8h8ZHFeOHa8PWFmg3yXgZNxjIESh7Gk2ITSQQkQOZhL
5nRBWulYSne2jhHIxhpMscp8zUzvIS88bJsRHvt45OWnB9h6/FE0ov2KxBaYmH7kpgbTCgpzto/7
2getlPF1Y2teCEXROGm2yjj1Dk7fMDdhc+I0y+hftNVLCIbyUEl4VVc9qrFGfvFx7j2Vv30IDnZ0
31w8T4ZL99ID0kuk2iDo5PfR0pi5NWUgNKe6CJzYMzRTyu3xk+H8NutP6H73FC7AR6FDGtoncYm9
SkUt4qEXvJKO+477VfYFDmml8DEK2SgsLoR2VnXqEuXc+XLjKrk3kNMUqLmwuBkWFJtapzJecmmR
8LaRrE+NqpdxRJ6xI1zq321gXCDuft4KBrtYaZNDTqnJoN2zDzCU7maKJlDBQ5c2J+4c4n+jfcdf
KWX++d/gVvppjFHmE83lVngDH000t+7jmn19YEN9pLo91Cayi3k3fA3BalSeCJCh3vrvMyRYwj0q
pvG0SRlDabw/FlriNNBMgk+3JnBPDioWr5CWKO1FK41Qlo76MdO9tFBwp6lZg9mcGexcm/N2OMVY
pVvQ01BJy0kUBCf8LPpGQn8Mt7b1zzAylfq91j2AjmW8SuwEStvU8UsMkW+Fbn7/PCYhyRz1+GVm
0BXRK5txB9A2xzAIpiuJaR1DBsLqWQQbTPg58EEV9J4CUGmJ9tf2aZTfsWUsgj0dQ5PPYynMRqBt
9k6tmGB00Hpvq+uQkZ5E8/j+1lLavovay1O8DQrMzGODLrH6w94VgnOsuDcP7XCvc13KY5eNBt2b
RAFS2JiYalgW37ekHwwsqbYlsJCLOf0IRx6u2FzD5wYp6UTwZUi30gZxRmuMFK/616topjWPTY5Y
N52YLqkbp1i0K59cKK/TlP/fpeFMSOsQMDBlDpw4lXz1aDvBLnnk/tf2kU8gS5EHugNB8otU79Uu
RKZ8tu8B1PzNWhMEN5qxLykR03bC/+dbJBUp4UpxsdSU3CX0e3CrpjhDcPIFJd17mYxJFLMCxohH
uwzkFCFi0h6VCURHJTDQpBI/8Xxwxd9XvRtq/gB2lvT5pqzByKB1N0s5vDjaPVceT0+8omC6JhcF
UcK5gT4N1frxxtUDqPT5brraf2I5eY852gLJFGX1MZMKeomVXLtPYrDUAUbXY/bv1D5p9xT6xEdx
XjybxX0oji/jqoTyPg1iyeaBuuaRZoN8381SmhyZgpI4z9UvOpS5Tuz+z+dmfnj5cDm3emachs26
NUbPZBtTBnVPlJPJbVsdYSTSpA4zJITGKQPU9NZOxsjqP+a3YJWg+4dhnvzKs1UzrOrsx4qc8mQo
POIcsK/5ljEk7phD7TlOfo2L9S8Pr1Rqh2FmHcMQbpkFITL3ki3J2DDcHhrTsDISQlzMAbM+hhVB
D0bgKhWg1d7Ue+uP18WUxDtvtlgvrT7lhGwpcXXkvHVuwUj6LHFwglZB1mEmfmAL4B1CxG+jUtGa
G4CLA92Sld5i5FjUReJT4JVWCbFn0ufIy44RPX+RUvYQ2c4KnFmk2Wfzn1c4NiNm7umyuMsTSH7q
LN3T1otZofL/ZbAaDFUckkQTPm9aUVqMmRjFajoILEKUQGlp0jFNJePHiPUkYIyRnPwOgQLUQW20
eopHCMqvafeS31dz3UbJ+wMo9Eo841A3JCgchFcSTrnCVTexPlRPIMMpQeGC8jRFUUmXm8R/Ft6R
9MZgC6pdAyWhUYKIhttHUYczQVA9ry5gS2v1QXcTqKnen9zOwyru4GO9pau30/1mzlp/ePw4jiFK
62/cpgK7bAbWXTUr85IUTnPWkDO+Y7YLL+HpaQfqy2lcum2HxhYhBOkThOFzTJodU8Jpk216aM5a
zQ2QIOM7vQkQ1oU0k5v5K/wy8KLQ4+1YKP8k726pvODelpTHMc5jVIhs7Rse7u4KxayDGMSVc8zz
6K8J5uq2gam/hzVcTYGBNHZ4LetMUJmw2A8tqbJdjJlYgpZDEJxc04Sjk53qbK7nJ/8P27GTTDjc
hr9VQ2xXf2L6h5dTh/D7Ofrl4H95uayvqYU9VESC+xuej5Yo9VCfSl9z0jaQ6AWaKXWz48brX9KD
geQq0hH9/3l+Dwry7kJn8/BKMdWBNZrsl7uta5CjqQturHVuon7NkY52eZwA/UctxQNgm2TnNtHp
91/C6xPV2mUE+k7YM0gYqX2TJ/2pxAv81WyZcN//O8IiWXyG5mdgg5UogIRDYJwWjIx7x8dYT3lQ
3euC3pFCmkma+E473UqKZrpXnk+eFMgIayazF9OWF26MurG6VtkywKmgLqmEDr7UUIs31N0Ike7d
sgOpG8h1dxwIskNenvQo9aJuCZusxLgQtesKuPCd4SGh7ZQnYdz0jVdWyMdzjgzjM6LKSXV5Jfw8
MuLvBBJAVpmrB9U+cjRP3OgCKx4xwoV/07ZtEQyb9bQLx2V8I+5nK+DvKN97LpBrmGjjJDmG0USA
yHaqTHQ4NkrrfGLmlSZIsKspdChe5aOkYFVLmoNM7nnfyD3CZTF3Sdpk65ZKFFEOmDGAtmbTr8UI
Q2CA/dpkoaMeZC18ptXdFDqg2gKT1ZRjjb0mjXqUefBOoNb19Rou4au/zqITdCj1YneHV7izaK7n
1cK/lVrKrQX1hT2Lo9pJF+3dtUodYcN0uTtA+C8jS1kt2z3mHkIb8RF6OV37nBS6hew6ybeCx+lA
M4VvUD7zWeg3sZd3LaID4Bsi23m347/GVZyG5/lmE8EAKVaNOXWbBxy+plzhIm8kayUChcWqU47+
GhGnlwdM73pblxuu2qBHVU2R78sz/xa70f3MYNI6Xz8qhoPOmcgE8uz1/fXoltTK/Hqsv2GbHxnJ
5GUwRSIP3GSDtjNAhLiAarZSJuPIr4/hfof67z54eFoajcQHDwqZ/wLyV1UFs/RSYThx3SHmdIqw
Sxn8+1V9NWTDPY0aFzIlmUKt9nZSGT+goXFlFBQE3kRmTjKtF8ED3XuYUDkNlwDJYMKD/noPmKNB
iezimudMUqJkNAJH2qza+vmXuSHpy5kn7BdBi1EUg1aEQiJtTs+rU5iI4FUIT6zgdzDdrOt2DU6n
l0LMJ/xwLwg81cAyLdEP2GsL564zzR+gDgRKaPrDp4k4LOpBfOxFVirDMrIgTRZ38hBszIdKj3fG
Kzg9VOOMg3509yLCyLWjQxtGAH8vgn9oIcYLU5/RBijw37HY2VK9UX3P/zHapxIuViVq4mL7od63
MumG65jZYo6uWrUfoyLGWgqdK7A3pMBjUT2RsoJgyY3TQOrRoqobBTmnsDyKqwUj4jykTela5WVo
ou7nRjZD7/dgW648+JNrmjYxNVyyU+8mtbSYbIVqZ1piHs7z2vT+kJUBBKU94sb3qWwuQ6WFzHKW
NubUc31rqnwKuHw1iUtx1Dpqb1xm4JoIJMNO1fgOY0xogegTOto54dBtoOiLm5/11pCNjh4nTYDJ
NJqKeGEfYbK1Cy2gXOQrFhESV6p/as430vx4Hw6tOLkEp2QNeomFP1zm0JM4MZtJ7HXK4WZolTcB
kTH1l/Kc0OmuXfbBlDKAlPgNQw3hwT41eqvsy4QFOfwO3FPZh4ZnncIYevqZro70FYy6jVaKLepP
sV4g1wfI7b3bwjq5V9yhZFekOC8nqLtVAD3tFGFuscz/evVVARx6rxI+eHMp7XjDe27D+qMrjibs
hXYX+2PB+yIYqqho2ynnnP2pHRungKHdyvP7V7XUIuIIAfop1wQ94e+GytpmtAmZSsBT4nUgYaNl
Ut1auZrdwIoegIDrg6bphPqcrtUunADSGpqGKwJDvb7XrzlwZpI8O71qAQdF6YoLtl/ODe7VF1q6
8gC6CjqyV+Ps5Hl0snHLkh9vBTySnta8fpLkgTUihS0L15Kp+YdEuHGF0Hx7T3sPwpSDuGkA7SHn
/m6bf0A3uShCpn5rTSC7C6tJjBU79WNnv2jfj1xLBg3eWcfYVQQkbE1riiQDFHWiPxZUt9Qt9FXv
lCyyASp8pO98nDEFufAs0HHl+WNg+sXa1VQfik3eOJ8bZhAwKVUSKkeiCe4lA4h2C0jMsGruOW5n
Q6i3XaOyO/24sDb0OSYImZi5pS2yETWjrgtLvgoZ+WWL0O/FF8nNpWAJSWU0/LU0ffB04P5K5bsx
Dq40R7KcyaVCnICxKwNU4JKKKtg/BQVA9bUl2KzcCR+VfebyMPrm/0KuJpxYblYjR3N/+BKcr32N
DegFZ3Y1D+p3C/y4YlK5l+PEc3ZjjVpSv6/iqSUZOKA3hBGEfJgwsov9RL4df1YH0AapZa1r/k/M
cQ5JhHhlNV0lZ+9ICI08rxUYUxFYEsMvEgriyGbBsLatIhgJ/t5bv7rE24Jx+tPJ/yjMhUPNDX6M
gzRvEJJbcKdviaHTiUkflTWu7HF3F38DFdHbJ+PqMkb1aa79Bnz0FBHBqHd174V5U1L26K3RkqyA
UYocQIe0WjYzN+c5YsFXN+wSsxzafDJAbj3qgIZwZSbstYcKaX1qhH7VCaKpmdsiOWAp5Fy+Quup
t9ybYyfOq33tsI+uAyubysyQbC4s3IRnpt0cjJ/UquCy3SyspD+U1weKdUgSPGTwxEpOvpW0S9ur
Aw6kIHN+wx8W1Y8gCRwZXOmT4By3CcYuQa8RFoR+8Kg4if8XE/Xztb4W6SOmAA21dqCAidO/1154
/ZfcIncf53k1ofk8jwdXeHGA9CX10Ny6b856HL5ffzfTb6moidL2XVkcvmsWcLvCgcU5iCRK3h4h
IqS6sDqMa0Bg31GMIMXOloJE3YgvE6O7P1R3P1k013ax8wzMY8DakzHs/YLkZBIlKbHEvoAkHW6V
hZ02VXpdGoPj4liVGad6Uz0OWrV/xpd9OJBbkz+CGmA2EDsz+R1ZLSop6Il1figBveezuIUVmQKg
zyqHlSdRt12A0HLcGBQlbHg+VMDhTD94rQBNCEzdxdk6b1HTgnDC65oFDTPUF8wJYpG50fZriBqg
x+YAPDB0l+avGlqRltBYE7CzxulWqyt6ntcNUDsp7rHKfNmZ+OTrXi1Bvhqv0dU0QhlsRh0iX/ZW
yh/uGWbO1LMs1PLOo0AD0W2Mor9/aX7L2wtPn2fctaeQ5YMBBNnHKecdDDoq9umYv4moTJajKkv3
YYKnx6tlR4/W3FPi7AQubv3PtnOQeNDxai9tZM3pzHdCKyNvdFgv3O5Xc1qH/Z0DzO1kUFY7i5P2
9IzJ8XLhqp/Wz0cbuNR5KlYSIJKL033KKoXKYsnoSx6F77/155ZbrKwVuHDqEtis0e7z9d0tT2cA
E7EEL6mnMm3qS1w6kIq0gpcpgY+BeQx19LNjRp8tzTB1oMMPUlFAyUBKNfK53xo7GbBK1CxI/NLd
IeN2ltX4uf20krsJw1QzkPaKFbnjYl1rCqmbdFB2BLKf4D2qBYQIHPPn1CERIhKI+7eNy16/8/IT
Xenc+KYv9Mqggr2qlU+YExGEPZFNxgIezBz7TxOoYtybWq7nQNTqORulGRGfjURjFDbKOeKUq8UC
vavSOpmKZrMZQC3Pro/N24wk7hy/iRH8wuYQn2FmoEopNxnAxbHRctzmSj9sQzjKkWON5dNzCXKx
7cHJu/68ybBO6e/sIu61Rid1/3YoQgd7PyG6hBAkm2/wjCzdaWWzU/qjHJkI7ywxqWk4JeLYLOe8
gB1MlpVKVFD7mfiLhWhOW8q0AXGCMDqYAcFJQcR+zlO7HQvNy1ibdOB7wHe3TmTjxla4QPJzHNq2
YX1spMr3zVSwg94PQt1hWc/vY52KBGPPrz/hnQYNthJesFj7+9qsAjV7SZ7STDGAr28zAuZYL0bF
fOyaLMN2GcT5ZSBHdoe2WXVvUk0CQs+UFwRX9uvOP1zlOnPc/3PtVjYahWajYnD8zARPMaacpiCo
YqW2Vb7t7f5JCoGT0pjPrc5IMeBHxXaeNO5ZSEF2AfqyCe9x2YgHcPbI8KWbLNpzUYxS8sHqG6iF
lnZLFzbxTpubmHXnz40W+rElcz1+eFFr47oQaLMx8/6nhUzDgxi/AiYlfvs0fsJJ7W+NqxBIG1Mr
8jVtT/CaJCRJUzqmJ6qpHGOVrqQHPwWbeI7lgTLnsZvr7wBJCZPKqowYMD2eHoBaW1M+7dRAElFx
h8uZzvLD5bWFcFmArwaTHOI3vcRPE1LFl0cRkqV2Kl/HX8rLTL6pPD2o9Dpyh5GY5rqdE+Pr5lC/
v4NmmWajFL9n7rUyuGW5YhIgKG29aZfCYBWVIkLUiwTWj4HbtFLqJcM1we/cYuglhzGeMQRc/YmR
ughXis8A4un2np41wXaYkAWN4naTEHIggm9H2vDWEFRXXnjbLxl2k5JnlOGufLEG78H3Iocu8+Ws
QNIzH0u6UbDXhfhIGSip6EMDk7+1lQF/fTGk+dpmsWO4KH6+a1N6KFuM9AXs2DGyfEW6hoXTtHWt
sqEdpZAVqcSM/UhVT0Q0n61ogP2bCll57mONChBIhUfdeVoT2Q0gc0icj1eNFPCjPs+4ADbXYK3B
Gx/81AUm96eY99uekjLZDrzCAT1BaBWFRO0mXEo+h6WV+vQYKcGn+Q0OPhdthLDoJ4RGkBff5JiS
k13k0GygjsrVbyFsFy1H9nyHRYxPa1r/uULSbuXQSuu0jZ970uJMMpaxgRCOjTidjXHR17s+Pfh+
DAWtyOzgcQm/H1JBb3CFz28xscvI500VeqZWEePmeokaiE+4g93RPWN/CzstP5XPCAECzjueS6A6
IdpHnt84YFloGFbjR8jf0dOKPa8WiKj1Ys76dRFZ9ME4eIRJaIddGc8BeduyGCod8kgQa1tQlAme
36Za4GzBFW8Qso3zvU4d6roQUl4QPA+mVdSuIZO+dlyAS92UJHJVEfzPGyBa2G9xKoTCQX1IFZMT
mAy/SUteVGU46lqjoVdMjbv+A96wEnK5i6Kmx+cKEtWTgk0A1GPC96J5kQcOPutVxYtIVpTZLXjB
5HvSuPj6hFdsjRyC8mUtyGEOsFtlNSDGPRESxzTrEJHTbVpclvrTh2evvgmvTRzKjulcX7Ohr9aC
ff1aKxk3MCNoKQgjefo0ARzICkkuO4mey0rDUXjdUJCg33cPWquNrUTjhDZKj/tCPnfa0CAaDrl0
kUc0bveU4gZd6dvvNaFj0qRre5tLHmRrZaePffPkWXkhgK42srvHnG2IvIiuMNZNlKr6P6yPcKrH
G8SJkJ0lAREBsAwPGxWCksLXPyE4ONU+193HDkZT+/DJtq5sNrcwyJTL9tgA0qoIYdjgA4c79Xyu
lYXvXV6fDgBHm84OFs2TSEzekRELlBHp5FQtl3F2iNiZ8BcfwZXm3m32NR4zdJw5YBRxPAFfOFeJ
Y/nj6uuc3o+vJ9Bg9PD7PZEjxCFs2BMu8xRjy/2BfJ2LzZ5R2KjrskgcRUbeKhNupmJZOaELoOVP
g9dGMGuk5Y/LPCjMd8lGhB/WnVbD5Zc8O3mHVemo0bd7Japqj9s4lCT+mo0f5M1tROcp1ouUq/yJ
WSco7Mjf71sdalhoAfYy/NDDlHPGrgfoJfxQ8WJvhwaPTGLXijLRTblk03HsEKAT90frRxBKiNYG
Rkuxhb7rcli0ITG2+JDkwltJM7orqwkqfMEiQ08M9sCR1jM0OrwzN6pfT9yUQ/7E4uyRlJYLff31
ntuVjSI8C8RD8XkSt1EMf19QGO1fIKhT446czYGx0GLivh4bVGVkKdlH+gDlZfjRdgAbM6Gc8/iI
nvfgBDB2CI+XH5KPp15w3Btl2I0apeLdTUq6GZ5unlvYyDuolNnwx6GkNo3R5HZnDuQEUPKLbXtd
s/8IBxZshO90+36l36s7r/l5gTGhuDTqjkFooSPs+LXiRmRu8u9AIs0jGIyoB39LgUW4HcZ/dBPu
2MtTaKSEjcEMbL2VGEmxKliXUr+6A43SO4eDnpUSOEMqQW95OqT/9QCEOzdtuG8BtBGxfPbcXF2N
RFkFm4dBYkTfmZ+t+IfKAMIdhrFXFaESyi74D4rXoO7GWC2AHK2YFhA+GNVxeo82OpRJB5Vw37Y8
IZ0mhfEZvl0ywDDfKsnoqetBXXvxtK4br6ff4nJuNos73obFY9ys+LGrcF77HfwiujsQ/VKtY9+z
B8L8Fkyv1ycB6S4UkBMSRFgDRPny+gPzz35U07MfxPrzFpvDoCgFzIChkY6e8b8YAwF+tE5P2P5Q
j4ZBgZpATQsCvpSmTHH7lsI4L5Xi/Qzm36XO4h7ADA18XsqdJ82eCg/DWk/VhX83V97KscdwZULc
eDzG19hEracWoB2OgtuEVnJrXoyGOr6KTA0aapII7tQU1s/h7nFFohYRAcvDVG/36J3a8JOrC62H
f5kMplnIG46q440NiM1jerI7/55z5oOiew+NKdvqTMe5vqt2qX6KsAu0bkdu3XWhySQiU4ndqyeD
fjRKa2hOWgndSiqjKtZQOrGkWRs4UtcUX46Qe2/+aeGcsRQr/r+oFC12wL86WJW4Bpvk+Kl+ccWK
88qcmyWYZwJPgUIxuPOXK77gqtciIOUAsuCITjLq41WenvnL0meTunlqNobiya7I/nI8/Iz2tpy3
VEr+NHydCEnUf5jP/GfBDRIQCWcU9Su/TwD49XiBe5P3F4H8QIaSJZIcFvixhzfR9YpnX9JLd1X6
CCNYUAXrDtpjrVaHpomrguyxbsooEOPDaEZAF6ITY+GssCMtjG+Ca7MKPZ7CbxNOdrte+B0GayRR
s54NKRDDPx3w9Ic0qyU6gCQKg5qiqO9ZMNFcWIoN/ii+Yx31ESW2/Xu7MSsKMeZpRebs+TjSpblL
+GufF1RVlOpItFWZgO3Pa634ERtItBWUgxJQ97EUHsbPZHk6495dfouxhGprxZRBVPGuIRADdy0R
zuUtB+gS6BKTmo8A1kVu9A+St+4Sth5bNsfhOpGvktHzXQOVNbNfNaRQi6hliJSwafslo4fjvT5l
QiRGdbReysxhQqmuJnMPznbAVjSlWbAyI8FawVp5Xot+1QH1jvc3HsVo5ADSVyCqticn6J4nAajd
MIk8yrvwxT4RJeOFPwbwx2D50VJSybVYIuwheuepmaqZdU03G89QRwYv9FzsowLxLWKOKj1A1w6w
c9gpBXPiPix+vTNd41N7asVHY3IC3YbJYfTECz/A4VOZ7q/kQgj3n2TFWnrU0W0CD+daf1mQ/8pX
etLoj9M/y8MEJakUjsqF5KTU8Gqnr0rnIDKyVxn+/K8vPMKpFu4is5zCw/60Ljwo7IZ1qKcJo0V6
w6HDvwk8l/txk3OtXUFArorhsFRBeo4egJdJxpqLgPQ7NwtwnJtesumt2xDiyCy7hpj0mBeWxLyG
YuCP6nz44yS5F7BgwGQeVEzQNSmwstSmtwEhWdGCH62jUsskjgWYkyvPVOcDJGipT+bw0pSjbzEn
hld/B3nX9kMePue9OCgk8TFE6PL/NyR/x9SeEcvmpVNUiEjc9puB77svbAaRgquP2R7IePx6yC2M
264rastAMlqV+QdjCvyiZ8FztmGYwvK9muzSOpi1rG+oz0Ru+IEv6pKmknkDjB4sVO5LXi98pY7c
G1YVSqMy5Nv+nCUMSSfxdFeB+8HNBbNBKJtYr/PeUqPvW0ENwOizHelTbjcZeXRJoI8cS0emdq94
xA7t86WJX/Q/o31+WTm3bEkLPLUKpTgCm1zUrt/RfkycksTm2Weyo3f4YG+hsuSJH/bYim6yvzBe
mBWNuvp/HSixBAvSZRp6Q0KXwb4YCgQvJozRfUgoIkfSS6WW3SDot3Sw3UIYY7NvS55ezWcDxPQa
mYG7Pd4hgJVAq9xBqcO+1L4U1gs360G96zBzll73/vFy1FKr0oug2E1uN2aqVkNquT3gXDwayqsk
17cOMNGfEl0dklH3zXAhU0jjitt8hwQSLyKSxkcpTkUM4NPBW5ijAG6RNR99RgR++Qy30ZXYgKpZ
HIk6vV1tR8H1LFIR2Xi2yoLs14OdjsvAGvXdDRRKEJaxPu8s5EYkAN2uXtjgLTu61BObp7fZuJth
AztAIUvQc5pA/gkmNfAhHDvY1R38YxXoQmXZASyHaALrrbJQ3UmQAIkIf3wpaxcAo6L6kahsjQ28
rS7ei3ldrRqzlOkJaO5UFGE0AbKlF33d71a7/WzYWkIcLNw+aKPUImKen/iqoEMfo0tcHq2jJYa9
ax40zaRX+Aj6CQHIsL2tyhwdMxD3VqJgUDMY+IscopORCKz0ZXXT8I/qjVpRfPv/H9RkY0+fV0uA
ZnpgfhbytuhjyvGkmNyEkuww6Teag0bRz33MTdNiJs7BT+ilcq9PdQh3DHDW/AVEFTHv2fBWpwnS
S+r8XTJOcCBbKOXkz4h8/DvGQu73wyoCl/Ks0yTlGetJ0TSxNRwMCNOOAhgKBwTS/M77NYCy32GI
q54oVPWOB1ybqk4IeQM9d8QOGoawGuUznfelsC1LlmSgQsgANZefaJjs+71FwYLyGKuLUAtnFzso
zpNZuP2bmdh7xAzEiQKRaJh7Uj0JLfe0VEnH09+Ubn7fpI1NEUM7WunT6797qW8SGJQ+dDrS5ZKa
/TYMBHN9mN0H+OME64dmEGrPV8lb7D7cQrmQOp6sYTh7tYTMo2YLBdTzggGtJN5hrCInMtkFGlwF
Ja6mjWx4LMwn9UKIz8ZRz313b8RqRPu9sC/rZRO8PDiUav9pRPmfeK2W1locR1HCx5pFDa0NsjNI
JFxFo8PtsD4rBz1QyuBi8dUTaVYQPGpVmT8nYNvjAqeWVL0/9YuFOysgr17coZupP+G3DcRPtmZa
MC95uQQd7jcqwRz64HQNzdlk4/MMCBbkEP/GqSOwu+jzlZr4PI9gtXLC7hrIHumatQuCd4rEt28f
uMZywxCdVGDEUR+51zgVVzhI092cLEhFNDQEboNtpLE/z5Sk2wsX0STjs/x4ON/hWxubNO833ONU
dP1MKFAHa0YutCGPCkV7EdBJztqrUHq70lEoQwwu25Dz8qp3H8roJFQg/SZ/8wTkxZRxGkYh0R7F
BNfnSXgvjCItNKChisDcO0Trayc3xAoOSHgAmHS3//rXvHChRH02f3K9fPggI3VTZGvfoj+gel/Y
NSCkUD6GWK2NQD+ok9dzmN+aqutY30xtTa+PIRGDrivVlFxl7020M89fnHtHmNd7u7PZoDF3TsdC
TVtkb41XYfOuoPAm9ovJPGh9jNiba0Sy2b8CsWFkLhweXkIzD4+Yp48kulwh7+E6uvEpV6ilr6FV
PBchnfo0GSm3VZxaRYpUtqg9wXbFxxERjSxHsRZejyk9bmsns56k62xhdevyiJiy3xK6J4nkgZI0
PwQbxbg8JhkF+fvtBXn7GppdFbToaxHCNjmG9AVQdcnMkvRLMT/mFydZqPua46kgCb0qOoKfcq/t
10NdEADoQvJWc+tLhrbTXnLQ7C9KooKfDRmHUo1e6XhcZB3KAPImwKVCpUOAgtgjtdq/QPSi7q8+
F+PZDzQTkGeXNAOnNIluVGlyRdf33vu8zet1IGIQLozk12+goct+Y0Ji5lVrHRgmZ5jWienzzwk8
ydnWwuSb0Oynbl+r2Y+2Glv93Y0sJI2lfhHUfo/666NGTirh2ksZtZYuMaeR0GZdghhnmTCYLxwH
/E5BVc7Cxs8nJk4O+VG3EnD79EWCCB32VtqOqSu8Jii2sIr27W68LjcXhwsg/HEdU5YHT5cm55Y3
I5cg+S+ol+VOfGC0BDlzw1Z2ybgfeUQhBvAw2AXKp9Ay5tQGT8I04iKWuksnkY22UlQzNh1Hlwxc
hzqgDHeCwfn3h5/9LKHXIxKBLE8ibLcQmZggqGA8E0OEe3rkGPmjwesnXf7rbXgaYV4f/lBXlqgl
LHg4OR+hl6xZsAcToUekdn7RTDyzuBHRw5UyVMFj81ZrVYt20hySH/xYezICXnGrJgrD5Ma9RNaj
43wd6YfzRlA6gSiEVZjm8S85zGggyyPYEhytI3FFbG1rCXHQdTpRKrM75v9XdmvVYpLATK9W16WB
V1JrWKm7mvT2ti5pre//Eb+e5j1HUSBwrUn65QxfItn1sLJ9a59dZWG7phZDZ626jv7faDqg4a0D
70/wML9htGp8enBSetrNAZuUD9+cWCyr0RddBEzVrNB7307aT0gNLP3hSillNso/xJxzb99IWTtp
SYaWAhd7OeX3t4a/c7JUttfM12ItVwP+8Hv7MeGt2c2VBNoD4N/x6W0wYhrofS37621lbhkPE0kq
2/b0ojS1K30eQLE1capAiW3agkxL6o+0SIi+PQNHME7JTd6pihXC1GhY8llP+vg0CR7NhcFtN36Y
LHSBl1A2kLiEjZrBcjAurtd+jypk7oqHKI75Bqvz1JWFQULHYAAzNxIBb/i7xp6zr9OszYQ6ctmD
sbmzb/PS7BCTBMzRZ9dF194gS+/mqIk8VFm69Of2hHFkFljwv8T6UiFekTLQ6mEAtjwy8N0mL+fQ
9OtvnLdEqXjkyZVyBQWlQ7m136TXLlQUKN9JlKKL/W5j7HMHiIONI0Z5aAzXSTFwMNwnneLEIWCo
qBFceyP26ZH1cRrejV49+pUxpbmzRyRpeqgHGA54QRa3sRLckVSnLGhZyn30aLPJnVC1ub9ArFL8
52/v3SY5UqJAMgTus8q34UFxMdb4rygH3OiX6WJXdSDN1oZW1n2/t6PKr6sVC17a0XFigJ/grDNT
ye4K1Qc8/Xd1gvf0zBSi95DSkBTS/5wq/R4vMoZlEgn1wPYWwHNLhiNf6LNJUW58aHvwaAhRM2Nv
tHJIxNl1kCQIDqYcyTuzLjy69Mr7QRCzy5Q6ig3FNVjGuOv2Qzx8zuXO6aybc556rxticLhmCk/q
MNVdKYiYuK2A3VJ3szEBlAYlYUM9FlyAOsaW1xEuKj3+LLxGzG6RO1jlLQcZICfg6Z6QQGOvD1me
obpc1C4dA8MBsY/pT5qutsX6DhmMTk9BA+M/QyBuKSW+4yAksLFzL9xnjLB5ab4PehGkOf/nYc65
Dslbkx4IX2gCqJHEk+lOos6YsOFkZ7/Q3sPiReU6ewPlAG9olDJHGOLmhfu56esEShWkG53B4ryB
pbpa+EeVOOStcfRG1kEHJot0ZF8xuM6hGC2D0E7EYZ4HZTVOs3uBx9Zq4b/johw8wDy1QFTMZGDu
GcwltHu+PKZNwjsk6520+gKc+RF3tZXEn0nLOiPrPMrcAc4+Pv0GExNgoFEvu4f3RemQ+kxwQ9Zc
bNbvqkHySFonyZ0W4WpoRX3B9NRrt/9AcQEkxOG+K0lHdRmRJWUznAHtG4cP3I0xohH6UQfQpQoC
W5WgtmOXnTVjmuvSXXrkm/ygM7qsEzXu5KiUTCh3hJDLGgdoCxTop2sbN1YtlCMBIic9WXUwt6R1
8MeCtCJsb/9lkXcQucQvgdnTiKtypjGUM1ya9muVTW9rDpnTpd6KL8ePPcvkMiWAXI9TOjNl9ulm
YSr1N/aWMv0Dg1egiwbhUcpRgkAOZ1tAcn2CM/DP4G60YuR6Ea98RNCE5WbASNXnkwPr4fK3OMld
TqF4JO7n9azOgh/Ao3dBYzderrCQpFLp7a3dRgaLzBSbIuOkulXss6NR9dDxND+DBT/9X6d9dgCB
OmcS4E2T+TJgJKYwyNy3TgewawXsdYPWlY1ewPlJdLE7kQz+eb3X1orOa7WoqjSWNGgBiVJnKd3Z
oPs/dAbGT3nSpH+zpQtEyAW0Vs0lF7fjzYlM4eEBqjmTzy5AuOPSBoNTZNkM+kW5wO2JA6J1etfy
G6XCt6g/tgjTX74yQ972OAFfVZPDtJgYEX/AQBkgIQpukIbNMd1lG3bhVp7EsNsv23YKszvXU/QD
9h7suEriCGKzuAaE2Fb7bVr0QCRIutHXrjWsijih7fiXBl+fwCCUgA2hrKjOKHvWa5knr6Qg/AqP
FanMSvcwCGbUK8pRbislSIMsjonxYNAIi9l9Wl8shYMcqkPSuYj7F6YPT2IsstZGb29LeSWGfh6j
Ql/zWdXEXb1xcKCj5K3cXd4Tqlx9tZcqFN+dvfFWMrWZADjePsDbkpphy/kh7CVXD0pHXrPX811A
JYVzaz1RmE59EGzZXsQHKQnZEMpwSbRrVgdoy8fDe7ZQJbu0xz79jynBawt82NiS9AvZagHyXmKI
QKioytGagp7yBfvZ9fX+GQukmi/jykpVV83XhjnHhf/E/b4xh7GFwbbcPY1PPgG41GpDEfayO+yh
trdIqDxo2X/9MiFZPZwzvEDpWFAWgkrUIemksP5vbBOB8y4JGn106qFG2W6YiIBersFvvqGAgHQ8
elTBJNotxxH3wxYnN2L9+LQ48ok+8EEkJoZQ1Uy1dUtbkN1Dvlctua1aiLJIF6l3Y7RY1445sU2k
XqHGyQwMCBoiS7+88Ftx0a0VW/3CUnOCtu6GC1aK3CUpmvZ1SsOgVcQaQWUN4+9f9Ao1I7gaK5GV
/z4ll5TlmPj9nipqjNJX3KgD5wDWizk8yObOoeVDcHbEhqZYifHjlwW63+6xGtx8/hHX3U8/+HNV
/tVT5SgMGz/tZpfNqMhTeUWA3cr/75rM5SArx5ZbFA7NBa1m91MRsYrLKM4U6WI1hkWdpj8I/26I
rjr9mPI7TTQqQLVlN1PzGZKPiEhsrTafCZh5Wq7k8st9Nda/v3xk7+fO/PHd9UHXgdg3wzbIvs7c
y7CPOJaF5sW82Togp7wj2ClcWSsueONsjGagEoAMA3lbZp4ymROKmrmvLLozx78cOv5Zy4EWDRM3
HSLUz3vovS+UjeYkrsYd6FdBPCV6nfu5mgFZAEg9/5fAPLeyQJ3V4/pCMModRWspSZdDcTUpGNW8
nv4Gn0C8uS4PbArgGCme7SXf9CIsY+zK839IX5enHLmEXC+Hpx+VA8RoQKkEOBOzqpr4ChZD8Gdz
YZW8wSmGs/24oUFHyypfK66xvYOJTve6mTPDUO7GkBF5uTWwqKcJXRUW5/dDmtOEKQHEnRTbbLGY
vy/ypfevFuGGHAlwqO8qhtma1LXOmqlS/x2JqAzK6RfMMiRpG9pto/G3O8lv7X85I3IsXNnWd1vm
HucUyLNRwfyFn2UOk0ASYGT43T7Fp6d49xLeZ27qG+gtc73NsLPY63JGLZ4cxjtkUWHCIJvX3fy2
V20hXiek+ZWtOKkjpwIXVnX7U3cgekRZR0BTT/wDmnX4x1oNl82MhcDnto60+FkDS/JX7g9ZLIbg
4s5npVHqslMxlVP2MDIqQ2np5YhXiBHquo1DNSQXJ/JVmYEwk8STkNO1Qw8zKVeD1+pJHyvfTV8q
u8J1wCZk37EA1hRs++6+goKHlnvEFYcHKJFmzqcem3T0kXyLLX/kKiGfo/hvkPyDxUiu4DH1Xc7h
ohbsazF888FiGITegJQXW5ICpWzNGS77whoMCcg4qBquL5FRQTBigKN5MJMtgiuo7JnsMlQB+PuU
XvJ+GVuql/k4Jm4wAOW5F9yWJyRhII+pSznXQpm872XvW265iV3o32YxSabRizMPaF1N4XeKRNZI
kFFcCPxeDei3BgVCesL8u8jtsn4Q25I+GULPVBizfOkWTdhlCBgcPBn+LUVpF4mgBuViA/nq73Ed
dOE85jHFsx/1u7gh5ucKnC5G7nWzQg3Ysxdz6U0B3g775+d1kYlfnFoKwzZRPriblpzhJ4RRMqGG
qgITVLA9FQ5U+UbtP7nB5iLdrcV5bRzLvbgDiJU0sSYD55Xd34MKFgSSgjrEn8EssLNTuaSWEGy6
HjSxOpK6rqxD/kBewmhUz3DZWdyb4UPRrwlz9Ad92PjF3kqY12A/+JX9p7OqMXHKN0QHSGpxC0jL
3JSyDG1ZglMEYHqGlIQzLHO/rO5M8f2vk9dakEBm5eVCp/x1nv/W4jvbZp2waDaMspeYyfH+uB2P
biP84OuWFwFM4h6kr5JF/LGnAg1AY9I4M6TE8X9Hrzbty47IoqnoE5elHzbrP4GZMGTr0IDkCKQy
uRGifcg2Rtqth8xBB1HYEv/iiJFIzSvp7cEmuT4Zo+zvx+VXVgp40pOl+/YJOwSA24gLBcsN8j2n
Ka518IBjx7wnq2gy7tWO6FTtMRf2uYUxxdqS47r/EPcsP/u7OosEQxZLolJK5TTocMu6km+rPKfy
luEjRZ5xPQJc1REPigtTWenTAC22VIfER4oDoVCGUwTcBTaKzillja01EmnXNkhH+uM4p2Cw28tg
b6tDp/fnnzFggm3VB4qfr0XNug9KFDXIYGn7t9Nulk0pHefdcIbKJ7AHv67Qmk/qPYG6l1vbKh0r
sPrfl7QWZwNQeVtJpSZo3X8TXKb+Iz+/ZwZJXyvN9M5Yz6pZq/MNTeuAJGx/jTUPnApCugdu7dWl
ZOHaUvIDoFlWv53totvdyEuSCJoKUw+01L60VDjx7jyNdFbfLdyquLf6SBuq0JNaofzwnH/lPg9l
hG2vU8jnBszDLtvHMEIxeMNRKtq0XYtf97iCKUrlx2D58PVcSfXjL2Vh0InhfzLfMdjBSbvw7Pv8
73pxjLV1LjpHctUradaEBEeOHU2fd1YTaQMkmvnQVj54ZnTe0iaD3u0pm1FeyIU5YqIDlO7F8tQQ
laEiEsPmxVChAeYerhXKP04YoZMD9dF9sRrRsHRYxdRUMV5IflJsY+/D4D8O+6NES0px+nyU67Zr
xwp/2Me0F+3yCB0OBIbC7uObxULg8VBc2yoeZCldKonx68SnCE5kR8LXVR9yXrhdTDr2u6fmjnoh
4X7NRJQJmehvHWKTlIwFaW6uob8ZR4rtSgwoBhabOcmHbejxEvZ+nk+Xdxhm+YTwdFES+65f9jzO
uYjGVw2p6jb+CslgTcpczKfaTaYfEe7Dprh7LNFpY70htal0MTd2xSSuA2rZqBdM8XTD/hko3OJn
5wJ0lEAaAdxzlXtG/fd82+QYbbORzGEJ0jv+SrdxjbgcQp4igXMBUVthU1nZL7EGGlXwUOAr3+Vc
G1ptQ6K+JT7fO1DfSo9simkfRi+AFmE7LYjkAJAORCo1lYcfyDc9pGSr7y53hXmPT6Mw+UMi9hug
O483waowcRm1cwzPM7zI02UxH7qVJUvNLR+Laz0LWgM2rbtP5UXImwGPc21B8lZNAE2gJ6BZUQDa
/PVaiAD63CtjPcJiyl7lrtWPB0gxLLoU051JvGhdZWTE/tdnNeMIq4ZtVj1uY2JgadbHH5DEEuim
b8c8JSWsktr5H/aYmGK62zZo4e3/14xemi3jtJPDsmXVufoBSwwFazciGO6G+dhO5BCYMYGs6LYR
wbgGR6vq+OmlnairMUKf5de/H5HyL7tQqSVZqWQbbAd1ebgNcjvXwz6RFPh/S2IHEZ9L2XLQhrwV
ODCwVSdie7hSqBOxRHCrWqx5Jix6YwCgrscU0iu4XXISXWZ34UYwCxG7kwZIfcsAzBWGGpSUH+71
DcFyZoYk5+0UCeCztWzgKWZqwPeZtxAw04W60sqstpVRU4C67LYY4BxIm2vQkWfH4X+f4olQf8ns
PShhtmEHxgWg/q1a/1VSgi7GcavF+zNv/Af+JSnjowRX/ut0vtHqFzVAHF6mrKwNh91rEMFffl37
Gta2eXwBoLg7oi4zQ4/umEH6OFkawf1tTu0Rs14UlJ/zZxENXvZqGaLsHsg1nNjXiSMG8dbHdklP
7J0fosOsyBlY+bjgskt3oy1GqoG74vt/78lFXOeSOCAa24X6cEl/puCTXD3mliUFIodr3fYpzrB0
wlfxFwpvVo92Bq3NnmHiDYhEo4mmTpwhe8uzrr0qatznpCmyawd4wVSztPNM3KaLsl58x6w6z8ph
c66aEtEP5b1Szbv+bYNjtQ+IdPxr/l8pgLb8nWtaEVQ5BEpFU4X0sj17GxBGesudKIAp07QJWLoo
BvPxLYx825I4EKx9H1JKYOSOjBAZW+jTdw2LIFNY9wC4SE3aqJoVORdtHr6TQf8o+vG1fcl0yPG6
2cRWHBkAE9L1k2Hvc2NMooh9JUPmjyGYp7OcQqt6EvgdibmCoqazrsO5FbihQrE4mvR4IQsVH7Bz
YWpWuePvHAbJ7Xz6lXHv5yF7sUhbk7ZU9wM4tRUVBVkcsKJYRwiZ0OmHWyCBDC0tG63c/G6e7/jj
4Psjlngo0Ltz7P0ce1iCCJKbXY8w1ngEYPfoGopnAT/ObdXgklINdCeXgIB1sAeY5rRt4PIXTGB8
c4BpqRun6p0qenl6201TI+kl5RMMWnH1E9T/oHH+6Nx7SmhAwczWaTw/3zMUzwaDuSaPsYCapgEC
9qvYpq/NdtZLUxsrLpAlNigYLZb8dA0Y1ZgLLAGfVzplWpne9n23XrXH/d5HLF32RZv4/2/a8ks5
Q/RrL3++hNaxuCW2xpF7iaNBh2EoPKmqqpW5dNwfWU7/OBRdk0GcvMu0B/BxaJ3GFR1jYt//M2rw
pWEgUfg6vG4xubzG/+Go7NZMOOieONbNkNIG0BPUJ7fOuXUACnjgU4zkV/G+Ll4BJEMvloBHoqWb
5pAh3vIltyQUhrm4VJ0UHvPMiuYrxdtdNiIq9Kx4n6rA7mPGYbKxE+rYVmbLB0EwZnj8klkJ1NEH
0EBwu1uHuryviavg7KB26B2jxo/YghIXp0zzcVgyOt2ab19RCrVlPWXd3ZPthc3OfXuMmROn1s8X
vEMv8hY7kMu3s6xuAtyL97woVWH+yynHMl6/CF/47ho5I7Q3GST/GVkT7Kv5m4ewITDTcvKnNMJg
6keszRYMySdE4S8/MdqTgWa8F//10pWgZNGTZtfDsdbKCFSoZ7YACdyY0M2JzOJ8w4ktDmLwLxma
5jOS9kF1FDmJOuXmVAb9fFW4WOh+4vLjtHyA3+GD0FPzJsW5zAFuMueeqFSEC46bzzbqOn43kCJ/
z8vv2Hovj+7e4AdSBvsy6XMnfOAMdyuuUlEUUIRVwORLCQYXq9BN+n03foLn1ddh2qznXonQsO0I
XsPozIBCU8YEIe03W0DEj4JLI+m9F3d2m5Pp4alEuFv64pqTxwakzr3DewumMB0PY7wkfEzx/hhN
5Bdu5pwxIHSIYz2yGwOSJTEaWYl9eSEr2jRN70Gi3lc+ErE6fe+Dujo6Ccgdi8jH9FwMUHi5A75i
fBwpc6s2kF3t9isFD8BBskAF3ZdcO3+MB/mZORdWpcVG3dzfQRUhT6nfhQsa3EeqzHzoaTvoYmmD
JJSah69ZJzQ3GNN6y3QAPHGp98b8EOeRamKFta1V5vHAUPDbS2QDKrspTAgs+oma2yew3PO2vtsQ
491NNLNR/tr4UxdE2YxIXbl0mxsfRgQ4MXw9FpDbH0LXqqXImdif7Qac4w1mtx//Uho6KD40lBcj
rS9EOSw6HmRzIw3zvcnqSlOKP7eMDnqpF1QHfAriSZ2I/Kpbasj7g5ph17Rm/jdal0qL9eDW0K5S
yCvCBTy6DPhn2vXHYJk1Su2f5i/TZHQmjVZNC9ORhVTvXk3GJx9AxZc8/wlaNAZcO4BYPcwOQpWZ
F2VADVC+GpvusbBkbmyVFEyc3M0uZivRB1AXp2VmWo7SFeY6jURBeBMRw1gTlpfjbrOcvGRPsiar
Wz7+3AU7QMmwcWqCPM3CnEBdsSjVmzkzr0THssOU0ce/I1o2bKFikmVCKXTXlOTaiZo2GEkP6jJ9
XqeRF3RfcQ+pF579gRLrg9ACbAg9XtR4Kw3O81+t1sYz5Rg74deH9YqQTDqEIZEmLNbc+EmGIdb+
oJdebYqTR5VSyX43fso4U5/IMvfF9MhTwxwGm7Mi6jh3H1HSXZM7sLxAs1OGNX3QTKlWCULUzBl3
h8by47KF/Z3FrU1nn6sCngP8CCzAtIzHkXPCv5ODVqLMeX4oP4U9gMaIoAJGQECpTOHYIc6/dn7e
5iK7lSAxYTFoKq9McNENnw5vWFY2mJ/1uJFFxeUUrJoL8Wy6TIpfI8hiYpZI5zfaegq9CnRdNDNa
aAGtkVs5FKQjJnZ5PTT5bz+qCEKQAIEt8VKztK0ucjwMEKvAcULO0tprHoIwa6CHMRnHIhwIXZ+P
xBDejBgj0WjAskJxEYtOAGV+3uJGI32eLGFF8ghVs3QOIVJEN0OGCaTc7lAMdqfbxsl40HrAkoAT
BCZ66rhewaX5V7aFkgT/UKFbDReECvJ/fHIsTI47sMLOoC4gmOLbqIzOZ9gm6B340N5OGJguD8Ey
xTZnLcLe+p/GDCJ+/iauCTGLJqTGx0JndSoLUNuzXt+o9cWsMqHIemqV7YSuwiB95Pdtkx52nbTo
q9dXbuWcW0jGQyvrKAUO91F4s/21mpY9t1xVBypEjZ2oxhScY0hddMqT+a+srNKMQlU7NxUxbaXw
u18eBG5RR5kBgN/IpzGGy6/VggkGZ848y2dzUMyzjxuBlIpq01vnxA9W83c/rm7Ig9OMXXekGVw2
/lme751ThNcmJF0hxYGGd24cJ/u9fTD66jjcIPxo6nwvtInqNCpvb2snvoeO+RgGTUTSXgsKZQhB
eh4oFZNJzlFMIiu7ibBOMM9CLAUzpIPRA7V4IIwoboB2noZ3MmRNjVkIAt/lc/NwLF0CH+G/nDlB
JW8A9qL7/1GHXc353DQlLGiefNxZt0NFTZSPlKZ0aHflfYXzva+Itw2SOahxWXdft345isIgRGBk
TcDhO3qj/OYysZp1VTFGzGeID9VG5btEndWKqp5sbvDMBtOCAE67dWghsotx3Szqu4vigzH34cL2
3wfl/GQXbKZu0cQ+PcuwS4XZuhYRHsWvHH8DjJnvUjzWi3GD3yyvVT3+Ni+BGue3kurIsP+K5NQ5
MsHaX3kANGWSp80h838s1MNL154iOlS4cKHgayRUiGCpkFy9oJO20WHNy+/vOmboYVYt41hDfzAo
olelcG5esXMwgp7RzrlgZDb8dT4eXiPXHJxhp79twvAEsGMlMmlZXC6aRIDzOlT/aTTq4pEngH76
XeY4EhdEAPygO2/y3k613YnHOBn0x5GME9h2HDmTSGfY1GOSEiypDs8yF1gfvyr2lfpDbAst32VY
Yfj8XAC906xJ4W2Pfzq2/hKvBnsAfDWSFCD4zttziFjQuluKhpdlRKKq9MXHMzpZHAqfWaKEnGB8
u5cYXG/OnOeDorI98WysU4cu/sz6Hoq9E57PXtBEKGv8/thZJ9Rc+7OY9t/SmHMwvo7ABS2IU2H8
JStV/gKYPc8/p/P2XM/amlW/LZw7GJrS0pegtBzKruDAinG2O6nA+nQFPaYTECoPsl9/D4mFceeZ
PEWLc65i/0rmhk4ZlE4/kku8S0b+OC33X8UXikzXOsp6QIzkI9jsubmiT/NQ8uzUJFVCSWbH5g5F
qN9QlgTKiRQ6VrvT8y/wrfhDSIQlry1lghiKZm4JXXNag6rd7EFlrE+wb5x9yz8qRu0evIvjEDiE
+didog9AQnOS1nRQzS/1btq1EOHSK7H+6tXSzoX4Z+inldTJpVheuI988lVifPYKfKrNBOekwCyb
mi0bcASwBqRkAUSu6PCBs/yNhiX+uZG9zE8PUR3PGKQIrD6Hq+Ynt9jANW/5jYn1/HNYAtEUF8hN
ne1OmUPYZVvbn0r2mUw1ZSVVYpglYTXsQ/wQYgmYCRXUswHT2rSP1ujZehrItuaFYR6315OMRrrT
aPwMcI/tCf8XhH5W1V08m6RY+AtqRwO9jfzH4aWlfpByZ95XQGjK7ZUmET/YZKzh2iHxBSSkKVVK
SqQPxvZ9l41OCmZMeeVOBiNsmwT95ejyys2PBCb8DjcNYGoTUJwK9Nl4soRYxiqJMQ4Ns6QnMyLJ
xnwC5lZhWMHnTvePkIXBlEPH7ihorZioJH/QtPfQiyBh9yrlknlV3synTw7uTffT74JFhhJwEFYb
QxMFgOlmJKPE/A6Odis5xEQD4JCbo6IP/oZomN2H4Y+2qEUyaUZebISs6arXtTAa65mTp6vaShS/
F14cU2I63G/Hmsk/Fo4YIUgwEOiYS6mMoEcbK6qjVCDAMFHxxYz8H+ZivcY4rJOO7CLTiZ3K0Buc
PRbifocD0pCRWmAoE/N24koYNAhqK+t48ExoQlGFeFSUmlsPaJS5DFRkCM8qTwWrKDfGcPwSfZdb
mAbTecxSiWfgUlQF7vg4hV/4x/iDDZ/obxh4hiwUjfjuyIUs+u62YXnVFKgId64uH951pkS5W/zM
UFiaJQNOdqu1rwUOMgjd9RIsd6ctxVuucQk2BMoUqDvlSY/+jYFBuxERNhpo3z78A4v7hBf7vyfk
qrlHxnA/nSvDVvIg9BASuUkzIUWMI45jjLL6zriy3/lrBX8Y1iIncq3xwGkl72diyE4RcUEocS7f
3OSOYkGyMcjE7/hODhLAQU5Km67fbZElNmVwypskFCS67Cdlb1JTAqgOx6gJFoH0Allb8T0+GqNu
Oy1VdHLcie4Lv0nKVH8tuKZFIUKZQZ/kKquIjyVBzO5+pp/rZXsjSq4Sr12C+HQ+tIQ8HfiPSsTs
beFK1D2OO4A8crlAvy0Uc2WwL/koMHd6Y1RtPSx3reoSXQfz79lYYlenfcaLsBMeSf/LZL2hl4UB
iF0ZxU+JJLr61ys53TtuS2+QGpG3TSTF9UWnsQkrgq0uR4vmzoLQmZGYM9hsfHa0s6JeJt999c/m
dOF6DN086RkyEFccpR2R0moeF0zYkk2ePO0yA4iE+5RuwjE5JA4M6LS3iE/N1fPphwQNrFJOamhI
O4tktLvzbnX2Wk0wsMwe+STkFGCOxakx8iUj7SCWpDCGw+/liqqwSc7PSRccEZQaZhNyRHV/X5Kf
SA52AJHsahjSK/7Dwo8PuOITdgHt+7U9Eoha9zvRwYZOw0KmoLPyL1672Vd2fnsJM2TdTlAxxKQy
3mh1OgNPltCuPaLFZQQfu8Gu/t6BhOcybaDxLYVuGgTSEUoYs4oLsn+WCX7nuBL5MPglqka6cB3L
D+96N05NqA9/y57W3yoM+aqmYePWnq1urg46SgzpkzY2BS/F7b5PEq5PFBp/G4T1lb/j7DEirsbv
qARBQp7cVpqDMCqtXMw0wB0M6fasBmnmEqUCXDupTB2kw7L5X26vn2hzMv2PoHihfiudYKNVRQyj
DkG+WF57CMVymBmv0JbbfJVLoNbfnH7RzjvuudsOCbKlC6hofxLad6FPA38/p3wssYweHPI7JiWx
6/edj6cd9HMW0U7pwHc5+Tr/8Xhyx0FMFM6XJluKHt3BslOKwfvEFQCXekgclmUrsWdMW83lIh/x
NoZUImW3G0UiGHTeVZq4ZBPHo7LxLDNV0L2xvEGDGhDUxK7XTnd8pUb0PLQt4TF0czUR9M6Ij7HQ
Z0EwcKHmapnPPrNNU8+mp5NxLEX5QHIViaRKniZM0lzPnteNMOJtDI5vX1xMydYZQJO6yDz5CswL
cuaQAp4RA0JsoZ9Q/z6flxATv/5L0RHu0yfbeFZM4jfQ3NGj2z2ZwHKqcRLHSOAPUFocdsZ6ntcb
OkoMDBBgPReiasQ/5cArl62qQJA+d9M9JLOHcOjjqtNk9ZyvrzJ/a7z3o3//YaO1UfkTksxtTb7Y
hxQSg8RrhTkLEUNwhx30IeauLBjed2/7/AhHgOeQyyi6h90EBOCSy8ixBJCNnp0L5QZSUjiuQ7yd
hHnDoMlyfNtGO/f2j9RmM0yZkW8AY17SBdIqbMBwxh2JiK9K8Fr1o1P8EEc1gRR4oEO7TngqTPgY
aQeTcE43tB4swxNsA71NiM+4pngB0HV3jnuKTBUCAgBwdTOj5Kd6qI+f7sXQWIN+p2Q4sTPCOneC
GyAeGTavszu28qtPiokEYpJc7ql0+YRPbSSku7sVlFGValzNC9DVhMQXiM36ayB4asynGt84rNmv
0q+8IVuBLvCOUfwpvESsokJo5cfJF+t73eclRSMETdtIrtlYELgtGFYB5lTP8FfOpClwxoB5TjK9
nNLB6ZYsC6Gm/9PkzF8GGVaREY1E3VoFNA/un79M6cF3J8PBX4coE4WjmGduRSOhPbmVwTQ9gskk
KOxo9ynrWwkTX2uZa0T8PVQncUyPsCzp0ssyY0KMvm0hvpou6OBCt2x2lAqKskexa8ZgNdgEnuC/
1Z2FwS5fKxt7auTA8wYuF6/vkcoTCdnDpmvAyCY4qMhzkSEVbKw6RREzuSzxg/ll8XUWerH4Q2w1
j0FF6k71b1Rvv8XDT/EFZ4dvRxKHdd/6860NJJT97BxrlbI57oFDbAPWuMCyWXJwRSYt8sa0qttF
+rR+YqsMYR4ENRinLSCwI6WLEzFGyW5dsaL2flnjZ/X2LQf+YLfpHZxwExu2/Gf5+nVGUBQOIheX
O+/2pvIIDe/kFJzmXtyzEsY+CpFgdLKx65kRKD1mhNNPKS9tohcg5BZ3DkYYdZ5Faan+SV5OViIa
6ITdXfOWaiEukKKucmnZwMtryb0fHhavpEPL7c3amqlS1e8YIL4fD1gu1g7IYd/59UM31BLyaqZX
Q6sm8Fnqo1RgBHtBHUgPjyGwlcqooeI77wkwOs6cd9UYgBxU/6pDWjYFbYtcIHNLDWPBSCGUwykW
Wsr7DEBsquK6HKRIkVGud2W/MZJGDTxneNKLACFZ2aMUHrnUhGxJq/GA7BH4FKlDHSp4ZBvrAP40
ZkX8JQiC4R/P/eG6gie/Fz3wC/58wHc8Eh+z1FwDaM7ZD5AgJusB/ip2bdpSJ5+9ekUG2aDStkSA
GzDO00N4HuITSDpUg0yMpy2dN33+1qucuRzBfYJHomwIsRtVLdSTGfGkV0HKD0Tq4Sd1zEwRiqgC
RCx65srdoaX8X935uKlNQzIMd3lxRf3+CD2hGnMvAB/KmxC8QA/nlE7dz9DDXFoD7LPR05v+gihp
/hPnd91GcAp0fNielypUUYt6EY1QT+KBRtnqzK6SXxPVngQsSx1MQgDQzvWlB2LTe96A3RvgbCew
qm4nsVIOO7OG0yJu3jOqpS1WyPr7gP1vrYvglfu9dmwl9Otv+4rM4uX0x85l5YpNABvFui3znPuA
nNSYB598hqB4/BR5PQBZoEmZF9cl5PEM3tpaNEcJKDylTQ5ZykzWtzLlHJ3RfCQ3jZ41PS5eZ4GV
HibG2p91aMaG4jMLdGW+x6nL+0kk1IRvoi7DEeSI6rv7GipXM0BZfn+1GVISYSFlETOrC762oLXr
MlWWYBwqcEGDhdc/Hw8DhiQ+KmvRKvVAzn5k9s67VWRxAakNI6KzyN67e91w2OldoScYY89J2Aqj
tEVF2+9ALmA2vXnKxmygcCe5mDfrofS7TGXWqm1e7lt/KW7uktgQqqLRaWuY94Qj4wWaoK6P4WHF
0jpVlBI8nrf92Y/2ep+jM/oA9P/B/DwQjnyW/q7VsoD9ykGtXm75aPw9fWWpdHUNHyCNFP6uza5V
z/4wZeWHgNKTwWXTQvXvDP3KCvRTuRGVnJzrXfBdqeRrZaEG5gXTLsufUN7SH0S4rg8wbbodueTo
R67KrKrrVURO3x2ReKW8MIiK+jNQ2e/SGeSji1aar2hjPaj5bmn7hebR0Hw7NefGRhXLgPKMjU9J
kfLgXIH0uawUATMjCdhDOWBq3dzsuRHDZcpidhCfKgzGqtaZiWeMTpzwFZlVdcMY19JIel+xyP80
rdPOy/p9hvI+k67YvgUZQoJbXsUHy0B51Wx1JRy1mFa6WaaXZpEXLESibvp/0nfWo+AvyWwxzbxe
KE2u3zKWFE03QkaGXpexJFmQcrxsjsfsoR88/m81RgJdIaW9IUHdnKXdrWlkkd2BMMQSRGX6oJHs
xddr5Vkgr/1m+c9kpxWsT7nbBDAHLLo5syzGupEcUYjb0NfwrywDZMYLC4pZ2y8WbvTP4yNwv1pD
w4gEP1P/Id09l/N7mf5EN/T4kU/i6ArVoawAlQAXYJW0axs2y4StoPKA4Nz9lifjCQchDF65g2al
7rBLOv7C+WDXjTOW5wsFb24NcfRJstDgDGqEdUAowYSJlu5qyve0EHbFJEtUcicQ/ATbNhYBdlli
aP1kzOV9ywTlv/x8tqaYsfgE5ygWVIIqnMxljfhxXkYzS3HuRB1Vb5RxriiCd47icLfG38RklPQw
c5ptE4zxJK8NZl9BFmjLUE3PKGDn++o8OP4e6+3BguaYqb3b0TjWXHO65Zvorhf9la4aKXdYNAQB
FBPnub6TLsKrD1NQVEdD6MerYtKSf/wYON1Zf6YPqlmrWlxDXM+cHRt1tFOaBJPxQrY+id8ttTXY
YTv3igpyeHK7lQTgNgCRfyEC6O2Kav52cX9wLZBSIfrztZWWQutUMV4IhHMfEzIfYA4/nA9t5uvh
zaeVT62mmKHsx2wnYloLEQ8LnZ95p5DqBxkaNP3pzA76dfJrRgLj3bCn5P/BnAZaiJ+CY2Ko12pl
XtUeiCMF/UiSTQPuZ7FWbgPW/TouJsh1my2BJDwD3G9f+TjRSXaWr8UY/Bz4v1MXIy5gKt/LQ2mU
nNSJvoaPHwepPg8pHYyvceeCuavcmCHNkC7culA9DdFcQU+NOjeg3lW1NqRdt1itJ0drjV2j+WgV
MQwoRM3nzor45KKfvEXptKNq2lh79W9JOSfhLUOWBm+TU4/+1Q6gm39t9JxV8PAzKh82vsUUj2Pn
7cLq59IZR/xv08D/j3jTm4CGyrE8o1nUepZKebh1smRAuzs5EIsEyZ0pQ3nQYSy1r88y0l4lBogw
NDlce4CWO+JNSoxj1BBQCZ2/HTlpf4ydMHZmaKyau2PWft+OQuA/fFZ+1MSRb3bsUnGHpjOYiNKG
ce9nAvY69Na1sBH0tppQNxcAsQnncoecH3FLpeIqA3a8R9Nxr3ybgruS6JqBJPHrubal50v7PcIX
SFsW2VJxhvmQ3yWkmnCE04Ex+drMxJMrjh8u9ixmmX7BIWrYpCZO2VthwTgt9xqGyfCHVLjRoAQx
KTpNKq26mfndNeK2nISg/VsB+odkIFHrHC6xcZ8So0fY5Bfm0VxfP+VhH+IqMLqi4K59oAv9/qbC
59M3a2SWhERz1nyg+tLG3P/Hupz9kG+RYKRAyISrPij7mdsRejeFvxcXeel73985VFoJKUDIVpDl
T5BstxD2STnFSdWc861Sy865XRZCRwe08iwZ+BGs+ee5FXVZDmQCydsHk72Viq462xoEhxNELhPk
KAPajFsG2h0e2qS1dYrBd//w9VDO7g+enxrYTvAEFjgt16b5fjONkD2XFmVrCrnWhAQylqVsw5Hj
YAv5TuMUFX3IC85Fqf3w+iEQfNdbYBtwQmhMG6kWsxfLjOoYje+ViR8YmdKqJKCrGCV1PLshZb5f
uurZYyIGmPp7kXnLDqXVANHwBBSYR6hiEwOsIglf9skY0aPMvwYsBBfgDDnXLqxJ8RUHrZifEGi9
Qc2tzz5tK9MucnvTBzSvJsOu9PwltGmK3f3PxSg8HHOSJJ1kIuRpFemdKi6d44dVO3WawKcp2dZH
T56DHGd6MyPlCZlNRkf/Sdi1k9BOWFAB2DnHS9DA9ho29C1DYf4MR4HWz97+lDJWlxkPhRgwrwkS
z2KiDU47zeD0/BQD3XFwZIwPaVOdjzXhGxIDhAscMXLfuMA+rYrDY549VtyqyvXCHCRBMoMW1JKn
lBDkAEdn8aYGTTk5hH8vuLdOUDTcOoHV15mrjaHFHikH6RITOXMT42CdopczaLkZ7JhxYr4bgTJM
uyA3XGIML2KloLbNFfk86JTcR8PG44IZ1JyOxl/MJp1EQpawTMpkg6qgEq2PRDxUBnIaLrezuY8d
42n8IwzusYpnYMyj6RL1PHwxK8C4NH0jECRi/cb0ybQTwy84YLkJuwql2boZprfZJ8k+nr5HVh2+
gKQxU9CETPgaen2IfNBzSuRmqBgBUJ70BmUNU5A6Wi44NDbfCSfh8y144UT21iGHug9Dq1nJBTik
Fa4R8iNpUc3kKYV9JrIuMt0MntKGlIWs1UtSGRAyzjYfXavh4YW7YVtQ8ZN1YXXKG1By3EDnZUfN
MdMuxcHlL15Oyv65jiaaeci8amDWYda7f8xSi5/vuRVX2Z3XZJ4ml2x5sIvYSekL9kJaF8QHUZvU
AlZOg5OMhMqW0Uui+8FesVlB6VqDoAh1pCclYikn0Z7NFCndJEd8zHaaCHftVgryilCV3nhMnXnS
brBPJuQMuRszVyWiIWpT5gijYBLfJomI0nOuikjPwClj7UxyAbTHRJH8KDTQtBUON/Po2NELye3v
GAuoj6BW7q2wRQwnP32JSa+rBYynFJWasx260k367cLFxnF8sCuMe+TOkFRXMjZ0ZGMu5xatg6hC
fJQNtaoW6PVOJexro/BRzPjqadXtN2HTKKnJEeGuzO0fNjD8I44UVwNw5Wq1R6PzYlGnVTZu1W6I
hmDUoWedWDCYrnTS9IAoBg2OHcsmlhBT5SPKOQlZXOOmZfubZkFQnvl2YdsCQbCa7SzJUMCNVwJy
hqSzUedV3msT0GTz0zPZ2ZhDkcd2WLvj+HbvER9tTgMrSxkg7WJ9ctoBhqZ12AbHyHZB/DH3lfto
CUczrG2E3LMRUMQeYCyBdK9wVv3ALd/RBVlt2JDyMfk0sVMqBJtShu9BeGe+RQDz+HjgXqNf2zEZ
Mv0oleiSxiqUjqIwDO09/tyRZ6qjFCqyaEYrDt2FmOd9LpWlbmcFw3lQxhw4f73FIslQCVKWmP1b
kadyec+R+gnNwTe3GDnkiNMqi7BdCNLh7FYFzQTcd2kJ4oUQ34r1xs2As2wtR7ia3AsLRT8v1dgS
OKAyCtnodBvMVr41GASWccrFyYeWHczo2Ws89g1XepRIQRTUpBqpax8KrkgJZCu0mZ23x69JWu7W
BIw9z97t1lHqpeebyZVTf9taQK5Iptu42I4mkd7mwnlVqh0mUz8sy9tAfvuPbuKQtMFyKQfLmhCF
snVMhKx5HRs3P2vBiJCFuJj60sm0lO9pUry4pdw9j6uCu3QwEnGZpaCbGbaW2iw6sM0k1nO8B2us
jVT/1Im2CDQg38qrAASgpHmvN+usOhjOWJkpCUn3eVexyQPcA8DUDRokyCenvqlNPc9dDP0TRvgF
I+siEyzkFYf7UVCaNtjoQijBMWA1z0LUAXwmKkukXr1TKVdBI4FvQaLBv+5RH0ajSDzXr2CeawXn
G7HYw1ir1ZAZPD0++TZ1godEbzFdudF1ix3yUQcy1pIA96HFX8yEmO4oU3XXdpnMm3dd2HuoGkgr
PoPadh7M2ygz/Dcala5kfAW5jQrnugtU7aVI27R/8Y9fKRbnzzed3/Mdj4bDJySc8yyAQZQFQTfJ
GXhphr1E4TcZr/b5ca0yM6Io0APBjyAV664MccKwvhttYkEBKAdIiMOt7rOTFGGQx1diRxANVfKy
zAG7eEP2gFqKGar53Zms5b7sds0KtnY+Su67uugyTan/Xyb9hV+DhAU7nUsjOAUNLSUaTDhLr+Nk
OdXhsCj358pCv1abj8HLsp942pBsItfPAxFaUOUoOgsI5ZHy0gfrkzv4qlTZ5QVfu117/3yeVVoD
/lMlZvKyVGV9+LulKtvDP2Z2XC8uVYgftqlh2z3Vk7H2PW8O2Ds0/8WVwdg4+1HNOVf1nOzj/V7o
bnlo0MDrw4OTSSHMap4daGdVCpXuP2pPuPCz+qoxCu+fj388AMgG6z/OeHz7KdfSNW+fdYWB+rOw
P8GNF7d73DD9uYOzvBrX6xiCu6jtAtYEcy4bjkmfH5xJscHE6nc8K0rv81EqNnMB2CA58q5nGISG
KibzllbBquUjYDIPI3AtHrLWOtMeXNCA1veFtVrg6iCPz6eKKQVA3+d6oLB+C8+qZRL7IMqxuC/3
mDomTuoLa1Xp7tGHT0HxyEfQn7+/FC/BLIfGcYAY2GUsnd4JlPHlkRMmIwo7SkX+T7xhJ80Y+1P4
0/dlvsnenFCrwpwNc9o3iNh/dRq2rPSezTzTY1vJXjvtbKRJ0BS7WMSzSSVNsWoTQotCKNk2/D9e
X5xj4i68tLLqcvE0YRibcn47WXxyyrMvilTYA8e9NT7QMjG4Gd3V7KA8hwcxCYPaIqct2UWT0Jqh
63mQClL9rsxOjQo1gO6zZqKbK+xhS/O7iUMAcAitf+9KIb6dd8nuAadIUTJnMN2lMC727cAEdAZX
OC3Xat44JqiVbsZH6484lHM9OcNAYTsNBVVMfemDd2z6O8cNecLbiI8RRTiWW2U3vQgQj+Y1s97S
JLlNHT0M0bjCjA2S2kQPrb+tqsYquhr5kIxXPsA47yzsQ/xivyOmL1cHFNd5XjQBIp7jLgYwqnrV
1waaSGFxPlj1nbYzVi6D0Ogm0MG+7yF5JUcJitZGIXo4jbXbY5UoI06EKhGtCN4q325xRIO7DDSX
nIJnghbItkYiolOnPXcwY/SFm+ACypxKm9Zu2hCRNZtwFEdjdaBeNJ10x+ZmsygOgYOUWV8E3QC7
DPOCtrZ1dBB02Z+gRYqXhKkJZKxr0KfFGHN+V8AipMufI1nQQS56QtKySmXzb/PlKUXZkYplYzgN
FPyK7Fl0czIYApbpfZZg8AVAo3+/BUAvhEkW8S3l/P9p2jJvfRw48gBa58uggyxRJ5jKSy+6tVEo
bw1vNTMhT1wJodajVr6Lc4YzCjUSAsh/khzXoKq2fptSHOHETfmLxgEU8XnQdkVeDgpjqId27r+n
g2SWABz3ns3QmJWfQGqGLWfcqtuV/U5AgrpxTlz8DqOML9yGzfXfRTIyvhL+VhKgfe3I9ODz8/AL
/HQYE7tdd/iT9jbzRdgC1bjD3WaRt+ZlaBhaZqpb+F2csI2+EEVxk/IDFKPLo5DpILk2SZKVgCGp
VLYmaDQke7wpfe1L5L79C90Ua8Njn1NsR94Vh4tEbOVbev/3zdwhOUc9/0VtrVKuTl5mfvYX6G7g
rmtRm/4g0I4lw5UV9M/5bWEQ1BQwvk2+GLDelhrJoBjqy4aWDAWrmvM8fB7NyutgQV2eHLmtlCuJ
uuf+wzKn3AZJugEtId7xzVOrhwzf7rJTM2BfFb/arNyOvAZDjNxDp6zwYSJKHvq0EpvNVP3YEaOc
+nqQ4hfp9UGYLUpWz2I1zlwQ7ammhivwuo35fHpO5Ys1VcsfqeHob7cly7unLU6zeT6Bbj0MvwF1
vHCorxj7OA3T48yF6bJCPgSEqaE5iHKXI/zQhT1D9kblYAa1O0k5R3WNd8Fa+BUFQU9TXtuMIWXe
qkSVI1aiE9dXiiF4/JFiv3TKEeqwWAXBRSfd0+Ng135EXq09/og5DzhOB6cARytIclKZNP0bAHH9
4hXEgCGT/aUcFc6g/q91kABPz0tRXEMEaw/b0GiKVfOkaXibp4ZHvy6rf+Wlht1vxBnbunVUIqOC
u/cgSb96f0Uzmbn9whA7nrA/rR+HS1gsT+IdAvGW45fyWPHZCEgz/kLlFyXnpTXT7clX6PnhtbkA
sUpTJECJxCNSzj9E9cAp/2FAxYnEvC6qlmRyuq88zVRZOIp9F2uYPqfC4Dw3frp41jY4Aslnj95+
I1LcWt5H0/t+yak75/otxyAq4E8tS+Oszz/QjKoiwUXhWVmE4iYwREa4bubiTe2oLE/S+bJQ05zj
koVnSsC7poFNxLkhDgBBNKmXY1HE1BDK3vsOvxOLz/qxcTxIysZCKsVyCz7Om9kq5MRsa15YOg3b
Iy5Qjua6uMDarvey7RGbq0hwBlGK4B4JILhH/5EeYHw17yQ18a3DhtrHKsyv3AjPA2o/9nOHtkI9
9Hey/Oh0GxdPnQqOZH5nDy4kBdsypQ5O3QdlaAOsB6gUKcu7oHRsGPakKNNTG//FZ9lwM1SvJsXK
r7AaSa1ViuCBx4vMXfSbqAn0vB+n0P1n6FYbuwf+R1mX2Er4jv5gHD9k61tZ9FGbn58X/zy7OPLJ
M1Ygxh+cXghRtfhheAhOKaZeSLf59cRXO6LgSEuR0xSyaDWxzU8cycnwu9LZMJWj7YRw0RJkh2Gi
A9N/ZpkXk2895i6ltfCbdJKSnSNQPVh4erNE1XAh/t1NyFAUKK45Y6zp7x7mAQvtm18i5723hHEa
OdtzjakdH3xrF0SsaOF/wvDTJthsumC1UZK7r8Z05LRPLCSa/6mSwLyp4XzQ0yKGf4ui5vIwG5pB
AKaFuyqLVD4BSWfrEJ3NvCwCGLlG8n1XTqOTJaSLFYEyC0jHLWhtQ+iLFuA/BOtxYYPFSIAHDFjc
IawlBUEjrOXsT4GTJL/79FL+/kZO2oNtopcDcW/vmAETMtOGW8SeSPtciDCYE++0dziMlWhORg8G
YNg+7Sbn1M5ecMZHMWHB6mGcx84Abloyw7BIiYSJuxakdNP4wxIwK7OH/4KJjJXlZn6uB+n6lomX
OCZ9VQD/K8/HQBaroVeo+A1plcZJv0D30LjyTftRRp171zCZbXt0tfgNFJtDo5S+FYBjNoCqIgeC
Smh3yHtRV+QnhOG498e0yvVUFBKIS6wKS7K3qg1rCx/6zZFWlDtXisCs7HhxFjrBQOc+oyimky+w
l9cfnF2VWFkF9MvDPWfUcZEBWWT9IC+YUS0V0N1c5zFc8Up/9OV6KGkcXghKYh1z/CQNjeM1R4VO
C8ScdUBB3etQteziNDwGDQa9Qw14sHSeUeuTBSqUvvmXMPpTQQh2joIlyINN5jHK4NqBgL2M8YrY
JaU4JjWDWBFlvamqZJJcVaSIZde5MVn0F0AapDG/i5MLGHmzuc0uq4n7jn+GSxTDEagCJiRoCQsA
za3ECPGIKjSiHcZQiqEV7sWDUp3s400lRqbbvQFWq9RyxM+kV0GwKfbm9ph+r6OUqpWkqpZ1tv7a
z1G4Tn9HL0FUAQGsFI9kAbhk3oN2roKLnWWt/pQGKVIcOwYOrojFQqnVuiw0ldNYpr3EObv/OwG2
npmII2q/O335IsxOJoZK3eZx3Trki6awazaL4gzE+3Yr8QjMXR3DFmG19Kt8S9dyMCkWvOvG/GEI
15k9p4w3DVR7v9xIaGRwRXbKy1vjEQTw/71ZB9c4FMaiQXwP8qBpAKxbisGbANbfzUh1q1o9KHxv
ouZ99QcftXOyWh/96cLeujgx//KZO2GTyTZsdUNaUV9FLaTF6/UD19ueG0CA5sINtaocqdY2YaUn
TVJN8GhnNiqz9n5jC03ypCjNXWvYkON+jlQrwsO34Vs9cJwUqXGfgGsV+DMKwwja3tv8CFby0D84
DtWYvspgLbYmGhkHmdtU9rBSZKtFycj/+ghN3gqr+sg9DGduWDRWX4watWKHQ2nBQs+arBPAo94/
8CW/8qRtmPMAPZn9EOCPZOmouw3YtZqOKRUY5A5vuF+jn89FpnsGkOxmp5n0ftJjEzOaRB7YxlXR
GuerIYTxGDmLUmv/Gvi5j7pqXtPYZ5U1gPLajzq3Eolc0Csf6mZW3+SFge5h/W/2A7/On1AAr+ql
0sDLR2ekmuN9b91h53jIshC4fGFHaz7ks/1lTQ9yx+1JJdN4nUqzVfpHtHXUG/0xy6iHN0s9DR6e
6qjAWxIZGqZyoEaPqdzwEdQfHhNt1x6R8sbLdgZGX7Gg3t+6LSWZN0bMcTqH/MWYfnd68D9XN2Xc
XolRSHeaUvSEUK5BhAFzDrkd+8mj73xGsDwycN1UaF+OgMNU23RANeQ9FrgcI/N2yCpSl4ubV0xK
Z0rKcSNI4vHNnfOhdICa238Bst5Xqk75VSAEoM8xJv4lA5MjUFrvXHH6an0upHMAyvp2yk8UkLVT
wCEoKUEfDEExvbXqcac85YJNfTZ1ihoeJOmQPnNae3ykRmmdhaJrHQHH1qslkeQg58cgeyEY+YYY
gcAnORMomg+8VuGACms065O52pgc67x4Fm2u3jE06DJp1Z1oweHsWUKgwzZRhgvqe5fzfv7fR7MY
bcaEWCDjnuGG07GUSkNSxP4qJMDbudiRq4k1bNxjThFKAHp3A33yeLZISwGkdP/hTqf2amYT5/J7
g0WmcOUN0RN4WN+Ccr1azIFMMVGTkNtZrrtmxZqXmHZSDwyQqnu2HbyDvFsnw6zbZbCUdhyMNzIK
ltpyvGKN/wCrcvcEFHP2NdZXPjKuYvxBbCOddwOh5SKX9foVA5lyqc1uNTOwhbzhrb0Rp1WVZCBi
ErLs3wULfTZkRp+9b1LN44GBvmc9xRsDE4L2tDGW3TveJc3Gne1UJgJRflZKzTcN9DeusckqprnO
6LhDbehcbLN04u9GDARTErhDb3pgJax4/Z8kKnx2D1H5hCxUgeqLykLkJ6eYeL44thG+MlEMK7Dh
i7hKp5xed6G50UoG46NTDZMiEC98IpXCPwb9/XhCkMYc9vL0HzXh2OiLAm1mnqUWc1TzwikoheaL
/FR9/R2liPoABjtW84M6rRK7Cj4XHSyhCOiTxOcHDXwoSa0ZNw102ZI/ysapGuzEmCeM9XNJ1ieL
SWTarBSIK1Jz+EvcDM3PeaQwtW/VLoJfCn4zyO85gfSSfwkK+q/icX6sMeJbPmH0uj5Aisvr8s3j
syVoemIwkaMCkv5sCxJIcXbGVGwrdWf6v3H15fWYgibEgymz2hpUMheCO7n9JC6i+euZzBDdm9Ay
BTza3hiiX4LbajwWGpuZSQTXH40afaVLbKEedPJKF6B4cVifz2j6hHOUr2GPorzX6RS+HeWZDthB
vf+PJDFlNEWNHy0rFxmSP1ZYrObeh7uNwKWQmB0QFaNu1fBY0qxt40vFf47TQ6P+q7GFng9mZjZC
1SBRl3oGGuppf+SkzAeOeuDQbZB5zLg/iUySeHw0z19x7sHXFD19da2hNh7lHVcTbYJcxqO0b9Px
cQPPD2SRgJS5959u9HRhOJMJMTaC8Pjki/m6QHHoD3p1aQOxQ+Ci3ec+fFxu+si6CUxzv+Bt8b+c
YKQex1z3AX57w88CllHKxOioEEZrQCLLLaqjggLrhGd2gIpi2OniYSXigEVyrPebfgglEQjx42H4
3BI4RwylGAjztt92+to6cIlHFvd2DfHHq5oBkG9R02TjVnmQJFjoV7Frz7gw9FKbet+8R6EgVB0o
eb7xhz2ZL1kRp/UA3QdcDZZ0PadwU1+RtZTwyc0fufaPeJxVS0NzX3DGHs2rtpy7fWX1Obx3rN6C
XtYwzufDip1UrqEhuG7miyeV9/tAQsgORKRxSWrqz3hREAkgjagY5qIY2rAuZ7L0NhQFqvIPr8tr
yoSAN0aXxgC//wMa1dOVk30Lr7+gTA8zTLRajJOo8yTWX39hP2oJCQH5binHOvb/KjzSC8vQelEN
rGABQZlIY4ergzjjJcd/K5gFXeRWHDi48pskBQVB1w1nJMtpq7tEgePl+QUM/asZ50vu/ctKWujJ
Naxrl3Kka8cWcUcLBM8omiCY7OCM+9ynFj1jRrEaWfEpig6ozQiGTc336bkzQPyKoDWA+0WFiVR6
uVInKQVBB3qpRkVD+ki3esEI//KlYwKgKz6tarkTb7V1+d2XL9hf7Q4NtvAlNl+01hzIFrta8euu
Lf63UQcssb7SYThzbbPhaL+inHv8BqK7dwk5xInexpqv+CmTc8tRLbfZjGsqLSHbeFpBvhU9vkfE
MOVlje/csaW5QoKlP7kx5ysGZjS0SSVRv17rV7kMYPAE+eLdJF6X/WzZugaTuYuYaXCW3E7o3CIa
IBUAEyhTXae4rMkBjdeiiBDPPc7UPb6wRBKcrot8AoyDv7Bp9Lnz1Djq2kRITKVDTr+dxhznMDj4
lONKCdo/hXtnfZnbh0pjBlR3f20QMzHlB7wad3vT+odeB4whj7ofp7KePAzrqgT33ho6bCdYky1/
Fhi0IGsYf1uFVBBzAQIAd7mGb8iUrP/e0fm/uVTzQP8R92Cuo1GD1SCt8YA74I+j1fz5ovtDfGuB
vdtIT2kUnehoUMIr7s0V+T37+dZfsctQIWbNsG2Ht1HKduoJoUOXIcWzko7lDF+0FuA5D4c9JGVx
gX/alQZNSTz3skRvHCXjEpho5ZZyGjXgLuUAtfWGuHc8bHSDMS41M2muifX1EWrptDetG7rF9Aa0
eZeNYbrcxgXaVK6CRYHJRp5eBRlH/5KwmL3SCZdV4gykP1JZ0PzRYyz9a3jjoN7ODf0fm24bsWWG
2xTxLVXilBB6ZWBhan0ClG+dyQTXPlmQM5jr1eNsJt2ACo5thLOgBkadCC0qGtKzldkLlxeao2Tw
hSC1HySTUPJrVIi8DrgWHMl5eCFgiZfO9ugD1ZYHePCGmzzDLVNPnIvufAl0yKGBd119aP2BaGC/
siTqFgtM++ftuxYf1RN1o9wYYcIvwFeRoKgBLWUPIKzipEujRyTCLS80T5dJ5bsawDk4n0ll5oWL
wCupNcBZBDtwqIB3uUMT7UmKpk4aPPdCmbshXlAreMbUIFUn3T0mE5BIlRuDdtHUEKZt7foTxPYq
wPNavwugCS6ylVEHuu9eSMVjwfVKRVHX5KorM7p7jBmJ5b31tdOnnmg2U4AbKUDsrHd8whKO/aLp
mHE6dWxs7GobWoTFuboLYvYMo+3GpJpfVm+fyY7R9L5ovBSP/EvDnQ2GmOABvRLOLdTZ9rVrDDF3
M0eaQtzY/ardm6It+67MVLqSOV2PkbH/0mt+YZH+WBrQKdb3oWKz9C4CWr3UFMFD9j9pgQI8ubME
VEePAswAC7zWBAi0WQoh5qbUocfRYflDK9uVsl3n2bZyIQuKAhg9YhNuLrvLCNtgkkYa2oRtnww9
CnhY0C+tlZ0/2vuctsFCZSZiZmeJrEx2PtGmzQs0QDCp+KBgco4cScR/1uMROvfW+BnQyX2vzwWB
AmlN3L74mp6IOQjaJjnuTGsz8sU8TdKZi3xoKZa7yBMgq3A6UHMZNx40nbC59h3AaIJN1FjChqxC
eeHEOddkUYDbzL+9RCMruKgt4xZ8L0KAx9Cgn2Bml9ulLf2KEqCNf+1ZBsZ4WJhmjL3TXAx3SjF2
kfo5vuod9Fsv62FUtXOy2M06V/DuPdx/zwoWWOYsHyiNQh0ZK7EpdTPZaYCBnzLwlrN3K35DtEdY
fCDBWuPnOFsC/wQPUj4k3WNivNS/ov69CG5h42qyU1VD5/rUKQEIv/9axShHoSztTbn6ldBqG0WX
F8mOeyEp2rhMxyYBbGJAKQ7/icqjy+fAea3VcVBUk1L0Tigi33mKU2rzUA+CPWMzn+QfeMAv0xKk
M0t+r0LkCUOwkiFWfkOX10msWDo+Y7o4A6SKHSaqx9gbVO02ufxr6+cRjsJ9j1u/Mq6t0Zrb2L5t
WviD3+yZF7KX3V+S3o8zWjWDGBcv0oo6gMQzfq9j5w6gIVNUZ+gdWHAa0Aw9Xw3JSHES1LYjnXMN
DZuZOwJV01QXN+O/A79zFU2rMBTHONhZGIpGxCjSlOd3W9QIjazPXKUPpa4KZAQDhGLG3T0xd0gt
pmfZ7X17BO9gGsPrxhLKA7WD75bWA+8MiMAQbFzzWL/l9GgCcuLzWgUwK0V9LLfBH8+OE0cIP3eu
T6XCM599xb7FY8edRvcu7G6Vh4Oj4RJeaWxB0cqu/yMsw2ytr2v7DTy9YVeFE3sFWi+bdicKiCfi
G9b6bRu8N6o0vwlmEvFx7FQa0kOq67AV6hOu4fI2qvDQMZbZv/qG1+GeCT78mmwef5FJf8NqSvML
Te3k6FsMeEZlNt+t/Er2NMSQZFwE25ZDCC5U5RC2j5z1JRkf7A9Pe2b0867NxiDoUBq3XphCFsWT
LtEdn08u+AOtNEi8XlluV+EQVd7ezBKVdn9ijflrE9GKNJJJvzE5ZVQtWBtjdvp4Cx/f34tPgmxc
Dr7hNH6O4h1EDxO9hF2NgjvQ/0w4ppO3be80HznLt9z4d1CzvaIOP0g4tBp//bQo8QfQ5YUXMlPF
YII5dDG5kZvMtnNd1t6Z8AuoaL2Eo4l7vUpn20IdyvgP5aYARrpBZjnaCWUudnfqB0WtVrGT0krF
Cg2eO131Szyyf4eWUIe+JPR0TCz7vUj58Qcx83ysvt2m3jBM9IK879groRxPm+s7zhN2d42jJQ6x
0fGLXULBG5kbnidGhzipyFnH+l5xxnaBTVjUiGE3ZHrF/Ge9JUvDlrAzEoxhA7ldKx2czV6wZAg+
hNHIaFFZO0eL7iJhb30QXcMJs4IxHG1S1f/pobtVPYivC4A2cFvSoZdbjLtyYXoFRHL053ZCl8xe
zxt+WnCbRy6YUBvn36DKvGpcOjlDZqWwowpylKrKNDaHYJZ4/JGE+FhmHLmsjHtke/XqU8x7wwc5
nQ5nC1ssOfs007eJS/RI2QgGejC5lXRIqXWJvwkxxlSeg4PDSkvCDA2ld2nxMFBLYSh5TSvSv9NL
84Yyhh0gQUe4qJgSUcXZTKZhh9p3eqt/Rs6y75GC/qqc92k8PAO2ftI7UNfvtEmOTlkr772BPUgX
K5TWhooitv1u65xflf8fgJXWsJ3L+um9y4J3GWqedyMDhnYOl5lx6tKncRsszdyszDCu8EePn5xQ
F+vd2/Q1AeFChioAY6tEQ/N7JLH8bc/T8MGTzi1ijRdDeyZzc4DhMn6k/N3fjH0D8XIg+59cZBHr
hxSwCvchvmsKwPgcdt4VmW+0GWikA/PuHmXp55JuaYdzByl0VhXmgSfhI7AKk4KOVDolRe1gIaFG
2hAEvqlpLNZersffjr5PvE6XmPn4glQHUF21O6Zs6tXOGfdgYVWMR0xjEoiCLRpKJr0CTb53qw8D
/SF9ZNU7RZUBGoBOiL2pGjeNDUNqdWfEuGhoNc6+kOCwKjCm3Kk6KnveSmwWq+Kg+3A8vQtfXhqS
YCT9+tpjcL1q+WoJnFw7CseZugLT/F9WPinhLwQTF0mIEzcTN5XiiNo3A6fCZH8Z/6U2OmHyamWf
We9mc7uL0xR3SIWyigyMonOixG23wjcvaPC2YZytEiNO3ZPwHsWXJQGxeIlfh/6DAqVIflQ1j0mg
fxsb6SJ5PKvWRAGzSfBQ7GQ8DKqF2uu4fPbKpoCeLypGecTOasdfp3IqMHp/eqdfEC8QzIt1G4jJ
js/gd3w0LzjzP19eminMCD9WwXjUXbzsWjiK2wHp2/xNc3xgwug8e372KrPF5l3LhSE537uAIjwF
j5vqLtgfv+ABs4RT8mXIJ0Mx7Ip/mg7umzxFl9RoSpx+P9mqc29yi4xuwv7s6r2tasBkXmeFpKFx
AKpVSPq8FF9AGc4KFQuv7KZEWW2LUO9oZeIRZw4CF9ni94PmHxuzRK0u8QCyj16Bxwj5DDByiQq4
1ivW7yeIkPBpChCPhzBB78+fTidV0nNkQd5TIt4LkX3p6LL8MdYxQn7swYGW47ulnFekWIpoFMzT
AofSQrjWnPT93S10MBc0DH2CxRLoTf1V8GWuukbvkE3OQm+ITUcIqWhsgEcbfA6yY9QItIX+HCwe
0ca3Rc3Aay7tEcP6dBCw+i6vuDg90JW6jYtPS2B03adyVAvsW1wFG4uigjbd38D0PUMYKx/uOjm1
TaO1vLOxd2istSdX9un+lYsuMK0VoY3DyzId5HHUmFYn12NF+ox0f+0G3TQNgezU4efSXIIjkvVq
nqlLtG3erpa6USR1Z+0QMIseaL/tYLNzBri1QtCxGehOpw/07t5ntiFIYPP0cTnvBS2FB8Renino
KKao6E1donPp+BM25GPWP+EBFfZmyJlyPBF9cDcXVFB7gpWcNcN13f/+i0l/3sHUvjzJaq/gr+xG
V6ZE8pme3saDPfS9YAMnFm/jV0j+iR72dw5yYfxw3EIrof4O9OZnJaiBdvmfF3wWSPgz4MhVcCwZ
evLTPDturTRPbckTr5xLXHvQILUPOXZrjylUqbNlEgK+kQNXaHTimpGS31AGi0m6d975pkPCSs++
uR3mfJcC3RL6eUOg/T7ZPu7x4JoGcK8bjB4ZIKzFMee3GNIi2LpxtCQ6X6w+9OkB0/MBXRyPHIFY
E8Ip6VWdhqFe4jOSTUlCHEn/P0YAkDX7uUlK8ZK++/VGBXQ6ePhTAzRRa+mQEgDnnHho7+nywp0U
ZinnFCAPHgbnfIZ2HkwGjK0y6iE/lWbCSGvdTR7ZjnBJiAopwLqNJmCYwsevaiLYZzQbzJCLDRqp
ehPNlfLkGgSkhjFG92i39d+2rg/iBEGmZo79FSLYZOwJvGKf3Lay+9bqt+LMikbG1UqDBFI5sG1f
/CbLPG0z//5DeZxr3rLr0EsysZy9ZumW5jt1ifhhnlhJ2H4ZoaNkAFU/TLyx73X8QBNSkrGC6aYq
SjwiDHlfE+e4qnjCiD24/ehopRWU/scyb2FLMZ3415Cc0y1u6lNnYC8DSU0Kk9oHzAPDsa5SQ7Va
0MZcU4AJ870A8CrJxzUltMln8BzdGw093iOw1vFOmGACyMrSGJGfKlQ65b4tqTDpPiWdpxQ2dQTf
Iqe12iU2RLoyxiNXLybuvn/W3CzIQv/XoGonbS3rzoTqPwrEBGPy3JjxgqB8Kmdo6HcprnqFFwIo
alKxAeoQEeUTEWBQG90iT0WJSNncD7+TbESfryiftpX6CupXHZmM8kyqBVmzVVVrEP04yqkmdE1n
ZBc/E4UoC96utYLUVpOhOFjl48WK3aNqEQ3IxK9v5Wc4uBpAdYDyuCLxsHyoggQrm6dTLnuafSIs
MlMJZMv0ocrBP6hMVoBybEPzLoEXpwXW647v9vCkx7Ns0K8ltjSfHMapMr14NvKvkpwhNL3ZHYHz
NApmilh8xP8usJIZhZRCJENbDiX+1ivSxtZcAO7a4GI9ggL/w/+6Xo5uvBTkiRKT+yQS3XffzemX
nrnOSEk5DHThrW7T6Z+jyiyuSg7+RduBEx00h8CL/zQ+rkAndSPju3+91SaSk3+mix5AKdYz/Ivt
n8Xcy3ittkNVbJp9NmyGs4QwahkE+wQNkhCQvDFBgq+H+k+PT3wqXxMc5RoRjbUrcF2ebjKgHBVe
uv1+ZCK0kpVto6clb/Npy3Wv//V2kBNAE6IOqWAoEdThjVdZR421JWk/zik+XQk7q2RjsVydYEN8
X5u9iRuwgzxw/Zk7DT9iMzbcTCA9P0OFt6qac8/knmRRT1R+2sDkr8bqnxDwJn+mjnnNTpKMULj7
rvKbOKBhBlqnapxpPUp1e8qsvMw5mc5BRVZlisahTnudlb3MCe85e/EshdmG7bRtKqPp5btrN+VG
xlZeM6b+5tnLt2F9oD1NUHwc2nOCH2fAM+sU3vF3mj/OttwtlvuJxXDE09KthUy8UOqyWYD1kAU1
REJlGNAdq42xTAnJQs1E4+ekKfrTfIN+9aM3Ai0WsPlveN5PFfVraf1dgNRWY5L4AfnVKM9Es5rK
cTGyiO/BZhsy35kFTtKZ3q716W75bhsHlcvul6Qi7wnBgjotGCInslL870g1qMMuKjcbHlvdMyux
8X6QLkR2Sh2nmY6X8KQw6J7M7on8T8T+ED0zQHleZuZ/Q7NhLCBzNGEhBjTsqdC/3Z+Fk6fO7S3Q
SFNv5bfkWGIQ4pJfoEgciHOCCajAV9bc8fvcyoyEanGZ5TxOYB11fyttyw1vdLPCBfAwvKCP2bXt
0Q6/vafBy6ZgBRm2xIu5f/EEcmzsK/wFr+HorAYgK2NFig/17l2+qfU8Q9mMjxDma/N+mViLFeAB
loADstsLMxyDHiG02AxCbs9B1BuBJaC0qD6zGPE/yz9mWB6SzRss5+y/azvgs9+iGa+zEVBdO8gY
IIsKM900aax2Eey1tA+dnZm32AMaeB48yEnrYoEa2w7BHeTsEfilkh42jXyJIlQMyIaCUk5r5qk4
GMB+knoxkdFHPbeixUyyyuQscmspw2MG/d4rz8+grTAvOrVTWM6RIBpLkUmGXwIyxFBYBZBsMsWx
RC5OiEAnYDd9vx/abJ7KR3XVrWC70sEtPhYN0xKp2DaNdkFADiD8yw5X3WnNkBuun2SKrZyL3Wn/
4Ov73TmNMafYRYnkQ9FUO00T77FK6RxcL6vOoG1hA7Ft3MN2n/JN9PMN2njwUjrnysusGF0z2kvE
vN6m87LHH4bhy40VA46LREWVqWs7RZDkpazvyszYOWPXQhMo6E3QSE+NtSq0EWXRztVYiBPjdmod
VQcZxHggR1ra5FQkzWG6BfNcmh7iOfE+MtzPAS90lBPG85cWwDkTvk71CyEst6j6fjQ5WOQRwgE/
vhDx+V3PKkPm3L3zRgi+WxMm08tAKC/fuJ+Im29mZ0rhCgk+G4ZIU7zkzMhkEVMlJgIS7d26d/0O
a3rvJD1na0kYiQ/bLxHKlbHvb6I30MtnIy7RfuLjx9JXRp1uyoVrPTDlHgF7TXvCYkxfgdUvnCXH
2q9hUz50Q8GE1wJ8cSAK9ly1xZxXRXNvFzriLinsPHaqGdb1zAb6pIgK0TSsd/LchPiOzpvVvGmA
t6a7ZeGV9jte1DGjUXGf0MWI+D6m+/Ak1yooYA4dYkovWqrAOjZKy9ddjzsQx7jFBk4iV0Z7UYM4
Qaa+g11vYRmA5mDOyeapb3vxeUiiH76Ymzp8AC9llvUSHS305qdldM9M7ms/Q7C92RxtsDKur2vf
er7fNyg8hwEPsAf6TeifKetsb33QhyUuDLUL+GRdwDmvWQuo+6l0YVgNBYOF8rOdBHyOc8tuUhTD
4pIhDnv7bNPG+a2bUFMTTAkFAGimeM05KmbGvTeA5E85OXb737IBUT1Ig/rHn+k091kA5AuzO4pP
dTBH+YFLPKWxlvS6Q0UuXmCc3QeDLe8SVoN3D0ocKSO0elA7U+sN7vkB/3zqlpZhlS558/7wNQEb
GKg+GWoB36Hv0bWg6nR4+fbgwJ1IrvnXrzGn4kyl1DzRKpOgKWYoZV4+NiA7a8+hftiKj3O6HtZc
TcQe25R8HPmJaz9W71ZqwzeoMhukPivIjsgCLzp4bBg/OSxt265d2VEp/fKTRlkTWdlgc0kFu7qO
h4cFxYsgnH7PcV53pIBVEsMXw6o3TeuFH9el5ggLm04foc412FaCcwWVSa6mPIe7qyZcrHNf58P5
fBiWm1OP8N/x+vjMBmAwEGBqou6Uq4zjMndgVfstgIHClzPjDpH5MDWRRZ6zt9fBj72AFE4A/19B
6k3aTlwy1WCdV8F/gxQyPiU2sI3p3AriOoM+mbG7TxE8trth3fv0Q9JVwChYaMtXfVCnmxDkGfj4
r0bpTJ/8jdba63LSq0PRMr3YovsS/YKzWM/P7sAz5xMKkYt/7mtT1UXvaW/PawnzWgW/uVBxW8lO
h4rmwL8V7KVMhBAqjX6NBgMjts9uE7+RgYlbkfa+GFpJ+SduCo0FPZbWEWoGMYTuBJAbvyhHyxv8
jRWWXMQNW1mDN7dCknzk0lwnQXDTQIrHMnxNRAJX0NgkN+WyJKF/n9leLFjCPO1RGugLMmHBZeRx
TXUSLyH8no+odkJBsO4APZdI64utzjtEEL78tZAeitx3+InQHDc91dG3yryU3U1tOv5fYNGLgw6z
y6+KdhtEstUDlurUnEnwV80Bh0seGrRoTav5Tcz92yhzMQ81hhaB0VqFfgvkXRuj1LsvOEg80v9v
avN+uMUVKtTRi6wDaYPv8G003n1NJxX/Ghf6TLxTq2TsyL6nMotPTd7+8xlIPjvcaraH8N2NHjIb
kzDEN3UdwBW8qzaNmmoOQmLWNXQgmvZJ/bf45tJqV/tVkvv8tgdX7gDC49/95G1pv/vNRkjughni
rRh/xV9Bq1UpdcGa/cgIK2ajw2vtxdxTBW3wJlVkIm1rTju954COn9Gu6iRT1pMcV5H+7zzrb0ur
Hx47V1NeP9oAcQ9Wo84Kfsn5+xMaTiW1Ms3pF5EiRoMCMwxZ3PPqs+hBC768QfoorFKP5BnqDfk5
jSZ7dT+x1uDtHh2cXMncz8xn+2GFblfhK/VZLR/f8IIR9nN4zTFOvOKd7A8rZrwttKGFC+NweBSI
DmlHXtoqgMBahTUIXmTmUCUVDwFzkVWsVrJXAMXZpcHeEBN7AcpwLa6NXzq//DcorTbVoLdeF4Ze
XUPvZnXbn0M5AR75ouE/TZJgITqkJijle4OdrJh/j7aYf/NapGrEuLYk/KVAmZ+3lDuMl5cFJXAG
sl8uQG2EzhDSThmsfTVYgT30ORNJsPLF0ywUwtXXYgucN0eHog0mVpsyt/V+EOLj9yPhhtLYfuOs
gYXEWzUwChlCNOCVzy3A0t09+mdNMrrQQs4DhV9oWqk74iRxyvJfW98qY4ztyiNMajq87kAsgtVW
oifB4AUh4Ktu7Ko7mZvHcQNFoOmJ0cSQCQMuonEzcsOHisBDfJtq619s7zN9XkcgLwzkbIa4m3a7
FA466tQXNW2H1SM+MTZyC0S2wq4ArUUcjEslN5SzdvuBUpkyOm3P5fBl/p6QS+XhIPnwRNvr2HXW
2c8uVJAC81j3nb6ihg7RQp3792XjEgPXCfdOKy4urRX7yQIXBwELzxS8TudSTPuZaCdS2zV75cLd
Il4p9ETW/Q/C3jkAHPhocIE+MXamG/wsHKfMj0uFJRQN73ZMcpoOBGt+r4VveeKCkP7US+qGPpm2
R/FftxnXiQuqbMAQA6vvo9RY0mJWKN3qnEhvcUiV98AxWPFgnDNJPKKscerEpOhAU68Mf9w8QAnc
rSfwiX0pqlDrVVLvKSNNAKnNRKw/DT9vwdJqfxOjwQgLiJ3lzOKSvR5sqn9cEeEhpvZkrH6gs47s
Gykbt4SmaQNJiYflNE4Cg5f07P+cAk/LoaCrMLho6qY5erQxkGK2bl1wCiYxaqCucbVnOM2eb+nT
dTIRVODLrjKyP/T8JMp0zipUJ1TJi6P+w74lOMQSd0Czh+5z5cSeb83QyxLfiWV6kb/pm4N4n/aF
CKJ1s1Sd9WgvJ55DC9x9qsPFursX64bJsBY9Zyp7kpvDm/lh4ILKKg0hLMgPV3YafCTaSXnCBBg+
KLUY0A6HgLtDAHtc96h1r6ubb/YzHMdxIiXnzdogrmXlQHws7XcICWszPI5VgXyTM3qNvS0DkgJk
0NZCznXbFWRj9fj/BYzmAyadegIjEuAmCQYv25ds3Fsk5BrNM6/L+69Rl56alp8CeoSWJExPXFQs
zM/H+oYK1CRud6czEjn/HjHj1OspPXzap7+ISTdVUopaHHu8mpcSjlFGKoN4UPyWQIX1XfCLDAcr
zWE0jhGirHso1konmkHNA+v+a5RSR0sSQdWhUWajHO0FyXwR3quXtv9GWjtu3NxiwBBrjU8n5crC
mAVZ6UhPrfsM+joo/KZ3ebN9l4OKZuqXz7M2s0zO+GceSB+qttsl+7C/DwAG+FU2DT/l8QUHXrco
K6o2KfeHJva8eOVmfwCzgnbKZ5g6FoTX3kbFJ2AyHrQBw1Fq/dGi/VfTARImqCc4XDaCJISEi5oB
vekveoQO23NA74DauH1L86U5PD0pXZ96zsOUdQvr4Q52igUyOqjRNM3Gpu4iEWnVlGyglzf6s8M7
x5K980yAikphiqSSchjB9Zc8axbc8apO7EvE41B8DHVvc+S7Kd1k+gYo6JMb2vFkAxvRJsnJJPfT
itrjepZZBfxZKHylSiO4b55b9vc/zdqDz2y8Qv+GxC6mcLkaHDlYx19fwqizC3oMsiRirMBwmm4T
SHdympNN1e15qibrOHoKMlOZ6NduTGhQ4Yx/zNI9KOyFarK23B59z9c73ZNYz7W8rdORtieYxwlY
fNQhe22HuiU3qXQALk0R+0Rqi42Kp9bDHpx1xD8m5iO7RG8W0/COZk80hNvzUTftoyeqj1cSSeBm
B70fgZ5dRfI7aAm848Ut/X61c1t6eBaN5MU1VS8YPnS4LoWU+bJnqGmuY13jrR/w/8NF9rG5abFe
/JnHj5Y6So+FcwkYw0uIyiSAtO4+MxgIMNzRfzi04yDJ5ilic0XY/7EQ0ks9Dc/COw4JoHLv64VQ
e0R9xq4EuEDw7nD+Y5DQ8f1Oodg1kwDKPICio7YVrszzMSfUrxVUVpRXcgJE9DffjXuRgr93DEfy
tm/zaiE9daIf0XgsfIktU4SawAEEFlbvZq7x5QGkWGBNWlsvqOSQyt49YO6Sr89OdGz83uBPpg/x
nwpndNxBZsRzh+57PWm9sswpSxNG+N/Ptx1sT6xmk8zDu2WT+bIP/g+HRYoGxrhINkgyRdi0FGUU
DibR8SvjJcMdZ/qYIB1yJLGZRfnoYYn5tOdJK2Qz4Xx36NejC8w4t9ydQ5W7Kueo9WyZh9pqQdR1
sAz8U6vQpC54nLVJsU5Qv+tHo6i33gZJ+5bsEkDqBzubj5noJIhJhTbcZK0H/8AFxGG4oo106GjV
+8YuRTu/DHuzT2WJCKQTv1Wmjg5AJIozzgsxFnC2CV+K7C7gg9VQvH7a2npBMEdjsEZs83WYjwrH
XWp+KreYcUuZLmllmJjvKmwYePVWaoEgIxvVlHyYFLToYsPznSeM5wZoy2OgFJNT6QnaBVISyv0Q
oiF59ixMdS8YAZpYctF5wVvRO6qIM2fMxudITuXcD+wqJ5sL3XfFoeED6I+q1l5aQ9/pTpqv8Kzz
eqLRynaX6YoR6ZYO62rUIsSrZvx+8hd7XaEauytg8BJYlZZ9p31cth71RxEGUVxuuJt2njiRK4qr
SUyc0sQGrMSiqWPQGhl9QBGnBXLZ33ObInTjdVDaGJXfmeUG/pIeKMSNpgoC3mNkqRFeoUS5s4yC
Y2oR7XdehL4uCrIw2KSSwwLG3WyxIKniy4tw1/It2Hs3umfzYpSe/ePIM5lDKwzGn5E+tJMNg0t1
qFmebHntT1pX7nOjfWdbUC+nSp3FLyD4NT4Ybul6L8sp8lKOejfN68HkI6e0lm7NJTwz+j1B03Jk
sjB4ED480NSf9DajF0VBjN5XrUenhPS8FuBbbTdGlOBgYDKmWo+dTDqF/BFleSpGEMvQRoFsGYi4
dQDDz2O7fsgLWQoZSITKWDwl2oALWRxJfyUMMrgktm38F1Q51TXfsCjaHLv8PD/vfTLFeE+8Eur7
OCjZTjcINUhmg2e0yG/Pt1ypMq2AsARm/2lskTIn80w0qpw/QGqaF3lH+bF97A6ioAuojw1uNssu
ncnWYVyIQf6e744wTRDWqHoK+OgZcYfUkyTmzeLtRws6MipfCdg8W5D4H4hdj8Y4hEa8ucWZmDR0
Zx0imhvV4N6E/JO2Wp+XXJ77JADY1Rlf41/RuW1xATgxrd6TaBOg/fDM6nGyz6ceUv8prC628CPu
/i+qo96r9CQ2IcObTdVPPJEjY7v/7hEMQsiX2/TNBVZqVXHTMkxY3RvMXPhFAa4kP5a2tgxVZAsX
+o5PgvzcTsXowG9rnK79m4XfuYlvbXwK8bhakr9ZxZtUi25URkNzc4JIxfzc/O+UTAK7LsxVmWp7
KD/s+KQxNchENLH26IDzeAgjtmB1Mia+UMICHaP4Hks7McE3VWJhrZLtxQjmKIyUtKmjmSaXXtTe
WH2fnKtAdMKcXie/S7I7znQ6XzYY4+XpxosDBWmXl/BgB9WaaIosGWcMwR4aO8wnnHdPS2xAQwLc
RWBkcyLlJuXT/Ky5BgmgrbTuSaVFDmlxNmkVpJ0ogMRgGHK8mbh5MoP7sqmqle5TdY3m6TtuDb/8
HtMO3SLNEdJSS1eDVHzInLL9XWnB6xV5At7xN8SUAWEtDrx/DPB3bdBROgC/wq7rm6kbR0ldfO2N
hwzVX44NcvXyH2Un5vFaICmrTBZ8kpDv+lvH7/bc05XsOkjvXccvcUDKltmckks/HnJDdmH/4g/N
y98qwUoeaELXpG6BEQrX3w/XNpdq5/UTwq0abtbdNuC1jGLN4UtBwfsWfGaJTQBp+DzYYJQKxTqW
j9jEsvgQB8CfhKY5+bSFQSLopdrGqAdLw/kMWzABo5CCf+0WbhHzjiHkSnUjs3CHtVPwahxstqem
zxUlQSbAfPdx7Ij6mRMuIyuD1bOP1e2wAM4XGHhU1GrpizXeFyNzoDMDbxyS6Y7aCtoqzQ0E9XRG
qgNUg3TuFsL7BM7LuBj9NUX/73jETWnKxSNL7S8y6ERlMxrbcvb6NL9dxvy39KooxJNpPEtG+cIc
WXSBLBJtiGVe5Lx+F61WsMAzd/XGBExFmw7y+h9i6G9rab7BhJPYS8JD/CdoFf8PwdoXpW4yXei0
F9OytQQdnmPij1DTo29wf1WwrWRX6yKvki019UBxtdvUipHr87zxUCkMDRG8oeYtajd9TW7zOWcQ
cBfmBgv8gNux3npdbWr1vJwrlq3GbHivqZzsqWr5186F9+x9yGY4E0IswwV3R/dou/GZwAmKHtZe
e0uuhlnO8WuSKG+ffd1jxst/l1pQ8IDKY0pltRRBI+GWNPQI6HrVQOEwiJ/8eAKJKkhfoIky7AEK
qicUV/yBtAwjD2bazHO1DhewP2oSt6NdoYKUG38jlJ7eUFGYM/2Ho0lVV1TpVHr49N+Fj7Um54pE
BAfmylR1J6jnMQ2SK0WLrb8sIXbUNeVoSaJaCVQMn5Lu7+bkC38BWWCbRGvLLaEUzRqAlrFV5MeZ
0hVbYWI2f01AGrzUYLdlw9EppI/mqXtkBZPE5rWAJd1vqFyr1HcTLkwML/U38eHizThTBJ5FcgbT
3AGECvN77HGKOEj0tpFqui/zPo4GPB0tY5r6a8pGmDvosJbTxk18w6v280NVKJ1s2n9xXqn0FMUg
zakvmcwDwUj2tdocSAE9hBQk+5Y9enbuVvEcSKwT3iBNzZhLAzJNcCmlXJjuvn5yYTc1OQKfljMM
iYNPibEZi5CPr+RETbTvLqL293WmoCKOqCMDAuEDcWMNeWWHYg0Rz6IqWB2YiVr7XJ08AfrZqSJz
qka9xwF4765M5QKk3V+JQ3zGLCKLDRaM6ItByXVDeTWLFk7cicNX95Y7LJ1fh7qTCu6Mgk0uIC93
TnA6mTRGMy8W52NumeeN/yX0z5/Q5dkcrgNPWfCSYEXPVJciFaNPaw3Z2CLTABahn8aEV6W+vIPC
oYniaJ6tH/Dgzgi/JyVm/M0CNnNSpJXe9ve7aehfjefhjq9DCYftoTJC4ici9NiGoYoRUhY5qMCC
BTXq9pkmTYgyEbn2vjpVci/REkKJ+4xKprj3tXxO42dSMPCv4xsdLfc5sfDqAM8xo+Gv0zWgUaYj
QkdONswgy1tb+UEyXJ3Z0678PrWkhzBDPnNqikAIaLU/3etp9wpftsLiPoxp8ZRv5LRKyh7RUmrE
Vx+Geni1FuPu4nKPk02f/OZDidAs4cUNtjv/WboNnBqybLhk3BFYOQFZ8GOU3nR5+G67QrM5bjkv
C0hheHQ2iWPkhGrraMP4XMH/CEgHu/jj4/0fBSMMV26dDxUUCantWD8q9cQB5hd5mwz9CCNoe8Bv
+t4AMsRpK0kv36DcwiiQrR+pO8+qM8cxDJYcdI9ILoct9WpTbRqoWTUxYqptEx6C61LNl88cDgT7
Ys8SJ2aDPx/11aoiEornDaFCEhOddsqRd2sz9AdZxFl4qkUafSJ/eU8j6A16eeLez4b1ezWQ9a6V
UUBeLFjo+oRrS8kgHwKI7+mmpy6Mcz1OJm4sqYFewz5wuTPEG52kF1w76vaplHYhEVBapoioJZbd
AyBGBco5Bep4RoVdX7m1YPYzYWUiad02poqphvtJ51LVXs1vUHpF0NqrwSJYL16RjEbghx+KZFUq
ayZK6WxCwavt4btesT09yBjokL9K3UePPpi5W+xEH98bnVF6zJ+cqZne6SYfm6Ngw1ppSxxz0yxs
a6GoXad4FdlSXDMP/61Ho3pdupGsLDG6LfXwUTklhMzVS9eqbpJGGYOerBFSqVRD03laXNmaYrW+
yTI7R2LoMGqhK/ob555oMns1wTPGMJ6Gx6u5bvTDRx0VUvUfeIfWsbm7dyIGmQEq+EsRcvPJDLzA
68aN1aQjQAQCDOg5vK5opWSCo+G+EDM5WVsIihsB9wpW66tpYDyAawgUhVbniSOVpWxaCxnv3bVN
YZWfdkWEmeTD6uraXUv7vpXja+R/RQKK6e8EoN08PxxoyfhOcYbmXCDBX3IF/N5nuftZ7s9gR/2c
/zJroc0X7YOzAwDtuhwcp8daBcNuKKHdPdkzKdI0Oi7KYiLwdRC1V5HNw9aEib1kliNH8mQoy2F/
pjPWBJNtbk27JsYVNtHIbD20UVn5/h1g/ecGI+5u5kR1o5FIqLo9pX5fj3YLQSqnRs+Pzm7dIg6u
J4UzNxhjQqMpkZVI8IzfQDxMRCELkwFHAYl+u2oO5Xbr90Au5Y4I79jMIwx32SRVdZqduXs+enGU
V1QWfKw03/FiFTPUyc87Ypsfvj3RF6ISx4Dkqu8XZ3ieejIhnYWT2K5j0GF+FFNmpJskBUzPo/Hy
6RXaiyLgxpofhfiO2e4SMEcxaJh/+ZV5vgPoSV+vmemuEZgH0d+X5WGK73fS+ldGzzW/Xs0rTD+G
KUbnOGXPT2YvMJZm9mxCGuHmowlMmEorIHtcZrVfqE37th842Se0PwJpZvZEE6SIkYqJY50nHkjk
HwKVKnUpqAP4bkDsrHVWpggLGrVTI/1X/w2wWK3DQrE3aw/VT5Dc3icKjf6pp6Ba25p7LN8qBxo3
v/G9o4CbQ0VyROW3vBD+pgQVXJ9EUI1jQtm/54oldMb+miJLuXqTfpUPvmr1PAYHZhRpmapj7Q2D
A/8MkGIffH70jqrxl95Thc/B3JsR2IHM8S0keTyTS8MPMEN2m0VsVV42Duyg3dmsFFtOciv/wrrK
7wobCm1t1OCuGNJ67iJXCKZ92KI9NmuKA+qpKGV7PYu+uMbKEvvE70nTIThhL67xC6XnIPyjuvgB
MusJPfksK+Yt9Xy/tmCGIaro7SfBZ9pZPFPxzSvsoaYMyzBgQwJCO9Dl3OjYBM/flzaM3xGKN4x5
qzVoRG0fCNR9wmmzwKdxnO9n5BDxGwlRgGtMNNLtvavGLiPEJ5EHNhQFA8lVmWds4DDiRTSj80t9
iuvNVgkFSCk1JdwmI6zkx9mvGjV/fCzHNjEn+ObxEYgh/8mB31N0AmcAREbgAPSss5yC5V29MuWV
ICj1hooQcJNhtJPmxP4ITwvk07tkbh5GpehGEYL3ZYWFa6M92memppe9VFQ+5ZNvIBKCPD/an6Mo
/ObkrXGB6URUhB4ByWLfEz+g+h0YqgTlqjihO72zA+cRqjgoIAxwPzlwq+6O7Y5gADkdpyEaAP34
TRCAu5PYzRPpkz1vc6QL8T/4/ufMKPQgEkLmj601SzLuAhnTwuS1vih+rHSC4BIdmmlTGOlYZPVG
SwvlOCMO00+whsOAO2WCtgxNV869FwJY+Me/k5ZlfReXJVOA7fV3UA4LTwXV0/c37mdXJ7RwIi/5
MAoTKhguCUvEIQ6I+ttVeHsaY/56W/nM9Y5CtXS0wK+at/LMgN9JhaBrkl3SJbW4AAYAySjZl6io
pZP8n4olG2f2xzBq4lEns/A/Isl27r75Bzy3/uwaQsx0DttmEFu3He5A68uleBwKh+WuaovXMM2S
LsBrSvRpbsouERBUUKJHHn51p7BWjjETpI9ar6nMcNvIdaFRnlFDUsmeC4Kff9ipqptSx5Qigno4
NgwyI9UFOCekPF7AmPJugwrsOtDpYMhEMJJRXqkAgNOkBDvLlsjqY5lVmB2CCk7abx65+yPXXYnN
p9GBzoSlQ4c9tNDDIX/jY05x3vsZ1IdhJsvZ+boovAzP1qXQIIMNLPSbOzJ69ssKpgD8ERxTN8g0
ifbZ0Rjj983hPwv0qX4pULzkW4spWZ7lF3dHMXYRdZqVwirWA03Oz9qi4KBWT+qPe3b2yUvaZsjy
qh+eiffuEIEoiON/p/gdhjriSLRI8u/ogz7IB3f1ItqreY9EycWxagsaqYQc2lnL9b/VhF6Fz1zs
m5cbIpL/wEosYrNLp9cb98BUcJvkGt/34YLL25MiBwSHfpN5mPA+Xr3CwZFDKCzKFaTVVO75W1/7
LK9ASBRMr3sLGA0uW7a6DwvUZjprnry5l7msfLM5bS3aV2QOdzy1UyXPXfthjGO6SiX6+a6/6Zzu
5m6mqaZA9KDaU8OVGt5m5U8e8IqeaiEAnpOlUwk8dnjYOVoOrNS3EMy+AffrBs+mYzLp1cbpqmkD
2PDvr1hfwjnobvEOwtuqL9MClR+xtjvrpCH0zRZpyLwEDNu46qc6RCoXwRaMyQExiliVrUKlHVGs
89yoMtEaCN4qwPWtCH/cJzNhxwzBf5QfwRWa0Dmc2SlMUmyYSvoHigNeeBlStWgAhCIoV6DB8u/k
AlEpgwwnAGxZN/1guiEf+Qva6SF3xw/pkQ9Ppga/CLmubMnF+077lfy4oaNAPiu/xhDfWPQqIy8N
b3StQqXwosR0o1D558Arz0ZjkfI53ndy9zJES4WbegQXsM4cxSEv4v1L9EfI1XX2SH31n09kDoR8
apnqHHTt7FogkZdP+apIBfoYsW0XmzlZRrL1AvmMmb1diGhf+JNK8nux1gNe7cEpLz/eehm0oPw5
V3BUI7tX9MujwqxtGXCIq6zbpOAfeohJEms1bXKSISRXYsgStZud6FcsyUt6zLLlnqE1X5AqzqVH
VkZA8o9b+izRiM17QA/AynOtU4RaLSkamyHaBjBIBnHq95/FABcJ4NT8KFGawjOUrx7hWA4bOzXu
ORviqrtdW6IHFmIvVgDpWWnC3P65BK83c1mcsJmNrGVhhBX9c6r691arTsM/dfvlJ3a+RJDcC5oc
+gvNrDz9FexTtfpgnxdTyzjW4LNB1yS9Ly5RW/Vksnh23rkWQqzm+p7vC6f4e8r+pq6ezShMkMUE
jay0ufKZCLyd8OX7ujdCQeXfi4CtUGVQmkNaWGiv0tmFwkNtWHDvR/0btQJBkIKJP4Lm0cHW3iRW
k1nJ/nioVIfDv+R8R2Z2aD3ubj0Qa0b0XIHqcbSANf0ao93iwN2W/sxVo+j/ZFtrfXEzT+7J74SS
gHiVg1Oy5AhC1yKD+AVby2EfkxfroAt4ncFYcAtHVNjpcdCLm1uP4yMhqCSkJ1YjqcJkYgTrP7JO
lH4K3xbFIu8/R7QnfnCEudBTjiMxtwdedwQxyKsCHhhs8jFgxzi1MH7LojHqi117Rd5/iU3GP0zw
svePbHZgFwq/cL/sqEaSLExjWSbiYcyh9auGHnAHYT5YPQF9sCBqOKxHtsX65Mc/Gen5cd6yudmT
VVxcTCQXp1XVdu+G3RNhCSUPc4brbnBg0PjbdEqT1PVlzknqO8HVK11M6Z39GT59BR5rYb4yfuIA
m3rYcMwwLyprgStooagyr66/0SwAgT368+giKRR1JSKOemEC4EdUX/9CTvtMlx1ncASw/hWAS0FA
Ge4XfCjH8MTrpLApSnOVo3j2I+jVYpra1f9YJBRMZMfcIgfJU5L2NM7epJJQSIFsgpneB1RWEQlx
WlSP/Dkc5gHNdar/wFPy5z8/4GAqDh7AJYc2K/k8C8C6hXem3snmkwAf4aL0HiKAnrxow8x3Q2BW
6Z1bLFkLQJpmftHaov4MwUfSOtYl7EPcEzWqvLsXvW+Ddz9NVPH2YloZ1g82wSRD+v0Od/xlMysH
VL0v4I5G6TtTQZ/Fnf4Ij0gVAJYgLmwkBT6oPn/6dlfO5GK/yykqbnQtBZPvXzMqteOBE0uroxU5
EA045gBlj+0ChvQVkBMSomBZuKEMMysv2i+qlUzT6C2FuvWku7sNh+IhyqcJFkUb1Ha1I72vHY3c
EXAz0Eml4cf1rlw6nSRysYB89gRkYOoEqZKE8vYytpdY30waUgZDsbgB8e6hd+y9YM/y540bXw/3
BRykW48YxTSJPUnB7cD9VuwpBe9Um4ujeRzYLu401CFwIRKj4JYakw3iXf0hJqinvw2ZWk2aYUC5
RS3E0b9IUEVmNkJiwqXQj+jwDq2AE477tO4KW7InUb/vazfisE0+YY05LGhHKihX2Wrs5qv7697g
gJcZiaZxGzjIlPKlmW2u88FyTCNqQxNfXdIhNmJ0Dt5oQ9YfhSGsqpvm0XFfteR9do2oRzWsa4tM
nT8JI7H2psR9OSRnhH/qMT0mzyJdzJAVdY+rLWIBVrbzNFztxsTbKCS97eS80o2K1uUQKzarqNUZ
B86n/2tCtLeCp9NBAOFOqFgy93tGA/wDhTVRxKk0ehRDKBZzNO8oPUWM2TBXm1qu9ZPQ/GdMjCnj
riWvSw0WcNpJa8kr/D8ZUuuvvU4I9klelTCpcumCePwf04UARdtWu4bXAfB1YM2XMbPFLhGzL9wL
WZXKAXPyl9RPCB37wizxRb2K8pwlNdEpr8LZMx8haT6HAoV3FM4owEL6AWCBqWmVgk0A4hs5gRKq
TyoNwLYV84zGuCNwRVvhkuzGNDVGZBErouxfJwCgq1MmKwLpCsvGWAaMFOLv2kfEhmsIPI1SuYg5
MxWVMpUcHONGcgooHIrE0tK+VYIx4jxO07f2ERCkmIW93NDdBM6yvlAkNkyNu7eT2IfXGArLUEqj
IFm//OiezGwtORDxT/EgIuPsqOTEY+nk1Mj+h0OGIlolqlXwfaw4pqTPl5+ssjN1uI5SHKvaV/ko
qSnssFVOVqKzne613lJ0urHajeVecZYlZ5fmbSgpugVz3Z4NfmFhMTxPMi3jeY6ahNxvbwttHrMe
wZ/nyThzaWbo5nMvObrCuBufy9tkThlSJ+C1CcGiFvrctlgaSgTDKnr5ToqWKZgjRTOgwOyVqFUF
H1qgkLZ7Dio1ZmGMf89BRUlwRyDvh0M1kZeX7q3Ycme4ygbCCfg1uK7tBueMTcLgCpE/+idTxF/N
rNuvQZEt1eYOi+97VxL1orxAGPC8z1OQxQrOCPhHRNXLCGtQeEZ79N1Q8HHkVy0MjkaPzyb7xE8Z
P5XAzO8go2K2HIiAb5MWSGhfCifZSZ2zOi+03nkdpi/T86coIG7Tg/vP05/mEh2jViZ79Fs8oMUj
LLwKc4A2HFEGAyICrwrJC48N6+2pcYPd/zFTTbcF6Rp6TElO4G+yLtI6adZ9kkbNq4mCmpWXbz+l
YItuEtShiwcYmN9iO+1SGtUJqR7MSDI3EokJoSuvwljWrLJkqzylMAL0WmwMajlRGWLCG00LXrZB
IQvdPIq0ihMZQ1rhMnqolyNrO//wmB57Xv5Cmh7wdkq/qvxRjz4I6BZrZIXint9yUptbQHSv/uOM
/NM2EO7b7rpaTqVnqr48WPvQHIFbH5x54l0JAUnc2QPZzY5Uh6dF1+y3RCE105YYOvT9arOieroG
32sd/Z4ILXuSVLbiAw7YMGl493lvMwitA83RNfbhPNikAXSwwBkZ/WHqeeNsVh+iO2e5WYH5FaJy
Q/FnogOJbKnrr/m5E2bMUqfOoxexfGsvcaJZuXdSXV0mY6uSxFjqGW6Ad9MkkQJjXnfIT9hqX3gj
3BCYqZoZAnf+xUpsJZ8CliG0XoCA7YHK6jQNkLgRXwDsZRDKA3+B1spawPX4V9PrzUo1k3FJNWX5
5M+zGS9jgWFLsiBfxsuMu85rgrtPaa10MOj0zSAhXiWl+FkZDgYXQ5bej/1X5buN4JjUx4ZwAbIX
dbNcBP6G26/k1qfuR5mXY5xU2SVUVQnoQ/akEClFoUT/4oWg20NYw2HzlYqCr8M+Jk7INnylyNED
5YQBUn/bjzRFnOIsdiy4I1aEZUGPF4mzz1G/1iBeTiyiBcJzhprU7qVltmZlvYm7HpolVHGVAMr/
mO1LxcqbeyN2gScBrao4drpYLiOk0wvhKy5btcwLEUSPxNf8O+WedZiJP7KD+RoQeXy/KKUNrFXU
3ZcfAY+RrWrf+aSO8tsnSWWI9oBpMKP2M4axqpHxRP5JLneyxo7aqu2Wa9Tc1lFL+d06U2hO8DNu
uB5QTETpZ/zJ1JflwjxRVcpQ0zbnypFlz8idKExqIlomHKSFl2aMlh+p2//+n8lmLfJ+0LqM91n6
OituBLv8oLM5IO2yvFe7enQsbA8oTCDzqy6bKwmoZmZDhdbtSkuY7q+32pXKqmAAK7JzITQj35q9
8d6ROsWrMKzBmICKVPpyBgK4fUS7q25AnXpHObuPY81Ew5SxJfKDo89wEVY5CsP5r1jPZ0zMYDhD
/pIZk6es+iCweC0ArzLQZIxArueLfu2tCozdmlEQF25Yafi9Jp4zd9uuOpdgHCh1xV4utIV4dKDO
HIuIvOQNywYJ1uoYlYlUI74bucdcrM0SjaiVjGzB1AZqT3peo4Q7MHUEGIOq5CFv1Tw1B/WlZRf2
l/xWLGe8GK7PdWItOeh/1OXTy+IZbp6lJIyigAMf8pT+isDPAwDFliqV3uxLGEeEU1IcIrh0/iUr
rNuK/znn/koJFFjbVlCADCVPObYNc7hutEFvKj/zwhdvPzTNgFjM2Qp6iVtEYa2rMdLE8BOdiDrM
6vKndPQ0ZZkJ2Kaz8DXxpsQcBql8eBDjPJBO2pQkKZDG4ZGFdJOEHjsXblgMtzqbTFRbQfhym2tU
Erct5fKpPyZ0rcYdp4tht8tZG9VURI4UwdhFymCN8t23iihF6ohFfsNUjWHUS7wQ/E6hwEf/hHk4
nj0O31K8tzXKxi0AYT+iAcTcK6RsJtALhUHzknjRadidlMYWMvJtnNqLzKkjO3v2CIY7NL4E1/Pz
iY3JVe+Obd1iwfmCV3sgZg68moP8Qh8GL/+5vnt+Iiu09CkRcy/1AIFZSehe0vSzXfJy60QSBdpU
8+TXcbBjSoA9hHbwEX56W4/YC9lcnv7bxSxhooyFhdf9eeR2ZTJUxrfNp9J6SehXKnER+lj2OAkC
dA3Y4cce02QiVgX21MKQ3bmbDKt5HNFVJhzr/Aeck68+tnrSrAXlL0MiVspH20UfP9BGdGPVqbNV
YluLYODkDODPo7UzClXB4w9K+9nrLZESjZlpVdNgdwJP7L27xDsjrOM8r1DmO/nQRr5iqLYQk0Gm
KccZDDCe8E9wFTA7toLRmahDFUmhAwIJxYG5QQ2EBKKuGOq/NPFIXqwONMNr1jzz16OZumOPyGFp
MtE09L4DF7v9JEZNmgE3ri7AzqRGJ0mYIjBaF2pVDbHVMu1LgtrpvdS8nh1bCuXdorFoBWQ/e0et
+lXqhvCDQzM1V0VDwtLnGwLFaFHVZMw+41N/4lLOnz07W9/VZLVBY+L3Ol+bxq9+oSgZDvQTjm7a
AqEI+Wu5VoH/ohwn3hdRj+uu8E18mUTOSOyiXxkjqghsa5KMyA22J1/VUhPeAPmm9oQ1zhu5U8WF
plyUiKLkCF5ijQSMAg15p8Hmzw5gyMcKIXn2tqnIEShib9CVxRW/FVQN4uk9SNNPrLwORcDkpMOp
ufZcY9vhQ3485gQ3B2P9JkxXjt0quyV8OmPKVH1j913ef4K3l7+82trMMEotXF/pLid4EdcnWUfL
2vKIDNNh//CTtEpv36V++gZTydC5QPWW8yeVUJUT9OPep9MuknXUbW74rfHHJnOl1vhuISeI+8i8
48ZfyoWCLmPF3/Mi1EeF8v2cmgYSbAG36Q5n/dVEGczUYlvjAGABIX1yu9u7R71qgJUTuIu0uc8S
5IxwtGSshMP0Jo1TILmib/72wySwIA44g6c/t6REflcUbo+cWl+aeimOaGWjPKDUOxX2LNbvr7V/
ywOVGsVR/ceyBl9rz28bng95/LWBZL33bR3Kef6Q/aS4OsbKYPdrHPWyRZFbRtf91FYBY83oc+Vp
BG8SRE+y6fjXmU2/vi1ZN6uXQeNY1dLCVjfQAOv5N89omrkmFHh5/Cf/XpUsw3FjUfdF7TzkYhY8
7Bwv9MP4s5J7FkdXfrk5AqXhyNgjfKeWVdy6yMCo52sWSzfTaEx8PjG2VbNuvyzb8fiF9qh3Q6R+
izo3aagO/xkkUfaVTayMsozLjAw2/O/g6aChHSOnf7BUPXYMyVBLFefvG1tW5J6pm2t3iDB+odvM
C2FMBT1QfA56F1thrtNCFe2sKchGKO96crH8WQO01C14Z04n2D9pHkn40FfNSWEmN2kt904SsT/w
KmgwYHVGyUimSNbmF6lzOeeMkQN3+esQ7G7P4NPul8GR3V6jkHqort7VvIsLqI6TyELkSRhIAfk/
zaf2f6N/vxdeIknAlLP+NxuZTGFp88c6r+qMx+6wOtFjLVqSM7dfZQfK1C9eJgm9f2lshNIDbzoM
F2xy1Fu6BimtZ+zI8XNzQKH/xgy2xR85lMNBJPf47bNIa/O3FHP77bCw/JRAFecXY6kPAOC/8DzT
VJvT9x3CExNkEeJ/qV9OMgeripVvp1eQyIEPrclBb8nyKJAVlKH/sIopwLweecAk/32iLdozUjwN
+wcxtYCdUK0Wy07L8bAl501mtfZCNddG5OwnDY78TgcD7uBdrsrhtSpzP/mikeULSTXWJlEhff/V
PPQdU1OgyZ/K4p7y53DLTxePax1Ys6BAuob7An1X/bXKiQGVJX5Se6SGM0KAz4ruMH8w8hzhBi9s
mbXl1kZq+72X0Y3rJyyvpfLf+xyg66EO1cs/+233MmVukyPCgKAsbx4ic9FoxyJZd4vFF/CxatNI
V/aB9jZnM9gvWZ36rmPkZzaKquTlStRRqBBi7UGLUFAUPXm5qgYNgMLHoxP1eGGAueDDCrioO0dO
7O/3CxYIPjSR8MHvjKS4mQ46OQBSNiE0NUHJlkK3c9MHdkHHimMKzdW2CUI1lqU12G8Lzx/bXuYf
9SOMzPjwY7UUxQb3JLGekhEtU4+XOPnI8ryRgwOmAZHT4ULdc0mTqqNAXIPFnG8dOXDkCPQUr9nV
Z69YdriN+SFltn/D8bO/h5kUczjJTEwh+FA/XoBrYzQXlVycn+fzvuQ2u4CSnf7E0vNWA5Mk344n
XxhyQBt1iX385E7/zpI+2m5T3kVQWntJ3cahueNeQNtXnvX+VKtUuZeo9IfiMcXfx0n1t+b3fuZC
3gNB6rsr3lMrzVQW2LdCb+PqDriTxSvLLZJ6qAOhaIHAFCik9Qggzsfu43vTjQP+NXQUj48KXzxf
mlBokc680n/Y2E6pXlC6B0cROfe06WiQ+O6FnoNa1+S7BXz5row0AywY8MEpT3wIJcO+ubl3HGMo
jKSc2HfspvxmTLeMEG8qtfqSzqaYtQlMXWvFe2IrhRVpMVzqcNguf8yQ1xTgyM7uLl6nmT+m2gRj
tXODL/iYlf2Cuh9LkXf+7XQFKwKjAoTdLthsPh1irv2nRgCpjyjqvShKLaNBhJe21gsSr6a9U0DJ
sZmnnHVu3BrhwmqXA56+aJDfD8hvl+05d3diu6ymrFYUuCRZCuput8aa4pjK/u3rG1qUo8vmxVSG
SBxgButyTYsS4aaQK5vl9kSRKrQFpiDIakOn1sWY1SMSF+uSrbEbBbJ0LmtEVlY/QjCiqwNziOWE
LLIJlw9l1gAN0RQQCvNoI4tY142W+F4Ke2nq2FS/z0NHEGDMn+cd4Pc5LKM6iQbvM5pKVYW9rZ9S
TBtP1vv/f273fPCNDS0jc08Fl6Ztlq9qosY2i98cdlKE2baUuwg7FO7m4cIXRaqNdLKIfzOdHoCI
kZRY7++pmXNOI/kI7zVx//6huRYbyRLaRF9KI2+yqmhNm3SUF6AECt5LkG+LjMucM7jRbv8g6wHq
J/jgJPUM+VRjo71AHv7rNixjGvMFLIotQ510yRIp/gc+hXuGZRvTDsOgXzlLPd1xk0yzJ7LdWX92
gMr9MCqfOFXINeoSTDjxgx7KqXS8sqriTQsoaDAuey5CTvWXUN0zf2JArkPxvQKmyPUGB6ghXuf5
q/lATytN8MVTGgYbjmWy0PYeAL5dIjdURPWseVpNVByFlYjMI3Ov95D6zINzXv9x/KX5p05d1duT
8WMys2gzk1UU3ynu1qRHLIpxFyr38nEfWCh8NetBdv/RUKAg4lTcersdMsWKVYJnMeRKIjwi+0Nu
g8g49cxk1os7HHbvjVxYftDwu4J+4tlc0+iYQJtuHnSCtWXzyjP6i3nGXx9mQfGu5A4ZOFK7as//
fj9Gf2ydmpzkQnGzXgtUz4vprFJ9NWXs+zoV25HpEP6gvSZu/Gun6MK1Plw43qNKzytDKywOrYD4
G4hMgX5pV7T5rUZzIwDyzqy79CFKUg98S4WvJEsVUKGSJY4frzgsO7OJLe4HqCW3PMbtepF+Q/Tq
NWJxVLYB4azuC0OZtN5F2jAFvXsdbcv2WODBi4jORt0nw1u2XaAgKGh11PlbK10KCuKkvrSftlev
Tk9vBKuCgTBmHyAcrEo47mdLG5mQ/ncB6P5n7AE+ttXtia0RvVTXKazwYZUDdUS6QH14+JfVgStE
Rj/tDx2x6QPD8nDpe6Egr4OtcDvB4P4fBHCILzVwzsgIWiCGuejWK7vBsxacepCsquDtjLXuHMKX
TLVQ7ay5AzINuNOTaoZUlmwJqlSrCeq3b0cM/at/NYmSOrr6u/YLmcLMoFK29ZxdmouD7k4XsCfS
lLyeUzN7moH3X8+J0ZWqWUqHI3po+xjDVrXvR8G6aFRt9guxzXxoHtYA+Q1fVnZDn/RadnkvHUpl
Yt4IjGGxwuslSU4+FDglObnmQkKcyzGKfcEnvZDe5mJWfjVHdhOxgvIR89O46IvieYtxoyt9e7F2
P0CIi6DrPPOXVBfyJvuYrO3R0T8wKN5NsN3kqLocHI4a5H0Zxw2KqUbNJVAJ06ekShPplHZVRXv+
A3bmAng/RpqU5zyfs+P2sWhCrrgwrJlIdAQHG3yrKTVfNIEK1TzTvw4jYA/Rg/lZ6+LCFjtis9fJ
Jj4Pe4qePwxuGEeIgk3IFwMMEM159NjZJ4ZgiwBr5RXa95WsgsRAnoUXEaQqMDk6Q/VQveoxLy4V
MiXz6B/AC+1NJRYuBnAJ4DQ1H1XIInKy40wIJzuKkR1H7jCyV2o2UfbsYvsP/isQ7ezCz+ptF++s
Vf2R+7udYFyAxUBbeN7s5J55octcblDhFu9XxHQXUaClhzJinT2uMCYSjSzvpqpCRp0eCmjvDZ04
s9AzuyOTssNj4iGENrNITikPd5Q5Npg+5km/VyD3rLUOP/9mXZeLH0kRJ/HvtT8tuYI2EqSaigAi
4u73bmitQsPBAZaVQKgc87xhTIa6qUGY/HC5P30ccYs4YAONhSkL8HhASe7ty4c8sPWOp2Y0DAue
dERCMPWKRI+lKokANAVWxgmXgRzTbh6W0wjp98XaZ3lOQgypBpnbDHyfoQIRoYZuvM8lIjlis1FI
/mBBdd1U52Hxu4B0DwP/i45wHWhSwLCM64yEY76ATMXzCFdwRCdn7fkthszVBme2jCy3h/hHxwkT
grEflouJyJylm/iuF03x/2A0d8Kz6TJk+OORM2AL9+VF9HhLpLZnk6DkTWrT5hVlwCovPAv0/oxg
OUQO0unjP3IeWLGFS2AvBZ9WXHIKyeERnb+4+XJY17HKd81PPNcHQOQIdizzNZFL4LwcAMo+sMWv
tXLQBecpbCb5exzL6wVbT9uMO7K2s1U2spgoF3wMW5RcjB1Va/CcIw6lWGUjhLG4VuEa77E1l2+M
UhfS8/gBAyUNwvApz7tgm9KK4HTO5snCQy8P/SnyZUinpGe73z04cug7iWYlMwIS4wzL8vFBd178
bVdcyqQ7gOHKhmgNxM4L1lgSxrFlaoRdlIWj8UAZX2zHCHLPj6Hy1d00FHSF/T45cZ91Yv9cSEdS
tf8RGwAQge8NGRHPv7yNhMCIqic9qjai0R5oyj+admiEmefAxy3l60nZHTINPpr7nZfTgD+DLUhH
t+83FG/wT0jJWMYlrRvKy4qIo7cpC9o8nWiE14s5vBDh+LAyvxirTCBLU4bKHOyaX8BNWKo5RVlS
lFkqUW39yyig4cm18AETxTHtqAYtcje5n5M88cAovmc16L9K1qKeOxERkdpFrD7GaY85+edqMM7l
DriEW4IsQfoI9j1A7W5Lk3cHHiM5Rc/iYGdFEJhRF1Ldb0HzJ4HJgGL9fNF+muF+5GapBN20YDmv
/zUAn5YdwXTx55g4JWezOgHpEM4sZylkKZ9O2xhAIrt64vZwFxQYmy1W2F3A9SojA57m+LgPup78
9a9xvZ5zFyM2tqH1VfvwbLMnA+H8HDdBDHTm1VQG4z8kVfrD2b7b3y+frQwVUlfrAr4nWu+9zAMG
aLBzaOoB7lV35Pj56TLUh8G3x50N6oHfyu0/RMfUXY42F09W5TT/xQT6z6CdV0qm/IENz9q0/nQ+
WH1xrJxeDL+KGQhWpFc2FR3WnWqeCkQVgnZfpmH8yHYLdpHH85/tY5CKYywPzsr0m121x9Q6j49D
ReGUHIKSMXKh5D8HBF5y1XYDLRkJIXlZODvsKcW/6OMwv4lEF0qiGPE7bDxXtKiQDCmCIvpO8jh8
5W4/e2kXdJotxJMSg4h1tCf1CYEJ1rJ3cWEV9mf5ag6s+Z0oFwDQqMVExfNZr5aoodJn1oJ7cqCb
n2XY3vlhOarZ/f1w008FxiqZVorSuRDiShlXXLJfIo2rd8h51Jpy0f5ddYIw+dW8oSlUvjIQUggf
l17ULrjJKQPyoZxDEz4g8JJuOnhQ4a//qPuRuKNAoPsx5zqD87DtlQ8+Hm6LLFU+TV9TL49jJ5th
6pGQNA7GSrm0wpNo1BwH/0n9Me/2AEJhuah/gZg2m3r2t7u8F1VscyiVYiQB8B1ub2N4lpIFfss6
A8PRYYTQgpPEqv2is121ci39sgJHrMhr7QqHXDHcO1RTo7DdsyHtBONXjjqTPpL78gaiyFS+kknJ
zirJGXBqrbEZbvWHYwmkmBCFD5yS60bPLy4JRqgeeLWxuly0eTbJ/CaURoCwHTjFY+ZU4mTeyICD
nTnNFTCn/d5U8O0I7uV6AZ4A6Iexat7IdwJhnKM0GOPHuRZM3O71d7KRSBAIpGCdjyzjreXBD3xQ
86GXyD9NNfU9W6o4d1Og9HaMxtIe/YG5aBVBTsXYl00ZqgDAYhCJ0+22QH0twQTx6r6/tLq8Ywfc
r6ZdCgzHi4R/sKnVpmL0NjJvcpQIe1lmQHwExEI8lpP6F5ckjycXTEKxj5+MPJO34+2N8jr+BqsZ
fubqih4J4VXjqREZYEiLHxneGsiMeXFY8Fj4W6AVxB/JiG//SNUyyFIaj7spfmjJb2KSCvEQsVNV
47+TCZwlPK7aJKAAoPjXWbsZgSni9tKI38rlJKfPN88bvPWA9NT2Zy5DJcyDZ6Fe0QpFkcEUwuif
XorC/Yax/l1kWomJIc0XUvKOAEj33kW9u42my+8XhdJLOb2aqV74Gg2y3ROlpdOPVs+dUE/fxAfZ
5co84d4WfsSwxjHcyAZPiw9nD+PD+rPKFD1jXOzsckjyC89PlZ6/qQ1z1tXQU0bc9KILr33jKbej
utxmwYKEGWJKnClLWyUwH4AzSY03mg+hYZfMujjfqRQuIs1twl3hbq+W5UJ49H8JhgsSnYS38P30
kS0MbEiwnC0QJaJtKPy/jhbBWVrkwwNKk1xbjE8IKl5rokLYrmVzRFz5+hXgJ9M+dextM6rfIb5n
ATbLNeHUW7JS3zaNjNWEgsDxJp/eX3MT5jCjnE3Y5AXvJu+CX0nGkbxW6Xe5QuwvEFhYlhP2U1rt
PylI0V2Jg89mrsIraRdBiDkSwIYCcXsd0oMVmQv/eXbYzFJCwgPdZMd1xIWpnFpfJu6wb7u7OTR6
SlGz/vv5W5aN2yR7Gb+QFH7ckRrs9+hUkYm9jB9WcY20y8ZKNPS3fTU+ShQOCFi3lWOcWdd5NSX3
zZFvI76N3nTP0QnkRHG9MwtU9B1TIXYndaI7Z4p2OGqqdJoM8q2Bd4q4IBs8UHRMK0a3PHWSyQIR
EmCEhmrZvCU9DuQaxCneGghj/BLMwSuEvTaaslUU2pyoWlIQRfaut3G4wzRJdUGdQ1zGGGlP+38X
jmW6U9IKRLsVLAc0fgJAyVKrCkwNe/b/IVdiJ8oRJnzqrGbIRusKRFlR2+DXuGBBpwAxwuohRG7r
VwyHALP/ZqUIehiMfcc8JfFKTvedWniTyAQKTY65dfB44w35lad4FmSrkK47bcAmCs4dGQ5aatFF
Xnal0+8dNgVa7h92actitGGIZnPRfAYBlGoHA9wjJPvMIdlzFvykVg6/YdERxtRCxJ+bdcvwxv0e
LZHqBkTbziKROtxmN7HEZVOXlu85qwfioglBf1Qsimd0xuJstYnDG8tIhhyVBdEK+LaN4NuGUTsf
d7nzE20QsEVb1KPUokABTr1uYlxlzIBW8MuYWIS4iT1BHpv01g9VnOm8pMPpdlTlXIuUZB5GOeZA
ibqPpfPKtBF8a21ku0PIEoVIBSwkSJNBeLR3K9uyLHrYZxCr+gZgcIXXiFe1vNz4ZDGwnrsIGP5w
HU8UUz2aGYC8gO8dNQR/hUCy7kHSRdxGiHE0LF6qItFE50xzAkahTU1PGXr8k/n+MYr1YHtV3plc
uxS0KdYy+S532hlXQlTeSPpKevb75MkIQgcqwPYVhv7oL5UIvSh7nEbcl/Yu4TyG8Pwh4QGxuT9J
d95xQxmAN7ZDI+YVbJqjGHGa6nmVVOs/xNB2xL3jz6A3coFAgFdmF7rgd3BrnlCrAfFnLXCYtf06
HODvpc0RDQWW8ck1qGKSdPHo8XQgAvIttbNv7RJRVstitZPATEfzoxZ5XWmWQS50M7qA0CjWwqwg
8sq5a3HtneHW/kgfROn1FkJ2f1ZOmPk+xRd9uRJ8hBjeBPC/LyXq4yYt6zaQVHrM78PCXzrP00x+
7wFqUQuo/pg8SohxCRq0BNjnAC8Ad4PSI74XfNewxQYBpMK9UmywVSb88QJ0U0W9AElWtUbORDq2
LwRbbagFKRvTaF91Z0erQHRXVIURlpw9k4W2JqnhgHaKob5Euu+NsHOVKCmHTkgfZpmHmx/XpFtb
7tN00Sl7D2/YLjyErkoZ+eduyzOsa4Rj+wqXYBrmNS7ZIzWpUpKG3mSkyYXehm9flXBEE6CieSZG
b8bnuH3lK5QNKYqr1dqePBhPkeyEV2A38L4qlaT4elgGnwLuHadRDnAol03Oi4j+eL5/nXMqyToX
KObvXwtJnkDJWhrXaVyzZ/f2/Qn3YLGhOdPbG88bjbJInOdZ5OAMHHQrTVTWcjAeUmYiFmOeCpHi
v6mpJ0xb8Oayu10tpIJhoAaGppDn2+DzIEAVd91Y8OHaM1ALGkA2GyaNGkep8bBn1VOo+Q2Eew37
l5rC6afRpVoi0H+g+dzZh+83u9usfnewLQn/9rLR4GcKGXJSNUbxER/xjJh4K3BSECHKFYSvN1Ac
23qRYN272tW7fORfUF1TuOagdcB1hoTQP+c0v7c+rNL6kZ9h+RbLCnszYAZ2vqwrs9ma5bLVFh8L
RQZYjETkMrP7yBe4F9se/3UThW1MDUgJcsuw+L2xaFCOLm/3ZgFJxrj3JzZECUoNRHUGLxHfs0OD
t6d0I5Tete7rwVv3YpPSMEhBvdy9tIyE2GuqXVTv6JojBdfeL2qx9EKudh9/8wIY6ayY2He4eqgH
S5UPWypCXVMugfuzKRLCnoIMtaN4a2c/iDwQDwGFZKb1Q21b98VItKKV7ssJ3ltgW1tQKAjPRdTP
8VGusiqLxs5rA0Lt+vOvAZiEhzcwiLgQQFH2w2Az60+umkLOcp6eIQJa/447leslbwyGx9AdAVTL
klDDnmaW/lvhTznDqneHdR5ER78/n9D9/Xtmoodw4fRdZJuqKkKJQSmayyISsg+OX3j6UqisdxVb
yOGbakVyh9seK+mOAr1b1YBS+iTOtKCHGZhciaovlHzfCgSBlzZ3tXfHkKiDhhH3XueOeYx/Gy8c
tqgX/BSWF2S/ZQWsrjI6AIqPeec06yFjRYeMvhJ5cmMNJU2qZPa0eG12z5MflMvc1zAwMaUo4zxY
Ro5QtHQro3wc47tHaxkFbx5efxjEHGrzN6ivoBzuiDvgT77vzcYsHlzmtxEr+vF9PZXZkj5rSO/s
zp5SE8vY9xFqQGEwkra0LlIcvzUJG1Lpis7UdHE605HlGwpxvYWDV23VKVD0Do2SNQIeoCW9asDM
xfokXyivGe+9jIgSeG86ObA4oMBJ61iaO5/uTX7FKa4ifOaWrHgEOT3alDtu8hkVEEeMx+hxXePO
//1xXuE3c237N5705QegmRP9pd5JtsIonr+yjUPIGiPGvsbGOMTQsPWc0H9D4O7R54CnSNps474G
3vAXaGUIRX73Eot/GKojOFiN71SBafVZFwOro9Rt/2i1DKwi16j2WVGJHoJleR6m++Mfn7IibYmP
sOFanjt+FU2a8v52mRLj4uLkko17+Y5cT6JvNlSSJlfQpN2+e+TU1utK4LyymPykRWYUGazD+qRf
TJcj6twdXLvt2y6BBxHh65Ouutf07tTmcdi+v1nfYBxGk9Od8JA6ENaDLl45U2kLoN5Lmlf9DfQv
AP6UgrOkY58TfvpP+7hh8wo/8G4f/G8pcjFJxXOOgvSUstfdhFtNLtAZIgC5BgUKD3vPTh6NJnbP
bg/NuzM+xXDJpBlQ6ZEi7mRqGDeWQ65AXcq4hhpmI1Umqa140n2VcbT+DTNAo7SQ+4GTBOptvf3q
hriMGejW/N5q7UH4ePvE/vt1J760sLvX4WGxtUMnud85OUpaSP+tdD9V0jrqlBMYie8VG2RFKNPO
MmDkKEqGygTFR0DYmarLSn4jLuXR6m4WJ7wd8qYRjT+3xErCAac/fdWGGGjTQu0RvoT+DVrN8/th
4AdJ8iveeXEXhMEKKUxkdCwyN/2GcTEviuqO2TG4d0k3K+BhS8X5QOzKoDxOYU6norx9C2evYi2M
pA3O95/q70UivMqdCNTcbnIHvDh/D97BGUBXrdTdx1jZ25bmdLxPBuqwkvyXNSVepxojpSMmhj+Y
DxQjZxGIUIUCFwyKUI9FpPwy69lLZBh4ZeQRXHz8G8jpbjXzPTqjE+e/72h53i10RRHpq3FzhRpp
dZwmDjQdsvLdOPnpP84IWsZvIXny3LcrwHUylnb6eUyGomJbRtnV/nVTcTiEjHsg2oi0oNDv3uUv
Vet+ym0fhss8PLHiiGqNx9207muDotU/r5Ct968cJkdpfs3gG+CwS93x0MlvKyuvcsUwE0CAo3Aj
oUY4D+QesvtvlSUVg2KLzWgOD489whySNdpHyDpmhvFKKjb0nU7DQihq/etzsR/LyQpGX2ya2qSJ
/NDOI2NueUP1o4I8XGM54wJs6/gHCwNQOM6roioZvBxIaBLUftGb7yzFPoiCIv5ocbX/z2c0juon
ToqdXm8/m5CLoy4DO4mHG2lfOo4FPGlLqTDE3cqTfFlQY6ae7xLajG3ogC9OE6PU41r9XnKMrWRA
cdtw+Rbh3XTaukNM1Y2ie1WWwbDP0paQrdFGqT00b38GpfqdwVpnjkfBT1kHdBKH68Uk4+itaae6
TRN1NbZJbhv1RMvcceOmN28w/AZj4P3/CPaZJ0LUvryIfxwPPX4X4Of/1r+89heyQyA7ww9iFm2u
daJ9VRyf/dt9g9KSJ9rZF65KKCtp0NWc7MFujg/k1O+dAT+FPh3fLp8IYdwEBBSubHrSa9pOT3Y2
FRR7JcWPrlmq2WKhvxioj6G3yUjZ1h5thh3+mdLELtSivuS3kUj/sVZ9bIPpmmYn919VflK0NRpC
wIUr94JQdkRSaKk9Msor8iRtQPteriepAm8Js+m3sWFnNoM55/PEDXqNoZDe1S1bvhsz+eainDbN
xgUnbQ9iaPaiHI6CcCvCaIqqo0tj1NNKL8s6jTkOEJzWGH6POgeK5UuS/TVTgAfmti6+0aRjR29c
UytovaKxRmxkcQpsM+RIctbmlYP4HB0VDuGJ+tAID+q+cDk8bwo89c9JVZG5vz20ULybTPOb632I
Yi/NXgAdPRUkWSi9NYow4LgT99FGsWS9JU5UKJQ9STqQNgzlm7iag6QxRKcih5qit5uBUrENbuR2
L0DBkXK3sqMMieUbH+EqC340Ge2nCeOPj5/UIESXDnAlq9HTO92mp6OjQn00vw1sR+udk92dYJTb
rZ82IYiEehC7csBX7feyirpZi9XUCPBxFVyS0eX6qFgkGHVx39liKwSrdKPvOMAChxrRh58QPQMJ
gCKJRCjvAKRFAz2ThnOt4v/pUSffQ2/tjVgtj1yeGRzqWGYBrlYlBNtvIz39jJuigGZzi96ht+9G
8tepNVG+wDvPgHCkkzcbUU0rtDl0gctmlMKh4B1N6qtz9+dxMV7VwcGjF5uLE36xuB3YXsg9+rCy
He+e13/7Lp+6nXFQJqGfsWoVBOrcEtlFHv15Lf7FvVBhAyPyk/XDcmDsqDo8MZn360k5KEc8fmGr
ZMbtPezFhp+nj2ZnU44xG013l82ALQyRj6hqhvc5aJTLcYIAA0gcIqcI4P/yA6FHku9YFo63byV8
M2h4BWMYCCnu1XVbSzQ02pE+SSXTQDi1/X7/ViKpQyYkaciw+/vNZ1in3QeXQ0l4kW6LGVeqp5ya
HndvVd9bwQZ1tblpR6N8x3XXIU3QpBsj4/iSU5Se5LhuXEJOYtWCGjL071vyC8EIseFJjUJz62Rk
C5a1nKSOU0aE7mtbNk6ruILLu6sP6dUPYT7Zx5ZLF1ipfJfy01NWg+NX4C5vYNshoIiRPZWgGxVy
9RaJOScUot7+QxXBJaG9OYw1g5r+2X07KPbaFOiKoHBNXtuzpG2+8rAfXleHA7SZh8s5LXsItvRc
oqvw0fWr3tKdnvhIDbZRjQ293LRNdBDmRCzv/EdqSSXHZTJVxyBq8N+vbYT/b+JtfZ2Pa9tIOu93
De/exVe/ToukvVuuBG/zWyA8hjGCbD09GIpfeasfPV/yHPlyQ9Vc0BvhzzPV651BurFHnu6Q/0Wq
OsDBtcQDhm2hjFJ/wrPoNUEAmg2138Xtp4ou6EHrbJTzUBdRHisvcY6XQe6WI6WjBrGz8kXjMHVq
modXB6g2/LMz1JdjuQBUNQ24M6PTd+WvnLGXfwqrIw43RNqK0dB5IcGgDv3RZ7FuT6g0FW4DHrzd
1G0x/TPMPvc9cH9ckI18UBaf+r58P4b9nsCPuA4Km2erLKshJVxoo9w+rmW/Z81Df+sli1J55Hqb
AWcMZLPyUDpQJVAJGUQds5fNaHKUQGtNzrJo4wip6UtkQAsDflPthTWV7jMOpa3oD2CV0mJR78kL
6hk36egZ6qfDRH1SjTrrDJd+uW/mN2lOX1dAR9pnbMn+qo5bYnLmeCVVv4+ZsDrGooe5VZ7IwDkr
JNkPzMlvBi9IRhlfWHpr5MeGhRhWMaNQWU54Bn6mXTdun7sZSKtMqQ0K3jFMJCPDNZCF6Pyou9U4
nZKaN0h1djPbAUjPF/wSuznq8bAjjsRxFCM1YRf4ur9WmFCBev7n1ppmNSNcvFFWJ3Qgyo+kH9xp
big0s//aOdFvLxhPh1CwDWIUq62aX0LpXJjr/KpCRXwSyDwdWnUtHtrxMFfKdpP9bFjp2DO/L+cD
LE0iypTgUskh7e5z4FA/YjKz1U9z8RG1g8U6j1YYYALZ1nhxje6E3sV3P27RsEhQdVm054GXbmHW
dhe7wcvcHKiMsRZVG4OXpNBClnfM2Fvgv1oUHKxyoaPKxdKIgNHn0RMvBgpwLaOYjZSdrOtDRKF2
McCbFTbs2rMGnUotaLQoYogB9CgRdAHNmjvm22qZ2jgWJw1S3NGNRCSGHA0qZSSKBKVejF0Moj6A
H4EymVKhuxg1VPDWQqxcKHM9dZDD2EiHdNrNdzaY7E0p/EnFzHAah7CUfVdVM7HJxPlsYpxBMav0
MiA13Pf8iz8H/mNv1nYtZIxvb44yPXNn6Zg56ZTDo+vohKB4p5p/9wb4QCJqy8Aa1Vd87cGYhbV5
hKz5JxamtNJskResVSHMAeSYU3906TfFe5YGrXf6aX0CEN/+TRk64heQF7TSBL7nyNakwZJfLRDv
yNblPb9U9iiJhqv2vVNh07P3eypavEsIC01Kuf2uYUtZq6EZYq+pBEGn8lSp7O8kIO0oBR4d+UHH
W3nxWX22tXFmYxUHd0lJt3dv9wTpXdX9jOvURmJDVQKC+LLe/TGUN8Y1IpWqeOOHgYJskrGkJ+g0
sG5AU4rTokVcrq2nNqlZxsTEp+/pZTXwPGbE4CML4GOE0PsPqUlKwizhgfQ1H3stB57ZqIlkRkIo
UvoIInIVHLZ173aDcALSqU8Aqf8COzkXUX1I55E00o/nYIHXoY6E8BdufC7wvO96z28X34kDy5tq
mdjRNu9/jWo7m5JpYyO9vjeGKtW1yOa4lv3++GVRnpU2TavFoUisdYXv5vTo4czSncTFZ6KQo28/
CLnyodWZMYOEaV5JdN4avOFGBRGYBB+K0FN37Rq9fSRHoK0AV5dEJrXxMUeioxxDNCgKT1eh/1aN
TklDiIRjadQjnV85l+lSIh4Sgs1AAmEmFv5gRVcLI6LShY1rO9mmhZjARVYItEkjQJNBieAcahzi
vV1gB4lqlYwHpP/gofuk3SAYxi1/WwvLHGYNxIRmJ/T2Dhm5ss0h2k8zGcMMIX1WY0Wc8xzValHq
d/SXkN6BA0wzAsXIHWXWNIGyAocvaTn0IDdSV0aGY/IRhJmCgdrl7JZbqWWZp8MjJgnsoRj6nPXy
bdxrq2305S7HTrp4mZ3VEhKS+gkMdLZN+SfYFi3LIqrRX9jM+y6R2zS6N1B+nDzrftmOmmasR/6S
Ov8Wkw2kviAOFNkEpuO/t7ntXoGPeZxPBAASSmAxSwwZysMtI/fCBvOKo6prfSq/o3rCYubKSbi1
uSvjxf+fHDOxaeDEJS1vrzjwbI+7tLeZGwvtuXyKWZGrRPXLC4KrecfVilL2TVtEp5NdaZeTXRnT
U6YBcNmAcRqi51dv2x1GzRCMi65yNjp6zOm1wKsKuDiHJqNFtCQ0bPAA+xCnPNWdVoxBXivVmKYr
mdod9hDLJjVcbN2uzH0NYziRpPdCI23r9P1WQbrwfe4cDx8jW4w1+XblQViIw4LPbK81sIExL4Ed
p+4KgCw9DDrPtu8kjKqakicHbTfEoR0BLdX6DKHmhGMbaD4IcHcTCjpRm0o6BcpJTNl0/UsZLfEk
gla8zvkOBzKMQ2/eWBb0XUa86u2nunSYOOC+94msw6AL+QnJEfv2spjesQyDa9DvgVPVH4EtwmPN
BmaeTRnS7ldWCZsBZqSi5Xnr1xq9rcjIHLwQCo0VyY4jb2Xhw0KvKHYOm3Ep7N5b/em53wjdwj+u
6c9c/15HLnvqSPqtne/lADLQbvOu+COU++Jz+5hZ7IR6Ewzi5WakafLWclROEbMYrfn1XEOJL9Fa
M2GQLBGKQcLwcxgyiqRy3aZ6aZv2DoTeBW9id32PJbDhAvuSfiol4M4feeu+cMU+SS98Vkg+zLEi
wyBUOWRym3ZfECbYtW3qDJjdv0kOnfOLkNkCN4iFeNzVruv4O0+FUa0ltff96BVhp5U0gOvt84p+
endgozyLBjALzTLeJRi9BNajrazGFJ0kIk4ZfFQH9Igp+xgjRZrV51tgNcKbH/iH91t9UqKVCPgo
RO509IU+yW9tcPpi/DsLizMrmgP1Nr3QPsb/1NmRK6gikwb+m+e2BLotAfY1aRD+MazXPWCiIINL
1CxjKFqLkBJ1rkUNgTWOPMNowwq53lvaZIkPMxpqnQ7L8PanZL4i0I9NVL/RXgIVQc8zu8lJGmhx
h1Fw5ruE5fVlCFBY4kUKuy0TySqwfsSqDJ/7SXhHx/vaTs6QQN3N46t8OX6QKLqrv27IYPteO3Fo
f6EBxpx90tl7bwlWT4GvYIekELZELZoPmc+xO2K6u5ByWMSeq3faDR166WyICfKDCjTDFyikpdyr
Tzharyr5VQ3ZJeYuFrWyjSKUWfefggpPB0gPYalMaPIerq+6EAK83aevw5ZToTVix/CN2pNV4VY5
KUqGtMlfgrlnmopIAKwx+BkG5eDz1U82Z3udMOu7Lz5J8dgCn6SKionhUZVNRzKjJ5ws22uFu47m
Q8EWBGy61Qi5C/KAAk4StKb5tjK/vl7XDu0KqL+l5WyGhT6FPkULfzHGYc7GCwnrd0WytXuLL0bd
hjJa6LILZmkhb0Gp7LUxa9DOwYycarxb8myNt/hDz3xHg7gjmhk1RWpwVLUpUaPBcoCAvMJJ4exS
A82yFPWb9IAC5hLBxWiZ4PKQdau0ze4D4gFzfAZttorlikvR0wKVyo8Z63rDqW6Np7hp6J1V+fsd
X6gLcPs5n/B7XBQvJ9qsU0C9qnJzIuwSQ7cAv2wPVfP8vwKsm1xIOpyMt9A6gXmszVfwFF8h9O1a
wY3L6iQNV75fsyzuF3iM5nuIkBXbPFyTrRI2f2f2hRoAWX1e8Df19DLcmF/zEDxtZ3wmNbDPZBrP
VH6T8oriNTvGA4jx2BI0Bj40GfG2z8texsjzXgFTNRXQexCRxb/iE/ZFU5e04LNoPlgmZLlT2NUV
nAGMhY1ub21MpGmPQCbaMsY19YfUiSX1Fakk8G7XakAG/X1t2W7mPbxvVfBY8x8fGXJlmyKtstcY
qED2b3T9ZxIKDVgwpZhUE1Z6UAjDXe/n82Xh9xPk9YZRENTKMANdqCCy4srSPSOOuADQaq00gBE7
GMdHpznMgnIsuFpQXmYUSMDSpEg0+JKm9Duh7bAey/eCX2pqiBpbs4CkbROXlUKjQHb6c7yoUe8u
olzdCRMblIHRxSeWy5yylJoX2n9bEXoUeBc2Htm4UO5ZjpOOcnbK9UsRU/Xou8V0DNzX+xRxQiFq
TNaWn9QQsVqjcCcjxkRz0FCm73nddcLE0uytqQeC4AnlSExEXrUeqJIsu72BmaL2RFdV4UvcF/LM
EKBn4+dqIvuzRH6YBHAguUsrYXakvnDYAIH5AcxHI0oCC9dUaVaMcuyQS1RnvUqnGfEkyCiGUIEQ
5bSF6vj8CFOfpBgx4yHzWRk6wp2AnCHyqtYqSKSsGqYySF+XxuwEVQoQSBkB9xqAELZ7pCbnXnuZ
qeURkyQnFPhJ5NHJDRHnsV/eh5UU+e9k0te2E12z9f8jj6Jv4gs76u1JL8esylcN32mvkD/PNGkK
mDXvfHqk1CI68H7+lqlP9boOkQbDdkeIdt2TW23JckdHTaiJF2+nTN/IjQrEJnseOyMMyw6A582a
fSPYhaLFZF33/jfDsINUvozGCenE5/4eb6cpPfeu0PlxOJSG4l9cPMxNRteYJI2fieaWzdEn/hA1
XOgiPC+SBa7LpqkY9sUqY3YYr1TNFi7oaTeX+IygMo3A1oFrurn5So5irMuizTlkxtN+to3D3RMk
5L/4Xq15x3iZUeZe8Q7hll11h2B3jm9ObiCm+EmcxKE1ib9mF5uhOTL+DUhMrCYGDHKyagOb2/yM
MZlp33+9LN78Ufck+6rlkmwqGefxTgEkMAuguUChTJRLi3LiYQreEp2ehBAwIFkjBCMyAm+fjJ7J
5CtMiM1Kgl6etV8w/GPG7JkgjiowC9mp+wXT+RbK2lgPVToNmCX9uF2/hCcs9oB3xvNhtLaUHzBO
xeG2G7p3vYAcpbf+n6bMLnjFlRid5nsFSVqk/VNBY/edJm3+DiseMyb8kej+RNCRbV/7E0Jxe61H
EywjQFRyMELO8SuD/5nnXUe1/C7FmzRnY3Y9csvffh+MMgUUZv676KEEO0NmHfJLRwXwmKWpt9GJ
T14EUQCe+zjZ6AEM/m2XWU6YUwHCWygsKLSo0KxEhEvVoLbIVM3WS2JPG27sen+9zxmBtLShjUnO
Gm4ZIO/oTBrSMTnGUSFaB7dKLebL7FRB3CvynjsyRPXIphP/rd9423Q+LQaLNw+F8wN6eJtU5K0S
zAvgG0/zfhrRz+6/fmByEfTIKL+jTOwE9CYn/oxAPVorlSSgtieAL9Yb3OMvSX81fyGGUPVnzB0a
vyl1qm+kO2jTs7bTrDXvkm7A/Xmykbpa0eNBhJrMO+sfkrEZNSU593frBuGuzhOkqFXLfme/Qs+r
Tn1mo7j8InwPTPbUYOgDWLXrNoONq0AAdrQcB4Z27zPVOnGHd02xcbTXp1PXQYOzJMpb6XKPN1C0
nUu746FSCy5ONQoo0Q6b9Ygs+WTyh/n26Sc0dIhyRUzPjg2JWSOCCAlIDAtxHRVp1/opV27eV3yW
kHcRZ+ETs12fF1NhvktQuKClMJqbhFjQKpvRqfDDH5kFNfsnEIhXeM48RYLh6gDc0T8qIU3e6rNc
/mnLU8DXj1JR1oXVQ5jucMCVixNhJcSmuZ6TPmKy9DwawGTBBsDmoeS74l4xiFltK8jPLdFsTk1+
iksVSuYyoZTkkna44DG0DRBhHWSpFAOT0R2z+4GYfjNW4RD4ZGDHGJcMj2pDJUOF0ROfPWkZw8kO
J5y9DraL5e5GwMzE0l4URy/DxTXtwAB6UB2bJJ0Du+Y/OySU6ymz8IaaH5Tk5de3dY/eJLYKfKdn
RhMe+aCdjc6Ix64B4T6QSLGe8vaOQEBiUX4HVuXg/lYaQnXbHL3JMbwqc2ulksPqVX5n5HjqUbUZ
TO5SlAfiEip0KYFuimiQu5cOU3dcAv9PjSo+UPtU93mn8our1s3KLPsoO0PL02pBTmvlYLcH+pGy
i8OsHTjt+3vss+xdOrwh6tt3AjoVPFwtARDrsgOLsUUHaduGylj2BNYnXxWXMJzJQrRCeqFf2/In
oCJFYx2FONYWtFBs/9/1kn64zZXkwTGTJhpNazVDZrl+EVRrfzuG8y+XoESzvgfN7uNvHBlItDcF
Ct3/tQCK4BKbgPZeXrpsXNtO0XMj5sFD5YhJwm7zdLs0GUAAM8UH/1j1mj4r3zeIVwik+xNGVcVW
+FXClgfGDkKSXUSCg94GVW6FBk5lsEQ28CXbIadFZ2rgD86sN/ivK29HDy+FMNW2796CvQsEgmbC
RA1fK61yb9v7PXEQonlIZlP1ZTRFKtE8ODk1UhC9ZG5/r16vV7fPzkqLwG4lBsisDaqlKatL4H5h
79HWXE7N7vpamJlPDHmUa50+pVIYtxugHQDjobf340t72lL8glHEZObdBGoecfRD291bm/IFQips
l0eWM+JY7cwUolKrh2+UAwY+uHsH6ZX/sM+Uq812VlrwfneTlnf6iA6XnwvuBKEinfTmWvtbJXLI
rxY0v/h69mRYNMzgpt3/XYR3v1T3+DNOphtJV4lXK3eIA2UT5IhF0TIiBM9r+npRVdkVzmvYdOcA
wCvdGbSclFkcZFSZaTQerrQUqJfce0yFLR28UAGjKHv1E2egCZYwK54mqnJt1sd066LYe8UyDzWx
T7HaHiatikgaP/FbhCnZ0HZvdc6uNHniToLa0Zdn8P06tqtBcMQJUYoN+cQO3ajp6S6hu/1P3z6z
5k0YfUqx62KgeVwpQQT1DvE4yvoWp72JNEZiB9umci/nmPC0qxYLxen9G4nWpjNMAJNg+7tXVi3k
M84E5Xo64ABbtUgnL7otyseSXo+H5JNqmFj+JQew9lffTmujzrtGme+GHphrXDtSWSZBf3dX7nHU
6YXHjR/q5D5aEYjP5GtG02EZPv7r7eBqV3cuHn9bVATCKssE83BqTXHi5NXfDyvbo6XwS8L2PfJe
QLPnld3NVgwHlqq2VaI81jNfwA+Bx2bTzGXVp15evCndO3Bjbz3u8iwOHkF8jyRFWczlEa0Ner7j
Nrb9x7tUcpu53rIj35xzs7i/+AhC90VxULarGYl6Ddt+ahVMXj8NPjxozR8ToIYibmPe/wXU3xya
T69INsGb4QmziPuPOhIaRr7lokfi8ehVNZArxoM+R0eqq9U03TSeThXxom003DFo3tA3UJ9sBzbF
2fJlNVAjL895/20RyV80EyjzKh1w+b/5TIuTETXdbjAMBTvC/hFkBKeYWC6FpVpPjiQu4Y8xaj27
CFyY4RtFUS463jRu1fiNrH5IAzoIaKIctWnm0M2bix03WmWBCt4uwWbBxB2r+YXa9dcyaKlt0bGL
xxCkuAsT0C6hISN8GUK5issPXZeilLG+zzv2OLfsUhLZXHX7NJe0VjBRTZoLOEitxRmrwmx/kbKR
d8/E/VHph/zlhkfU7BzgmOeqEXNWLtX2l7qx0Yo8YS989FxP6us7qIGVX+bczhk4EKO2814oMfif
AcPsur4wqyBAfVlncG4lwCTYJgesXLVryUURJtJAYPEPG9UVHaHego1lWFzkeYQFNeAmFJhoSyg1
8BSRhVewK0Kbes00x5flnNSHnf4doYt/xnviwKCOyQnOdGKGmqiykk09N6F4E8nQCmXgkuPT3ter
SCCpRCc33uFyiysrq7MlQPJTlswOx3E38j6/hciQOThupOVSFssw/lZfR4uiIz2553+6K2RbQIkm
jnTEvufYCDsHs3NIEpafmDZ1ljyxEQ8njiKRJZid5HnUCrBiKgkVbPwB2PzettAyI8+hAlaLXNvp
/NZAWrl1dnVt9L7dsM2g5cQIiMfiBgvJNlSz1PZUvv06x6BPTPd+C22AhQmfuBc8XD3Zjh0hg6RH
mYjh0CWgB+RfzKwCO5rCRD0xs7llqHCRtfpBPfkXNEzSL5e6CYZfR7pwRK4se0NNwSK0wAh3h76F
5yJ1Y9SsyZuMTU85AS+4ygGmjbrIs+NnxysNWkSi8lNCTB4pumhAVBUoxUGSF3qDf+kj4DlLGxaq
QjFMZDOLQHA9PV0/4SpzX/kCs3wWNnROT5WCdkuV/o9URxTNmspD/H1sa4eyNCw33wThkkhzr4X/
3klmsQIk4o8DbI18m3hmA5rTDmuX0pVO+6X+wb9SRkNd0tpePjkkpfQ1faiBIHgUAIWPo83daYsP
FLx2dh41wlHeIK/fI30YoZkLG1jsV7f3D1cI80yBn7QFEtwZZO8AhZTdGp13xz3rsINnllsGWFSA
z/cUU19rqpiYJ3ejzxOWCO/qFQcBueKtD00emyPerLmw29x+NZMc3Kq8cMPtgHlJYA6bkAHPK7hz
CTNQlaTN8g83B3Q6IZMm4ulTnMyyGJP+xcoEBb9y937rLDlJmuZad5YF0y87+/CvaOBVLYMPbXX/
ylzBRjQnKu2sAHW5k3q+uUHIxS7AT0PKx/TI3OSAxvCBY69DRM/jYiXJix427SELM2j/ckT5MqxF
1xkf9rmuK2aM9PVoWyVEeqeu9LVpILbrWwqEIHbJJSxH+cRBeFjZqX1D1ZwuKjzJzmWSQ/bHUGLt
gfZ+giNVwLADrvSWnUn+OdzVlm5G8rVIAAoWP9iubrnqcw7i70McuvvM3lu3vCMpQBCCEkrlfEny
hkiV6/m9ijpCvhC6iEGR37aZjotNqjj8s7mbisuPges9mvcejfh4oEZLn9zuNlGGuZJomdiVP5bJ
+fTFQfj8sgw5xo1Y22+OhtNTjnHJuNo0/Je7T+ly49K9Hu4XK93nCQ4mCCxu1tsL4Dx2wQLM+Htx
ZjHC482DCLLotqOhS//zNYoi67Ci8Oqks387R7LezBwY5v8lta7jB+2vq8Yf3IRFwSPuQ7VPBKh9
muMTweIrvjHA6UPrGk82ojEaW5965iUO/1UTKbpNqlEgY8RvVpQi4GMw5vKkdj+IsU5KbXuH0cP7
TORE7y3mSW6t8pjd4Vh7UCa2hFmd13hRFJ9pEQLBuQfPxO8h8OSKsgfewMwZqCylAEjQa6oEaPEL
Kr7MH16JQqhOphHD4VGjQB62w45bQSxM3x4MV/Is16pd7hKqirNpdtwa4c5WYIIu58C+dDtxb/2F
4JlUx+cw2bNBYA19k4tQyylNk/1olggO2Vr4fTXHK9AtKkLjBSMsG1gVJVbAEhpqGliqhBch9Utx
mPms9uEUGyRmiAUHjacZ4kFvwc2hHWUccPfLy1arasFJagGAmFuOWxSyZMCgn6c8YnrUdVo1Z4d8
5gj9yuba9A3jYAHqHl7VlYxn7DjosJUxG2oLVAswQDFBF/aJxaOqakTDgI+S5pWhFPodJAjEkn90
t4x+8fkby2Nv/u2elXaDai3SFRuvmYjo/rcKWiwLjX6yKe8Rhicu27e2B3xJHI7a4bb+6RPjBl2z
GVjD+ls7hEGTKNjY8bygijD/j8l0LunWH3W7HJVF8+bMzFPhL7cyXj9FNEjHF+hie+sbvxLZX19a
9r3eQjXJmIG1PPurM2+OyeQguFNaxm+xUDZNSryg63u09mbowoIafUGxqxprVTQh+fUSCknlLYbV
isGmPWkiDLmY/rsjywyxEEtZdeH5y0BPyy+d5Ds2kIJa+qAgdrLcHM47Y0thGsCdrjagQW3Tul6M
LBCpaXAbNBBCXbBewUx5WfZVSkpMMy9WAVxZaU70iU6Yy/AlQq99gsmgpFXMFGI9K3lBxa6FmLEz
XgZLqLtdI4djBlR1xd9LZvOFqCHffQY/FApdSr/RzSbWmZCNrVPoXhsGAMBMdZEAH4YrfL1DsVGn
Uozl4wwMMsWk93Pdfz3x/4bYNMf7cndHSLbzN0jBdFt6NIBb+ST/KQGKFUDA0lZNxVXYcOsEGBM3
K67Btbh+8XE5YVNuk3vhXdoHNi0bjinytQJ9sthvHGw1mNka/l1Z21UrYpufckW1DBqfXSkDvzU2
zUoEC8lYrimEPUOewNOu9/zWMMDFzRWUyeT0Lvsh4AVmeTdTuTYSkqs4RVrFp4Rdkc8Ikbq3DOha
OOR1jM60gm8Uw3Uyj8dDtK6NDn+G3QppahNiDAA1D+5qI5B9ViG2ffWB8S5SnGHFyHacpaNkGtSL
HKeJ4jqeLMAdX/McUdqqje7qwH9XOaA1p8ARohd5AhjdmAm/u8NJSSJJnO6ivq9Xz8rCG527z5Pl
7tk4jMAD76VWxlE0+j1XHZt7TFZF+mnVpQeC3dH4qtd/Cnvy9KclLy+I6kXsQvOCHMcDLhkZ9Y4A
DEfVDpx70VkaKGMDRNvTeGZLZiZY95lwOUS1OV1Q28ypG2nGQmWgGn8R/ynfs1AkWe4Ryr2DcdnW
Gax45XFyXAc6dwpEUwjwjGDV/6Onn2NNpDPyQZVu/CZhldSnXn2To7XUNufXWY5PLWu6PrkUmkbq
FiAT1imD0LRfU+EaGdRcgFJzjzRk24nsCbdMXtjT42UIbXpC4sGdfVPe2h/YJcf96jgHlm0v3X5w
khk9lyh/MLMsZOB0/rEHYZQucSsjexN8mLRJsFUMlnNI3zjSCph7hQ/B7ySJfuDYvgCvlOYHMUD6
uN+nKBsUs2NHLBB4PceMOwSfZRFmir9MgGKsWaKu/PbwdfvtYii/TyjqVU7+CZwqabNrw4po9GVg
ViQIroAsXExcShpIQ55IzfE5AUpYldqspdTt2s4XgNBmw5fMD/INU53X+0p/IQ2pfiYdztcGPCjo
kU0v/WV1H2AWQAzbsfr1VPaNwiIZi8ZY9fkXyxhmI/OQYeCf4Nd9mHo5ykGrqRA5K4/JgSHTes8O
0GUBu3nmOq6fA+aAnWm1zzfzvQRY8xIgE03G9RlSFc7O0rUVpl+RpiPGu5UGim606LMxBnKIxJry
iFkBWiYv1rTx5f83rf7qpQQ8nLN4c9TUcmQMAo6i5mIJ9W6wSYTkNycwdd80X40zWmCoCeIyjiGd
rqYGdylpDF5VbPlLQYa69goe0KiAsVrgySyVpBT78GvuZymMvwLgyZg3CmTQayALe4gKKyAl7pdI
aTJox1Tigz5zsktritPQsGCqrjpnWaSgW4NaIfLCStfDVc+j5zQxS7qsTSgEhg/2mY/El1zDWSjl
jKn0L0lQeIr/kpStOwgRQb+PMWmSU0bRGhzvhxjQysGFxQOVJOwq9FEt2R/k9W3E8Kic8ekrOqpC
MptzWBEUUoTRRGiFKWTKIdfq+KUWtHtziDdAe4eREVmfaimAe2BomWmQ6tn7wpNXaJpaGR9oOzF/
Tu7vRpSQ6ur4lDXDltHnBbJ/GorDFkv4f4mANtoHWAOX3DlwXuWgmS+hzbMHy+XzxppMr3CH/Bw4
uhbzPVcYFqj5loCcRzu7RxE4hw5F16yiCnNQAqbsUNaj2CbPSD0eL/47db1MTQX1+4QGMWA7Qoqb
LiI/HK+5Yb9uOnWf7+6w1cbM65hKQ64xZPazClHcUzBrmmSW6t1oGMiQZom+NMAnF1kNNPQHQDxB
XglZpBEz4bd5767FjyP2WJJn2L8rz3tFet7VcmPsjX2nZJxttvmSHND4aLUepoSSSn1PmQ/defjy
fASnUpBHM8FeEBnQh5gVt6pTC1KpgIWNDyDXzPtw+yMiaXpHx8hAZy3CULAvbd2n4ZNRRfLyFBxl
O+MuA0jXPKzpFkGocmEbNImJAidUOQRyQSo/1P5Zrh1JBYrIWLCNnVXc7HV89RXJkvr30W7vKiGu
DO/sNY7muQ+JXx1yfiOrNADP3A5b2DPvFaoIELrNSuz/nl7Ktu6hj17rFZr+AnkhKdQN7uQQVHay
J2GeZNq+Wdtm9asmHZbIoSaNdpNxvCCKJsBr7mA53gQNESkZL4JL5b4wISl5X/m3zIxsh0OSFxrR
OIZKZfqpYcs90Y2vTIcv92NBs6SvPcBVMLi+2rtbADd3YwRxek3Mw+/0RfLra4XP/sGv4QEV9nX1
HiOKNFS5HCiNPVQfIXRWJ40WDSXoxk4baKp5SxOIBwJhsmFt3ZbU15AATmfaobBwRJH1aVMc72io
GSpadVgCjZoorzpTwycaz4pIHIJh9dPQjaQb1p+wrYDlJoft/SrjVS2q2suwBqdaRhajecddgpzT
kMc5OE8uI4nBnJ5VvUanOoCmcPAKd5WWHlU1baswzfUk8qYFKznJwRbmZ/ebxMtmY/ixGswjbz/x
LDZEg3qoHp1771U6i5wp8jHwzCmnjetfwF++ibOP1ju6xySx4mDQZo26Bsbsso6CB8TYPspPo72O
03R1vxhHOjkMvUuy4GBB6aXVdTNNFz1NUaaSnIZUJU6xsY891CFXSRkJ1mHK6f/vdqYauxEer9/m
4GM+sN1yXTknrI9K+PFKSbNJxkpoFQAmIA4yZbxePaccyX2Vo0TR4TV3N2ht+v4UeUVzKbdN+m4G
ZZQvCIrNr/Rzo9pwRWFfbGyt8ze3aKOuLein69fndiHG5rr55P4V8Jf76Gx7r3oCnD6vcgPQ9wof
SdvIC3PJcNAo3pEgz4xBGpSOSrn0GXVuEhp73qrsC1GfqqqxwmApovdXn9MVa2cwz/Tt5rLYffyC
FAWYmWlhy/n1lT1vPCBNeSKp44Ph3M8o/0t0foWjF/IED+4iwC3kuvjhZkdy407U3LfiYCKORJEy
I5bpWQL5JPpzzFTVbHWI0VXNDgfp8gACHYjUFgfd4Rsx1GqJDYVDzdtcBHQGwM/1iM+EWbLuXHi4
FPoUkVpI0dqMT2+Kx5/xgEa1uXNH/a7HyNbtQv0jgzE2kg4bz2+AurOrHhT7CfYWaq8XbzadaaWG
JMqbcyvsnvPTl2Jhm1Nl40YXRTuthYTtUrEVlHF8RBuxx9dvC7xZ1EBaVuN9g4KM0XJrDaVEFIm0
RHXQL6ZRE966tzUBRORMn6MPkD4jqtyviElGoS1znCVVpy33NBE3lInkaUgN+l2C3AdaxfLsOXP9
Tz0RauCzBnB+/JM5Xqd4hil9psDmVxQzy1B98i+BN/AAXLKWbQsoQnLOa04UIfXklw5tI05v7JsM
+5Qy9ou51qHJftaoj5ypL6RnmoWUNgzmZ07cB9QWfy8n+eg1lndxmed6rx1k80IQEoNhqw/VozMQ
vKMwfFh2bzxuZa9l07uz0Jd5zT4pqqRWOjvg9VRB80p5E/GxktRkUMWPYKILxi+FYC9zrcDvNezy
vz986xWAsShZeu4dXS9s0mjLUTbQhDiBzP8oud823NvoY7HXfenpFCAU2UVakk1dHys73Uf1ewUC
kufDvBwzKw/OTS/T4Hs5PKfAZ+vxiXIL49Y0l7yjHSwloUqR3YL+/MPDLMcAPT8L35tAK6HsU6FE
kYCx0dbkpSgFKYkwpIxNLI44vrnqz1DRKC2QCOvlcnLvyWf1D30IMPT6jX6T/22SZ/789/asVycR
WB6C/OwbPRIHYR8XLlPH7GCgF+rjWKX1SS+8y8nYqduLpig+HCv3h221TuyyuLPrzpITmJqKVtz0
TT1APnVM15JtCfY8TYAOMKNoD35yoGCQQqE6q77QocspuxZ+CyIdTgctVGBTi4cvfde9tl8rslV1
xJxPGjVO3OKMjLmFRlw/RaE1EmPNE5sbPq/dVRKNF6hOrquk6LDLxPVMDb4U0Q2tFLKloe+7EIbx
UQxwHL8Jyv/5XzVLb7XCWj6QyADxfQtUKGHze6F49Y9JAgdqU6b8PUlQFoKVXVz7qY/bhtJc3XWh
IucQQTl61Np1/mli5VXDafCKdAHzJO0jd9LySiTzTDqQn+0EIAitA/hFhz7392cmcTaG9qF9VOtx
KRxr5YBCKKFp6/MGlRho4VVsKmjX4Tiz7AyHfPGFKwvEj+Ko3Xbwsdl76erZ4q187ri/ljtAThev
LKgOylsaLMhLHPr4qbcJOlnzbrM75HqrOn1yYGTsoXz/SwG6Ln8EHUdI5x/7lEqAmln9WnxKvta/
yW3Jy8yKVwYW1bo6pFDUBZvguyH8ZXDKWCYL4nku1xFQCEzB9xpbAKgymwtDiQ6uLvn6GWduLR2I
rplPnWm01QySvDqPW0cK+xG6td9IxG5olZeB/Zmgn2KEyz9w64KVkcGJ6dMOur+vd2gLtQISMCV1
SsfycGzbgECb498V8ucxhtB4OPzI5orS0EKIJ3rW+silMJhETZBJYVSehWC0zTZKbncCXAF3Btp9
jw3slHsjhdSMi3AexRInOyfiFHla+NJiFNU+big77gk08NH6He4YCjZJaBGzaM6MLGr2VI5LfTKR
FWhG5zKZmc81AVnnlxBN0UiC195tmwQObWzDCbAXVHu31gJt4Yq/ajd5t5FX+Wp2iwSntvwAj4jy
QSVG/7gLRy7MboWXMpAS+An8Jk9WobK+ruO/pXEdc8UXc8rNgE7TQqrr162kxeaMZ7AVb741eT+a
PoL3NXUA11oqE5Ix74cVCSH8zY+r/FVwMkLuZR5Gmz69DN8GbD7/lhDk8nisTVpP7dimI09PCaMp
jGW4BOMblI3R+EfuDccDN68D2a2S2tDnIu0BW+UW72eH/dFF/jZzjMNGZmRvb4DYtC4qB4KDrJH3
gV0jX1PEEn2bAFqL08uhSleTDxq5Y8mZ/CXY+bQ10X+vZhd5AXvHfy6riwe4Mi9pV4cKqZ3BCcA4
LOgyTfPZji9oqoMF6MV/n0yv/V2K5JF3KdBUbkw6og/MAFac23w40gYfiVb1VR2fnayi3B4C5IpH
7tE7c2hJ/WoSQS2e6poAKyI1EP31h2Rb1FW4FTRZPHbCiBAcd8KCwuRFXdimRF7mnxqncoUPZXnK
CSWHckUBvL8kdShTZSfqylWZyW61PxPB0kwnIXYV8e5NZLL8sKPoDeA6uct1l83et34JnTK42U2X
Uw/usHbMx659kGmrPKiRIoLmkBKVHc5bB9wyNbMX3jtityMAykvH9XMIUdzdRe0iO+tIYGymtTEL
UrekkzWVO6I5TZFQXSDhkeFulCM5Yi1NbnnLcfyNvacNVCkgkUmSOiLfBdX6VDH4XYNvxZDjdW8y
l72yfBXsuVp6I+rGONO/JAqJNArvjq3yDf0hz28/1F4EiZmnQG6BrIy7pJxbXx8dTSeVWYhwIYxd
mF6we9QdGgHT06SLEho5e5AgzSJ7yq2ZjZyZs5RgxcMLjTUgqaL7RAympiUC2yl/ja3JUQC7BJ+5
3aqHgkokaZUs4S1V6L4VTQtEWeS8l1U5ASStxdqP2Kd8ZrldNLldG11g02Rk4EQiPMlYjHlZmsCQ
Sm+8fvxTS4fz4GNJCVxlJsqJY/1LMzdiIILd2NKK+G29KbvOAJEjvjnfO1AbKvogoGT4+y3Pazjn
fYAX8O+9Dvmf6R4Nj5hbvCnaDPbS9jZf+IX0AE9v2TuK5dpObVluSqj+mYD87eXSyhl0Fb65bMLk
9XMq/Le3Linh6ny5fkKJHu4dFCIxoy6fVKPiKWC4OAckMmwQPvZ75elq6A6HPHLEFp37g95VmlC5
Og7wyswFZUmZR1MFW14lV/mjOeuigaJLTB1bt+L6xGvMHh6/cH1hsV/R/GkOL3+aDyVRN0KZKVtf
N1JcFcu38xmtCT10O1fG60rNE3LkrTAMBhpQvve673JrcVJyy5x/qnEjhuSHVyOHGnqtDMpp4YSr
eBkV7OTQap8sBSdO0xIfnLWrl5lzA5M7IMs8MlaDuLSEG/23sjEFftsNdKROqcGouus5oNwsuEgG
bgUpIZHsetoJdMSDi5i7dNFwFyzTEVqOk3nFBVDpNc/knU+qbgem7fje6tKrC8QmZVZCJ0UsEK99
iSs2CFceL/QDoIdgFxf91AdipCZWVtqaXg/0dAb+zHbQ9+iW+Q9lF1yeXbz2D85gY17M+NBdWItE
NtbHUVa6btK/AjSiX/rfKCivWQijx3tJO1PkcH+5BGSvtrZn/F4zHIaNfnvJJCGsDVjRHts6E59I
P787GwOn02hes5/LehrRfKpN2HVxInEdUBnXq7KzcAiMS55U8GfuHU3Sha8kQUuSNMigFdX7hcdr
kVqRszh+Xwk/fhHu2EsZGxiiaYDw8/yXaxYDk338Cm55yTfDCyYMSCcK5XEN+Q5cKgrW84w+30Mw
gscRHtnNXUNucYZ2VRhPIdBFroC1E5Y5cDhxqEfDRuf396TYBLaCnBsBWZgzr6+1w0gL2816+7v/
KGSb64kLNHMmLkGnuYGAJwS5VOpl1UIkNv25UJgI/L3+hNH5om8eD2MVKMJQMu+V3mbGyvYmAtDP
AXwP+q2KclHUOQ/1Uk44YvMsqb8eRCvuHQXSxdmYi+05GjelLXQXWNdeUdSFPZfVZPU0xP7Iyg+P
xe/Wx+yG60Y6btsa5IheyQmh+CX+xVcIgLJvsynYgTxjnSsD/Y2zkVO7uykKaNN5/KTa/n872lQQ
3KwvCfHm9/p+TOD4MlS6cRb7H+OOwzx6C7+KNmJPRgQi8nBuzVTGVkJwhht5euniXltphUK3DdCF
9+FCcm1H61Nc7V3b1YnYyoOVUGCfqqmls8s0oETFAYi6AR6HgE4+xF6fNdbWMmF2GJy7Ynbpynsq
xdvlspCY41Y1JLoQt63wm0ZAqzTo5HQoOHjPeKEkuKdnhyCDxMsCq96PU9v9zg10PgLSYtXRMNef
pvmDAe3wsUPuSfEkdyrYw/Pw9pOX28s37uGFyn69oLu4oDtQDGdzzIie5j52L7alwvn01f34EgGb
dC0zyy1QsEns2DjdzClq9eukb0H7QzAFDlzxtWZxqf94s2fVHD7RSP5vtw4qF71HC3lZpBBDyucP
K9oDLKoyhfkzEzzpv+xDuVdUWgd0W4qvTr4Bh+EwcTVWOQOPLkZ8Lz04Kd9g0S95471UR0lcve0m
PWGUJ3zGaRGU9KLoXAOL1/xJd9Cg+H+EUfnSAwhHw/HpACrvaHo2P9E/a/fHHEdmQLFH/p6S67au
Xm14484EXX7W3roWN2wvpFJ9R0LYLeCSi7gdfE4bmw72iAw654kQQdl3fzY+gqK9E4QzC74oB8w6
vk0OtFAz2k6/pP4tgAITkiC5JBXBfeRf1PCTgdPH43vpPDNNTkrcnvZtf0xSsYD5U+myEsiZR6CD
FQU2t/Rm28xCr6Gb20ZvhVA9U3qVO66cAiph+IUa+GGa+ObR1TqAVItGTrX2nLRdv9DJYBsg/0ZF
9CNBbiodYl0wWPjUci2nSL+wVnjj+5SnVnqHAp1R0B2tV4zlrF6thhMfiXFzYpBGl++tZ+SMbD5f
ndL7MVDhnc5b5xdiut0PfEzTiueBRB0XDgMF4y/mx09OusXQP1c+JK7N49bpi3HXlRG9xdT7LcQQ
M2UhWdSTWRaBvERonpcg9gdLkmW2Xwa8Z0fj+Q+WAipLd1Z47yecihmc2NQZUA4FZuiQCliFzDmL
Enw1cdAz/By4fMbgfJjjEUGZEHFk5l/uLcsWu3Xda3Uzc1C4p4wPuwc/TZZ9Q97JNkUWZ+fRMW46
Ti11ZaM5qNp8LpZXuT7K/aLtMl6/mHhDfTQf9Yy5hjGpvoRU36oCuePyvkK9b4bNq3WJ5nM3VX71
oouNP7n+jTRpD6XX5a+SHxl+814LqflPgz/S8x5qMBE3FBIArt1SAEQw0fTh7j3KD1EZPlC01l5g
29tISdyDqTeI9AZ1O6aKwQayQy9DDWUjtB/11JWha7ILcJRXJVnlymwG1bMvCzXdbkGOrJpxOBYL
GBEGrA+Fo3VtWb/G0ludEzfj49ZQ6ZJo71SDNvP7NYGVNqOdTZ2IYhoHI8cULZhwX4qa1ADNQu9M
Hl0RO2Vs6t1/wOwXMpDnK094aB1xKY5Z1cHSewNxbeR2Fnbdqz648E5QoD/blxB8J0MwNkQ/orc1
VF3D/G547OZWrpxiRVxhboSdmfTQlkHxkQgHqn8i0Rg5RUN0hWf763X5e10rxhDpaUmXdgq9tIRf
wxDa5bgo8Y1L91WGrc1rk8vCbmE3EMaD3Els8yOHLEOV/fx5XXjPW0lPtCDPDEJNfHORtUX2V3Vk
gVc1m6yNfJmgJ/GQ4+Rx0eviHP6ucNSnpyT98ipfuvp7pwoGxpyygC1w5XX0Ee3sXt/1MjU9t62o
cnidlC1Pq4YOFumxBiOoKk1UoS/++ZEoVmlcUFd4tybbL3yBh+wrdDbAwG9+fyM+koiU8cVBG4Ik
HBU1MItejs2LJkBv0E5yUGPNAY+E6jRquoJgnKOBSyh51CFk5yf/stLAIgoYDlAMLBDwjg56kE8o
FpcUDwUxqNlu83oBJFUhcPZHUCY8RNjIflGWQ9wgMD51fLzcgxxduQ/ks2fJawCO/AByVWhfWXPu
0XWDMGXmjLY0Nlz5bYsTelnLTdXBWPNXed7SnFythZkwXYhtFlknYGmHg1+ZjGTaH1krPKDiLNoQ
udQ/UFcIap9uUd9VRbmTZRLdeAy8ahpOrhMpxqrQpbjAiBTT4q2Wo9aWqyaRMZSxE1eVTd29SX1Y
va76XOIOCAKF3tS8zAHOmRlwgJHQ9b8cEco/pBpfDAcEMsK7NRpbuoTURrcSQPv6le9d0GG8gfmo
moUzTiYiBGzSxmoubunm2ZTfhS3dauX/tonEHieTSlnBzEZOal/J7eutBF/WWO0heozl4Ke2ENAn
2o++XJDM0sPXhCiFUjQTH6i85VCcYfz807r2NlvtnWyDE+eqSkcP9Oqoh3PdJ6OOKgC2sdif/3cb
pODtH18uGHktY7PNqxVzGDdQJ6wTe7ntO0SaOnyho7eanDpdHxuItm7HMfXjkQzUuyVTQ+FUgYBm
dhbDpZ5CA1VxG6+SKZZBiyBbXZVhloUSKZsH2XSbQzRLjdl2RJKq+3evlbOFjyZ5Z8PdZB9JhNBz
X7BwihMuW5Hca1421g5aqp0z4HouS9NL9HWd/IWK/l0qiLpv3d324/w8GKT/Kf+WIR2KBqJM7P9/
D90PYI5SWmxSumSpgA9RVfiSXwEfH1Mxfe6NKa6ix+s3O/UJzb1NHd548brGcugDtf+ZnJJHjR+C
gBiKu4rTwZBhxHUl6Wlld53S5ByGCGLrjJ2XGooDl3oI1nn4Y6KdqA4mLEv0u/P2sozILEDcVhCT
R8ETJHrj1IRGpuCj6Im2WYD7O15hUK1343GyGRrad05SGeOK+abvrtaRZYp1ZGi4z9BnRvE7E012
W+v7eC56sjIxDjcNnnaQw49+gpwszmdJ2Hr9uYsFvTP/FqwHy4IlrXBqCoNfhpO++QeH6zhJBUyH
C9sXvOssPNYQaDXtV0+0BH5uzBknblCzPNj/pplkkSCa0mVDnhqvIrV3YQZ5K9PjXr4hrayjOJFk
UF3vNhzwOdKvi84ps50kO5yz+VL0uLl4yGucjXm4y56QRbOsv0Y13ja/UtXDqt0KmzEWgoY3RC3h
uCJ/OL18iUM2ebgeLIyltyBkRniLTdso/A51eh/uo0gDnmy/sXo4mPuTt8mv8GClLYu99ESon78s
fK+TnhZPWVOTM71fDBFv8YicPHqXqSra9jX1ewDjTEYLfzAtM5atbxXZwxtvp8xMdi0yv3gVz0OL
7YOrQsLCPPXwICl5GjTtl9eMSdMpcadUdBW7rDEQbcnX+oeRYUVDngWti2N9DWmskgReN3NMNGRR
PhHAYDbvBZgBW37rSD3dvIUDp249Sd8XATI0hzmoF/w98SPEuQRZgfAw1JcK1lgQLNupSpMEmPe9
s3VqNykns/T8UPuXMG431+Xi6hOMqIvsjVwYJmghvq88S8ZG2TytEYMa1sP56lcYr9xJYpptvhKm
QC5bQ5HMfpt/unRjbieHyr8O/FIdPJ2o2wZvLnop51KJyUrpEv0uXV8uxi7w7cAQtK6e/mWwiLtn
8ZJ14vnPdEBhAe4POu3o4hMt5OLiMtgdYvU/GMj8ReHTUR5nI9JWhxxFLNz0ZIdrmo9Ub8+mWF7k
xDvOhmRjObSRzCIHhAZgEB3muIWw8kA3ATcI4Ho+GdSYay1elgK0aHaTKNS74Rg5XWq+rbFtJ+44
7gG+CYt+WrQtF6Sp9sqmb8BNZRcGWXdsWen2NbHHuZRhCVZqYuc7fMQTA3GWr+OgapxbcyKPEjvc
aFpD0Ffrdb4roPZEbjSr4Ul3Jds7ZXYPTGoAptS8sF8OO/W2pa9jtNjFP3UfeCKE2UnbuKbF3LLL
nQOxdD7V293dlpSvzeDWmdyNwxm4cAdRTVS33x/9lguFwVdxBINLI5oDcA2RD+0sYxX5hEiA3WbT
vHSpPzyoeg0/IzTeVK/p4bEsy/y7XnwleGAeSh0uWj9wP3W/abz9h2DQnIZwVrE+uIwiAP4URkz6
Hmw5T4iv0qdRxomN02qAkv80dlfK1fIoDW3TaezoesRLidiUTHYckwYYie1RqR8W3rY36SPQLpy4
sDAveqSM9K5f4YvCviWx02Arb376xeAMkmUR4zb5Hh5oORu23QE/pRBsZ+reK/OTnCKnJ4HrqSHe
u3tw62EM5Raet9if8IsLdRdmWtmx+Bpgdfa0jlLamFiGBpCjt6m4KbLDwmPJZKAQ4paN9xTvyUga
wbpXi+RHeOE5jh1PTWT0+TIWbIMFBBqaHogigBRRXsZl9GSPi2xdOXpzFO+n6rrVjaBEfvr86E4Y
fpLuz9YJq7RsjShOYlf7s4ix8xKpBzMAeFvasXILx72fD78WDJowPsgDXKae7enaMAgUGwRu/QbS
l94kl4a+BYktgzXinfQ2qGhPgO+SCrY5uRRpnYvn0C5GPPxT+EmcCJKWA32IB+rYWCLGZDLGybid
Os7+Y8MBcQx05k+M32J3rGIzLSlKTfCU2P/NOX6symuUrwCB+dKOliRk7xMOOAVlVEhQ68tSvicA
qCU4gUb8x6/Wu5ChTSujqGWxDzoN0U5TvVTOhpBEVjfi5RwIZV6mcVORbf+FodNoWrqLIkn0R0yq
N2UdSDf1lpSxZf843QlaTaGcXt5L8MNtmzytIrxZl4y6XPYMZru0Nlkprdkqhirs7UBI0H2UCPVE
UkQXet5kGLAm4iWFVgdrR19YbT3cyGAeO7OpsJU/2jYK40lyfVQP1lZ4uwpbAMZqXcqffWbClshh
48CnS8pTzNCOj9F1BhSOCZ4Dhjh91UXrWWeuUZPxyfUKKY+040oK3EhNhmc0v5FjflS4YU66fRhH
YGorN2aqbyrdilW8URlEjnfCFrJxIDtUCIDECiAL+Oo3Ac7ZzA+9I1g/kmHlk5Wrbe3HUENSl59h
tn3vwVUpB8CWsEMlKzcvVR/w6FqxX2Zb8DxBNDjMOTHcQwK0Y/5l69uSpytbk3aXKJGhIWdcSG/U
4PBCjr6JCLcJajw1VHor2RI1CBgWSgIQlaXF3BjplBa+eLqMm/8ysqaak9arfGwfwe9xo4MqUgf0
360Ogc1ccD/p/PH9mVam59yrDVQIyuW2P9RNDiJoO9dtCZhQcvBn9vCKLEfCpOMHgS53e1co2yQ8
RUt3JIxt6xcGjAT6eXT95O27HmMyw3w292xpsV2gvx7d27whjVgvl/AbJ0WmLsTnUCibqvoNyeCz
pveDPr5hlZ6xxMkGgLDCbkmNOqOIQWcWbFd9KUGS4JjVXz2tSvBmB6jpFduPRSsIAsuLS0srRD2O
Z2drFT7HXn6gMbLFmouEzcZKVnvr7SDCsyEl9qjCou4sQpiLYqOiYBHqarCzBz8LMW1uk9G454UP
VJzNzU/oEzkGdz839jR4mj5HOVVBcp1pe9L5qJ/x+x+xd4IAF23ZUVnd1iY0ES6PRVQHewGrVzlL
Q4dMjsYC/7YeZ7+UXM0UptYyiW9DG7OR30+QiLVb6RTMR5NLrrWXo+0nrsOaOVJUKNViDYAzSwBA
UnsHFV8+/wkGWeZl9fyO9SrOw5JVbVL5ixDfpggr00LXUkuQdGbwrgdBfLMw+92BvXn1Zeew2XrB
G1J+V2/Zx+cg2/8ptfLct5lJCqvrpUjoVzZIF/RQgIROBUcxoA+zDNilN2XWi6CN9pd2cbtlHcn6
ctY++q3kl3HhsEw1lItAkmwujNlmz60HALMN5eq9zEk1MWIbnB41iYGcl/sIAuI+JWh8U73vXQS0
24cH3EPVjpyX01ndNyRTpkzs/IzFzP29jAVhYnlqINOFkHyGOFn07A3dl3VKqr7zAvqIMAT+lUsB
1SGOwyMzHPnb45zfKN8xgneYXVM7DETCh0R5TdGe5CTHj++Rl2CS0CJ1mKIoeKKB30EEOvkxYR1a
4CGXeV8CELv7dpvUG4aSqP7HKfPrQ3s3ILNQiCP9gsfq47T3rJ+qH1WbywhPFi2Dnd3+4j50DtzO
zigSNSBzTygfq35VEGk8Qxe5OPWMT4nrovgFoPv9HbbyoN23eqBo3fntVB1FDRD0M89bYUpJhFog
8FG272EEj36wbwpNzKTZthJf24EHdSg3mhurhp4Qr2Lxpd4eorRcWoe5jkcmsiwL1wCwVl+VoqoQ
r+ixqfKBL+tgiev4ErN4/4aleVXaY9InZnR4vulc6rwJspVQ5oaFzmwKOg1CJqk2DjhWWoQdOu4C
rPsCaBueqz65ALuFn6co43oHdM6ZPqLjnuLaNgCbh0sSlPbZ5zm0t70W+XBAqNkHPoTQgKGwHmsV
vft07NNOhIpv1Knz/q4tmLq5z6bTPB+Fli/t3lw0WKG546xar+bXx34zdmNnzUVcJGE2s44TMNiu
S0OR58dsXnidX6JWT8yXcEhs7L9AHR10/WuEStJHqsiogqoCNDwgOn6jaTBmudLOVZaE9HAbRuUa
LStaLpBy77680zv30lJhyiHs7vyucjs53i/rXlkomA+mkjdFQsUNOeN+i2j+NhBKOAjn4BhY+KE2
AAkXlOWSVpAv9VfpeyUtTi3mZlpLYL+OeXPC+Jv/eaX3xCh7yZcgSn2qKIUfphlY8KBkVGAr2bqw
CKfqOUhGGZM+fniow/MHWvE1XpW3pqf4R+TrJizc31+dJtRA11bw22v83H5ngxXkte0+JcioSrpx
c3NpXSzfQWfOKFJE/9VutLayUtjKGlrXCZ0+j5OgSbJu5OyhHHLSIzEA6YQxlfO0nixkwlmqkekr
oCmdv2FnE2gOUvRBT+s7GSEzzF+3Nu5dEJkglqJsd0A+tORmlp6i2rHJChNJQIe9AYhlu2ty6+9o
C3l1iaJ8x9UpeDGbLYZjAX+0JlN3YPVMxWHOI+5zpOwXqA7JQlOqzwxd4yToo4HL79V5Ear2Kbyh
uJCFoYIo0OMFxr/nWWa9Cn67csz7Zc3vYbo40OmAfSxgoqQRMpvu6Mgh/IDGSFGdYzeYQIjX3Jzz
Ngh3nqOoeIlwyMPvysB6Go2/IuRKxw6F0I9Rwc2jL0GJ5MN7CQnkpjV9F/5FxafCGVNTq85IQhMZ
iHtvwxX6wwml2MBEcyT+hYzxHKoiaUl+/D91Ru5XzdMpTVoSL+85Xw2x4afj860iIyYvxVbxymjS
ut+7DIJ0oL1w4UOJgjQA/03W3nVJA9bNb9LwvbWkQ1rB2w9jgKjfhuAeXKmUac0yokbW38jlLjVJ
mWv6UFtlDQInB+VkTbKSUTFEmpVrbL1fsFD6o3uGFA89VuS0AWAzoL9CYeY16GhOO4H77v1E2nRB
Kb9nqdjXsnEfWHAB/uG5xBwK7Y/ZidmeEhC8JpYNWZ2RFG8jN8PHBraqKP54STdsDW4E6v/SCxvu
vNEZa+OB1D/mbAW6fagBK5gv0Lu2VCtvwMsfxFRvcrXzZdP4xHqOkIWcuaR3Kql6G3VzZy7bOz4R
2OpvC5zWVMDGpjBL4KEbC53QfpFGVd8GhL5PQnL4ZfWE6gbEioI2qKcjE+1Q2Ob4pP1adBX3o5RJ
w+cXHPXexvNp/7p+aHsYvcMByfaxfez8uB4kKgU3NwOUTbErr8Riu3putFWNW4LBpqrPNsXIzDdx
Fk1Nw4sjzsrXL5P5GLEy3xZG//WrHGr+n6NXKXaJH7H7umDeq2IDLk6bBhbq/LPPeZEgJS7hCHNI
fOf6b22o881Hftz33bgpbxD0agoUd/yTvv7Pw1w/1ICdjgS1VJElZJVWcvkIMu1H3rjeiNpIsbI7
4tJP37Jxu/0AJMddOGjLfiLKaInp2DJHMh++tf/kIb/qczsNXmBRkM74Vx/TQq8s1FW23Q/s1MJ+
OquvVsF4EIvtVPrTTB+pWki53vSUHRWr3k1Y0AzBHXGqQJvnlJWWCtcVvsgTqVFN4ndhAZhIsIN5
NwRr9fLcCoadTRJ7cOUVHOt8OS07twuBf5Y/imWB5PWN9xXSjFJalgd8LRz7rfbSnPtF+xT3pe6K
Ihu68gwcXeVnlU+mRnu/AI5gEIkvjNzO0NweinSQNR86gHs6sIVBk57QFjpkn/T9+Jkb3at6f6d6
Em3GjRG7eA8VPc72rzPLPOTu3+7sgwBglmix0HARJ6b5Mau53vOf9eFyLwUjhNNYeojUW09bEBJT
yQA7ShleHSxDSGwIWC8e8mDdzbPky3r2UZ6mDr41cinU8BFhcPLv1gMObfAcv1r6pMDyFeVYOo+H
ys7vK0FvM58G4vkvMyj+TZQa3MOYVsEOrDGh28VUMQOq5DHt6fE+9/nUgk2qBZgP9U254Yz54/Ts
qQBUvnAt5bdNOyZnD4oOd5rq+DWNImkCc+nUCHcHxT1DLuCoSfUBbXNlC0MIfiv9SkU1efk9HRl0
Ezg7RXUdKhrWlv1p8DdU4/tabwEZOmHdZjJc8SRV09SVtvY3BbhX6mBdZRnGR1x5pgOPyyAkXKVg
yT6Gnetwr8tsP+vVwA7nQ5YfAc2oJEOLWZSdeDuFMlY5dN2PpLn50bWCp/LLEBI699RxWn7tPTMZ
FzvGZu0DcznmLKpKT4u0Fwg3DITjclbs00QkhKS0zJhJbShF7PSRXfDf9YDLwfEgplVumHx/phG5
ZOqlWd+kAOrbtrscT3AVedphhMJ6sM8URosu4achXt7CaMbH1G+gj2EhUqTATRPHOfD/7WMU+VUm
Dw0IXpNCSko2EoILL+dLnF3/01cQDmpsy4dnUK9nFEFANgRQJaAx9sag/4gJHGe/NEU0OUcOQ5dS
VLhoVwUj1Z67cP8x/xNg7wgjVYXhooyElY5siWEeCAZdAHVkOegEq2kRIZb9AI4hwlzMpBL//zk6
38b/ouMH1EsL4ie9xysEdbahdKor9ZxtD5ikTKFOzt6x7fX30BF/2TcE9sx61pfO4d+Ez6UpifNq
l1u7wEjl2hOeafOA9VgADMEAig2nS3XDXJOsl3GvPDv1Pz+oeX6D/pTJndca9Inbrl/1gug6in51
1y45y6pqor5nDRNNp05qlaJrfTsKHflJ10rrUxB8G2Bj4rbnZawrwfy+Ef6Sx0aaIXeoTZkGNo0M
86yWzZt2ajVeRa8utQP5GeHO8pNssgcfAP+2bVVIXzk+50SEuYB4hyQP4BxqxgddAkMXGPHxaZno
LSie2MHO3GY7gjL6xsfkMKjR2GMPKGb2u9UuyjwZU5NC8DmRIXH8I3/tOE4I+SBl70XvI6Khnyzo
cTA6pBZROdcJEfVv8sM+r4aybgXoP9SU/6izVeMlJ9uP329dwMDZEBlDud09eIuJbdM9AvDg9dKM
B07lDrr6ljsFekR5O9/V6074IbrEDP13PQCD3Q61Bo2se1/CY+4je5yTDFfDYBOFxmnwn9rrg5Ce
g9KOb8kPoP4uDNCEgRCzM3uIwfPgBp4Mv6OEnKUXCFLOqZiDr1YpTBcgPS1xq6INkv4qMvQ0G/7K
iJ/EGv/k0sarEspAxswtECXRNwnbyMZzvksA/vMrqHYdpkQcBnuyZaPyUUgk/aHod5Z+Ou+FVy59
9JLg2+KItmi7yGHbGSBc4t+qPKeJL2DaomUJM077cu3BJrU5fqjVrUAu56oUwf/RZ/oz+WeDNoN4
Be+pDvfDhgZnhP9w6+y1bMSRCzYM6eo0YxdjoQER4M8aAmunuobWfSQtRGtbiNuTGpPXHQGFf6Do
jyp/3hnLttyP600n1z9dV1D8ZoDwXch+k2lHDJZRMxV6/yfIMBA00F0/XnxsfS38fjKlbDgNlbvq
kUUrV9yh9OeIxO5riBE35vEEAuG+TYDy8d7nEKgvEIhra2zByeNkun2TFxCYGZv3HZKLdWx6SAEp
fpjAVlJV6PhWUjGsalmeIefwhoQb9vWrXRdxYzwrOYUQ7f1ee4vMrJr5DHJyYApGgSq1TCBWp0bO
1OS6JkM29XOboaTWqnpdUjLwD2jPqI8iKZFEQQiCMpvhl6fxigIy2oJb70AYh0B4fVbF24OpsUDT
q3eWdoh4/KW0s2ui0q1k0pOIh/nS3ARjgXKTffAGXSpG5e/uBlz/Zr8ElNZwUNb7OcZUkbwJXeY6
dHg8+1Wz2nN3pKKbBS8EHRY5/Dwjo8R7vkx5bLCjuzsGMt1eyNtRZjmWaycHJJGmj9s3syATeU6h
Nf46UenzfSROrfzV/9ArW3+fNHwx8YBrXMLfI1sG2KZ36+/g4OZDuXAJzJw5eCAh0UwVU2BvrngP
fu9DmWkp116ZhOW+g3Bm+oNKyXuiXU8/SIdnAJt5rOjLUAZb8lKDDr4SRUK+LYH/MTmLCoRTJ40g
hrpTK2/AIrrEZLAE+kXPPvmdiq8tzgFjQL70ero92DDJ880ZwrpPsCCfLwDvM7Bqp3KDNsp21cGy
FHlvWGeW3itA4w1VRjycrxkQGt+6/pz97kwQUJRpAwGNzns/DFaSlNmyO/LyWwiuu3OznWQMb8aG
kxLZxPJiIVILkiahKWf9ileu4C8i6YK8hSVS/8ppc7Wlq0WHm3lccDDsWbOctI1ea7G5nq0Yfkl2
ukW/XS+y9AYp97bpFzLu0elYzzLKMIDKOx2UEXfigVwYYI6chSpMhLCXKb7xCTQb/ZBxmcJ0plZA
Dy0X1sgg6Qr8dAIROHYzD8ik+10XYmjlqD/uTIwNRdpBba5LdDXD3o8DWGt1dGPwRwee24dY0sGm
/hPZYoPFpup4tazZE8fk31p++mtqgXBNZxmINyXzXeyiLszKQ163iiiEdG3Okwy2dPe071gebu6a
krBepC3sgycdx4HcECTegdkVArhfkkVY+kepWFvV25J7NLuj7u8PDpDFOWy3lUnK6RkIHHtynmXM
AFOXbmuUxk/FKHukJzrJXkkZwdjVPnrrJSrzB2UWjKIhUafkLygfzyp09Iq/zY1+ULAUDjjO0q9v
/P3x3RROnXM77BR54+6otm7tEww/ZAsAYrVZ+1GlLLtmVE1mjrNtRsalsGuEorSeMwpDYvEs1RuK
bDvmzFh24Ztm0xqBdEd5YEEAve9nxhwL8xkA99NcYOrDYToRnoLUd+rL+T12Uj5q8IgbydjgKnvw
4mz9I1Lf/r1ig3y9weaF7WGK3tpjtWO4L2L0EizBs20DsayUsvMMSYpBFsLppXoSyYzTqQtsW38/
bv4etlATInP/3upn3l8b16ZnfyurwLXgPYOL2/ZKy8b2k4SSoE2VDWKJTHPZOvioQ3IoyqpphEVY
vZ1wcDyNfK0sHEyJq8aNnXjs/oqVX3dKCNkz+6LNvzKAJH8CGkM8CKTgE8uA4sy3XGmcH69HY6WE
s21W7/H9jpf7bJyAf/8kgjccgx/ZeSTC5HQkO+5NoAKoIPGqj7Bd5KB7/pdeLGsvbQWLzpNfc7qk
1bCtJB1OXNfy13cGLRQOrAZGqE7Cjz/fgNEsKnotN6pbYSY6rnTm/H3n8MdbfXoi4XqB+E9YDKF6
/ip6VvHXdw5xmzwpZs3FmtrRgXk8fZz4BSkYJzZoqEnUq7IdKOcWIzLNnY+qGrXiQDvg7YCv1evl
6YeS9U/Ct1n8/6SRIoc8dNTxQPaFYtzhXqc60UofW9MsrYL4IkkBSUK/SKc+EhY9pqCVWoqxl5uU
TE4v3JmR+RzPbGs1XK8i6z4XPxsA6g7t1UHAjmyIU+QlBLTjO3QWJu0AAnHdpynLWyIvggTUfiGk
p2sah7YigxIJq4V2Hc32GbjOSfABlLNgRdi7014tLT3186QEf0/sGwzcIg1dVnqZDUoySaYDjBGE
8OimjQQORqhdMON35g4Xv5+8Rxt7fh9rrcRO1Sl+gf7gwji6oNY9lBLaPZOYubwdGuaI4dTHIaJl
jTSqKL/leCv78zT5ltaiv4wzBCN4AlkyoU8xhqtLMQVjU/8XetD865ER1oGFBsKvmQL6H1O4Ic6J
dClhwNY0WmiQMzkQpwte/HV5qV8I63/K/6L6dKnnB0eA79Ypv2ERnGph+UVA3dR4aafni2Sb22Tp
sdFQoNM+8lYovAE3DUk2oDQE2HCAmUHurQpYy4DU7NJlUf7nl/Dw+llSdoHZgC44q/9OtJuY3VRQ
6RIVyyEhDITF5w5DfuMboA3jsaNlDTDYbtleWZeyyTyWLIb2hT7uymeTvw42HG2je7wPfUsg30nw
Vn2AJ/LSLxmsEMNjHE0JkfvDsYzD7IeDd9xZn0A7gXFl2dhCaV0PD5C2Hag2EkQyNnfKaVW/PmTL
Y7DccXN2UByPIr8ikCS8guwnRTxSRo58/ESOlJsszqqwvcv0FYAcPugnXABJ3QYaXf6/DS8pme4C
F8L9yT/+dAEz31jpbdRxULoc4fsckzINU9D3B0m6VxQibk/TrMp+kuwgWHeqWLhNwyQFmz4FRo/d
bNAuITaYbU5CGcx3mxItwsemQPJaCJiy6jGL8uchVUJMYcjXBq/dvdrcZMk5xlhRHzcPYpzMC5Lq
NclDCeqnTIQje720/SbK73+XAyZUnXENm/ncAhjL4ZFHrzwo/8zIGKw9TgO2onasgzRzg8vbSK5O
VfDQU6PHZSrRdZutwPZint/HzQ/Fuzy6YDI9aXWToveAzf9Hh7XYskNb5HozJDP8SqxsPYK7BvND
zaHojp6v6MQ24ATPBDH7EGpS8/Rm8s1UUfuMDRGwCfczH/ENemeZ6uQBlKfyPu9VJC/NVxgtwdKd
odr07+Xl9K0CEn/yra+yilppfOBSxzmgAE0SArv7DrSgDz+pke17wnrSo8IV+LaQYlQYWbRI1U7F
kaimV9OkthDbqdXGvc6WyjYhsopXRSAq1+DkuqqZz8x/HHf5M9eSKFaBvWUsLH6sAbxEsF3sRyVi
K5MW0fBx5jZrHZZ9xxpoxlGS1XgOJQaA+JzT3u4SMRc9Tqe8lbMKWC6KTybbuU8L5axPoeXDNIPa
SlnVzDZ9TGqV3hAqL0DJyxtWRmr3D4owzz6qCCMeZX0vPKqO15o6jqBDHD9RppnF6cecZUpGENwW
rgFGtDAjs+nHhtj2O3p0FrvfW5ENOlnxgXL2wFRX+3DZT6+wuh7tVHbSqiEVl6ftb1s8gNvGhcLN
tqxcUJ6PmtKrEffc9Ha1zU0MInrIhONj0EuLqJxHoWSiur6qOQAX7J57hKcDHSYCttyL4bh3YS0h
N0XaUHtt1Zk8BbPBcRKEsOOx0onKZ1R/hYidu++/5LT/D6+MY4BsJ4h/fRNgM53gJDxJxOc3r/lY
+wVUGHLE1RcrIt2tkxT5W4CIHnxG5SHgufJdnTNd90TJ0/7AY/09SA5ORbqpmqJQ4xRqxywkqaNM
vteUNkToVuM8RI8YgWVdCVP9Vm3fJq8rjn9tD8kpqUHmCvidzAvR3z1oMGEuKrcYNMN0ClG8wzhA
UX7p2cP3n57dyMZF4QWc8gYSveURMnbMrlEASy3VcFWgBvLKiqFttMOpG4nogz6rgA2XvkB5xF08
hQubloazze1EnqwtqUkZVEAeZk/WUaV2Kzn4u9Nzzurb7+yhQm15NUSS7VMxdGt3B6oWqDWrGf4a
0MQ6cLvYqRR9CjPKJrqSPJ/gny1ntrCIoswVci9e3C6IEVEGQyAQYEBOUbeiT8PLgng6fz8J7ljA
CSSknOF6RDE4k5NdfB8aJ0HVtSLo7GXNRLBz50tTcx9KGazz1q9LnZ59ppEpdUqshXv1eDJm1viV
yTts5Zs8VOdxzHVdWzVLpeYtw2O4z1CDWj5e4y2HoGTEYf+VsvZo9R7UB/8AEjm06lzQWG5T6S09
8dDUdbCqqd5udvjQS5C5ZriYhJ4x6iYyXIJMv+Bk3mkAOAjm48Wwejme4aM8KLPOeirBn0vculkC
ZqIzPV19AjQbkgKyiW57Tn+/Tbv7F5EQfSg+pU48dCLPSzsWRcORd8daLy2ONjRAtfsdoEr7JXDM
4/SWvG5bXFPSbL3qJmXjgwR9NLBpq31Vagyjrcur7SoxC/mdoxMPvJknNzqVrfNBncPdqRvCD9TN
H8kPvf14XGOx58Wj7kWbBx+j0MUmhQQ0w0o87jmts+MfeRAx+S/cYk5aJECSp2G3hUUs3EzK+Y0F
mY8ZDCFpFDTF43YNz39SBhEdH0iFN2tvlryUkAmPd3oR4wGSM2O/ZvF8CTaUKShq3IRW0uXECrXF
f8+sjdEM4tOpEAnj8zLZOatdDq7JnjhbY0lBWI7eX4SG7p+P3gdllHUT+NEzSfk/O84BJHQCqRYf
n5/TOER1A+Uo853MJT6WlT8+ZQcduEM2CN+GsvOCycNmejfZY48toOv9lgqoEn0oF1RoMxip5AdM
ZUyTxS/ZtimWpgJJkReUMalN1WPnXTHN2GcuL4knibsfC3VCtzbXavZu5R0w4hXgDJOKqWFh0xC3
GeOITdDRSXcbR2dHG3mwmFTifutHx/Hsa64m3r31NFQhj5s0dYnwlFtHG1vxtmebi3j57wijNvyA
PdAj7NPf5ADgXjeu3AaewZSK6PDV5nFYZ6tWobq3FZbRWnWiBcerDm+9k17dWro133UiS6svStEX
MuGByhernuN14D5saxU9ko83BsR5B99spAxeF424X42xMD0k9msK2eQ7p+qaCnOoWZF9ORW5doqO
wjCLNMHgONGyS2mdh2cV+iZUDiY7OHIuw+xeXIinC2tn+4dQPCD9KJBQjuHf1i3GEJJmD0GnsOVF
FZZhqYkPKD7AVf0Jf9JVq0bx4HwalkRjIU2jY4A5gPLmAv+EmL3OlMA275XcPzcqZo0sfYWBWfIp
YtksTuPg1HXJKgZnJQk3AWdFcZqlOyy1ZlNjqgUWafzoIijCBNlVqq47jukCeSUf3owIzSA4ZLp6
9/nLqA11D7KeZNKxHUqGfXphGJVlWsc1M/C1ZfnzvVauDj71R0sXP2+pvmDG3EMuhsJ7vE5BRrId
vu4+lUDIT1N/bZ2t1yWqnWe84Z6TvOBn3nixlZazYvYVtlHEIAqTduNJzHpronhYYyY0bVhvPw8S
LGE0fBsOOYELJp98uy3Ip9tU+xYBtHk2FD2EmobZGRpwFUZ4TRTGT2/1ohC1QfRSUXL3KG4YF/gW
P7atcvHVNC8ePnZM5BpP482zAmDlDoFQ+zWHTIKwhTrgbA32mJmyKzdC4962KOTgDuxlgmc8uMLo
q1Vfp3q9ZyOrO6R3rHYnCP4OfQhCcxnCdNDlK/7o/J97IDgawAkEz7NvbRaf/tG70SlUrzIK6MM5
dnMiXgdA3R55blx3wRBfuarvA9h3czlO/apEA35CvXkh0bJwNLk886dFZ+A3Ns2M9fWwLjxtfPjo
wrJNZ3qbaYVPXRYSpNo8J0VELOGmmUctNTyXSjEXuoSiqP8rvjcduAVnrvhtZbrNzPd8jT4WwCLG
aZ4lNnVTV8VjIPgZY+Nh/wVhMjrrpW4TQgp7/gKqETvE1RIM7Sa9ty+jW213St8WPMiQrPDEzNWg
/lJAXnlFfw3lzAEiUifRhjjay+DQo79//wD3lTpMmBxuTQB3YXeLCxulNv+/NpB6Sr08e0J54iXP
U28I/exg1mNlM+eadV7OTZsgN1KLWgRGt5XbsYjeBywf0VDUs21+MADmsFm1Po65qfHalMDwbWPE
VRWVC6wPMPKN4bQ5HAZ5vXguJ5jiMj1K9Zkbkm4SnRfMRhCuexzXnNSe7ofvq3gRysA3TSTv5cdv
quhMM7IvDofowkTv4jEV2q4Gy81TUEunagiYdwpB1Bn76jDYY8bSjNSzxIRbFwIVhcfoQSWyts0m
YcvDVnlXcHfiHnzZWp+SSeueH0Fw4rkmK/McYidOdapnHjdJErQlXEU7/2a3Yylj41K38NxIPL8K
en6i0ezbFVT7pkilcemvcMTETeqWTBELgu4PW5oN++k99ybCt3xce0cRNWjJd+vwdUDr6LJpa0lB
T/FhXW16Og7z0UCzIIsexlJamfCwKrDFgh5WTT/3TmRbndQyhiMS1lrWfTZmBK1ebCykMpkoMJTV
bF5GOT/x5paSGRBH71dJuZQCSJ3KEGvzf4WJMK4XMMB/hlBlmMWFnfyBNnj9+AxGX4kqM6bVxccH
fKImhjambpoW+BjVz2OmQ62OGmvQK9qI7xFtF5RQfwOMUOBFaNeZDu+AVdL6pga9Giw6f+ayRyjz
RnTuiEK3BckHuk8KpreUK5gbbBxYhs3uLeDfYIu8GGoD2B0G3EJLIxabpY+6t1h9FqT8eo/vYwb3
epPIETnludN0zsLBYa6d+W7367PkyGfDJ8j0WP++QbJuZRnlSEXTJk4pG5RAAq7/wimYXEtL2Nkn
zavGqQ9i3PWY2QQ1c22VoiyV2mP5kFrV6Yh+0NTZXbixXbv4xsrgu5MS/VPSK0ZWDdL/C+3Xpu5T
9S/lsiowA57CLjTVDgw15cE20nuZLQHlnJfMxpzX840ukNYYwjRvcBLS+yDYwvB3E+F+2tTT3IYb
KqBo9Bfemz3vUGvGO17R2LEEYn7VgQWZIN9eRcQ7AUdxF6lercroWWRS7iqrAfnxpwkhTduv6Hu8
thvwBNWrLcfkQKgdKE1kYAWjjoTnjF8cGMdFPGt7LRllijZA1q6NHnVXVx7ovdUUMBG/0ZjDUeRW
z2gIvhMVUD4bYNZc0CV8dXtNrMPh/0dXVYP9MbKjVQ0k+TGbWCt2hHPP46UIwU2t7zvdADQfl7A+
F/eAf+q9Xgs56t70TmlT9nLwuaB5ybwi2God4+FXkKURV18AHWa4AjvUrVrjkaPbW3O0qgcw4Jzc
4ST6XR8NYgkC8pk93bl3EJsQZHXDBEciphDA3O7WEi5hHnzkIBLTPI6Cr9VjuoR0dpO/uiEiYd5t
G0Pxe7xfpFUpuwx3ypCMwOCeFiOJwAEXKraipb/KdjV6ag34KerEw/xhLmx/ine7FGutkQvK70mB
dzEG0KqP4dYK/Ix0ZEJfGtgzjqpXIIrJj5jpzEGwdd6vjupeBFkguUVC4/Qo7KvUNjqd05xu6n1i
OQSYketkLZcymIndDHpC4/q4j3XxMhdJ6mkB875+wug90sqfLjdME5CL4pvnpr+aWOgxqcuYEX7L
YYzmLskgeQ1eNN0hDOG3HqSJbsIHQ29waBgeHrQjyPdnlrkdxpzBmPBSibPu4oHWFOYqKGfDspDc
0dB3ZVxs/m7/RJrCIFzNVh961GBS37rfHQ/d+bpKaOywYTo4jzubQsacEl9aNfIPtquJisw+8kNS
QbI7xxRnCZ8txKL6bBEs4Fq3hG9W+DfSi2MnKQKTO5wnXysCz+HihYMAGBdwSuMdHWPcbP5g3fm0
vCHr3tJ4Oitk27PEdE/iI46Y0tQHu8lNNK0nywa8srJrmReZjW0uBy0iTFxy2WK80Y0VvaEyXNnu
b2PY5QaaVEM/sZVs4fXQMxreJTPBDu+Oqzi8gg135lSmurDYuf+DRMPC73FgBptNSaHa34EjO9vy
/1oNlZ9DRtqxE/xNB5MN4pF1zq9TtSnW1Cx2DuHMvMvadS2gH2KGbbtmeeChrq3KDOHt9zlbIX35
xdn8jNY1PNALU0cvRI3Ac5a7XLlnWFkKnOuvLz9L4Asqbaz9u80q8ReqUdrQLSWT2zKUoy7qeMFq
fAmwWGpy8GKiYNqtvQwwT4FHUWEoNxHnSU+pPRnj3nw7cXxn9F1LSJDxzLvkbM/OCuqvFxtQVwiV
UTpLcfeZvMw7/7Cu7oX0+z9bBzTd/2ZBBqzKXsu/BUSLCUvPcuAu2zbsKJLGgx7O7gMOj7Hayq5n
SSJPdizG56yWJtGMNFyq41C84gAsYmuY0uHu18OIgx4SrrqV4uNAJuIwkRh35CCzGECHRvOaq4MH
B3idPnqQ6ZVhno0XsF7rced0OOKKFQZCykuGPKGo5kFEgJacgP3yAQeiWfdLo98JbkbRxkCJHwXo
7W3bpC4QlYQRMzN7Oz64p9oehvptrcjTHFlF5GnXlfLNgwyKfac049dEd4s//5JFA3sb54vdGuni
vpTlS9vJElcNOEDZztiu4WNblGZZ+/7qCM+tW96isYgeKyWoH0BbPcv1oknI1pRTB18zMlcgMTaF
2q1I+1JZcBQxaBK+sTc+Ihd6cwcWmWEvH1r7NoWEY8yQecb0/FDxozUPXvQhbLgw7Qtr7EF+TgbF
Ubz94cCbNsBjFG1OYEMVdxHCbg6FtmqU1uTn9Kzar7WBNz74Viq6DhC++XabUcnfn0AigtmDGKlt
Pd7BbWB6Nk4jCLkw5WCbL27k7xFi5bQxRQA9xLtxwphCfBZiLp56YLMV40NrLptWjZng+myDSO1p
iB1vloH+AoUpzoLMfD9YwCugvj1andepz8X7dZdGVjbF5ofE1WuvkMqjB/GAJ3iEFEoRj2J8w/Jv
UONVyQ8RsChOmMw+eMZG4h1PMM92ar5tV/1TZMWvBGMVyldSXUuGIIJxfk16hB4zASFSOqFOmlAK
YbvfoK9LSR+NHBsxpqpG5+DaHLvTdOwufGDL3e6gIRlveWnhVJUL6je6Khe81/vBYyX1B21iA4wp
oonBPePUEb50XLOOyTVpOLR1ShFCzbrHkRhFuZ2yD7PLWgUamIyGSoziyYwcVMd7Fm8jLtcvpees
FzAsI6VX5+mjGvKtBGmImvioc6eByaaXi3sQASHLlsNWiXWiU7avhhrQlZZ+FYZ9Zze+5wJkYDaL
qQRpCIvwSms3HUM/B0BOAG/m72kKHeQn5B/84o65lxxbJZkNLciZhWP3JkqQEQSb0OaheOQgicXy
xIFMM6r4oDb0b3dgLopM3SgXdVtiI0rq0TUMQnFCu2uQSWz/Nzss+Tgnu4zVrfj339lQkXfbKCS2
dhfjxD4f9CWuYGKXSxEpG3q7C6yhzt2BYQDKxUF7xG1z3P/qkI4/gmV4Valn3PRCSMjhb7TKqB9f
W+OJTxniyiJw1EZHKnjklQq8HMe/yq3AhL8nE5OKxPtuoMTYORS/bV+C0V38ZUD7Nj60f4F8gEdL
N4dRVL0DgnPjTVDtgQJ6+MhznM8ZrbZopfEKO68rn6pvr4HgbI+XWcMs0MKDmgEVU9j8dZqf7yQm
M/RPnvGJnw+9DDlNtNhlMJXnixgyfUTM4xcwLZ0C1uW/W8cz1kVBdPbR2/mcZP6KTiZ3o9eMdNKv
Qgaf3kRZjcze3A4fnYGh6sP1+SEueRBNV+Zf1M78FaWAVqYNjmp3l6YcovsLhByBOg7m043uTj5Z
dDc5hfADTeaIwF6UarjYI2F4u8sebPx5+Ep2QRkQwR4nG4lnjbmaKE5mFRhUICluU+0hTCVUdtlA
T2j5TtHoA3WxOtKQ9U426GMMXjepMugEJz7bvwAMIRiWFDNd+Scil7m8quqcyztS2wUZgdnxjbb2
6hU2BXLdNaWljt0HMQ5+HOgZtYhuVtjALNW7OhSw0w9Yu4viSGwmvlwo97kMar5zXUKpRMEnJQIY
SWakII9kMRWHjCv9K8MEe0JeAlYULLdeYDqPsKlZxnmFDoQFrNfpyRHNFb3tfTKXgX5xeXz6uBAS
Jzj0P+njfg3qdxH5p9DfROEqrF+r9fEN5c4N1Rq4dE8POK2WExOjbQ6YuQfA6KE3kVyZaVDPKcHD
B6jsIItZ1Hun/KWMUJEeU1jEMoAQngmfbKSenX1zczKubA/wfNuJLQqA0Sfx1U6dPW5m9Z6TIjuJ
woenpltzg/IugDSd3GriMg0c8X7hYLo9Qy5WEh//MKBUr5RRfv5jcX5FvqUEH/5BogOnavDhG/+T
ptgCtuIJDmUrYVDVEsK8XWBAFSTw8oZqvgYn7dIejsfbm9Hu4jrkTEcvS9pfT60Xj3uTsZOhKM9e
6AYAkJQpVZN3YGFwCr+8SAGkzQYqN+d2to1Huvg6Rk+HyIJ4C5SgLAGFeWTBirvGi+ZD5Ay/gE1W
e705jYncuweYBE62uvqiSIbmvYpxO/ikhf0YJMjKR9o/UW13unQVH2Hr2+ETYhhC9QvFRsjiQ8nE
nbnYp1KTtvOwgMkWMqELTNkkHgADm3Auw9L8nZMtYAF9x4EHWvT2qa1cEQzNQohW3rpMeiSQtsS+
MV4yqVDiFn/SGSRcA66FxGr3Hti/sm/T8MYvLNXOpgaHIW4Grd3eG/oMlNr7MRWkJ2DRfq0a+OyD
uh6IjG36kmpZ+4IJe4hbpvPDXuFOQvzq+WaldGZnzj5c+c3Pw5WtgdzvYLGYsOzqlQB4OTs4HX4P
1tb4fgTWZv/hwzIVUFBgRVEdPqnCJbNCTQwjunXs7IZhTq6gLzbO/O325G+6+ogpD5uwx5CkF6aw
7C43kwuPLwzAL0CGtiE9ZE4uwLL0iHFHUhjycwwDj0RuKJUr4PZ+HS4o9tvx7lbzTMyz2dl0pyJB
39WHtaAaylr7NH03KPW016D6XoIo9frvr67pFXBbvitY4Ulnrev1xbhw/7ruSUMrsKGuKUUsTJYi
FeNfwJbgT/OwmtNR4JrjXLctzQFswMKtx42cDUShBds0p8szThmA/0OuK0eEqB1pL2RzuwNZlzRm
W3aOx+jZPKusFlINFUrtXWEHc1pPyVfkwfL/VBRskpXk6CfTGnUOyxc3/ClKXk7dADN0g9wcsswQ
1XiCh3WraN4sFIbzPy0N1rViaW64WB3t6cElEysStizRs0w5hhYIuHUyKMmrurO/DmkC9EgL+57p
Pf2ndZxLmVeNsZLnJdcoJdzVmOBWMAKR3F03b9G0wvAvKCr5tcEztlolO2lZ1w2hHV8ie864gbMS
NUjYQGvpLZNjBjzisSzQcnyrFzWQXcax4dnKJesaupHpDQeII66HXH1YNUZRwr+4IcijF4tRgN+s
Le3VhOlIJ5noZ0rtOuIU2chTq3hd0WiVsKvt3moTuenSEpNMxiZ9s442ScEW98txJW3BwCjFNH6o
cQDXc2gX0VCos6a9brouLhHXvlWtWm3QbVHlBmzBx3iN9SmNwnYn1rnZ6fG0c7qPMezlcnfgALlK
7FWAYwd4loDL08W7r+Z+zzs4cpQiRb9XJOMURLC/yKYe17foJMKQou9TugyOGFcvgnnVreC6YGcm
EAM8ASJtEVgZDH/vylSKaFNIkDjlpAlS+O4mRqsQKdTS8ZP1Ll8yl+UtJE1Qeq3Tja0euA3WLhfH
W2iOE1fddctZWsvT+G57ibiTbCxrwhVnNDmzV0QDC9gUBXPn2GJsWRDMpEgcgJMJDAjSOEW5VtX0
BQzHGPNjP9wDyRi90soFTB/Yhdbsfy46SpMmuYhf09Es0iHb8Bc+Skzs5FXSfoFbyms3isOD926c
RQ7QASD8krYFiiQ1bQqVuJ7+RFQ3ko2va+mKrpNIksa5F6dP+t7EUnyIqql8XQWhLgzDE9FY1kIc
3MxqXlU9oGY4cJDWpboyA9/PSdmmyAOA6otKOgKxv1qb4fiMsl9+MNqESb8vYiKOwytyRiv/pwJc
MWK9osZSsZjmgAWQ2fu2noxXDFcA3Hn//0OMPVuX5zRdtVgtEo79Fl8ogvLUQaSA6IZ6P7zpjWqw
A9gcVpB7h5NHv4VC/5Q9fjck3Vhz5qtxGCppVVUP8rMaX6PjcrnO06Ix01D6g0AateoX9NNoA0dw
dqmewrOz1FYehVVufSbQ8/+hZpWKn7Mlrq+/9XItws1yJryNRVzpmrrPPnqd9RUOKURKsHZdjCQV
OMb0QPqQmj2pNE/F1emDYben+vTHv6BOQvEgyc6t4AL25kMVarSUtsNuXHqOMoX4afb+dWP1H6A0
ECL1R17CHCyGkh2xOl0zoru7jyFQFQQRU8AjGlCErqd+4kPGF+YO//LSl2J3v17p9vmzkW0jFHg2
5NTTISaVY0zDNGi//H9SUBWAdvPAyZVAHmYf/FI9MkX3AzOGF5558uneaWxl9lHPI8H/6yJ8qv81
Ylwx4+wPyKp17OXT3z4XtFrMsAn7VcdIdL1mFl809MZrcayGmnlWVf8rfUqJKoeles2MizuZIWI3
alHFeijWwgdXB4H6xK4/bHnoSBPLRfdIagvTuTk3lt0FQDefnHwko+WwZ8fOVN+QNHbkvTaUHqGe
QyFRa9yapFeD5YPDNwmeAVjS43YDkAfVu3U2cDbplIkCV3MP08cp38QGHDduz12X2iCY9jWF5MUA
Qm9lRKOs97Gy/Z9WOOlSyA+U2/jfjZBInaLKGopaLgVtzKwuGpxeLMKciTtWj1i6GhDlr4iVpqGS
ylyqMTXIPOOS7hxt1Lm8OuC5AHjJEoYW12MkhF8s2B1WUsK0UXGjYMUBZywPRAUBL7IjAhDpxwdL
zN4mbVdcvXwLsTTInCQhoJ/SnhXnEkV7bpCqwV8yg64d9YvWpbCjs4MIZK2g8gQjDlQHXfCnrQM+
mAGHpXTsQ2fjG1QAt1MudOxbYo6jeANtPSuTzDXC6SE6asoMEBPdmf9o2t8sZMPqWK0KwNcUoHph
afMbusrObtJfdJWztkVXk2u9njxArO0OggXDEGp3PBkWIjYctCTu76DFGZzjFc7csTbQ2WmFKNxs
jwkEYUgFjZ3O4rfgGJQv0VyQVtyrOD0C3kAzVyb8thMwDXxk4ynyl53BEX5cwBwbdz9A2SWuA/7Z
MDdEUP1vQuLUBwQWjGAMGbMFKDwK7XMVsVlXKGBlxFMV0NfOfrMkHly6A56p6ioQch93EP1LLHcG
FppykOwHu9fjKL4k4v2yabGJKQ21X6+hCAzJGQEQs3WKMfPtbxNc1D6ze5qb0E3DuEB4URWQ2a11
HrkZtavHw6x1lonTj7YbpKhOKgxotj5+ggoVsEbWtqVcF19pAPhUQqzQoJn0m0j082mET8102ggr
enpO+K7ajNat6hBg78kk/byd/i+Og06A30R1fz1yxUhXNvGw/HgyvzCHQTwdc3DVqnhmqztvo7SW
oOqf/MH2LlSs65xJtRVnGy5ieX+GHjL9heVIjek2qnGAs6edgh4aDJ5s1KI/EIi57K+3rGC22VwB
CI+1sk+MShkXxBdrtTHZ2hYWbF6DHDCpYqm1fRjS76vT31FZ9/O/7Hs3ZCQWI097TIpG2VJ3gJek
b9bomea09RVdDcoAaS3Z8/BxCqyaz7wXptOb8vuEX8sWRJFzuus23GBrIeGOeHJ9OYz/wSpWjRoj
WyAAbpFAnDRUqGQONZhAdyeqfsYjgNFJAHWe66mdcAiPIIXfv2IpR6qyL/Y1AAK2Gl9PWrmqmkbF
SLxQshH2O1guhT75mCp+W9ir/LWjteTRtpYcn9njqsyAYYKaD3kYBoLsyHZ4AQoCICemCIwbLzc2
YYBYuGtHyb6AxSdb5RPq4HqkomI7Li2CaClNobxmmV3aEgMhlxTo8ogsT2tDeLglcwzr6ekAnUXV
TJqJ4wT0RPTBfVES7P7ucXRl1gytOWIBs0fCDcKjwT4RRpGGc9wS9oyEZIt6o0zqhbdOY1dfjkEk
30uNvHBugv0UD5SkUrYZqa9PONPuSSdcFj7fBoxfTbzOG0GRtPFGcIIGungkp9ZBmnUP35VGrlWg
DiLsx1mO5F4lH/hORXgjiuj7uBlqy0X51zJSFQ2YNXjHYXORe4014BCbeiF0VyMeCZzvu2RzKyPm
DUsPcRK0Z/PUuOW8UAptvAZgjRvQD89oMAA09KRA2dh0Z+2R6dOlOmellHSpnopbhHsO7EyxD5ZU
bFhqjk4Im9crzoRPDLjtpa4EyC3wMuBA1df4rzRBYzR9XF6eQj6H8rXkiCcv8tpQ0QhuFskSHPTW
nU9iStaskZ16UkWn+Hka9fqEkOYOYqPvoM6ZkV64PUcAkKh7/u8ZFKNueUIBcDz5QUXy+q3012MU
h9MXHyRfIz5E1UOGBoIOAD/PTZKmxVvicmbURf2m/LRPyXaD+4R5+2S5+8V3mMcTvTCk+15Ivw0t
XeqiTp8O+iRxUlwrs2LkcK15UguqVvabLo5TgMxAbG73XrBU4uHmtMRamfV7qN1zXmoqxhkcj5Dd
aIckuzr8eiezLJcLbc9VBvcN87teNVnXHNkW/CDnQmLWJj5O9Mrb6cKoGxez8ilGpmKTV9rRORRc
gnqDhkxFYS+bOWk9fyIzmssnet2ioTHMg4fieBKcI0pFq2QiVghRyGgHMcrPN5ir1sSsVcb7g8SX
V+TPlUpWGIe7vc0kwAVW/DILghtUU+sq9hUuMqPYKUDAo/cQHs4/s4zbuadAhwE3zg9cHcQzFkKG
K63vDLAwTnRx4TzS0cL29jfELUTUlA6zWPw+0VmD3NXkB/YjHdNk6qke/fX4Gv+NRG/DfiNb1Su3
Aq4qzny//QxiCy68mFm5lSVxL4aufNq6KjTfqLitZikhX8gYJvInwpPlz1z9lFONTxsxgA4FaJLe
5cATKqejH+DyVYZOzie/Z/TV/gKnG1LOt8OlyH2Zv27XiHPN6uY49xbINw13lpAhqoOqqd0lHPB9
8i12KRQK0cRX4Ur8NJ3THmE4oGYKli2t8bUy7syGCKXpmUPhqjrDjnw69mv5zGHFkxgfvHEAPrgV
L2eDgmYu3CaT5lfm5ovFXeR7EMXmPnyc3wbBAZym6e7Yp5CRutGiFldWtVcW2qcX7YpTpJiBs8ls
y7fN7eTfYJ2D1rvtxVnMShUH3kIrvYU8bc1SLJrhUtV8qBrr4zv0HS6eAhyCZ6CLPcWAQIwCYoeH
WRlGPFMCTBSQ5X5JIOZTR48vxuUcl7YR0fQZh6ydvCm+3NFktuK28ZSn0PK82oX6iRAqPWM7rtzr
/m5CMOInP2AOgtHWhxDKXVn2U4r2RDd+Pa3WYEDqjtPz2wd4r+3P9yXi82mmlIttq3s0NlDsTUoz
jHVf+X5L0KoNI2rSj64M9ucNc5czljBYt0fBNlKcwcWTx6ZWCTPRK1GeJmOw+rjSLq2KKL/gVpL2
/RrIswNDAa8UZnPY0VuQKWBQgw8a13xzKtRkNNmp3OP3RZQaamJ07qa0Jmjqp0ZVt5rZfemIPc1i
3n+4FoS3/jPufLdPXxykms2oK2QwZyjL3Mb06yR82HxArzHe32K3CmBjSX4o0IbI4PpZuRJQzaZ4
OFTmho4KMAppWIb2fxFavhwfwQPMjKQTO26PFNAW7PEREI00AhMA44S60GsT1KRpX+TZy87X2cb7
kbtMoMAzY1JNiivl8YfTSxQ6gAOZlx7EP/55YVg5nLi+T1dsOo+XuMu3xhzZvlN0gcNDq0dxbQNO
IJ+yhsgmo7q+/PJqoXNdtwuS2SNA3H7crOHShShpHTjW6WpqRtOGrjz1EUogGnSO8YMQtXkv3ppk
Tl6Ah0Y2aaXLilgc/QvlPvI+QLVpvqKOx5AiKtPi+RlE0is9C9iWEA9equ9p07uzUU1N5i7KrNQl
/1qpP43YurSAlQe0lauvzAT2Su//HzNwJ989Id8k57+OxVKBZUat0eGJWJ/1lkNF/to5j3pdke0B
UKRS0WNsoUCxV3ilw9TOElYsH+Ssp0SuFJlv768mH8592GN0CtXidKFzfnOkcDWLWcDsTPAt1Yqd
2cOfD0nJ7f+6jCHqWM3JvSwYJhXAWMWuQtKM9a0cuo/jhfNG7mSfh6/srHDa6gt543U7d/YQ76bN
9IRNFoNbLeqhEGDqtQRRDavjmZp8o/tUo9oky2TB7qFZTZDWZ3sP5n0XD1f22SVbEVHWLu4Afd+y
9XnPDcapawOmV5f/cCBFY+R66i0krRfKQet8zCr0ZFLQLYHP9ZOU0tSzYmjIrJlH1qhgm0TNP7Z6
x5MX+DvcnvSWqrE1AGkKhVAYiLpxbtvDV4LDk0/+UIK3yIGR0H1FHjSi4DWf7bS2jujmEOaqKYxb
BnJY2Nziz9loKJXrVgqXbNnsx8ga6KkdrY5aJx0BMeaZT3Kh7CSctXrgz+/buQoNY4RpoRcU6SPE
G9FyXzLR48kF+02HdKd+ROPiTp9+GcONJOevytBEk1rdC2dP/af38mJ3J2f2wfWyflCi6jclYo7T
OhbXLgLA89b+6gGEgO5qNm0YhvCENtS5Nzku/oicARgbbEF27R/kGSKuYDT3Eut/ei3q0TmWyr/0
dibfXukgKd6tpybk5SDVxAvQFv6XwBK4ZMx+RRchzdNLN8ALKitgqn90NMKG3f/DezKACBmfeMGa
yCT3CPtg8XQEoIj04dA84LF1bFMMdg96za14HmWFwEvCnVQmUkOW0lRsn6EOGM1cDmGluSr7uIhW
5PcGg79U+rlR+MmXDwP32PjnMYLiEUF1hOcS+/lLrniRB1J8KMsgWObEQ7l+onwm9zuLVn6zc4Ck
3umCa40XSJYawhDD8hTmVx53NMxHMmD3brPuS/kGfr2VJ5+SXlLumGg4ERS3VavYtbsnS4egR8g3
GVmhm8+WE+GbWwv+++2BC0UVzmv2ieKcT7tUul21HAiXnU484rOX72GoylaDssOyLff7BJSqPpaZ
t+7MEfSCwy99ca1jDUqJYqkHth48wQongEBUnCSb1femOm8Bnf0kFV1AwIB3rWncQrMW8KN+zQ3L
3ze6WBxf8V6jwIisHvWmrRUbygVel8yC/TXA6TtmW/64vlK3ustBe0xq6JJcHKoFizXW08nIm7jG
ZZT2ogzlwqEHob7BX78AxTdO9V97PGlbNcn6iTdMk5r6sFJPy49yyTJd1KL9JXI6mQ+OvK+UtptS
Fj6kl1oyjTuFlRdtnlhfLfxC9OX2efVVnkMeUTua3p5t0nZKajQAYOEVP2w0J3gMM94PHya0cK8D
nvBZXLCfOzO1K8T8G/7TMFxi9Mm2hFF7SNGzKnYAnFrEnPdx07VKakfexQ9+F1bwDJ7CjGfbFK78
Ho5CDJb/gnoiYvj1v/U/wA++1N/KiUAMilUC7OA4JYOu7n2K+sEM9WP4ANTMXsJliLL1srP/S/Iw
4rcOatxzJAV9fTkfOtk1F7FShSFTrmKXGQ5ecNDfovJoqoGvfExwr2nAJpImEgjvfhY5uQyY8csQ
5H+KoS+QRedH2yYAGeDyAGd97IqE59FPFGEfuawn4NWjeWK6RHrvsKguSLB8jSDOshW0qNW8ZjYh
Jclxvr5XAx//08xRbeZjgfRzpOORyDs9ZVmqN4amOBl0gmDLSPGSI5NQQeLfDXYCspoNo09kj+QS
k97zPTEBTcHpSdObnTZ1O4DwVyVlT3H4LKNwSghhOjU9YEKpq1CbtPoF/INpj94LTHVcyPwD48Ph
tUoDO8w7BmOFnqj3P44jssb2Q/mFO7ELsWwXQkO0lgW4D+MTpcvgjgzSBceKLgRx401xCSywq/r9
h62y8vik6uHJr/u3ghZ3MbaeToBy+LGTDAqT62lIvlALhe16iPvbLBIhsOS5gCJeuA115thTNEq3
CF9/PWXdUQTA7mPoYe5A3cj8Rh4xAT1VUw8WGOj64LUbEEnwi24neJht9NzGkftHw/NmXt0Gu3LP
4+0WthslxEasIxk23T7dTInHAe29TnjR7OjlIYmOc4KOM2TVA7aZ8CvLzmTYdSpBrm7xC+0iWwrg
5ddq9pSdgEgm8XWxGapteTKMiZfsA++wcmb+otgLL5GkrTN2T5Uayxm3Robk9+JXqzkGiMWcsTTC
rXF5EHPxdqJE8hA+rV5xbHRVMOlBdf+asyJo9rGUSiULisqt41x1ZBsXexgONjgPc2/aMm7GOxAP
dgIJ5jHXD1GfhLoatqBFnEMDqsDZdlRJZfa0xuLhEq4p+MqvJeopKTkGFMb4AmRc4rcdD1OBKGyQ
0aAt3zRl5NOJZftFwmkfx4mAXIIEXt9FpuAjDzZfk3IaQmp12Mv08GJ7Vrcv8zR5eEgg+jnGzXUY
IllkfoBOVNNi9CRGOdzjC3bAq//hzaZ8R90AAxcPjtCVlm44cYIf/gYc35EWOd2Q3Ifaj50NCK76
ry9rGC6T6J6k0n7/KihgMnGElrx2tb8Xg0P2PgJA4xTm3T5pLn4LEjarhCMrxlpYWI4ZJysCvLO1
Xcm1dXLMmUduFYao0/Ay1m3uS60aPan9dbU4swwxBbqsnxFvpnWmkKjhy4GRToroiahLcZ0mLtHE
WGw44MRJ/8ZzgtIsaxo57Aq5PboF11a2v+z6bcij7ppOOzx8KEhbcT+Nza0om1rhW7/kP1/71o8u
ZeMK4T+wVguLEMKqKDU1bsnfqudalwGAen3AFDaYAX8rXDK5VTDeC3+w8WX4r0DDJ9MkG4TrEicN
Wv0muTSDbAwbOrJ1RUJ8VL0AGipNKzbBBV/D874l8r/eXLXafMlnDFWxuINwUqfTbffz1Ohz0e8F
WZU6mzWxo6w/4soqE0tReFw2mNlGrqtdw2XyR2g1CPzvnyTBaWwNm0xGYolFrAlmqcxBudurpt/D
0NxbIWoKPm5duzZHrvGR7K6ibTPmd90yjSzy9piia/OQjoOWbeaF4mB7e+gqV+Out47qqpMem+rz
eGcRWsKoWIUwn3MTocMRc0k6bhGsIPDKTOTozRvM90OAm1M/j4yhByYGntbcd0EVFV8QQSwGudFQ
0ypDz5rSrHyDWU0d6plJcTLgQYT2wL2E2YUzLoZACfDpTq7Q8i1lzU6CoDVVgKyLFqLWeiiNw5vu
F7NLZldd75PaLB+zJBRQM3GqzQM99mcAh9wV8LJDKFH2R8xeskYJDAGD2lI3e6BHcfcWwvxRPKIq
SciGCHbNjnKOqkTyKY9DnT5voxlgU301QrNjDaBUKFE+g/stccZ7atNlGAU1w0z4h2bmnh0E5WzS
VmUV8LkJiyYLj2PSDpkgNCd8ykiUgAbFAVPM6xLmX3FHEzj1umcDqw8KqoSguLWkomnkR/G855QQ
unG+mb7dUWb4tsAkkcxV0rLa7AJrEwAd+O3UWxzbqx+T0XggdKJbyFtDR72kImwxptBXTSkTNc3/
B6Vw4Yv3hOCK8I9pklHSJuN7tqdy+8zjxenMm7z2TreHifDqZMxvR6AmCXX/gYoCXMiy109AGlcG
VVGYcFvhB5XVQIGn1O91XfJqez8HVZnUVzSf8+HADbGPT+NSOnf+5v+jlkkSEWytxsVCP5aocoId
P1bEv4iFjtDDr3ag2CCe/s1f0BgpJncerzFFuaQAqFFHorVDu+ZyLDOIJ7ehKBpDzR0lX6qz3OGH
bzXBFNbH6sfVHuYywnOxYMStUdrjb6fyFur51OCVX9/YU6i2edDozRElwA5nSbAewiF6Uiz3nS/b
gYMv1RFZ6VQAXazS0MqnFYPKIRWvhI3todDkF5/K3iH12jRoF+2cltfqEy6AzOKD2B8LqptpJrl8
nPH/OT93q57DX7SjGHB6Rr4COJdUmYRU6PZRsKiaahs1W55gzjGPx4NdCvfvxXgeR66n+Z+Mo3sT
r7NCr0uS2eKaL8fLhHidGc9yWOJ6ZK9rAQqOS+5W+THip1Xo/Iugdi3OxbbmteuGqixocCiQrFy1
d4dK/AAzwErfwbn2UUl5J3/pEzKm2fwj3Khn2dlF+Co2IuZTHZmutJXV5SlouvPCWC2DJgOEcmD0
m8suVxhDhyPmJlCDGSbVa7VklCKLoglH//2KToNPK5pyP6CJo5GAY+jVh8xoIgr5mWN/HJZMYDBm
tncTubgSOPa1s4LPcsOiH4UyHza+9PtI3PHZQxRoYzYMPXQZEEeDoVsqh0NCBB8wvWYJ2wO/3VcN
t3rUALvjcwSlT2wW1QuF1mdmxbekVnO0da4DHOKEQ2LKz1qSTwljJeY6avn+V9AYyigxJEE2LNCK
OVCbZjUWvV0g2RcSOnfDob2dfN1i4I9l67r5bDRDj0qBw1fTZLAIvmFhxT143WTIpZcDHCPB4nNT
BisAYbMEuILpX3A6wGSHeeKfxvEPbxUNRg7/pKbYrZOpFwwBsA1kkuyZK1h/9UoAkF9wf2FN3Aeh
DjO2XmqLtnI1nt9vU2A+GB8jE6YXgR7I9+2bHfab30Gc23pEWUtlOIG014h3Ll3+9u6KZ/unm6JE
Yawf1f0LMP53w/zv+o4NhsQPih9ubLYMxkIU8sPXw43F/kgg4DCTLidsuzPqxBKzKMVyJi286T8r
4Z0JYzaPZXHakFHiIiQYPdeFn4G7cyYIk6frIFihgvrmYe/Wv23u413VjdzwJqChmRPkpza2XAjc
SiaWu8Cp82+n6aUaeNwq2/4DnSi/LBQimhT70CXtnzGEQeuR/9XYHS73DMteUi7Ldpw+AG+ErrET
wup9ef1WhE0hR4Sjz+U/1uW6nE2G4n6e4VMsVwZSOaFaLJUawg6K8IXXbmkr0DqpXLofCTUc7VWg
Ktkqs46SEkgf1dXL8kceVDuDzCFaX6LF6B6/NlBdFKEwQiJMTMXPvxRwgiWIFrlvBqFeBW8OH469
1vdukf0KjLAwaGv/dE24fF5qEUdCOB0u8Qs3eLSe8Y8CVVghW1s/4ddARxb0/Y3B0r8A48NMgVnY
ds4tI/QogkNsQN6tuYh2c0rupTgpffonBaxPKTCnAKNJwsgO03zgv+gChInb+wa232s63Y5mOctq
zUuV4MZEhnSXI2FWjYttEWnYqPnkTaFRbRAwkf/BhVJMT1jR2SKJDuWRVq3fWOJZ5JFAeMlLjhVC
hqgUuntxeoZvO1KdAlNyDQ1OZHWiMPhsUO2FjsEbvDixTJrKAedcKCvCSyT8993fpIpp8MHb5wYj
FNfHoSmwPGqdgqLN6ukDiRVIpUID8mLwKLYa6T2MZjamRWD/KmCDGBkmY+8bXx1rUVnrN6xgJKkV
XE65b/7L5Di1tDDPF+bRFdFE9IT1u4+FSRjpdKAgqXFFq9tunKjrPPPPgCX3ZvTSEcWtqG9l3mOy
bgPRMtNwuCh/RblxezSQsNSyv1IzK4UxY+KLfzXKyFNsF3r0AWbqNzaGFSvYMnUi4mmW2rTDTxK/
7aRa3MRjPke5xeXL1bjC3tPCSgXBaptj8VWkP1fUlOt0eHil+NycW9jiuuq211uRcnm56q+k0vyi
dvX2hNEsINSgmYwlkxCKJ764oeLmrnhBv/nNWat/Nl9v8I3AVY+NZ7PWwLxt2mCBOnz1sbh7Ay7T
7vnUu1q1j5Xgnwx1mDrEFdhGST48J/pGeyx6r1KdBgEWB1F0E5Sen7W21z9PGC0DG3+Us7j4lofv
A18bpXvu50zH6BkJmYRq+IzYtynkOwDXUhyc21IHUXSGK3Gk6ORZ3b4qV4Y5A5/rqgn8y4HDCY7S
1hW8LR2FbTbwy3sdr9B4qjKSsM6xf/U9pyIts+z6Oo8d1gE4pXXhNnW6Ot5rall5iXHWmJ6+dl/j
T8ekCRacn/yUkdVWwqhcdIjwvHc7RrbwXv894v1b9AEcZ4w+To4+Zg1dzQiOv13sZHq6PWJVumCg
NDMkJQ5qXjhVsf2BSh1tOkraI/l/PWFBe/qc/XjFmwCrLI6HbRxMzxcSuOBUVmTBGOLoqTEDR1ih
acUo10NEHhrnnxECI96vr1QrQX1PLn4SQL1/Tc2aRLvQK9CIvz3FdZJARB8F+Ya5XcaaJUJjyEek
+o3OH2U0fQcOSys8nPn1hT7l1kH6iFdWuJoQor4liXaUA9QevXqC8KQZLsrfJTUBbxRZJOZbjDAA
gzgeKLw8MyKeHSsOQnmVx5t0ol5Qw7w0vumiBePiYIdb9OuYcq6/tBKKd5nOUBz1r+hOeiX71Vc1
deKf15Jn7rH9yoyLx3k44nJtOTy1fyAmab8/1dNfivhk9EHnZ1O6l+jsGcjc+cS5Zn1UcP50WlV6
Tt3wfHsax07p7PzmE4i+nP0d6xfceaj4+BcB5et9UybE4GJSh1+p2Us2TgLQT2u5m7g5+gHPBhAp
lQjffePEPTY7Pq7xTu9Dk2mwynsuv/hptRwepa+AnZKwjFgG5cHEfchbCBiIoRuaNJVTAwELC4W7
b9r6W7/B49Agi8U3robMPEI3dQGdbbw8Xgup4jwX5a1jzpjWelbGqKKeEgN0zT8g7clXG4gmXFdN
WpZP/xe7Ogxs1AE1MiKldSavEs2qtDz8FukrTZfg7+6ZSFtb0waazPHuOmM0lCoqvw+5wi6SShBn
IMhPnZGFmJbGPDLVAMQGVQc/fHuaZwcRlNyrGRZ/vuiNSl69Uad5HEh1RCHR3vit5MJ9+mEPNbP+
pBQ2l38Tj3ZR6h+cUfrcEhriLjJnVZr0C3SAfxbgVIpHXvAaBqt8FSKENPFvTt2gtj4yVS162Rs3
t4eZ8uOuNkSTHbEINp/uL9rIdO4afZK0UfEW/2QV6B8iJImVymNUYy2fjaY4P/6GrJNIXV34Jgia
97jkXPlqa6/DJeSEz5/ahIjZeA1Gs4n0O2Nr8weOvSRYbl0ntveYL/eyTEWfYqWSlJSAvGs5qCZE
oQ4AI2OiG3oyEwtyQmT1kGWiwXtoq+9Ln5Q23EQ1NV4E2A8YKZOJyGDM3wrGdPU9no4QG7HL3rXX
aw20XRfT615Y3NNijXRg3oNu8l0GSsCze6QR+0aetxAPQywAanPdZ4pOr6dte9YFbZ5xh4d2IlMl
vI7NaR6vC+MkP8OYElZyvx6ccilt0Fybv2zl7Owd3DCsW9HLwwfqbejfYdBQ1YYxKYyFiIgpuZPV
APuEsBRT/gEpv8zY5hVMTxjfF+L7mG0N5YLy3gUc4+8bJxcdFmys9L3VN6L8SlAkTvJO/AjLEt7t
fREn2aAeVbqb3dV3OR9yg31++IhaKVCraLiJzujKfv7ufzmMz0Uq3v9nYbfma9QZBj8cQmBe7+Xy
+LXUyX/UhRh+5Pq7goE9Zrt+i7yLIW6QH8XajMhpY88xSiqVqQoEUpLZ+IpsrecQqfAZ/AwFR8Fr
gbwrr1C92ymI0SaGidq+p9RDtgaWmHoG/qXGKMDD8cYLjDXqH1e8U6dWhqNb5KBGZrZsdqgtdpcx
VTvjqXtDPY4ek7e+VBoOfTWExo0/+JIXo2RcKuBm3m8FApUZ8tdJdqurO0mghycKm7tfh9ePFT02
eptS1Vhw/NdCyHgdkGeGOD3PVYt2xUVDlKJH2rbfZukkSzrqbDr1EChOjWWFLsQf2NVq8UkSz82s
CNeGMm1/eu0stTWoVfgBqWQDZ9oiVxBFvQgIpPoDx/eYfha4wJpsoUUvEkhFe2yFV9eQXJOHAdQ8
HRo3J6Eh/aPVe5Ma6VYPvbsh0P51UV22vmcuJxD5Gz68toxgIhyi7WVr3nLXY0Ah3cxHZ2DEskj3
o/l45OeXKR3oopuTXQjrHDV33WLGnGQnBtot6zCq9ZewmMkw47YOe86fwESS2zNppksOmva3Waxh
6AomPm96zrl3bnuX8KcY/BbOyy/R97TWZnyh83yZ8EaUDHVOyvzb1HHAV75wdyVGF/pLAitI4eFF
TCVm/nyVY6S7STVVeQfGtBUxNFUNo0uYFouNkJJkCcahJcGePdIHv6fhKz6Ry+WNliPSG1ZIUhd4
xfdjYy37jRvj+4uu11ICSFYTR6ivKAijt1d1bGT+H2Mb71UIVH/rYIzRkAFamWQEAXH7arj5BM9k
jy9ib8lGi/ucHlP6xYgoBffnsFkuff7Dhjkn1H3n0khMRqmx4yKiy1rtlxTuHNb1233jZiP68MMp
M8/KQs8YrzCmI8pUlO/N5sAxrdbt2kbuVrcbST0yiHb1wMxSPw9Ukb7iawq+qH11/5AzkzDpRqoZ
hKbcCnTMV2boJV7q4X35aUUojA6XFRTiP0Bf3T5GbrUHSgEAylTM/KWGMk0RNqdLYf9wQw2XDQ6I
nFd2I4SQgYFybVx/5HC3tQwmsi2p/WDnwQq+NUcWlngZO669ukYtkudnHLT6qFNvnwFMitDmH5kS
y5SkDDx/F6VgTutuD0C16ylV7vzRz7PhnqsBlUN/+ZfHQa9w7jyiLYhWSk3sPIl+nhovONEyh+e4
zX2ELTMh2Hr4KuGigT01u1QKT7jRqJeOXz4V0oVfor+OxkTdRwtuiOkhknR3frwdhJ3+bdJHenqF
E6fgSHEC+Fnjz7OIyt7D2JbnbvH0N+mmYEbYkkaKxgxHqTYEr0KltInyFpOzSHyNKB7yRKGZvM7e
mkXoA1ZzUx+c74I/MIsRD5hCX1UNv31DHqvZGW8tSpOs6LS66q5jA0pQJZL8AVJFjI0qECLtLwl6
BgrVMHIcomIXafpQzokimcdwHH+WhKVDeTFMov0FujEB69U6HuE809a8N8D1s2I9Uc3Ois9nWrlU
17qOAHYbyd0YWGCDm3ddIEzDbzBotdcaLOoCkcKK66iD4mGTI7q7E+O1r1aAk8gXmgW3UPuzS0aq
t1dTU5qJRC+A8xUAh7m1fy6EOfnitC66Yq9zvub0Rt3SWbK2zNtRua35iqWH1B9vmfq49DpXiaVD
D5keYT1Of29wD2ylGysAH6T1NmMh5ybSYLz84SFdOhA+XD15jY8gJOv2HmFeFRAOltIdHsSXgLaN
P07Bs8mFkUA4eO5TZTLIB72a6DCPqqpQzGUbZR9da6yeHbywix4JpLEQ4Nw1mUWmgAj8K2DdP3Yz
lHBCyxqjAn2S/m69DioSngpsdo8gNwHCT3OhD5OIDflLOVsbnceNF2RAWnttED5v/abpRn9ORQ0n
UDP3MCRqIzRhq3hIac79GnomANPDKypCAqu2HZt1XCyYnKzEknPafi3p+pfRW5OqPzvy81AYdtQS
a4zbXP8qfwdx2Tbx3DGs5nn2n9y541P/gD/WIj1HnKhhuyEzvKY7nIComJJ9OzNM+kX9ySa2Tsn7
OePQl/wweyGQOMLahyW8q0vtAeNWFVE/GHAdjSAap89sGZIJNx1xKPmngrBO3A+pZ/JqT2EL29f9
inKLhDu3+5flPlx4W5Pve6DDnLYmmTGhS8WMdaG21Sq3yw4z7tlr46g3T+nG4RphrN7IhLIleBjN
PCxfkw4m8zlDUFjMojAfXN4cU1Ofr9EbvHzPX2ajBBGuQ2XIayaZAn+tt2HuVvkSi4nwSZ5vEPgN
BgL076nGuhhN7lIuvm2i1Vv4uN4vndgbhpi18trMFI0CcwuDrlX9Y28iMFVeIA6MZ5asm9yyYaHG
l6Rrb1vIyKNEoFux/tXo3szYPkwON1YaYfoS6dJ8Dm4f+BUSWqomqiYHsaPeoUwck7BVfEq0HPij
5mOJtZYaFwZhhvCU9nucUm/RpHSPa3JYufDqI8tCjvCoky+pQ/xnkKC4wA6ha95CAqjtQGhH3gfN
pJJIRYKCzDRCGQVqeXngG/V1fRAdLcwaDR363IzCSHZtFtE5GAfvYiF7Wojz+X9m7OrEen8q7La9
gyfQ/JDfQ90bJeD5Z9D22tqPDB7w7cLwiLgOrzHYErYfcocv1ItyhG+7qJBjl43AIvFRNSiBNyGr
lq9ZQ4FBnhONjstdB0ocY6+CLR/P/HDvF3gr18hkchJ9DKRoRU7CFGI1Ia0kJEnnZoKlusk8/XXe
5I26oRfrQRoeR6N8ayLpSvTeYP5uIXbKbZssUCu5AFvqVnN1OVvl6w412NWiDDwkl/2iN4O56ur/
r9eAk1VEOsp3I9Kn6dKQgLZ/jhPY9PlJ3TmvIR6BdwhL1XrePAqCqHH9c+Q5dMS34bmFsEJzVTei
aXJCY0uuuUSn9hNXKx2NI1ZdKTP1JSptqWnPUiHLcDc/3voXAXNaW/F7zmj1IHmGg5ph3XNJyK2t
1azHztoNKv26UiwejeB9tazBpGxBa/WhJFhs+OiI40KK5ezvO6wLsPbRmO5Rxx5RB3u7lDjocVaw
7JPJV/ggd+zDcOX/yrnsPD2r3iuk8bFp0Njrdy64uI+RnlVN5lapYYWtbz8HnnRcq8V0ZauCfwTw
JAiuo0sQ1wuXrbnpCZ7p1Cw8iQHPCG/SDF8W2hw+4AW0UxSNKBpE99tC39ZzCaBCWpqUJ7ukJ2bg
T7abG2lcat24kzWH1MYaSXaacL76741AIrVfya0ZeBe1687uQ1DbgBiF3IQKLw13ScH4K4or9sQK
dL2AANd1C45Dbm00dgBPPfeHWdEn077lajaKXrEHqCla/DgUNmao5TJyVIHfDgv08OEP7/IA1R75
h3y0haQnbnj0WubdOyyHNGjN8e4pbsJ4m0YUSNPR4RCQwBAL+Txy9IRMQHr1/wm0Ef5cPtYwIi5A
HHRzHPwbZRLfrGPzvY56aA8P3Xfdpzqr62vsJtpabdYufLHwJ5oHOPOF1/dliRi2jTd0MhW3CyCp
GJHDsuRbVjr2Sx/1fNfPumcpsvO7BrB48NZyr3hiLu35Ue4pmB+bbPE3fuZ9lDDkMZmtZxuaBBbc
gnoTy3zrM+tOZS9UmOzYLz/lX07Dhf+kr0p4NbsiRtqg2K9zTM5/snlX8TP9CS+uow2JXBimkFN1
Gd3IMElKAWBcXqttLmbaDqcmIfUjg9XXMdcVGoumAMHcfSV99SYgSdnn1AnXds8+kDDhFxYrjAWV
rIMnj6iv4uOb7lJfBO/gVzNjU/JqGIDi6I5TZe6d2LxZO/HOrlBngRtLut4+r1agMORaoeKQrPdq
mqrapWtNg1qmQnBY/xA3kgKEefI8bwM20ix3l0JmXVgmZg5YpPE1vGa/RyNvccmgMQHfJe1Mguoc
xBzno3X+jaXqxg8KliAYeFKtcxKhet8ufwXzScEeV/L8D8hHywE3ItEdfMPg9+EcJWDkb0u4TfP0
NRk7Sz+KkoatjlfPmx9kgE74pNnQLHSzaTONHZbHtKebIif1oFxQVkm1uHOib1KFh3I/5DGi58hX
+uaBtTBx2EV2n8lPAwgC9ysCnGcTpx+cu7piBqIaDcYTHzlIqHy61v7fAJHrDZT6YTCAzWJb0ng9
I2bbc2RxS14zy1MfmUTrmrEvRmo2hB9xuKjx6L6G+miZsDp2lANCZR9S6mKUInjcH7V8ilNXwSNv
c+VB/puD6SvqugEz12FugvtsBtnClWVloQ8vURxH86KYzIl9dnJlPgt6ldjPjtMwg6E6YhhWozON
7ysH7wEm+hyXhBpLMefa1VfmAvAalBZ0CioJ7FqdoGDlmn36yCKdA789h/se6wR1mrgno3VyFy2V
MTAoj+ppsffr/x1rftNB2EDvO76YV6JTJURjvEzKYfaBE+/UTV2pItzgr3P44kyGCfiOkefipZqq
Ase8Oe5JU7b62IqUc2qAvrzvuCp2eHqndBgR6DYUpVJnazCXPe3LY6nka6bmt8PVJ5ElPJaC78lg
Uq/0pewISP/WY8T/oNjkVhGIaLP+cbRwiJO4yiVBa/KMTcZIKzavxSE5CmcYrXRSJ8sY00jwNvCI
V60silDkl+jOBN+bKZYrcjUgrKXS4NthddIUwAG3xlxoELiOMJNcaEKw/Djlm8pYlMOypdVNn227
/sLhcGuUgkIErpu9/x0FKtOzz43zBfEfTYoF2TPaG758lW9ud4QthjvxROaidMZMfw19c/7LnPxQ
HKVgji+L47DaWLjQDCmJjB7OdLFwo/FgvFADRlRYsi/upyoom6j0p1gUOichw20CRg114cnX+9vi
DIVLL2OFyQq7N8n/pC78ZsAD+gMEzVI+8nwC8NbBHe8uWzBHoZAczhHyGYcmRG1yLj73vAOTMhQq
iWooYe0XctZr50VjjFieOuANwWHP5cNXMy9UIWkzl64IbsOaOAvv9zt9wdfP98g/eCVad8JAIEO/
HRAIvzshZSzDkOOFX47Z152Sh9Qaa6Aznbt/aoRq+OyHiA4wbu3pG+oIZoVRucZ5tJH/ePHxQKyQ
1xCUvuRTmoseWiV7NgBFkztJHs7TkHB1WHYkT5MtY3kx9gfLxIGAeV4uy+H1wPYM6TvnZtvwdHCa
d58eyS05e5DDYuaeVxif9+tUcD1v8964Q8xX8HkUOF59Xu67W1NEaWe3j3tyqnEydu3Wf542XpKM
PvpQAwDnZkXVJFQsByYExz0uJOgaJNhVyNDfV6e5DHyHfHo1h+RLASzQTN8jQSEZSawel+8YMFtZ
ncbFDkU+rQrbRs7MX7sfCwra4xm610DPtQ8utBg2DlYXjpRCN306GXzUeeqY5JIxCT4lHGD6YoM3
7hGsElTq95BKPkW0TkO5aKQ3KdUSnl44A1ER4O+1z3n7zYw1BNCD1I9Zz/1SX/mU1KIgMk6brhf3
U+XQDzfOpeYKd8GOgqn1pmMzfgbP96Mvnjk1f4o41pz5omEbzcq7sBpmKmeFcnjuDEaHN21ukK87
OILeRp2B0B70HMHWx+R4t8S69EMInKMNP5TjTLppMpIKg5d84EaQ0olCHuVLurDHe/ND9Is0X81p
9AoXyOxpRUJCb6nMX+3MCLQxXwhmB2866l9qQ65UYx7eE/BhKgFo78meAwTAZ6UQbX0x1dQAzIZ5
Vq3MYE175dgi4KZW2LVVACrMmJwPhlc17T/wnPyY2D5s1AshKyriHSsJNBHdBgdOKbpghdmyZdeq
p+LUSl/jlcKRMIeKhKf06WiCPAOAY1hrBU4ZB4xNIV9nO2w2x++8sUOGtiJ55fuENLayuANKHx/m
lUVeC7hq/i3861iEp+OEOcnIuKS12LeIupNdHDq7pyxkN0V3sKgggC0kF/6cUNECfN2HLlpBxW4a
k3HEs0Xs003lTSJadcUAPkeC4FeT+Fq0L4gM5LNzL+4IjXDJ97bDxXEubscPO8fjjPmozHPSAmg1
WnJOlHv8n3zqKThUwCSQ5lnZJgrAIjMsS8mHs2LHkNU4uFYb1ytWzYXUx1bCQARHSr2jmwLVRvKi
p5QxrbBqOwxvJYkx++3a+FcrcnfxlcSdqKnV25wnJDTGbWVEapxDxcjVFeRUHJmh7jf5lM0T2XmB
dT7VKFpN14B0t+t2U9p0qg8UKUImtKFG7+SAu4HN30+VAsA/vf1lAJBXsuETh5lvIo2snMAmO/o7
f5hIdFNimF48Tm498uuclUfKv0MWMiI/eSEH9i1x60jCwdEbg7OXVWLQCmHfAnniX83XGbdHrwFZ
MTLyPx3tkFWMWlkQm1Z4SFUpeRvQcTPTJUgQzP2wOLLJkECgld9msd9JC3eh4Hds3gsv4vDLLf+/
p0pbhNCdgAo7wI+9o29woULQhkpxhfXJHFQrKis6w8VRHCmDMzWIdaqK7AEizqfnNcpD4gDiMfWk
cgjQbGkPun3TfATWA3I9ZWaaCGLyFdYt9orms6symN7tvpn3BjnbpRTqDm5KnudWUCtVKBLoyIr/
C+rXyFsOT/NVh3Ni0diLpXLhHiath1yMh/3V1KX5ZZ3UkVFe7osb4DvQmHygQ/BQ406y91rQ4Cd7
u1rN/tYymuCZ2Qd9RcZ0oD/YyOQsf2Jl8kswTrRSjCYvMEKLiXjpU/w86oy2av+oBg1n7/vyU29E
11GyTNFMG0L8VzNaX59zPp0GzHLx6krApI4tv1EPvF6o7CfecKLSSX6jlNZJdumkE+/ysB/IF8Mh
yGFFAhBscM/oxsRb4cp2nm5RivOZhRhB2VH8GjAnCRzN0v33nSMUUGAygtet2xgw6P6IBAVTJZnL
HadtQDdZij3zL+XYlQfXPUCctjW2jZfgegL3qsXxC8IlJLcHNNCI9beuk93eGaCaDm3XUL6UPFZo
2Nwr+KIUXoBHpHGzhf5G6zaDFy0yWNLP05TSlMDTbpO7Ag4Pbv8cy8RXVmBBLQxsV8yGPs4G3Nvm
YC2X55HAf/a5uNBI3yeVRCVmpXUGngw7LXdYPPwXFVWpHCn1VAr+/DvDf+JfsUmjziGySZ4TLfru
FddaT4ZyMaKOC5e7mjMvm4f2La5lQWBYaSWh5KuReyvQ2MCs4C7bPRQuKn1GnMss+Hcpkw4ZBWk0
Lt24hNJDCKdnUFCLNcm6lmkDj8QMye/izBm/1yQ7ddkCNS82MYKvvj3vucuvR1uEmGVbwuR3OiIN
3Nu5+LoAUVN3vuMATYzf422yRwPvxlJELrBH0IEYz81mTk4tAGYNCDgB75HcFyvb2R+a/eYJsD9+
XUh9o3bDnCuoBclTxkK2LVt7aQWFUQlv0yASrL86IPJRV3I7cv4gZlMgHy5FR95LACAcy1YA0MHd
9vO4GI/NUtqs2eprEVnHd8+sJ42ywdnpFIaVVmg2XrX8oqJX1pCvRznrxE6a+GJEF4mfGECUEEwu
8kYavYSZ96DBb2AhrK+mByjtQmWy8DqTCtM69ZWRmBNVE08Ct7GT8pKvOliOuzWGEnkxHGXIRpFH
Y7rIhGKKlZD4TW7Uo/bDVLShiZutA0woyaQNOxvJe6AihmAKMAcTXSh8YHHHIagRqwROeE/45/c3
BI2CrRnIK5tiMeNbkvhh1YbU+2X6Z4Lsh+DNGxYGB2hMKEJg2fkDcCVAvUqme+/LkahjmY2omhZR
vyOnrcFLjl30/0qkKDEtTGAeLexoLJxMCU8J0ymLQGUQiwYmalUfn03e5AGwc97njI/GrmG2TR23
60kpchCEh97EgXv+VYWb3bNIo3OqAHgK5a+uMaWjHF70D73RX2IkGaTVlj86zTqjId3DnonS0VV0
7kSjSAKZgdLYWr0yuQm10GcZsMw4AmcF0PlVzNTb1qUGZi/VCUgCYEXgQ8CFzfQ1ljb5LZ03+r41
LX8DBU23LltgrowDfnohnxv+vq1dX5fdZy/Jk9Hc5Lur7Tm5XDHjutkDgnMPbZ6XtmNxny+oPGbL
xs5M0QPF8Lj6rIysPv4iIoKjTV+HJKPYuZVrWGTSr4uwEssbDt/Yy5mgPKrKh22aZJb08JQnC8EW
phAbJzY6yBmf6jRDmIEeGqTrST0ItSWD25Pz4FaLWsQ4VA1Ah4iDZxU5UxjkzicaGhxt9lB204t+
oTPuKqzxIehIpsCl1m5io+n3ZakvvaW8gezjZjLfhckR2xhRX1RF3LXRElRM0MX+Q9pKByYokoIT
Jha02+YbDj32/GuPC0q/YSGbROAA90QegLUOhX6tHTMzQ74ZM0L6RZhLQZaJPtjxk60GfSYEHF6j
+AbIgHqZOKxnbIU2hBezUV0m799kzUy75GF9z3k3rbKM/LztIg2wC9dk3flLfl1Pyzis1UOyCS5d
IeZqyNYrT+oKMtzFB4+iNoHL8ADaHUedrWK0Yv2cQH8JqC+HV0w73bab9mtC4cR/1APQ+ch/B1Cv
S+T7QKgwQTqycKjP3trCzBUBaBe3cqW6xNVNSle7pWlUCFHp65e9+59MFZES+Peae2B0QTg/14T/
v9jasYiSY337MAeEbjog0OOmF7/KYCbwQ6SA7lmicfIfLymSd0545i0LTZL2UdhcC4pR6Z2ZT1+g
XfbWIuvYHgygVN/N3IbZ7lMi5t3F5bFqsKZQnpx4n0mLqSJKC4QbZu4QNowoq32C8VlhzA0dXLyd
Nh31r+SFKmj11sXEC9ZHfivQ7Z52BH5kTpS4/UelkR4fGjpD0yX6J/AVVtw4jEV9elf5vXREXULe
P1ymngUHP78/fWpvOFgEIr4hvshMGdvo4ehhDJ6DjJ0BWfudKKMBhaFv+h+Vr90vy7EOewF4uYEd
+Qvprm/XVD3IDJu2WnpJ6lcHiIW2zw0noRz2VuBuiDP8h4RS6F5SIxROv3F/Xgl1azfPsf2k5pRf
xAbSemlHQjYqhN2DHGXNzcyab5Mq/JLjRMNzCHgcASSUXBW9qR9+ayw8kAc/L6hgvTKncl2jwHzJ
07ISkgpgL/xSxYFP7KFSxE1ahrd2TzRUKzzkqqr44+60Ux+PwVa0iP50wJFPori82YumZu3+m1kv
L8UIX48MPOLtq2uliACqvZoPbCj/IbTLZ11djKosAY640pv+NzQJOgiGWppuUbobXBWFGXuRIybk
Rt+kbbPHF14YnIOw3H2xktXp7s1YlgtxXFu7kj0Wkjm3evtpBzTRfWOBDkjoCQcGLKbhohijglEK
6iPJKxtLCm1zMqgTyjzaPuk16NkDpc4VK8bfxbnOYoxmEDeloUlqXsgQMMk2CfdVQPo8yrpoLKeV
f2PKpB3D6LrfrHPud272GtF+k+136I9Mwo2Y/0fqO7p0MQkRvnepx3yFQm9oyiPqwtk8v15OHliK
RJu3AUEg+hIkHrV1slSje+PvyZK938PGGliEXuSygJCKbii2nScjonEk0Ua0mF2R2cQVlQAkh5vR
+PU4PFrMv6Qv7nuhLqTUnhJHHd6+n94UFfL2K8uoFav+OjOkBth/hR3ibTe8tVpJEiDpCWnc8Slt
x+l+CV754lLUCIbN7A44UdEHWqBycJMQL3YsAdLjL/9GBDUCCYmpEqGPHZuUg3Py4wMv+a0u4Jhg
ryAcgSuTftlBNfu4CCOMGQkZPBGm7mqSkqHtjPaPbu/V9UEDU0Q+LmSL0eB/5SlguYKE0vSO8x7Q
qPgKGZL/nwf8kBZWvTG9qDY/DpVSftrlAp70xZHrfNDt9dc7ielYXOEC0Ybt6EO0AYEKvDNBLHO8
jFdfzbgZ0Nl85t9OFeGcvl79oowEPSx2FXq770ZEBKH2fPYqWIa86VP3SbkdqrY9cARtx08332na
rs4HsUceDtbiYVt+q1l15VsJQ7wbfx+tFMWPrZkZK1tZGn6LrHDLFX83kWCQlJAVBspCti7epJ7Z
2CRfOTckjrfEkd1ek+4xow6EkneG2rfJgGDA6H8EGJ7M67IYtVpeKB32TUefrmWfFOrXyZ5s2Oqm
7SXh8dkfUOS0YOyyqNT5bdd30wBCmYS3W7hZcCQytGwzOvVtPN1pMNQ3swtv9jSS3qSUhQCKIYGm
Db/hAt6AyA+zQefYo4eDTb+FL4t+KZGKo+tBDtSwEd6KHK4U1aXpA8nZsqIXLfchAvagZZvxdD+C
5NlWO6ANH8Pmm00bTJQfLp4Ir5JnVEQkJ4r5DLj+XrfiS/FmsYaAZxbhHwFMIy/511DGwQOGCXQn
r0zf/+xsqIfi8N/nVdQ6KkR+Bo85xwXpIMmD5bnoat9/M6f+AqPfkBPdAKl6eou85Gjt0c8Efm3n
rgQJtxWUiK2dxHX7bNwLyHihikFsQA+VhlMd+AxX5FyG23TDBAdfe/zdYzSkOdKL9SKPABgNcKpG
GMqL4pa+TOSeYuzVrnqrPqNL4i6g4+XtoMaw+Ix6vhMWhvwS8y9w7ZJd3M8Xnh00wz5Movnhpu6i
gsleaQ7B0EWQMSsT+ZzB0RHndT4R8obhyOM7ncXYF73VVO/DD8fQyYJee+p9IiOC8Kw1aGW9VTWO
lREICxE/I10moVQkEEogO/rFECvE3FUL7yDL79+cMuRYwIvzifduoqZck7KGAyHtCL0JvPNRB67u
gELC3PQOh92M3zaHVx6huWVU208PiCuipR1Wvg5683fYXjX0arlFKCuJSb9JVpRv6G6aNLH9HrOw
bp1YWKHqGt26ofA8pJP9eF5pWsGJgX32sbgoF/xis1aZGCZSa6ksK3l9wtu3UJiE3kqgZoFx8NDR
BarJj7vKp06ss9hiWQ4FP/GMcTscol2gMCbDBKeIXPlzWjuESBBkVYHeT9bRx+HGskK2+6rIUPsj
+OTJ3Qp3qaI/chlxaO1kljV/HF599CjwFWPs+BbE0V1nCs/Xz5rmAArRxqOutRaR6SJr7OKg+cab
rFDcg9EiSmFy40w24X9uzflZfRTSWW+Avmot9XfwGwftr2SG6ViXQ7ee5K6j3ySCfVz4UyaBApPW
jtc/T18X5aL1BdYHRgliCe2RGyzR0Lq2VP9D9Zqvdj1f0PJ5IYTqxz8hflB04F9OIhmP1avyncop
to2uU8qcNbnTz1jVsQkPIajBGSmE4coItISzUJO9vgHxafIzNjfnTPcNgtUYffD5jOJB5zYrqj6z
2UmhUwkO6hmnmx4eFj9tspWgx8a4COe13da00y8y5KZAyVk7osZbQQQTceGc4Vn/TYAWRHQq3gS3
AGzMH1fQSoP9ZOfryIp0Qa5PPc0gr33RuN8bQpz2fTanxZnVAVq3pbTObhYaEm22/vWSCWqM61Gv
Ow5UcU9C6GM91Ca5M4JguZAfo82mHesdn8hKJ6xTDFgla76mYT8Yd6lmb46nD1M5oj1Sa2CQfyG2
xd4s+T/rmEoMYQRE5Nu5mnAieCN9MFyH2MgkZX/qWLayQQg+6Hv1sV8lYBF57f0dMclCYe7oHOXe
axceUH1v+7oGf+XgFlwxbOtxyc6HzUfjHRP/St3GWihBW4YrTtwKrYEcn4aL9jz+cXN2Mva7e399
2wSR3QbY02Mf3S9whYNWQg/MaXbnbr8kLruUbTIrGrc98ouYZBmR9rIrfaZS7GSJG/aXCxX3yQ3C
yb70Xa7PvnNUpVIMChrhyi4Gjq5yrYXgcXDmv0AQozinb3e/ZvKuSkMalKk8mD/9d/u1XdUncmok
T/VP6CD+7RVNjChpvePB5+2vfgZX/wfl1x+lA4YqU6uilaU5a8DEb4A+33dwzLIWG3yWqaZwuaCH
TfHPJt2ouL3OhSMy6lO6qFLqkjOX1aXw5U60IXqICkTU/7miCjq+AN2uS2FhoxUhXSfQ+QxQXT/e
q9maEfkfqvnJNVuZ/jdRyEMDmk+GcriWsRFxBuBK8XqPns60ikdgGUQcXmRmkAaP9uFd+rcihOUX
UBk1+Mo/Z7tjhgXTYeHShYmv65G64VkIhgxm1hD4xsgRdpUntWpNNGU3TxsLDAd6yYdpkoWrzntv
pxw1I/QbGzkI2lx/wNUJK9ivlIqCCRyP+c0aQRA7ufNXrAgENnOV9SBQQnezD7T5aqiDbOAzOhin
EGY0IdAnpgKR+UCOQiyIKZI7RfedwhE30JHVs9Iq6Uk14YNdlTjXUB8hIgrgGryCJkk7Q2WVacRO
rdDkQIvLvCunHyHSTxlrSfEFa8p6c5vWRqT047upktdNu4+if4zRP386cCZaaqVsFY5A89So8Nkb
gdH92Rwre0bwjwbyFMk+W6/e77DWTrc832ptXwW8/ABO7evCW9UAYYeC/VRJiWvPZryYcHFOcLSG
ftH5ZKyfg4oNDC7C/BYb/5iiOVdaL2fvrhZJPGHAkqN0USwdTfM8c75YyL20da3hsNPpyeM6S5jO
HmxFw2ocH52B45U97uD9v4ouKhwRKwVDjZJ9hDoSPT28N8BoNWUhXTwuuUN8RrRXJfg+mIGD+Tz6
96OPXi1tL7aFi22dF6MKADOSApbZNEUiusXmk06pY87EMcm00q70MQKCGdsufV4wjIy0Zv6aNkku
dZRpqaFtQ4FqB7Ob95YxxwzUgpzwLMx1YEKTiyxokpaqfgekTOpibPjDbFQvLRE1b9U1o6YnF7rA
yq4JNzS/c+uwVVmSPnN3VSDx9GzVMNEQqGxd00V8G3xNQr5+ONs2yZiJ4h52+IBAGKdNzQOPzoBO
z5eB54uNIDmctT96SVDvE/qfDA6HL40HzChRQXnxPi/Vah1JgqUqeuyJO3MiVt2FbEQrbrFzo9Dj
iPymlNtuw98C38BoKBcgUi4mM4abwCxyPG7fTayKx/esEkWrXpt/Z5Nwkg41o+90Fh0hNaqsseQP
pe57y/qLUiwaf87+WcE9hb9tNK1HSOqAcLiO/G/4PGITsKl2jwJYfVlwjdkUCY+ANbmNagBdxtSY
XWz5cVBKobyecqpvm74vwef5UZoDTL6QhIYHF0cqljauqRVgB1q40RFlqAmL3ImXay+QkNuVy3Vo
8gk4Blqt3ihC9Ga9YPyrohLEx7OTic2C5fifI7Mb6xhnnoNoIGquY1MF6DJ0GwbEC0shdzGJ2QXy
t2MKHFUxgbna+i6KtsSgPylvFNTyjb/WGnUDW5RcBz9oDSNyhfChflu6RRpU1jS7OBYuz0UIfxvE
xFVa8bG57ccoqX57E2oDbcDH0uWI1DBb9rwBNp9zjC3tu+98nByLbzSffyIXuNBncOZMVAjJ7Mx+
YSwwnj7PQshXVv8SVoiMK4fWVTa3B924JuPnq3IlL4GgjP35erVPRZIR4Cbl11R5OMD4mTcWBhvl
DvCYvU10Mzq7BMo0QghnjUSzIJA4iAKW8SSA0vXO1rjRNTyf3NxNdT0cnhu5yHyqO3d0wjP6n90r
dMf6731uNbDuJc9jM9OouEoTqifKC9a+G1voE1k/HnaT6QU1weKb1Js6RjPPVU7a2aAnK/4fjdWH
edkYOxp13pn6t9DOx10n4pSBGkmbG0KfW30DWgRtMO8z0tjoT+tXPw5xOjI/W3jdJEpSCrZ9DpBl
jRsxfd8WAxO73d5DsL0DTtNEJS+4u2JIuxEe4umAAW3KaKCtOK6Mq7q/eQplWkt8oXT/2hgxVFp/
CKI1DWvjDt/4BRwcMK0Z2K/0J0BqHr8/KZr30F5aLMSE1ZnnEs56KKOT1acmAha6AIn/FcRYcBwk
ZoSNDke5KYptbIfnvGYfX+H8RfWsAAVfDPNHbnZvxZh1aH/N54rxQOC5Ax8eR3Dy4FumyL6PJ/Su
pESC7u/zcOPmTRvZ5Mmc3BvHQhV80J0W4+y2CXrfz75sR2Rigt7oUExzEYpno5BblTo/IVOF+Z+x
OE/ftCUUKtVs36ZR5AuMnhTfH8OAa+txa4hsnSovqeds5TJ5IcL+j+w4qWT+V0Xk07XjCeuiBgPM
VNB6qXuyiMAa5dWgSMRyP0RCjhqe+pR+Te85vAvS/TJKJtg53Fv63qfqC94ikWvhTi9YqKCXN4SO
M6YI6YHg34Mq3WBleQq6XN/YvN4+O8SR/mOGNQpO/R1U2ieSzwtvfP6q95VfQ/dd24qOM9050BPg
zo2aT/0M+56yabQ6MZa9HGvgwaMOG5t26mnmL4bywUEptrPoLUYrQOPNzXMLOvlfdlKbqZuisrV+
1x6bphSaocVn6766NXtH4gdWqflGEe8zv6wJCJTjCesW0T3F2zpl/2Oo0Y/SnJNd+W88eed61mC0
8UTBJ58R3ICsb4NNqURoi6koH8kdulw/rDOWH695TMcNXkQZWRXb9E4e00/Fj/Y3DVHueHxeP+Mb
DSu4sIxyEtJUyCTL5N4evSnbuFIWH7ySXCIRu4G63vOilUPGUicGEJ5chwvfZ1JKg5PnTxDshTtg
LGTuofIe/msTrlj327afI+7Zxc8tqLhIkVSqZoHDsDtOvPyU4iNephyj9ZEINqPjBDkUBZ34TuQz
SNQ+DJ4uwt8GvyFsBtaeS/wDQICvgvGQh5VJ1VdmkiGgQghy5CE3WTIoSAHhqBaD8yTOwmwbMHhb
nx72Ab0+5i2wXW5F/2yHGiYQjjEHEiPah5ENHDCpN6RoLDSDDYlaGohl2Jndgzlv+XMCbYp1HF7k
QWEamm20hfEc5KdnEAuqRh4WMJuXOZ0TX8sWX5sZB4JrP/RcpN0f/l4SFyVT+8BjHOQaFub8Xyz2
5/RWHfcQVBr+lSsZNbHon3J0HpIc1T2x/sY2zKjbf2koVbnTcUzCBYF8FVTE8lJ8yd0j51phsEe/
QpEzenuvcSn/q4uTk3N9lgf4WPrBYPH9nv/W6RAeGB+0uWvRsxOsPznWSukREcFTGX86ER/E0A6a
Y6BhDhzl91O3bCII0rCTaf22vbaMRcUBYkX4TupSDOQka8OXjYPbxrc7hkTMVY7QCpjpQI8bKh7y
9B63cOUUSPEpmGDDNuLn4MqUUPukPqhpIa3CjYpuslXF98oAfkewMod3uf++1f9KVEn/c6o8v4Aq
xgRVST2OkJXfLtm0NLFHtt9+clKSKCtgD6cFdAFnAHbE8+T3kclZ/sZrw5zyUtsh5Q/Bhg7K0QOJ
YTi9WYNSAnNkWQKhl+pUExd10QB5moo3jcvL6jb6dRW2amjgNV0L5AAoVr/hGeZ5MM6ACKS3b7PW
yIFwLOTPbgrrV0buPneYNnrVMk4pRDWDWwnjuR9m43WCTlAndu/tw50fQOKCSllRuAz4bOg1NWmu
X19h2yuaKkZLP4HYdaeXIkwkoo1PYvacQZqt8/LodwZlhmRd2H7DkmYwDFLVJ4n3T3bVFOLSIYyX
7vGsES1MQpfPoXOmO7iHA7yf57GKefYr6Q1b5RyI1nHxBr02dFyW26a0aY1oOpgWjzmC5H6q1OtK
o+H1Nn+38SJ4XN6Yaxpie0qRbqmAbx8N9HzFk6pQ8AVRG/SIBeu5IHJRoXDFXd1lJTDi112ZSy7y
TM7H1+PfLTlAffjEsR9bgeXaecZWklT7GJi/eg2x411oKZRcGLuZLa5yLmB9m4d+wf6MPrrw5IBj
rItKpxM7MUM3m3IW0yNHUtW9Od0DZEn4tYBbDQikncBcsKpQPWoTlv9u9sksWJ35Dp+aXgqbzKxQ
EL+aUhy1SQrh4XfKc9nUM7hwtn2BUSL4Lqzf/5jpllwoE2yvRkYo5V35zp5rnWLnAZDKXSDdC8Wv
JZU5J2Pz4qTx2Fc0iWu+jx8NpxS7Kl8WSRlf7gNYr0z5IjlzL6RVt8SOiBrHSnI9vyhgzeqdnuqC
DTkrxYeaYWuOXC97fACENuLk8e55kVgQRy8QMVaJ4hiYqpc4Nin9mOoM5QoHfvsUONQQ/2nPCeDo
HkWORM7e9ujDX+skVKySPzxcoTkXwXXlqKGoIZSgC8IFXOK96zQluMhNlohL137FmBXfL7DaXMm3
6QdY1htKaRUiQn22qQxBNLbSC1JayCOwY5gSiF62/IpAUdhTrcwikFBuj8AltmDXOXEavKhHLpaD
M5W/d435Dlq9IQkQQAznuwmLidO2IH46TRYAJbmXSDJj5VIKvPyYPiZ4b1vjTnWZ/deR0kyJ1jMr
hLsd6w69LHCvLxXmEYdt2IpasEvADLjiK7TxftApJTw36onXT5xhtW1EW5CN6P/GDqXV9bkuXMgB
JpQCw3/WZnXNJ2jD+9ctUgTOVRVZiOuIwijfcdfimi6a8ClBrA8sINe7LnNNRQG7MNwl6SZzJckz
Iw3XzA32BtdrGhpLi7+X53q8KXROMjQNwfAgADdmSR6vUelLcsifk7J1BCiMUJefqiuOeNux+GE+
JeGAPmL+cnIgmWyxXli5/wq0a5kUdvWm1pNpiQIcZ4k4mH2hABgV7JG4N8Xh52ke5nhJkaww/A21
hEN7yqFaL5MtaZiNWmgz47gGvyf2gPv+Thie5eiZiVIhgpw/i6WRX3uIMXD5ufngI0kqtP+cEJtx
5V9U09Ffe4nK+OZI4qgBeCJjae16lXoZ1U9Q+FvUB2hWvdE0n1qFxToilo+RKBDyYD3HMXriqRHj
1CxBrq6HpxS3G/NtnqU5fsrRA5vs6svFAkZoF1Wz4b3xQqjIoV1az19u6xUW6DgzFX6o8pnSPd5Y
QLeqB6M7Q0Tc/Q2LfcF2dLx7qIG3wMSqkIVnbTVIQaTQqhUua+vQXfdyzWWt7l1QaLg9FOFM7MFr
IWCH0+CA/VWEsgwapQsS9xmjVc5VwEeFlwUUkE3s9vyF0nKLo9SpXaJTbVdraylM6Nqf+u30gHAQ
5gaYDQDMY2R/5x7vfy0NIVgOe0uHo/NCS0iiOwAkEwl1KdxTU8xm9SYuCTBinyamOZMU++VfVIuw
ZAfybHNjyIfR9dCNP2OZen+cJuLw3OaZi1BsZULo7CyL4qW0GBVdusFkKuRKuSgBbwGVFlar7fRi
2DehhES4Y0QM7OJ8xVwLFY40Ze678l0AA5jmQXg7hVOWln7VJ9QzJMtcD6KAH5GgtKJ4/aU0oYNJ
B9+anBo6YfETUn1FMxq7fHOXzrWbLXC5GzzEd572AZeOEzGw/HC4ohmjCEv7VkJeguVu3FpQbrZi
eB5dhpp3Qx+QroGNHxsbkYYbbmazFkPELlqShzyB1Cza1NSu+zr1p0La1fo8jxYTQvkXGBJBNA39
npFslV0jlGXU4CvD0b+eiQ0DnS/ic5xNKjXUsGeAuWhMZDMhcoqpK+npD8vbWerLn85j0oVwOCrW
TJqs6FFOtQ3QVUKJoVLqltL7r/+rUrQoC+RuSMUxRePtyW6f44Xv6LD3XC6nlxh1ruLKpkkpTNo6
W0a0Cyel2sWxAUHQXTavdDi+G6Gl4bnzx92tW/roliLcZCfssVpQR7pifT+IMHRLtRHCcnqib9d/
vULlv0lJmyHDS6rY6Ws6FD8xtR45e3QICcyif2JG6KsyPICyPUmz3Si+MyhK5MPUy41KMpUCAVOS
y3Zh50PwPiZrpdC4US1jJ0t+8MGdbbZ3ccPbnKrScQvcBDfYC8haZm4dbf69+mewhODhLPQsAoJ0
9BbhOuDebpzcL6lRxUtgCkcxbZs1Nslmqklj5a92mLhDaebFPNCQFQETBiGqivUxKh9F2189OW+O
Q/SP7GMU1ugO99ft3LxTJ5rKrj0mSOuthqfdoZzKH/eEvU5+5LbY9n6N2f6iBfv2Tuvc17/lJdQm
G/WpT+xRjSTM6thNAOKcTlSKbJO9bxmvNHhyAE0+DU5M3wav1PD2pYUj2C5IgxBgKFWAH/UAgIMg
kBeW2oF1xOOLkpZVy3H/n5T3EtdktLtPBdyx0cFTS6qjDNhh1kL9nWRcqjU/KTXIO2zWBgK+32O8
B/9IKdrOqvkz0q1tSHcfsmAyRGHNZZDNRPBreEhP3PXlJrXnGB9i3bmRxxpCzS+t/IiN6LT1vy0e
XdVOQSR1ufcJSgQ3ZfIf/q2d72JoDp+STOIfZnh0/DGS8OO3fZPe/2Lpku3JJYHr/xSJ7IYLE8mZ
Ic1rKw+OE4Tydq1NSMYMRNxGVdR2zyAITZRbU3utvcC2onl0no4AyGM5WefInpjhH4izkUZn9K+c
tTcym2a1WsK2FAjbCWH/G+1WD9N0z05CBHtqZTic447AD9D8ZlszRAm/IcGzepMRsbEou5j9fqpI
EIDj0zJ8epDMp9ljknloW2+UiNYrST8ySokrnA5ZN3lib+RJAjHNtGgoW1UeyPnlDSG3FNwqByde
tD5XTLZMfgp8B85JcaS4SI9dxjRItEGmZ62qV1Kn28Qcv91cw2EXRKfDMoLudA7iBCRnNh8YauhZ
wxCHKZlptnjqGpJGGt79tibh1QdwkJgZwQmMiHGPyuxPuLmaYkXzJ4QMiAN6YlcnXM8NWom4VMet
Xal31JWb9yv0hr++rch3E/dYwUNSVJBAJ2/KYBUKOR0hn6oP9A8ck33GpD8d0o1uL+MMyX3LhkDU
4ZH8f23Yl7sa3PbEas2vpeWXLUWPXgdRupHpWEWtC+SzRI2P1Mf1QkLgKaX86/y/rvTLfyBgxuaa
NLTLqwWY/mpwcef+cFsqIaTAoQc8+kcfwsSxeSDW8eUD/uiTW0dk2N26Ud8dC90X6SZXp12y9jbg
B2qFs63MUufK5UR5Pq/mIEjXhh70QOUUNAiFFW9PE+rikFjox51VWYkI4lS+c/6JCiotQQrXTSi5
lQEQEPMbtmV35ebmpicMCYvQBJqJu0m5WdvdlaC4v+xt7Nzx1BAgo+e6ADiqe6eBPDMf7Sfu+jf2
F4BSGfqfKeNOcbL5g5yWwnerywNSYKx2e+xaMtv86uAzX/owk0yDpK+vPdxpC/DrWDz78MIpFjZ8
ZuM7W0zgvu9FgZH4Jh1xU/zI9QW5IWWKroSS87CoJyDVjIY6TzzPeGVxzt+2dl+F35yl84qWVijm
IOAip2exzFW5+6bFGiyaFcoZRWwDPqV57MrwOwK0nVxeLcPvQDNDxl9hwJLkzkvdhjcZEv94TZdI
iChDbGR5QB5JNDfS8w0S3NhkfE/24MSDy4Ryu61clEFeBwQJIqY2mFTygxnArqJwuJ+N0WIbKKFS
DP2j7ak7RvpIHbqiysx8xauqXMlpVq2+wFBa988XlhJReMuX0PYbio8zCOcF3/0fTGiPQ4UaazPk
JXAMRBl6Sx25LKe2iARdawXOSZNQeQmdefTE1aOnDG+fm0aRrsVAx+9ZfLNdw7h1p5LTGAVBqoMz
igvkQG4aOVHFYQWVliMyd5OdxJpBRznQx3fQMN8Vg3B4yupAM2QG1IymT+EPBFB7G0PMqyM833lj
lv7yUSYeNc2CANAh8grZooG5fJC7cTY2txgUQ9bb4ao2KlFqzhaEXc4cvh0SP5SaayVtYLsIFhUy
yRKELOgQmZH7IqQj0lhuQmNz7Ouy6CIPLqMWgAeBWp3lNyrrAHdBUizMNgPGWtGvrteP+abzCLlq
QrgxXUKhv43lxiMc5sFYPBhy8OTJVhgzg15LDSgUGHc4By2RKZu2+Czk8NUdbarkGjrM57JikmeR
KgPJXxItSVB8XcBh74p6Dby6O5OPTSjKEYaf1DEQ7u3ZcIq5Hnyx8oNcnBz894edbve7bcXMqWD/
E8tBotgNAyQezaTicSDOv15zfFa4d00LSPJo1w48fSbrr4aNitPgvf6d3OmynzhA7SRHaEdMK7aM
1671m9df6vVActP439B3ljA6U/nzSecYpdQ/fsl8jeIzE1yr3wgfPvPSs9QlasZz35j9MymIdmQ7
Td1QF2mpwORwqMVbiebU0ncBNXkZkmIBlz3gTlBcPpTklcwoeloXf1DR0WSkWChttMXEHYuCKUWa
4j4fhYB5Tfc1WnVLxD2TVdhmy754K8P3rrZKDHANBUGEZ9XOfFWFgZa2wjwfwnOiDtql2MeEXZJn
C0YJfRMQZ0rFwIM/MAP3Stw3gHBDFeLtNhhXDJhXvsjbXnaW6WxR0WbErXb352z1LrLQDVu/bYvO
jfp+cHZkePBzhoOvmDJZUgFg+pa5YyfzH9rE2T+Zx9rMdmeC3KkAXU58vRpJdrA9XdH1j43j4qXI
6ZIPBdlcjnfp2ZYhc9ZeyZs+wXAHNAizdVkn/A+ntY/TTatXKbm/mRxhuWxZPovNRV+mQ5HQNsYV
FVMPPrcxz8KqtBDRS2M+xxQ5BATHeCi5iDhOJ/iOG9aru20ev5q61D+gu66KiKvnlBTunmsFveqz
1hk/toR9ITW/V3ooUNaJweLQdxdUiwPjJXst+/tuhC5zTECLElpP2OAL6NixHtoDOJqSiMDG7t7V
lZjR7jqeIpa2ebphoE2Ffzfc5latPJkbropWLaPhJPSNPP6jalEw3Tyg+q0CbpffC5tvl5xPKIQl
3i3623XGdQUjXb1P6UgiVrwiyPlp/rPiNwYbT7BZC4sFrrlFpnKt+LQsCP0bBcIZTKOey+v/Llyi
dasBhd8Nxdm/tLKkn3j/8Jfc3i7sogxjjCxuHg7uyIdNNdjZJdgu8WTHugb6s8LCsQh53zEQ/XYD
Ss8yd3uVUXvAmioFgYoysS0l5UoPs9/kznqOzgaSRWjrUhFeP01W/OLhITKQD8b/NGJH+0yLvIWm
iS++qO8nK0tLDXribbmtYr51+qSbkQxTjF0QdghEdTjo+7W90WoyCrxm5Lm7G48I/U90S6mxY4Ne
wbZ2AtvDPpvcuVDzNRB1jAIqftvzxjek4Yfy2glSYR77/QavjkWI4l0vmmCGzNkpZRBehJAOJ0LF
/Il3jQ7+2NB95JadKXZSZqoXxvStiXmEtG7dGd4rl+oxERYkpERQmAxl5U5eLyhipKIbGVgO7bVw
cmDFvY47Dtj5QjBgclYcX3aOk12K4xSuQLwXtcPuVV5hSUzDhTc99YlEDbeh+KEFNjVtcVbJazax
VGhvbrJKy86Pwd8lu7aqfae2TY6BKRLbOnyuIo5XRoSiSrGMDCXXFmrUODFW+q34rhmQ5aXGAdbh
P7JzVkJLMiXouOkT2WSU1T7diCNWM3eWNrVdmDc3IfVYJxWt1Wn4qiVUUdc0cLVvcnkwHSaCskP3
TYteB7Yc3f8MJECtX3PCqmWAgv1lczeCj+SXupxDP7/0+46xyV8zRUCvngm9qYG5iLxueGD9AgZn
pJPyNeT07NM6OsxafBUQC85p0xRmsSGg9dgy7x5vGiXkC4DFg4I7t9QdSK7axBr8wmfM9yPR24VV
zHw41YALgVjRC4xbzJ/AjOMvXCTCSOIo6xUGQIu271N8O9wGdUhrI6MJXy92NZA6EOST2ZvOS7KR
H7DSvhI9998xh6gGCZHYy+5ZzUoizJjG/AC+zzgd0dophDJasoEjcmCNhdAYeqvKr6Z8urL+dmDl
X7+U9Pws6qOEkse3MHaVDEoaX2pl/QalDZELlKa1JUsL6jnTXydG0n6605rcc7Zpe1CcjWGv6kKm
TE62Rb6dt9bcT9+bkyupvLF3fEB5N4Vv3c2hORITS2EEirj+xdnvoMjgol80ZwfTtZB0R008G0+1
OWJY6O8y6xu+6joPJTO5SdPutF5+AqOz5grC70daAS+RzqOLMHFzWbfeq1+pOoROL0l90zqEJARZ
tmK4k1BOekZPFU5xcRnOsCEWkSRCfQQI0QvSd99nHRJqxRRtTrzbbeZeVU/mL/CMUQMxSkNr1g8P
NJYMDj2fZ5yeIwW/Vl9KZ3/P1wKb+ehmphXaz9mecf9FQCzlEyBCDejvK4l7zo7/yuWHNyiGWZTT
L2FFaw3qrpSAravu3/LPaDusbwJU7woJDXwcfNTcr4nd8F8fUg0ACh04YV2HpETYfdobYC7CF8jS
1qdnfQiO9q4+3pBUsJVFA/m6M8aUuqx9GaElvbr7f50umNiZ9kGRzUhpYs0qKPr6WFaAqkn3G+wk
Jyta7gAmVhnfWivVODg7ofdSf/6HkSfh4oFEd9WAzVRmuH8ef67lUWAbPcxmpVtZplaTRlt3J7AS
KA+zwDldNxnZn4lfbR5O9vNIiL9bZpK8xvtVv3/kOCIWxUx9USV6YQInv/VrEmzZTXWKcmA2gtLi
dymWs5tCM5/AjhTSqypTqVYEIFWXomYNoFGF4JapD+VSr5PIigfdGYB6O2Cp/RY/28YEl+OezTEb
dmxJX/HAn5JVohsqCODKo744cohPE7NdqylYP7UX/52SSNrlzzvCqZzgvKvdQPtVfD64V8MzdFSR
XrjLgMcrNeyFNKJeeYlunHSsqJo6u2uCPl57ZIN9EyJu97LBReyeeUOra7zOevt13vjeoTxrEFHI
WD9pNdxsJxooesyOad6W9Hi1qEpbWEXPT1yWhdeMkkP99RnPWwLsNVqbFejKGcanjFcSJxzWr2Ge
ivyR+cpZTa64VBhv06j+XXeGiUtpizbFtX4O804hUp303yQpHK8mzCIt30BJC34eQskNFkI8COaV
Bs86LQxk2TRUC6LgUeDZFmK2J0iTbvEHZ/Rhmg7SB6n3hzOZbhZ4Cz6nsdkAGD8jGXgI87bqgrbb
2BXxR1s5vbW8HNBWtvd/TYGRU0D658d3z0QUEyUps80QNzByL3FSN07hnN/tPxIpla5sqRPeUWCo
9YgwksZvs6kGOjmyvOdfX0q4gCGyr5bVM8yFX0qdfY9mGC/BJx3v+lnKorzi6QHsJs0VEq766zUp
d20OOH4nq7ZzCa6QwSSjNIxFnctL49njl6PYbmQ+LaVDXqZUEfhm1+H8GkxPaPejI/jX6qKea5t/
mEu9JSQuP5CLugACvkfbgGgc0m734WAVSnSh8iLhU0vPMnOzrajHc3XV9lf5EvYSqDuemcQ1d23j
KKjdCUgPrQ0W11JiIGgVn9Aes36nO21IcIZqWMgOBbKG/sl2bn8azVnX6PTz9Ejg3kViy7eKD7XL
IbjYQstFIDujJDvvAvDShYPzR4AF0PSdfbrNMJPkwLsMIHPW50VZOpOG/mIFpTb1HK4xnyvinWT8
JYnpVhKLAq4prJ2lcCuiZ6Sh0pzifCUc2HPuQmaEXaXC2Nuh7aU+airjUETCpKj+4u/bh1HLVvRg
GFPHrCqCDm+EsyctppYV36Jd89UwguMogPAkhj7+C4h5vlGsv25yCoLp+GW/3KnrdV/lh5SHuknR
D2ppzdD8nmnwzyPFb95pxvCqI8liWNu3XZp07gBXchBJn8OcvBWISOTkIsOo0msWuGmm8XB7KfJc
LQQ8efac3tQ5F0Si2dAPASlYyCEprnMNoMO/K6JvNTWyOgz/lj7+2tbaeJyMI0pfWPCzoVOO+iRR
7Fr2crGSZSWFFrWjPgchl+d5DdtvHZ/hY88pYfkhDH7uLNpX1rzFd2t5csSvvTbFBo2zHjhWCHZ8
015kiSRbvP5VhvKedS8X/hULkxsZGL4Es6S2TBtNmrzAYN6fo5E/4d75NxCS1cxvGCeWm/wVcW1A
PDK4z/gZysqb0uxkgLguDFVbagEEpq+6IuPAWkFdm8UPLVevLYAqAk44uxoL7/QHLVaTs8pNCICk
moFKQl3SIZaQs3PbeNkn2VwhVKU07/4tzxBG6uVdIMn4lxOmf1EuquZImTL80bakYG9Xe0oHAbv9
iAFMd9w4PfupBZ1BHCtihLJWdUVTsBlOUDr2DsLSJf4VReVXKJbO0YATLQmOA17epIJlHZ2iuV45
MvKP58NPvl1INrTouWNX8f6yI/6Xf7lO31DYZPoVqwWGyBHkMxf+akQbNFY8QAOkkBLh8y2PW8L7
SzBjStCo8WEfdKp4kV6p/IiIQUl44dsNNTCkWdM4wLpB7rPjZm/n4qdRlblh3Z2Ix6VzGSX0PcDt
LEUtJdq2WmvcSaaUqknnJ0mAadc57y6q2rqwwV99pPUvP/7D0GOAH7Fc+ReEBILJKyBEmYPrF1cY
oOhkaBzVI9j2QKIXUZly+7YDs9OgrGK06qxWLaiwnXI6/hC/2bLdF+/xrtvYr42YyCay89FCkoLU
YUaCH1Tbrue1SY9BG3Iai8zSXbLe0zqhLdrxyMkZBo2sr70sTSSabyrsRH8kF54ygiUVBE8oOwac
WhJTxWYHyGRuGKNcZ4f+IryRmagdKaQe70jgzFQquMCQ2WGdYFJMcg8w3XndY1/Dy+41+bmftyzV
957nMkXzuj2PeRUU1rsn72cNV+mXXmCYSsJHH+KExacIe49fRvS0hVlVzyiPMSUNVCOspeUGQSJB
OvCicvpOYlFT9y2ohEpRALIljlfbUZQDc4IA+m4aCuMwUubl3PIz/Sch+WmAd+wlMhlrbdZ+K/MN
COJuxsSae/gJLSyfmsAsmknISz/6o9XP7NjjNaMEGNxhrsEU2JMMmisXUzlPoNe/s8BrmFtrnLSR
i7EcCwUDztrA9PpjXmmZAyzquher1OunGE7aqs5sHmingZcy0wfCHEPlLZ+qolZZMW4014Ah3ZQh
aNYGD+brhCjZcgizXGt1wtiWSSe2vdLEMvFnmQ9wqRh7jhbJlll9pYFcvMFaCEqgapvjfUKbdDhf
IM25+Piis4gR28SKkG1sWv1fsM7R7yPxwbZ9WuMTBzX03+RTrYH6jGTvxNC0ymquA+r81JJQG2pN
2TB8Cdnk5RM20U3tmHR2EISGyKu1W9izTpm2+z6VX3vdzNFaGaEFz68ubvUEVM5a9MYmDFVICG6g
wL+X7vQCKF05LcsSFklsXfHiZ0RO0v2tbYBqffQqFqrMfymYeUyLZcCBgxDbB6PMoellARr20vCg
Kz5LOLpVicmsRZqw0MhhfVLOt+1XDZvhKKRLoz3vx8Ec1n1KM9zGCWYk3Hkn9eDbHma+0vWjn95l
Ld5PkEYeBYZ2HvGjH+1zCSy+wl0w3dXayybmVyN9w0d1PrkYv4POOt3MEchkUav/nRc4Va3Yn8ze
e5ZS5+NSQYeuUcEVvZG5PklSq7b7AytiPXSz8E9Ogn3BKfkYRvB/3rF4sP6IYGPSHC2/6ziWLFhI
flR4lz9nHHiJ9QrrTPTV8V/7Fe4eXaQwhJcsb6P2CjCNwvnExP24GgkaNOC0rtlxpRuyQvGFWZaQ
QBhoUA2afRy+G4k5E74zTeqOyPP4hbgvTILT28YOhYIkhwBmVIuJBIk8o2W6i1oJQhjDcMhrAS0H
DtQcxxp3rJcF+QUtjaRZawc5g/L4TdC9JXNggCPILe0yRNMxmEn3W72/7lb/y0oE5SV6Jrc9tUhm
Sb7BFIVQeFG/A4WHMyiFCHFxIUtEuhg+Xle3w+7tVfdMyspLlYh4Le8Hvqw3/Rt/RhTSK9Dof9da
UOPUmno0gUgMdjkLpx50LzpHHpglec1heNKEzUjsKwc1tXDu4CzSX647i/ZLSE4v79ArewRPfWmd
AwpVDV3g3GOxXXPFwFyP6D/g17MomSTIk2dD68S5vHpxZPD3qRwhHh3V1FO2CCNPO+whZM2iXvPg
FhiK8+WzEtSqr9M7xJlIjJm39V8qSPBPN/TB8erpCsbbSkUbz5dm58YxgYg0M1CSHOuGjJ5Iv0zI
JzUfsroxpsznQUAlXK28q+/mYK5PxdnhuBN+MflxWc2eu8XzTfSf5Fg83F5cFCEr4NOQDW9jNkrX
nbDu2wyXqyBpVa7Q6m82bj2YW3qYq+vOzyUOAL0Y3yxd41i6IynZKE3hz9deWzmT6iHwh4rvvOVu
zg56KVsxQBkDe7RTuB6LCrnSWKoYE5/wMToWKD4rXkPiu4ddJIKs7DzEFW4yYyNpLPNmFkTSxm9C
yy1ARCUlF3wJx9hW9lfq24KSB5N3aGXRuwB35e66tJmnxjORk0+ae1uxKcNEtZtQuye0KhghZX3+
M4lahmaS6y+nilwpIkg64Ipk/NDtzhxALYUsE/V14xnBOJdr6O78nGthDSNXgL7RCDhFqCK+X5ou
U/7zPPGueiIs3lvA87HJwTnS+v+jI18G+hQV2BtVo2IQXy3zYwwHHUqgenSb3oQ4je/AS4rojWlv
FvwRxWPVpf06HOdptxlCgcYw9LvKH8TLUFXKPnhhQgomrvDSiTyX1b5vh1IwDrUptgSuPOmEXYwF
yZgTMXIEcpEPjZKi5GTxx86yY9jWm8rNydWSc3IwqItBopQ+8wgFQcrOZIJG3uN8taUFD+JQg1s5
uERDA1XR9r8fdLTA36Cx6My6Cq7sKGd4B02E9UejHyaW45Ue/hVt1At4lURjk9jbj7/vLOiRvnas
a0oQyFlogoKrmG5i1vfsyUfr8sT21wrczui3uGeAPBvLG2XHY169yogoWRhiahGn12gdcJK4BFPB
onVrBJ3QnZ5Nk8IGWyboUybIQkhfCPCcg5iLNBaKJHuBqjKYUpdsAAwKE2oy9goQKx0EaChsUUfa
3/V+gxbaMt6kC6yzgwd/8ZsodCkJp8SJNaQnsfXTX5i+bm66z9Fhnl4goMrXIao9wVtk7eSfBdez
EkQ71czaucSgbbTuWuN6MJvjiMECKfbt2uSTdmQ1xiKaDMhIMyXMcYOvF++FyhmazMAHk31w+XGa
IQ4cxifR21UfdRZrkp0BPLneGuSQy1W3CRF04qkEfgAOOnTzmpZvpsFii/KqOkmN7tOa4bw7FdbC
jdqtDg6REbEuG5pWHbEOKqO24K4GHGXMXeHLp76jGIMqMx/WRaFAasNsTz9G3UQIBldS1/bnkWvN
ZU8dAvABLHFKLZaBD3qpSwVFWr4sK7JQ5SKNY7hpVutjGem8fv6h6WAYCjRwO3LwGaW/Lo3F3sCP
VNYmOq1qby/kc4i14UwfCxFFUuz3SZxNEt2QZXCV69OEEMjGN8g15kJYP+Skq6axIkajnPcsSbc4
8tDzTNnj95wAUlA/x7tUer8P8eJuy+sBjv7klf3SpkXaABUyT1+bTjNKPGI8KUTpyVowH8tZiMvm
6dYGc8ksvjXOwlj5TtftU8FzurK1mvOIe2CN8gb7cQs4oq2ROXRvBfoeze0DHqZiu8Ydap4oyEWc
vd85Y+8d0qS1RpR1ce+UjHWuXIeDkKOAmG5P3uqmTWkoDf6Sj2gGBYQg0tjoVb72xkm7PWjywRV4
Bzqb/O1CjkmVLU0KtP3IiaAOiu9+Qm26pBKFe+w8Qg3ocr6dt+p1V5SuqtxqQX+Q9nxHQep74vx5
lmYbdC83gpC73jV4Qd3ZmxTPei+vVCp8Zkryn+7Dr48zjjC4sJ8Lvi0OWUKGONpsuboeOyB/PQEy
KLq6zsgqANCADnqcT4xv3JTk8YXSsjNiPfBT48XNpeT0lpTeBqVJ6v+qk1GA2QEsMSztGa2GaStE
Qw0t7sFUQvaRHpGtLQ66XEi8ylkE+0B9a6YBQoM7zEAvd0vw8DB6N9GNfPL+gt+HSeCZjGFnBkOW
+wMXuvmpnWIRWeuoIFh6gh7TisFeZaTxbD3OyM5V1NlYMMvs1CwjtTwI4Ql59XLdrv3ybMboTfr3
eNjrdY25N3X0O6ikh1q5IVZVnjLt02914+G9rm5Go2G75vlj2B0XRHaliykM8kAggO1QLqvAqo27
NJMOR+W6x/Au61Ud1lqvYmLgOPL2E9l1l4jNgH5mcePClnrdtfSlfp0aBtXA5jiDik6z1K7irP8W
TdnnGI/M9G7gHBkA43nmok5XrWVKA5YzO8J9QmEOugNoA+OJiFKt/jxBM9dycLYRCzaUfmny+05I
mphIU2pkFCHE9/jqWojWxJe9KYWt6JAu1ZTipb8gCxlt63NK90u/dsflDyRBylB0tZ7o2uLVRLkN
bLht4mhdwZ4PoeNRIhFKvezsC7ApjobQMtZPXfptzwfjosAlWMKuG6ZDZIya3tmoYABFSNM7hr5s
HPNleGW0FUpgeME55x7F0T7TSYVe0Z/1x5EbKg7NlMTWcKzLraUsRAxXnE8bl4ujqUhc42PZHpit
l2RNWDTsaW4xwd/4bGnyJ3oMHfYzzx714Vthq/EFpqz/VS6WbUW9O4WyxJXw/PNLxNRtfKD0w4/9
O4H/Jxr9lRyp/aIGMsFW1xAMrMPJ8Zs3MWGsWR/kEKflzW9uuBXt4BgBgcFX9wMQyguUN5dQLcdU
RgjQoaqCSnHKa09gg5HdvU3dTWCNvjxu3H/1tksad8ws5ZZubTUVeD6V2WPW9OUAUf7IWZSVbK9y
aYRuhrHH7O13jZMcDhVQejVvQBanBjTd2uV2mdEsebBVdKYJuOgUcOYeea2LT3MKUqjYdoOUDnDs
FPF9TBWTY3Py1d7DdqqlLRh5S/VfODrHuKJkHHzqvL6J7ROKXhphx5yCI7I9o8cFzJxHIQCpPHdp
ORHt5UsmjE+d2uEX5HYcl3ZlIIPTb2xq8/wa4yfO8eo8hTHwgeNNL7C6p7x3awIurJiBy46d7xna
FIcByoJhcNH6KMEKMzvpgFnHecNHFrg8aTdrDdGt2tqmgQty2KHUm2w6QvgYK6m9QgqVLocoumQm
tRMZGjZDSC1tC6KxedzzLCX+AF0c1511+1Tvj8g21G5GWwCu/08ciAC/d01p1TuYMDnUfn+T9N+V
gcNe8I5YfVPTHHgSYPmtWBmGXDUGnFsWm3vmMESWFrpXrca0rsfyaS7pRlryG5KCjcuOWrcRXRko
7phHtvkujpdfs56RYgCJBpNgbyAZmqssIIjiohjx4WtpKJz73IzB5IFSAB6u3ion4FgPZq7/n3No
UYv0UfqFQh7njGnLeJ/7v8Fo+6PvSN69IGQ2+4HZnzpQsS92q1A1gUJ41G/+Zg4WtB76QlLRaWrA
MUUccFqa0dz1UDDmnLUalWLFNcEq2h+l9OOEfB9uGuaWctRlffrP8PDmIqriQl7SRC1/vUN9PLbL
h7eA1N3Der50vnanPAQ1ixBT56d9W29/EhjUuCmvJ0E/lfLiwRca/BwhRDRiWY8BMPHiT6qEUp5w
ylzusiL61p52sbMyMY4DaTjmt5MyJGET1FWvqAmgkqvjWzUEdpcyJwPQH1vA7KF7n3ajSHOIoCTS
mhUmAgjXNR1xupvE8SrVkwyg3/sfupx1G1cqyJeTznlgqWHPYZt6f3ozV3pYfapXFkI35kXdHOV/
XD2jm6TKKIjFFYZq2gz3BobIBVsYFHq0AEKpLgf6xcMWSVjwzaTkiwR6ldL0tXNNCmnbaNk9EHuu
XEfG2g53SVpRvXkHBOCQ7mpAZs3dCkO761jxlEdTfPOUqgujONfhXCAhTdKsAj4eo08dQbmLLHeN
mWee6vJGoUo6j2z/vI58qnaUKTEhRxorcu78C/JfWEG3raD9WbIGn0sQB680ug/ICL46yRbkONWM
ha7Em36TF4wQdODziruj1cRZXI3vS/GzeRPGUeTCb7yqcB/3uU3uiNDOr/vyK1aL/oqY4uEdJ5S6
txUYB02VC1BfbKMnLrgKHfv35Y6m/DAW1B4NmyDRhmIj2dfNlTgIEpI+Tl5TkYFGMf8pMaoSmOEv
lDBWUNjilHFgBsp0xxGzFLGojcaoLqyZcdQ6DN+o4UwlfDGapeMR+LjuBdvCcnc+OVJSviIMd3hQ
FFrD4DvEjKDe6DBh66/ald4/nP88F8DqpZ+l02up3MgDHqo+K2YJsTuBpKPtQAU74pmNuJMScq0P
PIVCQJqIgTa3HNHF53PEaVAi6ivqkZvVz1nj4t68BblKD3Jh94VGi+5YK5PFvo6C3vYsq4AtbDBy
O9SAxqeMgakV+ce6iupXch0rozFoH1MAzqy8Ac+I+Kt5y4RfysGpSh+mOgBn8SE52p/maNMOEPF4
+bhYF/tOuZ/bub5Oe6iZyyKwLkgRlzqCSrtS20aobAJFUIP2tk+zHQpE1AhawB9B8J6xI/TSLJ/7
1piG9tVSz8XMB4C8G7Dg49G2NLgKa8Qu6O10Y0G0pTJRp+WOfIWCehn9CzV/1SobhfXQfUWhW0wx
IpaTxz6eIVCfpJpDciHRqLqo0i3B4pUF8FTPqXDTpr2V6Art4MiPINlvG+BodavoGX2qEafP5Ewp
e5H4+oiy9HVbCRdLCIV9Z4qzg2yJWFpdNU6SyQqR0SAUFTeyCInczcWF7MI61eSPS2nUfDzMsk1D
8yfBFCjzip9jYEzxgwKgFeOqiiWyBIs6ZEl7c6Q6tcE5z0m8VXEaWm9f0E4BE+YPs3KQDAp0khCB
4EHaSZxOb7Xo675tSwdjp8XHY6WYJ1R2F6t0Q3wqKkmRiKj9PXxRLqBVGmXoTIVLsd2jzdBR8lPY
eaQHUV0ve/pdsNEImts3AgQS/909RVF42XNwQBwprE34w5ITz1lAqi7bTtOid5KBAOEfX16Es3Vb
BZ+z5PYctqIzTFPIrE4qrm/YBR4O1zoVA44rQGrOFrx7OVdGmOMbZGzbcAoh5FWKXB7eDLTsveSd
WxFGn/74c5Ga2HpowDh8TmkOJJs7nm1Df8M+HelSR8o28k9s9KR0297Qi5DT1yOGRL5XhIPbLC+e
RUPvfzqqokaPcKx9d1DXYyyi8k51oUnD74C1qN1j4ByYgSKg/Hkcy10alt06ARuQbac1YbmK4/5s
/8aKvc4EgGKG2jQyydWpmbJxtM/zLh+dNvKWHsKNH2jB9ehI9XJIT6kdaw6/2H9oop9Fl2X7T5ns
Ys/HKcj1+gPAFbQRGlLLQysVlrJ2K7FKDKWB3L/WY7F4k21Za4KxJd7VSMtxlApgXntOkBvRHQi4
6VyT20wbWXwfrT6JjTqSp6epoDxChcuyZNIM+mDTOYtpwJmhlA5kFnRau+dPJ98BFdRRDRFV7NoS
PP7t1fZvRQTEsE+b0f5lHO7GzIIq3qFyit4D+CLgKIf1SdFW4QV3bZ7013DLbu1tdAbFee2HV2j/
zkh37QUt9EMM4yRwrN2ucH2C7Pa4iC7DnZTPGpTI2/SnnO+RM6J7mgJ8i5NWfGyrThrF+JrhtQyO
dtP1/xRf5cRxCESjoN5YFSTYQNz3QHQl5yvSVRWKkynQ9Xtkuoo2pT+Io5DZ4kUlbJCeMMFSFFlN
wZLRadcQr0WxJuVhXFKLGLrsuHMfGC4jpi3tKCOYLJ0ljvEUVf5NV0AdEltQUz/pRdxXBK1fGnoL
Gf9hAfaIFbVsoCVHt5Eg5zpXUna4h8+bKRiKslX+Iv2RYagoe8O0hA0poQj592CalEJRevUcESN4
clh+2g9r0LXJRVXq+AOGQ6hNvHXcY2cThMVAIC4gJER1bp07QgRvwdszB7KTkTKMdRB3UXdB91d9
qum3qTi6RjFdqCYuD6XhBYNfc3+hDF0cP2HTAXfZ1wqDDiBkvhjMtzUO5tiDIBCec5Zf0+YeOCiA
IidQ0BBpVXK+zTRcJHvMEVmo8wSTrBETlqXaHCTYGJY5TRs9EIiiNs6zVZ0rkd27Pv4xA0Ur0pTt
Fw9xBenGICYWKSSojIvin6DNG1Ms5RdftCAfepxJox7Idu50eOCDHn5mlXtUaiOczOsTAfw1hV4v
aTJh3cFWmIq8aT6lZubnh3IcioGHMraP2BB9RmeJ/e1yqJzHXgIw3YU4pPsQnFdWzTZsTSpXwCwc
i1UxAu53NRk6soKNYO8xKHfnT6lc+rDXWY99jolQ6tosFvC59ND3aMxuDYtzHCxL/D1joJRM49Y/
oJfreYzXhPL+7FI7PfnArkuRiHVoB93zL4KoaPzufYt74kKIxkXJriuxAOeywO6v2Y5BaCyJsLxY
DK3kJxFxan99+dgGI0CeG21yt1vNTO8nb7oGlvagKSTJDQu51yE4SNlIAgpWjhKqakQi+L6PwmrS
KqkydQElQniM/T4jJfuXB+QQlymYjkgsnt74J7oCAghdbatGQaG7pAJghH0zGX6SnfmszF7QavFt
MXBmAa/WmzV4rEQ6kKFFSR/kSCUF5XhRAM7vZl8ZCZLIhtI0JKmp7zvjQriRt2ETUYn/TPF7ax9K
asM/Xuu1D1fT1QwkK60GKKyZjcO20lFQhCjCHVnbryk22iO/N2+EBvtMlAWd6E51qWpA+fsQTmIr
alJle0NUgxCYA7/F8ivSrwLUS/6wTnjVFDYtTX89eWC1sW0nNoL0ZmhJds2gn1na5VDqT2QtFpPm
oMWi8Ym4GC/miCg4pn29O++tRVjxiFZCqQxr9y+E3mOsyBJt7kJJmbnyDOZR4MHyE6cIjEX70PcH
e6wGRNzqTTDwWAk2R83HV1pmqio+rSCn6Jt5C1I4+xaB/oFu/Ompg+TJir9GR8VE/LI4aC4yKGA0
B96+dQaaR19MryLPffCPsfkfDtQ6YaJ5IATU7ep6Wo76WGH6+LL/QlZngBVIRVf3vJpZLPsfXcS9
HWuWpiZ0S0f7c4J0eumkoI56Q5M3R/eY1EtZQecBwNOAoqmlhvgDvlmipLLWe00Jvqf4xSpH1rtm
M+drvOAlupADlseiHDhqAn6gnsgK04htDyQsW5RYxF6VuMtOL5a/ZDyfBLhRWUwbBc0ZMA6ZozZ0
M1N+Z5YEp/Q0gJCQBE9bh8X7P5nwsjCxEiiZXtvWGp5vPFN397Cy+9v61AzPMBzVdXb7lFqhGotl
rd8a7TgebcadsRsbSFBXb3swasBWYZrXXatmyA53wjA/coY+nsyiSptoMmQ0/sap3DeRDzBF9y1c
/P3WqqvdjanH3YClQAIAzZVdyi6mDWOrqy8HU5db1ooDdVYgGa9UebSxjojlnRCyFiFOqB6RiiCI
u/rhsJ40k762igeNNclq0uLCZg0YYznFCMds7IuN7ozHYXxaF2YDP3AwJN2UWWpSxrawgC5c4bDd
p5CQ+Wy8kvl9YedVIX/2MwU16SH9Yx6bGR2v5mWGZJUjQSwXbOB+w/pN3y1KlDRGLdI7/L0haazw
wEB/SkeKUP3byLvUR59FH1MICHZPM3KdEvnHZkIxpjxJ79N7pWnffberSB6GN97V69Sk2oqRnjmN
9llpk+2UUFON1RNhS9LaNtHjVO+Nt2j544CKMgIw9zpL22sNLmVM/BEzCyRy7pBt0wHYSSOWVPRO
sqlNgq0oskW9E4t/QDmjvOeumJjZ87d1MaMw2Rr20u5muzvwERtHaSU6bpsBmys7bzklCam11Pb4
zYlW6eVapppIxBTXPuSYJTdrgrZPhEaCk+pRNthotdReOxjilgq6PkSLr9k1Z5IIUuL4sI4Xh+Ea
K4jXcZM1d0nB89bKokO0Hh12Eo0VIonLBKMvH/lBgDgdffM0mXaG+MKPCAS3Er9Df3giosCIPeTQ
4hXQs+QJwt1wwCF1IIBJZCL8/I+/fmjCrP7jFpphGaicI6MM2DqLHKBr+CFlyJpC2kQZhQdY5RoK
rwyZgRnbrkGmOREGiNPkNaGrIkd/0UVswL/SYpBM/VmAXcd4mLNw+Grcuz7MDB/WbXyue9lrFEUZ
uSAegtkF/AlrL7eXgvcDKIdAY9sZvdJCTKBNQKjgHxEhwEUo9uMGG90I+cJEvzicXmYKIPmlCC1a
FLTFJov7oykxmGnpJR0MG29LuY3152BhbDKXC/RzIWNBMolBn43i/35GFAGlIVn4r37bhqgrzhGF
hSLwkCYULvWsj6SraFqvSq3jZqitYTWhV/bFnajvYslf/BxFMldRc0KyV5a+5uPVAYoEvWZIdfcE
ANzHl3u+Z1VX8kYwo3nrD2LkIjQAbjaTsS/LWraTAzmZBV+PDF/hsPWF8IsHmmmEyRTdrqnWY5G/
XyHZTez3sYB79YjLWcqHJX2tteIjTcXNKJTfyJidnwgDVQJlCM40keIcbZE/OB8Do9kGxAT8wYgf
/Dl0wJqy7cC+rK/VodeSlMa3pu49Z+7YpU2KmyBrzca72N5usksEQcB+upU2DD9v+u4/Rs4elKOP
cdQYS4nGMNlyOOzg8tZNkUZHLLxImUU2rLCP5db6TFou8FMQ5tQ6QAuaNs2UKusTK82yB1uEa3Db
MJWD2RzdX4/La8NOjMVgou75aFkzfGr5n8RiQVB5YGi2YrMf5l28HBEN3HGNE96yQSBCj3cTuQrC
3LPReJJT+0gShpCygi27W6psQGZ2kb9r2Wh+vAu1ZEqhAONCmTqpLA6JiwOUhI8jKxdlPc6E1ES4
mrOP/+ilFuFLJa2+5pjbhoQ5aTqildpuDoBG1Xapbzk4X6yeykDA6vsbdSXFi7liFpKXWxbNfmDq
1dbcVjMvzEw/Nea4F82Fs2I2Ge2wmCEiR64KLbRGrYgYiwqEX4kOPQOX9XjSJaJ3KODYs5FGMypS
9eJKXCI2dcIlZkRoXw9ztFEwXANBdnfbGOCIOiQ71Eug/kHcvdAJb1PdSFiRCZsh30R6uqr1yDrV
jY73LPtdj4ZL2e3cKZvKccrEt5oL58s8l7ry7upWUzEkZIIWQ1GKaegT16obA7hsIs1Z+QG++IXt
eYZGPNjICCyy9+/mzDOQetJVCj0CF7+08irJl2GDvcI0K4/z5V2HXRlUsom1OoBbm8EweI29J9dc
+btjN2dHngsBJTgkHQ3fO1hNQXHI1p2We5iV9JSFuC3FBwI1KonE8Ee2/fwLrgcpwjm4a3vefYQn
zQ3KVMy9bGMNIeBtoRqey4A/XEx6g/aQmfpcUNzhH55ASoDMhWezlhWELMhuXk9G1iMMgvM+tDAi
ONrp2IkbrgZgSA2FbMZhK3gK2wUrdbGTdz7yudnfVhbH8X5WToRbezNsFc3PlLkzfF+IX+tqTl/L
7MjLzjyk05/UTBuikJrxFxkxrRmNqiYlBKrejsv2UxeECuQP2ZTdTpEJr3HnJkDHkIirp0BZtGlw
cZUJ7LFpvFppB5KsoBoyW/VNlpAMntMVpRNT/AS7+ECxiMml8rOYopwqdWt18Ee0LjTcONargONq
3eU+JkpOvs0EJ4+pT3JEklIxQ0/sy3USFoNf4/29bLQTAzVHKRRdXZyHZoOQM/z/a3akGda+u2eB
k52MUO1voJBCkREh0pioQGCR6WCyKgwSmGl2rhqmjZ1Ir+clStpVNMdMAi957tTsurs8/FeiZS5Z
d/qFSSOIC7WaW798VwPU3C7QU0U45EsAel9xUKu2pFk0xFKPKgezCpkXRc7O9L0J6DaKMqtwLTwu
ZNh+d6Ga65VivRTlWeih/WLmO9CTMHY/dhgEIPAqzwbEB+jnr7vmLvFbWk9ysM064RsQOJCz3+1D
w8pPYllqhq2FY8S4SA4FTxSVzG4eM6DFfY4zz9Y5zSTNEr8Fol9kULKqmt/pQsYwHPi3riErOoLr
hasyVGNZseHLOydGiBaNIpGX3VUlU2SS9TuZDXgQgubcSr8XMOCQb9DWm18cGaFgRDkfaOlCkfLj
NZ7THXl/Jx8SGH6UDSM7uaBS/QWYVLbYN3JzvWQTE6CHpzYEQ7ExGXiRdnZttQsQ58fzaqmzHVT2
b8vNnCFDkYRXBM6EP8e5Bglw5BPxFVgJQU8oUo4QArCbTw/5AQCF0cJoH60vI6vxHRpvVJJZuxfh
mlQDx5hRsny2w+6mMSnhDNFZqsRPS2hyIP/ZAdDL65N52qiYqINZWRtsHbVZT/JW4V1l16n3FDVd
HpgXOaViEh2mufpxmurAskDnzccRnZNkR4BZGgw+EoHmhF4KqQhJzCraAABitBlKs7vuc3BPdRaB
U/XbBGZMXVGp2v7hhS4yslRHOdHC1gmq2SS339TZYL1Z2eXifiJ2YIwdg4T+UpHINnFCzkyodMOq
xyRJEQ73ccFNjbRlMbdwzBbGIOYxJW7awyG/4vPmJJVYcPDjFBKOczJPS9QGIlLi9iBzlQJWooBO
gbbCpEZRbKYVQbUmychYzHfhipc/pt93bznonWYr2AboVFEK56Fklckw4d4QUSVTDSiOhbn97uUL
9qiTiPAM4OsAHgx6dVboDxKR1PCB3Vtb8v8URxnhkNXHPXwNcqOn46xG0fAhQjhrp5TEFh+WFJFO
eYWNWRpCFuqbCl/rRF0dHWOs56uZwGd2l/T1iLMstQO+8RRakzp/MwYzgVGsCANhPawASeNKHZdU
j5HE8oW+CkjBsIP4vNfiBwMsNVXfiXvVli/oeK/rWx7L+DbELThM6oRxSr5k8AysLINfEqmD1r+B
wSZpdfZI3MaA1oOxPVrrASdUbjpqTW4u3h0TQ4Occo3vI5FqmfXXzVn1ezjPg/HfWe7i5AvIfmWf
+PEPprbcj4tks04xcuJu2a5aP1bb2e1E6C4Hu/WNANvHQOuowFVUVV4NIZcsR1No5n3OqN3/2+EH
/15QyIXcsRhz+6Pdhfk3FGnPulBsxsI3m+WJWeU/xQQf9hv2abgud+LYj9FBbBjzre3WX2V8Y4oR
0LJTqnPjb8C4FmQsMUEn3ids6Yw29dZ0HYNYZ9GXhiBnSs4302fJzMnzysskwGdxUv98QFL6hrVw
PlpH5wQsHlnAB0EsPECCzbNbAIroX9/G7sxHX3Jpk4KfwU1LKSNMQxCLsS+hnv+kgdIfyREKaiPO
Qphz20WYJcVDCOJuZHzEgbvG1RB3xLd3JQ23qo64R/X7tokp+N06wJFTzwrc025C+tJxF84IFPub
nYySDShGUEJkcctHgG1byTuhSGfAaiYqmMVbUtDymbCUwchG2BeNyAfBMwqKWsW8Zzj6ejPExln/
U8WFlbl4O9K242BEe/N9Q5rNSktgGD4diXli4Q+h+wfpbGHH/96KnqGEOYarUC+82wwt5biVraGq
eTS5MPid88NLbnWlfj4l5gI/GVXH7mqhXKOOnAeCLJW7d3KGINPUAizT1Zdc7dX+QGvNIXc9E2Hy
pUAZ9ziPDIhLBFWlkZfG8KCQk0asF4iHWUdIvsA9PkmjvYE36rlEVvxV+Br0+G7Oi0pgANvDnbr2
D0RSO9UI8ogVvtWXcNWXNvl6TNKHvuJ64BPrr0X6WNnTuhXlOZPyaVdA6uB/72wYydneqtRjMc2H
sDmBD3WntevTCUZ+g2fbWzxjs4GFFszDBjnrVKRL19VKMRLBbd9lQ8KvYwcW1hjZ7CS8cAfgVJX/
3xk31y/JFUNcllLaomKWuoq0d0YHaLJzmkFEZy6Uprz+gRzGRpdF56C3MreLHXFDOuFjUAdXbulN
EdmS464H4cPce3JDOakj8Fh8G7KkkCp7CBrokJomcoZKjWU5nuRpysNi29uHXDErEs3T9D+OtEqx
403DSJBmTq95jxyZHUQchd67x1GNwIxHSGDPGkoXf1YSV0PrGd+3ehyIqnWeOtKheNSPQOLRgf3W
vys35T+pHvT9eGA4FqC/KVXwll9Q96fPD+4xIjTwfto5Lx8vQ1Uf/dY9/Cb8o9AyIC0aezITy+0v
pnGpy3mh+49WCit0txKth5Dky/qvtqTz39Tuq2kY79OOzBouEMNxmujz6pW7cRaHXcSn16vGC3ks
ZLXB0DaslXJuKDRrpWOf84VINJP8bsdxMDNUwackS4QuxBHgZrzKzVWJmWs51JTopSwnZeFkge9R
7Zldy4QRdD3JT7X+cTpPu0Kvix27ATHOQV4+huKg9zpVn7yBMPtdYxQAb/usoBte2+sFqU9c2VDa
fgK8ZE8raxnX6RM0ACPbGvvCeUUFKdnKROVlIbmUXdI46t9oPJ0wPOTTwtw9I9u9Z9hBqNbMCsjn
A88iByghKsPgQpeCHj8jMzhGaqOk8pCyYrp/mFmAYMKSFlCvIs0hD4EgMNmFHwwHUPlqRG36JqN2
PCL1rYZmeUnzhaw6Ioj98VKfJ7Uq7SxqwhJ2JVqZmdcx8UZKx9Bc5BwTzxeF5HmlTPQRAx6zK3Mg
pUf3FBSHJ04mNXWnxSepcvbcWt12KQUTZSW1YsCkSXaDDg2XL5TrDe2FEcJXFDElbCrMMIL93YZI
KM9D/LrnL6vPUK0Cx6ZwHh7hP0vdrr3p07NaiVuBmgugt48LQfNPQN0G2dURPTas2Kb9/Gxb+jg5
uiT0oECYsGxdCjHN4akHS9JdLb6kunwrrZATZQItLfH30+x5liUEkM0h37I8Wq6gMN4e6Pktbder
Ywe36GVisLGNiA7ksHXplIkezcQmv1lh50brfLG3QsL2cYSdqQXTRR6KeSH88o6JYht4LUrVWwwj
QEb7IgWsNzALmjSKIJBMmU+ZwBi+WDbFm2nvlvwL6X8g9r/+oxSUIODMyAkkIevP1iyBddcW2wKB
f8+6+XQrU+nuRDKbxvCfgFlO2jGF441T3x1xVAB1UbGU3X+GFwzk4ZKkQI8vFzUm7Kq02jFIuA2h
CLuuKI/vAlQSEuK1Kn7cJvUzgO5PZUhRwG4W9S0jpkjzTpKdy0qKduN2Jn4jf++cq6Eaz16BNMnb
5OAiiXP2A0c7L9kAAJ6381+qaievHdWV3JUhKqZnSxo0yhww/z5kErQrZL3fIt2ublOiQcIYAVGu
Egm+VaAZPg9lz4hLkOObd326Rsv6PBjZGa+fORi75zAgl1cEnEiBhgxGladkq1HwlxmyvylfcIYt
CrufIK/9QDvAYX95B7ufGloIDcOYKMJGBIWqc1weIeZ9P4abMfNOdWGw/89ATmEGgZlpo4GgQ43N
Fwgm6Yg0FLCMXpKnFaCJfaVuI9LWN43o4KDgc/VVGxXFgxOROuLDVuGdgJMHp0lBGBE4EQ061zWA
ap9fVnGKFnCOY/oZ93vDyn+wXcmYP9+2Ijzr4u+HCCCpUOwUUKWAK0H4isOsb9MAW4U6FrU9YO4z
vQWExAPgn/9be+TVdzejJbKK++xkp8gU/LfS7S2lSy18QodX5YbSsVVctTm+1c4jmFtqj88on/vr
/fa550ZbFeifwII4gv6DghR7FX/cchig7PIPXizhNR5X4fN8b5P5+7Q9kfNG27fyNoY2whMrUvQ2
x6Pb1nRkCBrq4HS/AJUGyGczwns6xXFqkC6B4eG1CJ6gVeUmDOX/EW6/RfEhvwkDndPdBWJgdi1l
FtoV3/T5NFZuOFkPZHFTa9yNjOGP5p7uX6w8vgS18r2fISVcP/BgukoHcI+lcD8TexNeXbU74DFG
Hqu7rdwFObkiTsFnDUPYK22nCAh4nuaxQzg+Xe9NthhOfJUwrDBtVhj3jLGyBT6nTbx0hB7Etcbx
aO3R6CIkJFKzKd3gVj+93xwjBs8jtehv9w9AN0wSwlMizAyEjw8HaEaCIV7/K7DxfR3X8RlQPgPL
utmiC8w10Di1rqisriOge+k82exMp8rfTR/WhemlR9rWOAdqaokPY9o00IKUpKojHgU+tMzNJULL
lMFW21HKDMbtH+Sk7nV5k6jxThuo1RoQrW7BtOaIplCjZMnsUA2rU+dLwL7VKVr+KnEdq2hP7cpP
+FNm8m5lEqJrq6ErmtNYwZK32AoOnLS7J/Xi+I3T5+N+PFWJaL14aBbAGHJvaqfPTftr13iptOMG
TVUfEfJIVxulsF1nG7iF5l4a+KPoPwkpFB31urNIUz1dGHd8Zjb8OCiqeWG0bnAk9EIYUFdwTCDe
l9EaVts6XDRIJz0+e1gDFgYY7AFgK1fKwIZEBwNa7DH6R73p0kXzSttbL7pxYUV34OO8goES3xnt
6EF0JNuQCWQT/JuttEKFCowyaPL7eMPVV8S9GDFnSmtaceI6cM0B7OoIZkJn7tN9kal4j9lnhOqI
hdm8DovqVRyGLk/JuBXy4TuTkbShH2tWnSoWyV9bOkbF3+nz1aytTcH3GreTN3QxeO1PL/mpYbr6
7U88WrQdI/fPwzyi0ocPiEWJrGZAkHCmyu2gVdaz8snhYa5VGq2JMriAwcZtba6K0wSek8xmjVqh
4GHlaGNKfdg/aaeiTKKHWu52Fx434TD6qewAlL6ZCWgORgYRz6oZ5GuwBbxEWsuuDZl1V4pL9azY
XYxkt59c/QIIOCs+TS4NqGiD5CxVJl3mPojBvIdBToawfK30zFyYZoRZG/0vD2qeCndZN24JI4VI
8dHVGV64lJ/hLbY6wjoGjG6chh4RUPWX3ivWsSJq6wd+zmmZyvOG9xTivfncFPbhvauIgBfJLWlo
L8nlA8sCa8bekdd6qm6iMGzRD1nP+U7H15scfkOz6jBrUd3sOwVBunDDdCybqUyHaH1Y1I2WomU7
8tx7gxgpXLfFea4fbN6FaO0mHTouFJciC9UGxsOR1hJGopm2S4GZUKsIXU5Q+u6eA35DJkc9NzSM
ZeWo63qlZS4M6ZcQcOCML4bKonSuvDBJbUv/2fiEhM71p4zL9pe8ykOtCko4G7ddCbt1EDk9e+M7
ujXS8IuuezUzD/ITjyknCQOUfwwNiqIqF3RXIMsJw3kgapQQsqDRxRQrc/e7ig+arA4ripGIpYy3
NpRDtt2PG5l2eTzxfkqehJVXzAGdIhn4FleyBSMxuNzMnQDv2cuqz0mEoCV84chjRAnM2X1Kgfg+
4O78pTZScnPKcuQP8ZxwWdFrXG2bz2ov9reSyKT9T8Cbi0XJwJwzCMyn1ssqiIaQYtKN8KF9f6Eo
mwn/ufyaUWlBDHlAoomItTmXL9qbIB5ZMhOmYh5WqRJSW3ZtN8lS6NNT7QsB34T7fYW3B6KLnmKg
/Yj+ja1sQlF51REP3cQNtz5OWZ09eUUcRvNlnZ6Th+ovkN4GVbcQawqWLIpHNfPut9T0qRppWQ+K
nCu2Eh6/yCLUJewce9tuKeQPAj7hh9cxDtPNPBVYAlDyh1eFRoTLfsD02ZAGTHOzjVb4NPrgGtw9
lvBv5ULf+A582XAt4XVY03j7dI8NU092HAV4fY0LITUerHQN0GplN4bmwPavj8tQ5uIiFyH3J4ad
E09l+SL5Y0WI4JnQd4E6kUhKCPNKmdAdrlBuUdh0Cji9pw16sU+33JITMXt+R6lq3eg6MNc/sYzh
iWYYfAWga4GmAF//S2WXA4F9FL+EYq+TenP0Wk3fsmjGm2k1Lx5Eft0LCBvAPVEHf0K2Ao+0JxnH
TvRxQM9ofI2KFD0Fc73BYwztT6PN2TA776F0VRWerk32IZIPTfTbThYnkhxuPMVBWavuMv3DILRn
3/GSITWkJEq02F7wL6w1ExyzfwB0ATs3vufSHnTbC3Gy/L12s62et/qSTulh1jAOCnLuRB98VCgB
70g852vHsxgGSrqOc+EWwR2kUjwzfqJ7vDRhGQkjua7MjNTw/YbZQ647m3Af+7jZ4TBQBDahG738
PllMNZKNxohGoFjRn8pRn9LiKvfvhlPAbqvYEJ+K/S1GMbU8LsjodX486FQCepAn+Upv3SfRz9Vd
xc486vtx81o8gvkTc3J51sl4bp40FbysZND8oMDs9HDsfiUWz77v8f90yuTeiN7ibOJZodG+WPN3
FeiEtPeo/MBp0RleCGkIChNqZVN9086X7x6UNcMNO7g7cXPnmC0AwtsRE2OKBhxBr8H7VYM3DeHB
IGFo0S+gYBNm/c61olaRvAXlDLH/skIwAk+ZY2n39/uF/iQh2lH8Wcoj5lN+7Dp6TgnHZ1e0jnv0
MkThH6F7YrM+qEGHR46HkwQnw04aKsjqipuZw8fLu4SNpu55ccZw5FB0Lftxkg5oGowc8gGbE5ni
lVv2YMFyVM/Dy3Jb9QFFi/vqJ9BTy4witF7wfI2hxXq7MyOfsXOSLIk77q4ZEgYVQSbemjRgPccw
ECBeN/Ad1oXOTVHN7f3PWMMuZtGmNItwE9t6D3b2VnZ6AbtXne9ecseyzqER3qOHeYViB7U5pxL0
uffdi5tB9L5OGKD8bif0MKwprr+LnZG4/LXI/ayN9lcadCNzwdlmmqgD558j+TaasdeUenPmtzNw
wHKZlqBQPkCg+uA19I1OQ5plVrCni/6yZdqEHSonyarl/SrsW/Bw0C3G3LInCaK8XIYCuvdOVnzS
6+tilCU5m7t78m8V2S020ifKVMTyHTB1/DszySj3agVDOklh2nBPIT7vigS6VQ71Iss25g1lo54P
LzqBwBlUPg6ynNo+ILKNY0ZE+4gS5YAvB0bhcG7v6t8by+35sShiVGhrAxnZuT8Dx05W2vFXeo7b
jAhQeYLdM3RZTSm6JEkf8oEO/x++bPOfPC9sfiQPI33//3heOLFwNQFy0rrC0wmgpLm4pz+UuPtB
C7t2HbFkto+vPI42OZqV1Vc7VvxnEVKXUuiEyNgAuLM6vLoHNT9gT1Uucz+TXeuUQ2mBfIpCKL4Z
vI68S7iwuCwkRIvKSQGvycgLkmUx0Bayp/ZM/fZPdOdreWgXTqd52qyECuKVI6ndbmgvgcJvLAEZ
JCrcrxZv6CeTDUtYUCSndOzGpKAVfJbnqUZB72pGBjvt4zp3aGwO24NB2W06KzpJug1xkdqTqkUE
fyt5ksntbDaeiZrF09qunEs0HAdGWovbNw01GkZv05arC1CFVxDJewTjnNEtM/YPwwpwr54LsjOx
g13X24id/XRvA5BS7trbRdQrjB0N2vswTDOafa9HmDqOLoo47VWKP/OyMaZpyBRb6Rpty9nBEYir
SU7hNxLWhMd9rBa2jVHwsJARGtMUdkMeBgFs7TVtqrROCKlwCVeXiV72UhB1DLzJC9C2xVcU4NRs
57FTWxaaUt8abD+pu54Q7F13LQsfBoxB/mTchjCpuqJcN5doZJAF+YE4s0DFkGGr5JKRwpuCcwVq
37Xk5pc80MzcTGAqsYLM/Vt8oIoeLXmBHpPO2rMXAzUj6DHUCFAosldE3U4RVxkBdQOvUqrPE1NT
Jt5A9bOVGLp5oetJzjHAwVaBvzQR1wCwLH8Wrz5fI3P77bLz1V8RPpNjBrtFd4oFhkHLRRjPV/hO
TG8A7HVHRkDRYT1yHw7/rFqpopCYAe7uNcicduTu9f2DvElVwqTpglZB/VglmSgfnfvLc+Juk5th
OlzrVR/3AkCWkW8KfsV8ND9qABRaHWCMnS9RlCGwTBAv+UeXnu6VRVK92zz2Pb18Mq4FQX/PxttX
1kZoabbg04CEQIl0xCqyZEXiIaIwfwKbF+dBAypkOcZ1DcTjFZjTbGWIkqvK9wo0Hg77rdChv0E8
9sKXXWBSG0lyfB8bxupcr3ftdymU52w3Tr2jtETMiVugBCtRoBZfPrfj+fhtHWLNnDYUqyplRFvg
MmDPNTmbdhDlPhoFzNtGhMOqnyFiCoQQNH4EFeAECk1MDfS5/19dFYiUhoE4Rck+ziekrdlDHTmd
IaOLkB7fpJPJO5H0rLVoGmywbVSvG2DGYRNdTWPHebd2JtC+UxYszm9CNiPYcR+rHxMZyGHZA8sp
sZB7TngxkeiMo7ciPWr9TNejq1A82dJMnQRK6QKBZWXk8NCEp2rJJssUK4Wmd9z3jnvx+vyhEIa1
YDK2GdxgB+zskHZdrDNgcg3yzOMuK7KTKoel7URQGdrOdxoETk5YPcqTDuJJU1e8wS5W/KZNd0iQ
YfkQpz34c9jhysrV9pxzZH1R8J/4gyDcfShJwtD+WKNMIiX7l4V/kqzD1oc1XNjwPKWEmZ3fp+jZ
9A3dq4yzgVxjnv6HDjyqx7WLVTKDT1NzhGDPtwC7wWE8ftWt5FtTan58Qc4i/mPlNFjsrGd2whLZ
O2r1DROubEWyNCxTOJn3WOmap0gw87KpVF03pwNCQmvzMyMc8aZXJo4DG+TtXj0Ke85G2E4n/hH/
EjJmsMaVP1qf++EMAwSWpkjvlBWBPn2wt3mgqlkoFfmyuLmY1EcSJLqTKlL8qyLs7ln1OrA2N2V/
3nAf2McPCnDV4TzlBmBUVA18eNBa9rcObAQAiSq2mBg0zleFfJ3jQc75UlzN/0xIBlWk1YIdghFd
AwZfHOYvYcqWP2Dn5AlsCWP5NnMQXaPEQoLrUoIdT3JhTENUgIDTZD4r7ujTfL5qwds7KgHIJ/aI
SkwyxvE6L54BVLCuXqh82CMHZ/2h5LlM27XaIRfigoCxBDR7+GNLzLW8ZVdGdx/gmau2iLJW4b2I
kNRVve0+Qfne6mM/K+Syot0XskHmYLs3danpSE0mrN3TsL7D41x0egXq7Bh+YD61sGL1RtT4y06y
EbG3X83bS4CjQCdUx0HsHHwesii1SYJBA8T3ozDj9T/QSRs/+ojc+AXGKm2exNBW70ngdqts+zWC
LVCJugF2IYdQt4zjVt0eiw6vC2UBBW4Y3lDkgDCpK/qq/sFqNMYx75h40bHQmjSlTOC9Y5fhfLuu
+XZh/6JVsxRzQp2PzTs6ldgagQokWuJguYWiRE3S1yTpsPTy+59WnybslATgWWkICVzlNbgBNdqH
WtiaJuZASmBkweNlUN53SnE5iAzyx7AZU2TJudbJBgeQ6xJh85/ZrD3m4wj95CalMeX7RkQ3S8ML
JLBEJhg2Qdl9CC16VT8JRfAhlSq29qbUQxKTQ8KQawZ+PENva9oUYubPBUEYUoKHszjgtTc7LwV7
Ri3IgqU1ldKgVhjVDsaAmlrpgg1t/r0GdDY3hQpdse1zTjxfcuZIZo6JVibu/CJxlbtThGSIhQTC
F7KE7ZDdGXdtB0X+AO6CcdBY4cZgpbtYQuhgVpPAJ+wFM9+xBSAm5FIqtZyBIDtRpKZ45LbapqFm
hyKWEsoO7upOd0wqIfhWngrAj4V/wsOnGVKx/F03IS5a9KyoPYinq8DmXHtlD+yHE32F4rcDdU5/
jYWdyGuFho52kf1IoyEF119Hszr/y4g5SzJWzu/OG1IqsFk3ftsr/rQP4lLshL6ixD4HigxVdbSF
kRNnkavMve6YRcuFT4PbEKqhghSI3db58SIVCu/cmyxa/lK5f42RQ/09vBhgSXw+JcL8Y03s38r0
ujOn2QWvLrnPOYMRl19b6Gr0MH2uOHSFPMNUC8+xT8KAAtNRJtt/Xw7XxD0NptMnKusI3YhVVpQG
QT4j1sAnsYZDPxWY173JT+UXXKXu8OoQNyaQuM5IRuno+jVvb+hosGZWx7GaM392bZfq/yCgzdBg
Tb8qnbFs/LQYe8DfLBpAuEctCAyoubRz02bYuPmb0a/QrCCqeVWe/eqPva/a5dPmb4RJA5lK5/u2
SIDemlOf+H+TiwI8FgZRFMZcwF6PVg9mMXCaEwJHxg+LB1DFLqoWwmdzWWWOZj8GaN20pYfTdrjR
yGskVMeNcCeuMoDGOE5s63gducCWjYN8+lQMJ73VH9fcgsMgaaTtRRRLB3efeWqr5Kciq45OTkSj
nQeNt8ag8ZXzfHpfMFs+oPnn7PRNcgfoSSsYUpRQrJk7ZpPJRk3M5HxI5W2s/F7Ofyj7JgisebtV
LNRGV5nD75JYcHrwNzs9taqre7w0D2FPhyWiCL5wqOBxL1b3U/SCskbzTe+uwf1ICOXrH1goFM6H
ZKmeqBfnr22OpDqeEsacKMkS3uTl7lU5rHUp5UUg8OzEOVM5n20XvR5EOKgqxN+dFHmq8IJFYcgv
FbMqWdlEMvgiBPnDQf+s9QnZM0Beoya9Exc/HI9pbJ7lTWx1dMPYcArwO/l6ScfUeT+spHbRFJ5A
fi2v1CUsOMXfSWvFEyeROQSY/TpHnhAGnQuLRQ894m+gAYVDd0lc5eLEtLSvLCwTvs22ngkLC9xj
udxI2B85itTF38ayNya0IzQpa1fW3Xyso55sg+QnB1tIufU7qFluNxFPvqM5xGbBbnypvRxSNmuy
DyIwGoS6D4yoQfyJXNeSNald3qDsdQSvw5Mcs2Ag88/x6Cm/0QAYzQYDnKSgl+eh0JXDHO40J4qI
TaYzhqfEOoIE+V/dvwDCuFpskQVNHrTDNp8tb6+3AEZJMD8RtmMyVq35lpwzgO7YwDqbAxnMKqx6
BPvHnRZU7tEqR4Wl+ej4mLK5FfOiIBzN3kY65hZXpoIl9Lsocci/cuCkG1QfCKtZ7YBArNyti6Hu
Vw88Y8FxjhBjl+lWv8t2hnb4BNZF5Tp3Pg6appzPwx3SyWReU5OBWdNhkUVpMpu1Sd/cuLaNP8Ns
HoByzsY49MKbfA9qLG9chiToUD8CaRtlIiwlzXB+Rikv80MVL69Ym71Vkzkj+MklIGwGS8tsaMbx
TeE5s99Nqy2/p7BHen/GjSV0prh+MUfGDr5Uofk26z699694VX8ZmVQYqQUS6QWODLQT/HYyQpBR
D6cTKdvhHglLm9IIB8QCtA6XEmhW2ViI2aJajTcLQgSLTyK3ftLBJL/5pU0WOTY9kV0042HqmJWY
RCSbA2x3XTeb53HcnSBZE6WoYxqeOQaZibsr6Ci/7+/u3NRwNWgxmRvG3tSiQrDBjvX1dibtArD6
rNxR+JtnfciiGg8Lq5HqJP1Cu0dfnHWIXpcUY7Cg8n93puaCnT1usFVRLfv/pEKIGtYP1w69LeDL
rvWk05Ea/92vZv3MRvejVubps8Y7W5BJUa4zHl6M+8FaYWqAk02WriqsDm+lCaiReQaFju5/q0Rp
mYN8t6yAmnJvhy3lnhD8lqH+XQRRBtVLRp1HlZez/AISAx40QDNh7kvAXRJRJb4twbAce62tucNC
bFGPh7PsVIvHRwij0AxXfwcAXWgSo/FX5XIKtkBJHZWiGW+F81z+PpvD3wPivw9KLxAbSCmDLtSl
TgRBVrRoN5e4RYuIryic3jwWakxrYUBc8kQ1FUdy+kTkEuNlIDiEgRWIXa9bQZQCwB9DAbBYVvkt
cH6gCGul+CwLB5eCu22UWvF1X65tw1/LNUvZdBUhBkXDdXxXsnXIuwqe5mb/x2ZF+IItbxej8kcF
CVlehNCtfnRn05QiV85q4fio6CiEiqGYbI7ut6Y/qKR2s10QcE8Mbr4VIJ1Wrg/deo/1exRptOF3
oLcvrTCeEC6+1qiXzDlsXPC3Sh0EmNymjYx+34AWSTW+qLN/sXQligHu4xWdL5cAmIhsg4oSB/hi
l1SNWFdTi9R8eSvq8OltCviyIknFxP+HTtDgBLCUFCCXeX4qYz541g3M4bdhUWVMTbDtvgpZBrL8
E8GB9ciu4AtmZ3q/olxbraokbaUNsQuTmVme/OUIfQZtSsxIh8ZNTcF5P2v3zrKKsfj9Yx3TuJtM
PWGfovvBznFZIo/X0wXF7YoDEoHPWztbA+rLkE6IjPRtJ5izIH/3aezarSw+StCA90WyZFYG7S1t
bKfGDE8j+0TOuyGrvXXUW6P4UX+AO4yaiCRB+JD3lEkJETwd/cW2gmq106m8JJ7sj42izXeYhooT
98MNOVMGd9DI5/5VYM4QuoINjvQxVB5cOpj//iVLy/nfMGVOWMDZGru/B5XwhSVu5WD1BOGgNDjL
acXOJ7MmNPddacIGvpN0w+Vticlk9eY4CrMcrRZ0ITy9XKPWa4O1bwAy9zZ1Uo5FRk20O2CsuBye
kLnOuoa/Md32BrrzgWgJlrt6bY/18dLsug+xVLkBNt7/dNDNbVWPlLc/+EC/efpFJ47+Hko4++DI
B+fySZ5u7ru5S7bgdm118fo3/ckKaWlR1NsQ9SEvdi2SgBcp5/7SYsW3wc/V9OHZcCg8sH1MggI2
JeOl0HZQQ2SrwFFn8XQn8dvdZRZyxRn9sDmkpL/DvDEL/Cv8DPZPIMmKXAlflI7l0PUc/hfKXAFA
iEBSztz4VoQA4J01ZpfPgUDqxNFtOzmhg0zMT43tenslpwGd13/TiFobJhYAtqU9VdY5Sxwgs+i2
CSIgRsYOiwXQF1gh8dxkhIH15mnGjJEb35j5WeqaiJ+NJaQUi+7F1pRej2jbdOKTW+fUouCtaXfc
UsJtDP6epfM8fl0EZd0L89XUd3VJANbDtPWw7ySSkidIZwRZlg4zSXjA1+JEcgR/PXmJ/EdCYQ+O
N0wZ6sV9LQyeFYaoICNx
`protect end_protected

