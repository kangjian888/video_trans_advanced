

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DKaw2YF5X/sI0l9aLdTgbK/M5GUdtEMTnIFmxvSMohXCNpaRunL9ipaA59Dc71YrenIGtec5QT4M
zCoGKmFbyA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QRHRuF+/6jbJdc98CuDuU1RSPkw4Mrd2rWInSv90clZq9I1OTAA5/xdv3Hk99Vg2prXDV3YjNqoB
pcpnTJxql+YZ6VAzN0qCk+oUeO1cCu3qiinofcBjVXCdgYxomUKUeE7FJeYz3Js2G/kJGoeHFW9U
+zAl6jadwyF9Jbvv+i4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Lb7wQIOJLuT7MorOQ8eHbXO7nLYJ4w6DRb/CRc0KXgD29tV/pKu8nH2e+iVICJbGwJJtQ3k8P1j/
LscOU8Hk23tTbvsi/KP4jYIAhUNpSlUfm6H0KJ2yht05tm7/nGOSq+YwUD5ni46LH6TZmw9wRjLo
RAHSpBohLboc3y/hVTXta9kQmKPnqAmdZWZqkVyyS5o93+63/fdqbFaxxtwx1mXeZDQ2+2zbTCKf
tbrO065IQsNhLqpQ6GmWS0y4Yk762FiY/PW8xLoCZ1V1Fh8ocFk7LKyATUlQjo3T4vsNks0JLfh6
k4wW0gpjLf86zBHim396ye0D0jCoECOhPpGtaQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZXacKhqAwgw8zLrWO0Oej9oQ1uNqsfSW24Ju9AdSqiO9hJgeX3QSs/Auka01BXmxZF02hREfAK/G
6uXtwOuytUDW3C0vu69znjuzfKa65iqAvitXfuV2wV2SBDUohxstI576S9cHfGPfoJ7tVzjIg2t8
+fXxMYGWVW/hL5Dt3LeBc+ul5BEG9/vwugVmMP2uMG9nGEtDEQeLb7bWAsdsP6jyz5L4K49swiWc
6TrDCW/53r7o1y18s7qcumMrH+8e09lZWlV7gV/qSGCmNFjNoXkvbq7X5+RT29nF6kaEY/1Y1wcM
sqDv/0rI3Yh5PZatD+o2YnHnz7Es16C87EBZrw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pkb010SLYsAhKXcWm+QlAA9Be33Kx3pWG3KQ8c4OXZxiNI+ziOzdNGDZkUALVJhYeeODAczIsICK
xPobg5BZJdmnFjXMkYzJiVNc7H8OtQ+xwCOlZfGQy0nG30bs3aCt+0ciZZz0ed8EJ3QfOUNUrA8S
ACDctQvzk535zqal7JGqVOcbax0rksASegZXl9TYHMAWSFXsQNDtHG7HCq8QaEGySiiJnEz1Zygi
CXmAaOXrSZ/75eRU/jV0Zmfl2uX9M3RD4WyT2L0mtTPVI1Jo5riNKDciMqi09G5yCgGBizlVK0Le
ynsKW0Fvo5j+TrmGuES2+DcsvwzxQUmrQ9n9YA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
saU9xQVocYCNVhmm+/jaIKt7f7lGDiBCwD7GUeN8jk+fV3dDx7VH8BXnwqh3bO2UtgQTq4TYazR5
PsEJU9lk5Y+2uIztywixaUOcY0t6PGvi6DZ5S1UapcNaqz1GzVDJNMdFrGWeodfXgyVpIeng6Jtk
EKceFNW0p1SgbLjlCjU=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pbTosJ4LwLIDFDsIbDQWyryoCwFpua23V6z9HaJa95eQ/VgCaYwQRc0pJmp/UgRFI8GxRIcCfLjR
nDQiDTQUzYsgXuFi39wSqyum1ybk+zJc/c0tfa3zo7fAh7WEKBR6EfegxJoOfQ6umn8yMUOq35ku
5cQGVgAH0mV2j7kgcszzSTcMNu1shLKlPJejpCdXAsAct77F4/JiYgr35R62Nw5TiOPHxLGWKlD0
S4rOzGqDzYI4jb5eYbnrBMtpHWXse9ybFZPj47SvpsioKcFIHeUE7GrNOvNDQPdNPahScNll6gSb
fa6tuXH+3Q3DQNGg7RW23POGEp2w+WE6Kef4qQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74224)
`protect data_block
yMYYqGgeVsQe3maRM7bLX0c2N+asF5cD0d06OXdkHbgxOuw/Vh4aCYtelqhgXhb6c45qtJwEPVwx
WZwp/Wm7JtYZtP5hT6Foz6Sc0F2JjJccrWr08RQobyWSaoNn/6Retrd5QHoO5URgsyLeqxLi5LlF
k4pP86cYhA0Ap3IysHnyNcewxldPiz4Nxf6IMdt4MXKo+nX3XxWbs3Gxt9awPY1cAEFxMOLXVZYE
gfrfS3bvX0JpdnYx7V0fn1RGwhAFqn7poFrhf2b5AP/SutCgRETnJHHu90jAICP43KP4d0i+SJYU
sQX6SPkVn/V24z0ZTILLNWKWNYSMGsInjm3333qgMcnHwODZ3tkuoOTVSK1AE7HKkVWFQS8mUTsX
qce4Pz/zje1n2TbpAqWg3DWpGTblHryaD/LVq9sthSx+qZw2q0VKIIPltB15ba2LZnY0Ysqc5jV6
PLC7MXZao8oqhWjXw8yiJMBYy6x5uFq0MM0N/KJYoiLwxiXw3+0l1bSKKMY1gVtH/NTSadtz4SZt
Ix+uQzYlCRPUK6eu5V2kxcsq9u0IGHNzg/ZSmFDWDQxfJqtp7rBeNdxRPMKnbgDuF014q0nICZN4
CtFhvBP+k1m0Vn5qTeVBn8+sL3/TMkWvl8ci/dbaAf33JH6ylGLOTGTv4Artzc6CMdnAnJIaFG1t
9vsR7a4LaH5jnzEDZqqfDxvk1TiH2CwF2ET+fnZnYpQ0Bv0pp67BkD4CwS1nDfQVLfRtYP36ABzL
SYcgLgibzfSQfP/BlYjFyxLlIPJ4we210bHM7nNysQOA/8aTYib5TpiZw63pBuIhdIN4ghabDuVc
7yc9lxqgvnGfiGOzJc1MIquqi6X4/INn60rRmdgy4r1xskU2M5UOmVetaTlwLUuI9iG75VeJL7IP
Cj/ugDPGf/qcJrnhMZPXNiDjf1Ni2Z4E/T5fasTlntEIJdtT0RiC2i6wd2qnq6DDpPpC3SAaheH0
WKuLhcNSWJAe5lHgZeRYhDUi7gq2lVU5tPz9DgFEkZtam7DZZCUjMREFu9LWa9cvKXr3ZXqBDxKH
laIG2L2JXr+nM33LUbL6zdrNPRtu5B5qrht3OR7Nq0JQWHH+ypZbg/XhfcwMrpW4X3Xzsxf+85o7
szSx/GSO/v2whCalYLD0jdhRyOG93uwGn8BS8LPyDmsKmWkB7lculy02cUyxSmbqmAbjfCUJ0Ix/
rFZw+MoplY2PZSpA0lezL75E6fO+uwwA3hl3ivp4p01ysYWQlpFcju9MkDJxxms2Xw3HPg3pZ1sV
/97JXoU09o536ehXkyAvlEKDNqj3doIKMVt+O4+dQm5qqA/EJg/EMjD1c+gkqOTCvzybfY+6jo9Q
6pLM40JtUdgyzinq6362b++BSKoH1MjVKkAhArWLBONWuieshglxXCM9Q0xrierSc6iYD3VxlVf1
lWIGYmde+SamCmyoui7eS4eW2CXbZTJZsJLmloDrXecr1IgbGrtgDpBv5sewJcnfYhmIMCiAVidC
+ebAWLBM3KU0dVDGLzBLDjurpAMIc+yAuTN8oYGJeohBBoN4pIWtJ06DkUftl4gDZuZg0vWteRZD
IaNHMHUzssuSMc9RsV7xV68TpWLT9RH32e96Wex15adrkWIAodQfF5zEaEmtDEyl/mleawXlVY/2
UvvU8/RHnooEf8G2oZjG6MowCjN3U+geA2bipFuzW87JrLtVSBwvHa6t5qmi/76tN8/pGgq22tWA
M4JO8xZafIw8P9iixTuKeVyhSigc26IF0oPFcLpEFWsU4G6XpyIxs6MypWv3jRhDYb1MvJZf/RmL
oIhrHiWnvwNR81XlU+fE46Fe0S/cXYj8N2mnkjf36Lmsl4RmiYeagPhd8Sy/knbKcvu2hcO7YcQw
5Hk4SMQZ9QM5cnWHx5xI7LRFDJgY5RJ+tyZViYPhmyVCufj+9Ps6aNxVPK8FjY87gIm2Bh04e+ml
/ghdTstmbaLgdN3ZT8fFxjgKJeM22aQ1jF0iaXfPjzcgrxy1E+6v58A+mpxEjJFEmu2an+Na1FLC
YHXB1A6fZQOBXCZ5CNqd3dZ6vpqBrZzQbk4cAmhQ6t6XP6Jxn+Ib+dV0TePEppb7n0eW58lqf6tI
dCd+B7CTLoLIf3/eJeqitJXa9g9VvuRmH7djrZz+2qPGPFNtXlLAkpO8NDHFasaLL7X76hfXcQ3I
1MwzuD1cqxAkYiParPt65dP7qM+FSsTqZYZsEDez9WkIK68K3V8arm3vAetN06FopAK/jrEmyErF
JXkJlWNWPat+KCvTKdI5Do0eiMF1Wze8+AokC6cE8N+FkgDzmVLViqyzSyYedJuyoB+uEasDkkPb
km5UWfC3PuZn4/ULlwjDd8UnqQqS+mWPuBngAk836Kp4K6m1nM/C+Q0S7udYDR5jZmKaS73Rfc6e
8npkN6cRSYY1rIrh+usTjLtePEFfyU/9Q5NHrO/s5pMumDWT12OgCvhHg4B6n7Xt2h3jt7wI9NvI
VDFnzmyn0mdGkr/BmfKjWvosovYmPraKCd7SKq4+ziYnjHDx5Jm0O1bNdhaE9zUOsxCcwmVL2tWG
NAusZRA0sko2aIfjKe6PupOIJz/fpe3q+aUYaPg4U9tpfxs/iEdhNR6Q04B8D+u/bjMdu3CAzOJS
WBUY8VGM2fU0oOUnTYsbKBelyzpU5DbgI34Rysw6D90rwuoqeJHZRhaLU6Cf1SpOv7pH4rT080OR
wpxirZeZZfjmfwEAMk0hOw0kbN/DbYN1OWnvjio7cz84d4BtkGAEbF5rmJELsgzADsM1AvzvdMLG
UjPAF6wmolL80uMO01yTVhKLlYJXCt6PPMJTetJ66jWePybAfqo8SjVnELU1IjcoLWVVe+IHdb+o
9qkQ97GJj2rWjJf+dFH4rc6PWl6YoSLE2jo9QD8PizMBG1i2xwxrSeNj40Hzwnl2GsJVzqHJ+qXo
pbJLS2nMhGA2lD0Nba44G27d4o8stRFq3i4f0FLx4Ge7B/0Hc1ixzo+4f2HiaEcpEKkEMw/0XpIT
P5pY+w9eXS7uceW5ZXy+WMB+PLNB7cRe14j7gaPjAbkHsg4oV/pBogaeHXWZ0XhcgYbdidw55AUb
RN4Bqkm9OED61euw+jz8ug41rAf63aZzDbp2sWMeWx+dWToEDGWr1MIJ4msNBxVWRksSvvOj6gP3
2zfXLME0mvnlEOWN6Koh0TE++Qqdn5LFcwoyNE3lgsL5pSls1FnV9I9tah5JTQymqzB9vvgPiZjG
BbvnDpPHvxvQo/VpIIbPwzEYvFqM6cv2VedHWyaxOQOQUQubgoEBIrrgXiV3HQQ75bIcQBGAHGRE
2/4K6H7Cznc9gcTYpdontXt+d+gtXSj65LOBEnuvQvCVj3fiRVM2MWg/+BWWtQXprj0KAeY36ec1
EbanauLjKCCjtxaC0BiYcAtJumc7wvz9E7eOS2y6jadV+SZIoMgeRI2PMlDRtCUd3PM66bBImMv1
otn/atdBYuKmtgLNLSS0m5l5P2cWSD2rKVptcj9AMhM5x1qcgiUPeUSa4vXkoC4yS0dhq27EAXun
mEvM1TOvp4UcZiOEySD2fi0NcmdQFS+hFfwaJtQjfIXrTgFVS7F7B/fTs+VNhmPjAvQM5iXWZe88
0iOXjPYSrB4mxDkIUzn5HuHpkNfWPN15s+i3DXMlgutmmkzyAwxOZL5rPbnPYapzcE36sWSCPP78
hy/n1rTzerRp4v0yyxeIc4greZYr+/STtsO0okpH1L7iqa097Ml/kZL8UtlvFQTLXLMuuAFGOdRe
yq1SlSr4yASLbiR7OVuOCK92S5tSrY4TK3UlePUPd3b1XKQzYUPjxfM/uh4XWfTxPbqh0oF9an9l
kGRk3uMRkxcdGTxLnIJ5TMTYC5+JCtKcD5RlJMTJJdy0Xjc0EjKiAYuq5VxujyZ2k0RoNMukC/Bb
u3IDcNqKJsdW3Gw2vTBjYbPZvbV5dx1mRqLekZngMV9sSd0+DirgR835/j3auI8/+pq1dFlSq51R
Zb8Zk2vcwKu/uHbpiMaepg/I5QjXzA/88gYTzpI3qO5hfFMGoVAuC2+hynzvCAO+vqWl2go0QxOQ
h5jAU1QldDoAbQCiOuZaD21Iso2FsdMY3Q5Zjws07tJTcGhQ5VVj1lFWOxB8yHNc0l5b+M4WvIOQ
vuLJk96BJOvI0oivqdmUgYNNClPTYqJlhLd4UNmOEjsVFTPwZA3QJEcGdyVed5iUt41O1yUlamRg
rDaNuiCBfLrl8mJvse1+VgPir1zIb6kFTmY5K6bX+Jg+HpvCLaEaNi6p6A7UlSvfCldJIwtaFijE
Ua2EDcO4S2uCuHH3lXNUyhyR3ljfvz9rgnNauqr3/yHM5VhbBsHGtQqFdBgYxZSBABY2bPNJnVq3
0McfTsHvONgnv8dHZh9c+p5atHQp8VcPNrBAa1hIi50VMiXI7ISW4c0hrdY7VUQxMs4EMVObMQG0
mcMsXr5xx6+HW8ySnINKt1jZQJpvm9HjB54Cot9c6mRvFqvJkkoTHQmoi/DgyQKMfBT6cXx6Klhk
AzTuRGsJYGHro/jNLogUVjBeqJsBO+FdMt680XFmvjUQb5tyWDy9IMOsUZEQgvas+yXg4s4qbj/9
Zm2Pb44Ol14R5s7nVDQvhuTVXXiqShsVFxGzgaZyxeP80cn90eZKhfulnQ1KlPRmZUeT+YKgZfZh
AospUn3/9tiRfGw4umLsrarC84G15VcjxUb1FQVw7ZckHzKCVtUx9kSrjTRUDpoEqPBasLG8w4WD
mW7KgNacg9AUOg6L78wptO7sbLYWPEhkZkvPiA9ZclBfwyVn1SUdu/j19XadC8hxJiAMqcViLfLw
2wqB3nF7oNzQRbFinqvKF/xVpZ/5crIwNJl9C0nawGR6d0v5smN+soBbfWBjnrpvLf6TlC1mWPf1
wPEDqLEmCCSNBrFMfh27Y0aBHrNzVOuxNyo6YiPSuTtMaGPEI3TTzEylA80AZ9okdzyDwrKzJMhO
b180ezX6KO4I0tsA4b5wmTCMCRqB2RI+DFCkQlP2qfXJRV27uiXNVGq2+RE41Wpkq/FTmsnWOpI6
bo5ZAYZQ7h3MkvOf86CXsvpi4iTtYW9Y3futkcRQ82I5x8JXESWOW4VEWDNhaqgz3X15+TDCy+BZ
TYinw4aXvv9wWBM3nCqewlDkJcobA7Nbg9cpXwgZiQcShO3DjgxwWF8PwC6cgdP5dbE1TTWdMx+7
S20bjohMSLsjRpJujG3px081xOExq+s6npphzydRGaHh/IIq8xvmMyazVQvsIHBeO4B4+7iklBTg
/afKu47DiLfez5WFB3ElmaG+/aARKVCbd16taPMs2Mj0Z6nBxejBFrmGh/v5zKR2wHaXTtyixYgr
mt4ar8fkQ4xlhyyE43e17AS2kQB2m6HOqh3I2Q6s5JRJDbos8tYNp67B0GaXR3kzxKRVaB26BLDX
CFtuM9PJ57Tus22jOZKOlUSBp4A4mtSjyT2Yc7JgiwlPHD9hskn6kGMMKAgZYy8ILvqiewpSTaon
WqWb91eslQKvDahGvduF/685GBq28ecdbdug1VnwIC2CXcauyhDRtrtIld3/1g/iZZh12H04c4D+
sVz6pjLMw3ih0J9bjwq/5i2RE9i/5JfbgPdWUtlDZx1d0IfTRCNICsTeDGns9jboBDo7idhCnQN5
78LdnIg/cxHFdArtzNEksGzjmm3L+zIc9EfiKvLd0rD3Isd1P9HDGj1oup/HnsD25bASln2Chnnj
IxWOLLEVPtL9QCFVTDWyaT1+2EKibVix+LABWpfhTSEnsztElIbasJW4TtC8QBjpqVmOTdgM8T0X
+fZOpTR0B7kUD3GeZxhWzKnR5VNsjuvNTFqMS4Zupvv3dEkTn+yXEeF/q+U70/InZGU4Ks1iGimf
kdZTVUXPXySNS1TpwW9X33Yo9xye0v5qRP/I27kjlwMuDMHYmpkf2+BJUrFYpwvzM6/JgPOtcSOo
vKOMiK8zpZOvQdKi6YW7htSjcBJi0x1DnE4WHeHMX42Y8P9Ggil7ATP9yAQN+e8BJmZqJwM16ms5
eWuQrOzdvhwa4l0ASwezKmzbmhJr+mgCEYa0Ge2uSO/dOKBNUeEuqmqgqriNQ0e4F3MZRHIZ0+wf
oQckqhr5eRChDUsawmVhRjL88ysOuPdF2e4Xt35oPP8Uyo1Fl2vNb1cQxHDiJt+NC00xcEcFk3Q6
lX0l5qcxghhJHvKm5H53HUVbqF01hc2rY0J6rOWJ/I+jdqTh+RpQ8sruw8aDvmo5cC4bPMSwjprt
h/NX14RmCfZpCjkni6fry4xNNkq8cG4I+Y9fsR1jsyRDhyhHLRph5ONR0OSokUwsWQunkdph3MQf
cT5o8ScPjMoyKZfnD2h3MqcbiYIN7+tu+CnSqYRuMCEN35kb07X2Zjq6Rko3w4jqEXRnu6gwUMcP
AkPCJXTjdVhbqZ1PI2tH3AoQtTv3Npbw+oJeiu7ZE2Bp0m5FW+blhryqLQEcbsHSRDE5O1D8y5XW
qZcGLsZu3Kl84SFmDA7u1GJaWcF8s2F++TusUuHti/cC+7E+Uo5MyZYWhv2vmSKgztBTbjkP2W6M
f7ARL5rAaiAhfRsLgaJvPS033Wc6TIDq1n5GA9XrjSWS0XrJbrHfKRz9WXQns1QF7JFoZhnCc8v1
98Gm2qlEeNCAs7qPiMymBXnYDdiaNpAH5S7svBQgvSy68bvwLZn8fWT1Wi+U6NFcMAHC+6lwujOZ
5OfWyPfgn8CMUYSPNfqrhIhAvg4qG4aoxq8FPkcy0GqaCtrRuwNXGy8euMkrp/nbPi+9dgrMTMNt
ng1mvCFHGASNOP/Z7Bw9a2myYfEvb6XtL+Wabo5B0if9MXVb2mASzoe6qcn6blahzcbHHTeNxN9K
l/8Jeuq4E2cMNAP2e0je28+E8pOhnNJWokufDrWGLoxy/85E67RM/YnlMHZKnCV80bXJ2y4QHUR9
292Ghqz7zWbFYg87mmiji8hrqCikAS5Vn8QrT+mYiB3XVj2k+OYW76YMM7hafDfGkMSJJBl7DRvP
P4eOhmJ6Dc3HdtphI/r/BUo8QPQVoZl8AkK0JpN5nrOJlXbYMwKXxnNtH5cxGfBKW+0bRRKN8Xi6
/gpAexeWSjO7BIpUr5oQVWfMm/udYhBivAlamVMLqwZl90ytEQ8C4o/snciMFKwEjzMpbQXZMpYl
VX1wX0llFwdPTF9DF9WYDfJYDlHZuGJF/ET1ZyJ0G3+qeND0ogNZ8htc7LN/u/zUad011EqQqWA9
6OS9SrZ0haQWp8x/TBkCivfiMWZkD53wegdVYs3ZUP+2rTNt/JWTozF9aRs7u1xmeiUmM0Za9LeH
9A0EqVjiNUMXjuy7VklGDI8CzYRn+thohBv8XRc8L0FUBRcv1m9iOfxWZk35EVdZPbwviJCiiW1g
0BZTcE3ZHz1b4C/ZyVKp+3MASmcUrucwpSw+lWJxSSItLGpXfoyAyr9h//2HAzrnseX/r5Z+ctDz
acxpzAN41ErQlVHcup/ctfY9E5gw4yWzMXATyTaGDm0JUzO24v9B8OUNFyPD3xvbfw/JE1JWWDdp
Cw6QR6F5+Vx6Je7LtLZJR+qn5MPD7xwd/oJUtvRIWlqVZkv1I3JELY5AU1/LVhFn4ZMN8HGhO9ev
0lQXF9g9w+pjSg3wE48e73di/iJ7HZ8XFh7xEoEVsHUq9vSM41axib2v6Pg/o6DT5eeLYgDIE0/f
WqKA3/OJQH4RocMkPdSMt5tDwlT/pai5U3Fz/gBfTERLtvB5UTLgRo2T8vrLMC69LPA/Kxv/KeU/
8Fjc2EysVEnFh5uWMjKNoF6djnxqi4u4pCqc74tY7Lhy8E03ymtKFWmPlRAZMmaW/aZFNwv5fKoV
nkMhwETv483HwCkVg5chb2fTVhSUV0cue7Wa9uLE3yTj3CwKD6Gp5GapW0AdRbqxj/2v63DZTaAR
hq5Bm8syA+z7UenDbNaEZcHmrZcPHixMpCQLZsv59iUOcIqQUhld25VxLW1LxDbVkJNBue9foQ5B
yjpv9tE5nOI8MYeT+5e9HUcL2DHscNdDreLU/CJb4TxGLnHU+0dqoRorf+4ZYgqT8cksXXbr7WBs
udWAspskhoM/3uKaTpWdTwtjEmz/9OtcghFnArGqhpWqjr1hhp15HDYNrxf4/nyuu/nLzh950TFM
o+XP+zy0OeX+LVNHcyRCvbRhdRjOdtyxFys3aHNA09TF5yrVv6rub3qbobJ431mUeHRKe0YTTili
SjLl1Antujwaz0F3onDqG9K+9SqVWWThcOq9uZL4BQ9WQlXoJu1pvr/gvY7mLCZjPdSygz/VIwLq
d7EneEC23i9sXEh0bwnOLz9zSi7Anc3ex/usgY+bVbIed1UzFvn3zrGewPieSOWnMPKLhOam7kfH
sHqjw7+Nzl+NQb+5kogBo/Ar/VggRYm8NpNYbE6sqDn6C3meXZiKSySETL+GcdlfXIoY3u6VaBn5
iE+NftX2nUEGquIRLd3KAREOfteMGVMED2nGDCLihvAZxp0/iBccJE7P8F+CnLtmeiDD67c8l/xZ
is3Xa4EC1vhvUsgHZsqDaYTmtcihBglnoHAF1n+8sRsdUh8BWX+josOLbFKyXWAsggCOm8PA0RrC
ESd/Qm3QBCOK+y7fAshmREDM5Tk+3UL3fgLC3zIHAHNyEJqX4sliEgG4JaG7pBt6LasaYt3cdoMV
aUtCOi3pR3KlsVFG2dpbKl3Pkb68cPnUE/Lu1kJrVXRpj54N5nCl7tONB6FR4atsnaRWEbp2nDc8
wSFEHDuQ91orm4cLFblYvKxwBCbeUQTELUU7jXP+T11t6IhMyeQFIgDw1g+IuR49HqELkLGZyPQt
YuB2uxWOpoATAZvp41n1pWQ++emhlEINGqWv6AOjlyAJNERQyPAHwzf23PbXhChf/SjCa/iUQ6B3
sLtsKadFQ/ZpFsmW6VRkDysF2uyhYUoEd+YlPUbnl+0FKo3YSf4WQ9uWroZa/xqHg9/NaQZ5QwEt
Z00Z5H+dki9e8BTtyYEUVXdqciKE7+fPDx2f1ix9OOWgnNuQ0HI3u4rpDrN2aL3DNo4EDx2a6mAv
kll/dTd+anTr4H6FI3Wl25zvim/9aLwVb4P0TehP21oPcHpC8Zpgi9LyFq9l4MDfxgvKQW31N/Ra
voT4lbUoN+cbhRB68G5ilIdw1UfMBhHo58GthKUqawGtfj8LFiiAz/IqbimD56ijc7P38XTFUplI
51qRKDqr0KG3fjEOuIttA5vJWq17no+WWDD4BOaz6165Q5NIBI67yKp/d4WOKRA0Tpa6JiyW2ccX
Rpzd10RzgesOb6+40KrYwgXutsOID33LXvMZt96ldg+ZivwVHigJS5JwpH2soW7h/c0xpJdO11U8
eiBjPDdvh2RU+D/Cgw6DM1WtxffajYEAvw87afjXEpgis+411LEWH0WqPkGM5ZSnza5x2Ht6w64I
3VHo2hxCkOL14djQqnVRi4UW3WBmGDj0GZ9NMYvmzzTJ+2EH4+KGdFKnpg+5+PpaX0tpiSBXyBUD
2MF8JHnT56p9g6ekqFCZinO84LivQOTJnYL9FkSLJ758NTbKShy3YPj/zH3V8CrUyU6ffWjkEc9B
Usd4jze9oFerVEVJBeJc0zhZOXQeZirxGrIsHaCSPY9uVwPxLEqOAL+IlTCTHMO/+bcv6e1DQu8S
5Yqi2MbslMQxWVfBLOA99Tr8eLcd+wiP0wbZ62OOEzCj5hskH/xwg2mux6fmXSuWwzcxSuqeTror
AcObuU0kZnFypCdvdY5GpPpCh628vU3/eSbizoexfiN91E00kQOLVX87TcVDIMj4XHz4h4Z+jBxY
nmUwHDahATSzQjrEvKgqza+J47lMduVfRdiuPPSpqIShjw/b3wo2UoJkDDdsSR9nqjAZWKdXnt1/
eItHU9UhgtBE4EesZeCSQIcU55JyGr5FEmyROJfxSchtcUU/NzswRBw1M9IpFKo7HbszCR246THU
gqY6DtGqge1MC1eMHpF2CmRqNjj/vwxh2y86shvnoA2diABIF1POUCpHbfTsLfjbHhcsZsIBls4k
Iqe5fILxqLDEIkWnwzaPPk3/JAIpX5GtK5Csebed7Aqvz3hgT3vs3sh4W17BSAeRgre7QczmYWm9
Ibqp2g41pfOiKzAPpbtQrsV4xT3XdsE71+Qjj2XdWwLBlarben9CdTlbs+1y7DFwgXtCjG/e7krr
n4l6x1tCb5MmS9pFdWQf3lJ4K/t+bqzjBHSiC2r1rOG11lvnqOMjgvYOlX1c42j+YuxCAcL1b5RI
HIFyfihJ2ECQ4ZKcCrPClqarhJ9Twm/OJFirNV8+mIlOtTc688ZzY58Qj7qV6foPIiIFkpqN3kGO
dtaptHU6XoF/wue7HOnkF7HnBMmuTQOet/iw67BoaeNn1Zk2N54u+pLMkEgfOIRIA75czyXunkFm
T36HEGJyAX2qxRYpzfqYfAJWaetp/lGu9IvcwqLT21/oLkG78Jwk/D9oNGpWXhCXsVHl2Q3HrHYx
4sQAy4u6K9TQC+RZlcAJ9r9X8O5UJZFKLgZn900hzD991H0voWQyGUrfBiUll21Ib/rv/g93cOE+
6dsxfw54SYdQwTFZpLuQM5uhe/Y6WAcBT64VL8iJqi3Uk99kzEtDPuWgD15CtJyUWHB/QqCf3x2z
jm9CrZw9iNdXeUvGYHUSTafbxUc55VDwgUWuHsbfO9/SWHHWXeLbbJJvZySReAE4/6muI1lN7TGT
tF7/f/MmYsqBrKiQJ+IYAswtQPIj/UecziXwWCg/q16jrPGESuUPmdz13M1htMXWzk7GNdf962ty
c+HMVUJ9lDTwMfqPHMwhn+SL0367c/Ukp826732DIaU5rkdXRDU14u+CVyIRcfwGOWZSCTxB7SWE
geELzTA2iGIl/NhhFBamR0G9FQQUzFxhMufses6RrqAIPY/8WxybtC+BnlylHWnsOM8GhY9eq+rX
jJL2XJ8h4gV74D07qAxcVAgP+CvM37KoxUqX13yzZwJw/TJUnPcQfSEiOsZD4g1h0YtiUsBCIxRV
OwhgMJ7BmAUny1pX04V48gV3ZPwicdePSmK24ZkPZzQfCDmX0VXnXzXP8c9fiEBC2DsyfLY9fEAl
PfQjrmxzNyxHvDcb0ky7ctCwdEm5TSvMw0pEBogx5uSJwP05gFrB62k4qzznmxmTjVuCvVmEE17l
n/RbFnrmBB4c/IR8XZxNZLHyLGiC4vUlgoke6RS22UGAamcdTTDD2cGKdtWfY0Uwiihw2bVUiKKp
A+RewEos+vWQkExIa5RHb2fY+5eKe+eqcejoEaC5FbeFTnl4OF5h/AtJKH/tDHC+d44shovqMKzK
uki/Y1gsoIcMdz3cMnRzdA+oQL/mW3o1LfjDa+11frEVTtU+02dBaVOLmew3SKCsQgnSDLgA2g07
evOILVSx7ifpa5pAde1EwtjUw+82TZ/EXTENXF+efILrZtubA/nsxJWYVbV1rbgXEdd+p73en9Al
Lo1o1PAbtboBdaOz0V2tS1KiEtMU8FEIxvU3mcSP6vz5I70hUcCPl7kG2oxBrtO0Pi1yLcyyuUfH
aKDWTF3kAJrutAuit6UvNSp/Avd8gMTb1zBnQS10wuc8AGlfnbM6Xg0VR3XhXFBssRyvnrK14MLx
3ILg+q32SmMFSgOBOBQ/kzJ6T3WoZ4d1T9Ps5YvvIXXmrnLErb0bEP1VY8d/MTHRgddEMX3pWg04
3Tst6XQxXgvtxvvR+aHtFUuTydisluHSiYPERdqTkbh08d4S/HdKQTjWR6WMKFm+Wb0UcZg7bfBk
G2DSXPyx2nt7/LW9MsvTLZSVBan/UoXYZTbZKIOKy7zkrY6joX4qCMZxCgyVJX5AGJVaY4k8sg10
BqfQ72LGG4LhY9LDeUDLd7fqSYKlNl/W/4Q7D5RV2gckFM1/q8xZKgigG0drKosRN97lIrBVRlnj
VU9cMePMjwIUrcl6nbQRseReRCP+ZOvRKlOnG5wSTh2V6gGKceLUmj+sqpIDaw6xTT0pyvizvbkY
9+Jk3SjjwCVGhM2pHDK1B5QHAGnKXo5qlsIUYsGbrOvEOhNjClrRt7X+gj3isHkI/oLsWMQQseip
5Xr8RQF7dQdB41IPiJbyxMEvBPeFkXGaXbvkXzfoxeC7qzcH5j8XaisZk/mURQIWFyKLynSFREcE
wt8SepoPTVSHOFjqk7sJZ2BywVVF/+VMjpmnZbPw1g72cExsQnLEtszu0S9XQEwXk/X4hX6vBp/w
pWcdPMiAyU5dYvbFhtOQqexxOvDunb/aDuV2pFoFmCHAyGFebpsrYaP/T0bQcfSdq38O6ITTctIZ
PQ7BISrXJ34YKYQadMYL9rFpIOx7bJhBGICjc67QXpisl0WYwf16NPQGmGt96nj9zUFQYjM5BFWu
3Zf+KtewXD6hDuTVtcVlUtN8G2VnbMIYS84usg0bBwKJSRrpLUaSPzSEcQK84uKwVNg6dkOHKmto
PKAMBx0aqS5fol+JHIB0cmrZhRbjgCcaoCQy5YNDIbdpvaW9tEJsq72zaNQx4zBPUH5pE31OsMWJ
Qu1Q3zTWBhmeYhcBDXKvhZCq122Js/ns5Mz5S/yx1rEAnZJ7QJEFY1LJ5u2KRyfg0iCnDhHxhnjG
YFGU2uX7DUkOTnmyq6MPGWM3ExZa/J22l1mjyXHYknSuSWJY3i9A8XeAA2Tcup2MEwSHcT8EJJE9
kVN7FopCBBxlE0uX+g18LJu5DXqGUuHYcMGGJluqSEJYZGhC1QZnzxHhJQmkpwqiW711/bo4cDrS
GJjXM+4bz9EYzN4OuW0YXiW1q49kIhsxtqT2ZCXVnmfLBGSefz1LXd7ZiyTuAQV+rGyQmtCPoVEZ
hR4FGkPLoxcpt8meBDI+1ZkAMKNCB/pWfFNC/rOarQBvMYrITl7uNwqlGTvumBjjuD8BkNvq5oS9
2hen3ieTDRJv+4T9/RBxHK0s2PoMMbNmB1AObbgrM9z+pC3aQCWuY1t9M41apwLsRRnUl39D1mt/
sgK9H1SJUKvyTmoRAlVxNi5BhdW6frsxLCHz/kg/FjJIXNQAsWUHJhSOKYVkL1N9B3AE3DmRZAcO
UZy5lYpw3/pJaYAy70wd18XeezLduKsuKvXiuvGsMs5yc/SUZRUTaNLUg7RPHrc3Eis2YbetvGD4
5I/rMoMgkPm2jvmi0CKYbH8V6Jw3l+ojZnPQEiJJh3NzNucUauVO4MU9galHlhcPDopl9yn7qODL
4Ysm0I67qRGr4TgK80AoZoqsEvn/QAo6tADMhh6ZQRBJCdUD7jNbz1MR8UnvDLngLiL9csoK0q/W
Eqh9wpP4yRiJtc9EFix8evIL+A0QTQkykoQPqHvu1QM965m+ojxsXx/Jccd2qcwJ+teCi9om6dvK
Swq9Cmgog1q6yuKCnRclWDqe8ofMgZ2GdfWqhn6lQRUacZYUW5tE1hkH82n4Gl+VM7Lwl/SQUrnI
AKQf+mkpvzdGeJDLBfyjAWpMa8bnPVuMaUsa4qp5DeP+EkiD2CCjvNCOWMzXB0WDPKuOSx/lIPs6
oXiMpk0lWXidvFNsO4K4AITs19Ul153Sp9I2hSePAnXRBoE4ZrYIR3qhCkx3Vnluw/CX8tUUcjyn
DKU+oFsDYFuYGNFwRKVs7uleb+eI9fcjoeCOfPw45nQ7s6TeWu+9NJBnHjBvl4Mjkux4+mzQfc2v
DalkUhZxVv337Sute7uKNfr82gNFv/5E2nnzOY79j9OMVaGwMhYW6APSQPj0vcgf9e6Gypex44HB
qr9kX7Su3Iz91mEHwDU2YaIDxefo/VFAyaprP0ETZO3g2jfcbQRQCY2OiuytfxeZAdK61faL8rI7
gkGFjA7c76yoD+NMwNbeSJ4PKqALkGEBWWpSZa1LPdu5UKn6bGOS6FsGWCNc/4ZNkd9DqMxohxla
UoTBPH3hhaTJA1lhjSRs554BO3xLIj9XFxljLgd86aDxVkxEcD8Kbf4hp1t5FFbGDueQOExFJWXW
HYut438iKcZjOXf+yU2mBYMm4qLGlmpeBx/WT7zMzhQqaDJqSKTzNXee7RRBeWuWVAOuxfxiYzg9
rPnCV52DMxytE4AmzVXRDQk6suFOJE82EkT8nqBa0hFMVujLSvV33tvIvJHSFIc1mzL5nvOvC1bZ
S7W/pPU21lucoW0aEGSLJGoPdE9/p1exAdlcqFuImMu9wghLa8oeBjuxgZQBFUbqy1IDrkbWz2bK
E6ElrGgZt0oWdE3wp4NhWtyVRwerQXIWHZiI1umTderiSkCxGkPDnB/qyC8ctEe8JNTVmAm2Pxaz
8v64/GcgEK+9BPXcJ2CDZ6DAz+uPumHFfpQBJLj+Iby1TaRN6YEqORJUd9T46fntpzx30Y3SHSIm
AWwTrGdHYRc57JiPpOTnj5fb4Vd1nfe7O6DdNDoN2YRQGG51kihx18XajG7hsLrM/sJKKaFwByWh
nlA/hf1Tb0dthiI+a//VPHTNfeuYzf9H6Tac6D3cvATKkSAYsZR3QPtv1rvv2lYlRhH1UhvxTvbJ
iFgC2qu0pXpsYYG1jff0poPFgIrYTJU8rTsKHs1svrzNZSLrfleaGq3rNipd1Qb6P/csm1tSlyNd
eVuZRwK1eruEEEF/Zh962uJGLURlFW/3qioZa2Gs7Cg9Vt3P/2DOBPzRZW3IL/MFBcVgNFUqI/Go
Sq1dmjZzYb4mriFiMO1zGRIG6mm+aONREjKbGVPvmDMfyxy+AfXFs0MUuNs8oN/XK5D81c5z1dzI
CrFgPHrbNDFFnS6t4S/3KpLy4I0HwY/xIS/SykepJnZqMKrdmkbPMp48oPKH4k1E7nP8USIYGwwQ
OacvlimIc9TdrMYSx40XXbsbcM4vGrvFhmyUfv+RuFoXUxZDscTUCPztzL1kLOsqJXEyJqcA98Ze
OhEgdc51+QFS1kXnxODD+9YYbtfvd5bylP3OG4J9gRU1KdKGVP7yyK+Je1UqT/04Mq3mRMQu7b8V
fC1kZUMmb6kJkfgU24aQUMt/Hqx39xAu2OTezKRS1Viap0xoce/t2PmSRZP2wswfdsR2kA9p07UI
012sUfHf5klGhCB7+U9sIyqyL6OhKmKCvXiFTmC9VDXwZZ9p5uymTr+Cz8Pam3R1hM7c2FBq/Dva
QJe0EWq5v1BRivPvLq4p0640OnWRefm4AfyN4r9d9Ge42mUz+2/huhlF/MIncjYkt6GeCTyevSHk
fHoRCyb6+KqjZeG2bhlLTZm9kA5LKxSZ4JhU16VyZkpZiXp4pGVjMGxF5U2vOpobeT9oekFPvTO2
ZQowsfE9jALTG9A1gr7gOXI6JXX1rnC8ucNgbvtj9leY619iXgnqbQrg3ds9xfBJhmYvowzu9azF
vsKfubmBIJw4tLJHfnsBZIVsx/+ypDtHVV0fB40AeN0/Dj97l3aLpbCQV4FUrKY4DQrxvOBdnRpx
uxh9ZcMJuDCcUmpHz1PDaYvivJ3XUraUotdZAMvDUPRXFTxC+nJoQO39tSBMBd7yt4L9+/i48nDW
zAw30FOK+UyZK8ImyP90Z3gbg6FHMztuErxiYnAAk3dOqQ8g1wfPSXnkUMD1oAOsNAHM4ibXDgjf
BPvQnF/XUyggOqPoS8SnAcDk+jJ8gUVOGIEDOwDoIy0HLhvf9s3mXZXdtz3mbxpxQtuRFvI0hpXs
m/v1b6sVQnWODjAp3omiYoZYo011nfKdSrhWyrq4zv378FNR9fv16MzaQTN91UWBGLO2UezSic5e
8XCpG1L+vGViMRmFbBPeT4jiCXQBs0Iax7wt+/9o4mKfG71d9NpCzZ5yK6l+nrHXJV1AQN6+4FuO
E8tqRRuI1uwUE3v3tajDL581ZXmN7Y0qIYZAX1MJrXT2PuUGglOpQMkNnrzZK+91eAU+3MveK3Ni
NnTkS76/OE9qeq4986BRzH9FXpYPtGig05arH0UVqqKZ42zwGCvDT3u9xvLFgmSL0XQA2+jKTDbE
Tf3jJeYnX9bWwSk48qclUsI18WUHFG0JjTF/wghwg/yY0k0VZciqRDNWVcin3hOC4A6rkAOKMCTj
KdP3O1aU7UqwjgUjC1LIHL690lDQSRHUnF9MgfF8kvC/X0g/GvHvVbLy5vzWrCemtkXbr+TFug/M
k36vsdoE74j7W2gXAQkGMYfIH7CjRbTtvOuZDv0Iha98Nk9l5v2QxwZHrtSx3XQBB6VlWfUePDgs
jQS5A+k95LCb/E2vkCHz8kqtNnc9Bbo0YLbVe1TzUB7Lr88xfKjK8W/1iCMdwxNDNOIIoRG4fn4b
rbAOdXRE5mpLcwk6zrZjK04BGuoHcyJycQMV0sELR59lk61vdj0ygCRwefWjzy3nam7WRBDBHMYT
OUQDY9iNRLMgfxYDoIO7H0/qzEsaf+god985LdWN4ho37fNSJEJgErvvIVwMBFU/xOHyYbpuIFCa
o645fBnaVnoMhC+X0/Iqpeqrt8joCl4w2ElJInmZWT8lObXR3pwwdI27/xazFxxh5HaIK6NqIe2D
CRJB35LDoTv4i+gsN8yGoNwk54HHoGCrfo7Vlrzf0aUi2xasubzdsQUvQye7i8/GFfPEXfLQq+dr
11tkfsT5IdvPYOGMPbxQ9A9S+DpfDz4WYx/P1otqsgbil9gpsv+fWnNDaOQNRECvD+WSJXFQQLWg
o4QlaCpE+a7XreUpL7hUzpjx1C0pNxqEb9FHnXeeWFTPvrFD6DmEfVhFYe89d4hc28KCfc/mjfRP
WFsdxSr+Yc8wQI3oK8ELfmIpm+1sDqF2Cp1u/+2FNr/GNfBO4lcvjOlHnBavSCgK7TfCTViT5PuW
ropX5Fw/EjKmZCf8GtCowZhdNVOzwYFx82mOQ7qUaLfcej4Z6veOzNx+3Y/YACrtjIkqGrEtQErE
FfW1w3aI2xWy4ODh1yjaXT0myqBfeLi21JcPj/ELXLp37TUjvY4/SR/EworqgvAxK6m3jPQr+IuS
rPUwLmLidVezuAuOndolNztTSAsJgVqlW7BK4mQj0RjqMatidiEQEkT/3uwKI2suBjfM5jf1EHUB
2Zz4EDAM+HiaVO1l6um9JA/pBXDrYRTseLl6V1KfcZYk0qWGWTG94xFbqJClbjH2CKvkMZq3TOr5
aAEZUU/T/E+BMK2kbJz8wH7noklpfGkn47850kx6ZBTmlrjXyo8JU91sfcM+rLT4uYu+kymipqNj
pggj0DkEr6fN61SpbIlt6nRPNMfkmaQyr3SFyz79Df1tUQjQl3v0dnSNhnX7jxcRXt1DO4TXjA8p
TQ88V9OZg5ZSRALOFROfOaoqZ1+zTU8fJysGcY9dKPfQLnNWkFSdHb0TTXmnaVX9vfRz3pnCvQ5+
eRPL+t3rx9MXFMYqK1vKggyIVRHe51xOgjr92raO/ANR29FGluukvWP/gr/PeXb8YNA4TFoK5kPY
XNstPFuVuNrcJi9WUo2cCgEtUr8yMHCj4z2WFejqKahRUkvkd4ICrvHeMJfHZ51ucKef2GG8Uu1g
m/M8Qes1v99T4IgmPSTElKIOxbZj1UZ8LFdYu3P3c86K3mo7A9dQaLNNHrLmJvybxb6gF2PqABRB
G5aBa3D+FAb1q0k/3zUnDeclW90WDeLsnZRlTOuXOZ2/5sPq1O5lYPBo0Vw1Khu/HatRGGJR23GI
QFlvAKlYvhQV6ng0L+V9k9KaMKotgTitpl8KMy6Z/GR4ov/QmuiEOrh6oyFsGSVaRVnazvmJntRf
FEzZVZl0nJpeSF6YeDG5mfD8tjipSA+Pr65FFmL6zgsYmMEcYy+ToIPuEA1fPWxCr/SkpGmJioDB
tg6aZvO1uM8QaJE2RHP3eWlDMliOYo0npYD2UYq5fRPF4PAe1YfxNW3feQcBMevxE8UF/0+E7xss
Lq2bipRXl+gVLcmY+ABU1B1LLrzMyA9Rdz8YIKQSRXpGdVqez4lPsLrUlyI8yEdsNV00+xunuRjW
C7K7feVbOCh3P+NfaaHRbZcJgECLVgu9rgnHzfNAuUf/KgiTSPp/20JQ8L4r4sdRJTNYzCLjQQan
q9hhfOVxZRPeCTwfSPD+8vslzAjd1RBvdkk+K7RPVwc/2jKYSjFyM1tLHPc86+/IMQ7k/Sw5cyH4
q2IS+ryJngqAAumgCjfRaGd4wlvL0LogyFNcDcOFRcG6wFqeIFT8nRvsOSlaaqLDBqshG6sF9FNN
Ckm9sP4M5gtsndYHgU5MfWXEjwrhHqAruC04ZRu2RbYvYeq6qjpbpMzR19U+LKd6a/3V264V70UJ
uP4KI2iMhI2YIYv1YcLdre8LgiOwEutBkAUcn6DWkmtdfyNrc12+t1e/ag4YJiEU9GPbG9o+UxpO
fVk0rBVpu9xJJ4rndFnjp4fd3IaR/2WGY1PiLGFeCS+BYyHRgQJOQOyGalhoJKnMRTop6fjVdQ7S
H905T3k0XYukvyumP1Vf7d0Ir0UsOqtJw4HhxNTfJAEO0OkVszmtjqwZLbTyIilGcBY8XLJ0tTth
nJbg9AXRZ04nl2Nsd+iPtNxTtPsU5d9U5GVSbjgbXXs+unYdbXlUEp8r8HL5mtbqV+q/UAoq6uCE
dYaIV4Zh2tGy0Zex3Ykq3EzcYqs6J/OLsazyTNgZRhAk2EpxGtt7vHYxDx+vZlQCwiO4KX0gGW+j
qFMqVWHiozuBg8E2SFWxUXyRt3PMXdfn02cGDfjPDszpBJ2Na4Z6pMWQ1fZ91li+bLoDyT1kF4xp
hDzkuDmzluP/8jiojOTrRzM8/Aa1Yj7SvDL2+sGqw25UC1UMEwClHlWsCXwHV5TBaZybrV6LqmW1
aem4CrUmj40w/ZX2puiFpg6fTK1lzx3kt130gHBz9lF/iodRnwIqRbQLl2I9rtBmKUbEqCs2BUIr
HKKoZVfKN5p8J1Pq3IS6QFHDmWhQ9gzSoUP3dxbbr8lqB+4o5Tmb8CCBuCuk+t67uvJg4RklXlTd
vi7YetusEGgKKbSQDGZlXQVAJ1zKxTH2ymKqebf9sRM3JZabYj0nJ5H0CR+q1KHwvQl7XEEJotBJ
PXfkyY9mJkkhH042Dp5HJjiXH5VAbMik811FcuASjJZr0Gsuwem32DnGC9ASEs1qE3srTkrTAkDo
LwvEv5ltF1Zsmfgy6KuqjmqklewSZmqUcsA32DSqbHz2rop04RmksrM0/MHN1qBYmDCB2R1gvFiS
SnUU7ucU9ybGAFlHxZ6glc7mcS6/cllGNRMM8wHJM1g7zMGs8/+8rd3gdCj03b06rnyGYTG6pYVd
LELqOCgczCWC39L72IqpjZgD9cayy51Hvj4SkA4mikRwSLhA9ZssLf+IkSu93UMfY3QOtFxGnVaM
qsz/0teY2GIUbxakn7u0cT0P0g7AFkujwP2k1r5sduBvYsO1k96l7gyIMQkpSWd38sSSQdQRzr26
6gRE1CowlOZJ7p/ppEUZ+IZyXvcx9mMj2GrUGFUWp9fdqRvWFXKdCSw5aMlsBLyW/qUK1WHMyblQ
5OjimQ286y1aW0ii4tN1JEpDcajrFvAzdcFM0Or9dG89GeDxrYJBXqXMDYxS3TcUD6rhoImD/260
9U8Vt7DsDgel0q0RpxprBFPj9YJuWPft9WnA7FCu1EamXIIlwuosg2ZVvbzoET9m4HwRbVvt+Qbt
Zse0gcz2sngTNIZQV/fbMXEk3FEXF+KvnfJug77SFUWOjgHQVVw05lVqVxDsyzBdqGhlA9Rqp4c4
iBhWvn8zXNAggRbO6LsB3Xx/fXk26PUD9WpwpNYAhkDQn/etflBY/V0LVqOAdwJoWojeu8sFjepF
hkNn7oK9/TZvaNtmmO1N5iqkI/OGJ+qe2f91i7fbNXXtiK1wVk0hDOSd1fZlF9vb58Ly92qraZh8
wEHid8LL+aZwXhxnvguNgKqGNwiISB7RBCKXJdIiNCnnSp38iliMEZCtHM7pDySMviPv95Qrv+mf
nhCr0QRmRhkJDnvjXHY87lcofwqVX5PEyV6KWeyRQ9+hownscw2GEjT8ct544Ob2EMPxLbqhWLiL
uB6KqbPqdfvLvRVda5vkhpT1GjEcccUYDMbzkOru7RNXaJ/SnzEa+CmBhIcRveNjFysTb43aA96J
Uo8HGPxa9KuNkSpYBdfqJl6QUyD2hXUm3lqpIWolVGL5z4LcChNjWQFo8N7Q0FTnCq74jPo8GpVg
HLVQYGAcKB+JN+MVZQMQvXrFZ+ro+5GIZoKq4Bk3sPp1NnJRKu3hGHlp52nsiaxC8kbyd6ckRDqX
R/31P0xfo42PJu1DIeyQmj6MmnoQuovDwggveIgddUMF23YVa1ILEm34YBFSIkTS6PyGz8fCJahx
+ROUAP3TmgEJRD1UteYO6jNRUnBkDhO4XAjfNCAIQCDDBrIlesOiQ3N2nJ1b9anmNKfon/hf60ec
baB0N0eDspWbYVwNG/c9208zNAtMCSf8akZUDSSzMtx6HI7FxBVShZy/snP780/KZw2o9FZSdRFm
mWM1bHfYgKs/Ryt4jf64SjH6enbHO1zjbYvTU73MRT4Ccj05fT9cIS0wDkGnPJ6VlYOvjYXVaG3e
w3CEgHhD7sPWvAtu2b6aZSAV4VwxhpUT0AHcXmcpyOd3kjmsuZQM8gLo5YUbhlk3KXW1f3edG9bM
ePxJuSUe5tCR4rw0LlHP/mIpBE+7kpGUDGgHVkBkpRfBIOcUL1O/7A759IVR1z4OrSjCBjk4fef6
9FoLlvkXjp1Mv+yo3sHKwjC+9oQIQBYn4VbSjGW7iGQoxioXLn0cvvXXFFXIsjQJ2p99TTnNlNS3
J6eOTeMS47PudI95m+KvtyGufBXkSAOWqQlqSDwxV53WnX57KPHblUOhmX3MvkzPRMGZWXOxOzYG
C2KJGVylYJxbqrznveB6JhKyCT+vFp+ic8QczlyuzHF3nBg885NtvdKZR6fFHndKULTEU2HlNPLX
5Tw0JZhC0IJuoJLmrKWmpTztLYNMBG3tGVKOBL/ko01OFbXThPddYWWQMYcwZ5fqcWZvQLsxHjTX
3Bo0BYOZudMNG11ilw7o3C/UNt5xfb8GeJADQWBhISmPIslaIxe3TY0+MiEIVVGnNgmRNa8mz1iu
qZlMzwwjm9cSoO117+z9TQqn80sSkSIGeix59GSBbD+6e4OcK0El2xiXQOEPuMPE8YXoik2d4CjI
hCM+aiDjJLwlq5332ck4q7FXFz1DCAbtLfwU0fKR52Hv0Y8m/Un93YkbkcZI7I8PMbDluBg/k5ww
zUs6QMnZO4yhCZ7N0DmVhK48zTMZ7iKOkLQycJB3jKMB0tDrf5Wo15LpM/5tpxA1m+QQ7Ze6JM5j
GseOiBffR5I8/KC/e70MlPu9S1hB45RQcgxJfWDHy++t9/PuPiEevvEHJG5oY5qQf8s8Q65L7Ctb
bYtBbIbQjFZZx/F+075+I/hfidBvJJ0msH7GdoG2iwqDtzr9EFX4lo3GxNhvqecLi2YfPnfTUkeK
XX+St0Ggj3OOJn2hwSmyI0n7ciU4nY+2YVmuGMAgEYbOo3K6A20rI71LtBmgVYSOtq0g+dYmuEbW
WQ/AKC0EDkZ6/cvSBJpq3MhI7Q0APLYOpaO3Fhdfiv24QssBm9iE6rglJmqKX4RQA/iadDz9ZmRc
ArpX5Uvmo1x627TrxF8RiN0X5BT8wlWui1E5xIa72rgG8NsKyNldMZwR4/UpIw1DXhgOa0XHAtqA
ZL2Xg3KMfEoRMjKtdxL7+/3af8bP18+fnRP/p0bPrReyAXNCNYMohShYuA7phduzft29CD9UotNT
pEfP1+i4OKtDWtG0u2zN6199z2nkzDJ7i9kURxUFSYFNfr1LpSeIdIGL+HpuGIgj1Yjkqy9DlY01
QQnXPrO7vzcavuouI6ChZJ+a40YjtRTPE20Xnm6WTh19uR5Wr0LMshbNix7bSPTaHby0GYMYVA6y
EHTHzj8RkhlGzqHoyL31mnKfl2OjXhU1JazKtXz6toPsXrVJBaIYL88h//N/g/MAigaiGbDUoEw2
gaJhP9tYWKfKZikeoa6z5eEc/m5JOhHUpssiBOG6j66UPJq/C0Gv6nD1rOoY13lE4001kaF8Jx4A
XBEpYZPtvByQH+ZFGzMorEMMRygkkA6usFn4P58DEqdI8hMTYmpCICFPLK8VVpk1ZYWNNxqLVUEK
oEbMpMW5v/b3LSQyXV5eZE5pHVZe5gVv46gi4i3S0TOhVHYKEdXIxnosv+P5WxSJdFtjkSkZjFAW
RsnzKfHPRte/uXwRf2yH34tFk4Nc83ohl8TIfDT/o4BjiSNAdfOfnw1e8IS4rQPnO2wVqTMTZ/nV
dfGdUxmnD99V60ZQIH/EvJdzddWxdewkWiLkKvbxepmSEJr3xaOy4GRnKo6aCV4M8pG4P7099+8F
meFctZKYVPa2iyRIhLenOGU9ubbP4c+g014q1FCLCYzQT6wzu5g9VS6OMGrn/XpEqk6JOsA42oIX
RIKLaK7I40rujDIOO9r18dQkig/bwj6xdIeaCobe+KBcZLVEjspLH+JS7aKzpUFV+7PeUG/KjXBO
T1Sv3mwhlJjGG5L6JBLWUajttbRcavAlxprJtK3KqpIErduzI6bymsZTIImGmIU8NRZyZtZpBlOE
TkRVcW4sFJbjprLFiRbWDkSOyAnaVsetyguhWFpO/yTV+gsYlzTCjIUdf5nRBonVO5SkXrkL5d8b
exP7tezsTeJ/Dlwa+hWdFbit7ksmnL6igCEzyPX0/qAkehzriKkXKKneK8N+uCS2LdKpl79Hu9+4
D8z6gE411i1et05mrrj0ehhv/f74cCfxqaIombLJQZCvjWe9jLyTaGvLANSil3SbO6dkeVOQeW3K
2ssO4C62U7czH7m9J25G5GQI4gygscBFrVVKiidsT/XmqAnVvZ8061Lo3fe0e4RUs+ASbrRpI3qR
4sIWxSRYOk+SE9E1gGTWxxq7wdijyRiyRazCB/U3pKpcJ9KDu8dw57Bphfjqs2mlYVFJXdn+vHZs
1tdA8LsxxD9thumA9aV2LGomcGwCITlycSp/9mD7VLYYczQgpLgP0XMEB7TZkl5FCOq9YDSZM36C
P4c+Y2O12zhs3DdlxXxnSu9x0ewf6pp28ZQAEruNHN/OyDsnO8u/r96RlVGulcwEUiklAslj0oQm
LTrG9PHwj8sIR9Tkdh043WKDATp1m6mGXapxS8tgHrQI4Z3sg50KjbP+B0yphgOOcUQCBSFGQao/
IxyQA5ZTEoNHGId0tCnqWUcWTyJbfrjisj/rYaS5vzcN12tlU3U/0YcLVZ2yPJVBOAumLCGxoZdJ
epfko+BGbSYE3oLUW1Opa+bQb5Y6KcOwCd68/LrniHyvTSSFyIH0g7n3GQwQwfwf8UYNYGW8aNFV
YOwwrldr07gDAp96exo4buwycCCzzSM3yuFOw+KFfxsiG7l+vxwEblWdYj6cYbopiJRq5KbJFPzD
w5oiTCazR5mSxO70Y3JuPpCZfo3CKgjiTqmsRlAEtmGZtrXtz0sParNPFHEswf8GlfL8FTDAWLjC
HKi8YlyRixF244vc1xAHgzB+lAKhwpVNa1D+w3rwirV/zLFtYsBbcRSTdQSOrjddJdFYe0HmMVfU
yVFG6k801R8z01uujYT54MyV8qcjwJt8i8sB8diQEbw80LXQN0IIOFJrYHrfVuZAQpE/el4QFyH1
8jvaeT4B8M4hG7hUZ/aZ1ZrnWm+aYO+2F1cPlGx26TyKIAzLzgDDYe1EUz3CDluOmOSBUsNZIEXT
DZt9kH6yWk0QRZSIi4xEeYMPBTAZir3gjx+95J1IQ2z5fhRuZRovNYoMRXbVEHALx88OAA5pF3eg
nAZKIUAI+D4pBFw5WPW+750CalL2a51wJDAzqVem5B221uNCCDGlyGl3i8Z1LncoXPeM4SlMG1sx
981mTRdIU1x2Hi9q5C86cnp2XvBbSlbLZxgz1Ahx6hoBz6vcj67QBVmbvVQt1sE1+o0weCkap3FJ
sgLTn6zkWnua4L+oRiIpMxN9e71CWFcDVFqm7Pl8f3iMwme2hohl8K/5fE1Mkde55eDQs8d9DimB
2gEQrkZ20fVeP0Z8Hq5/ApTd7IKlr8MTSWPL5JZzjD7YpUxrX6YeyQMEiD+arFGKTP4zs++g52Fy
rkUK++15vr0G9DoyqXLeQpMyqGr/oUBcv2c+oAGr75WnA++MVMfKETtbrl3wR7B3z+HkZyDi8tZk
TDBmkogbLRFP0bBY2ooguoEidGwGCWgn5d6fJ2Du2BzAGvrJwv+SaeCLu7zfJOBjTd7Ne5uoxPEZ
BLtRlaO4sMpXvFdgg0tkHPQ49w1IpP6lATTYVkAx1afNcsaF7wU4081QhpSaowZklI+JpG3Ds2n8
wehCZpCwFyRItxc3QtlUuCYGJMQbLEZtf4udYRgsoRKPrLVBVq4DR/dxoqGlBO/9G7qJhHZzt6Z/
QiYMv1NcW0bqLSCmeep8Cwr8VBG8hg4CcPykZxY4PuFqvSbcqK8W6rI0H6zrtHpBYPn0yd/n6Itv
G5JZqqA/QVs4GtJxCUy+QVGSKJq65UQymsvQC5mabhnUVTbdh7PP+I012G9FvHxCu0Q3QLMe4R1T
7TUVe8TpiRH2Bod27e3xUe18N7BJszGoM10HsmvJw8WI8TQEc7MbtpkUXmb6kG92am9ooN9PtAaU
IgTjTTFYUzqyBEvbfHbmKgvdxUJ4LlYF2NBT6ab2V52biN5YKmOWvF0n4HAnxDHI3G2hGSHFVisT
vYiNh//4MUWjmTEB9n7wcym9o9UgJ2P1qStSu+jiwEUjcMayEf4iOry5iOLYrdsNfMwtiRMcfYN5
1PrYgThEjWjAJ8QoY5m35J/QWKf40liYtgBPjwBBNapJSv4lGA+ARpbxjuKOvmWCEbczX+NOBDi5
hklYqVfYRooWXqbhUDKvaGfTqxmEgtMN7x0AM1esM9uRd6YY3fyAYdyutX5PPDzUQ6BHNf+NeGz6
b2WbC1jmOmK1WMWgpS5yAShCsKNZsPj4fDtSaouDo1hZrGnPKpRHFs+0lL0d+Q/dc93CrjE3/HED
Gd9RS/7KOxK4Vj/Fqlai1IO5ytTg+DrylHLyMJt1pkTja+WJD7Ufymr9cBRsHmD/O2z7w9TS3zab
Poy0F9xG3lJUGtIBRFxcJohQnPimDtCDowMtOIfZEbEUd5n/e8I2/VdArGxVeEIHmEd9uZ7d3lK7
lKOsrEDZ2355xiaQ8MSHVDy3py0NCtuWkF+R4uOEKxRjgDoQ+7g29hFEFaUy6nmdsrr5ZJ09BF4X
m9L+zghif2KLYnCnEQ8wY37/44aUNJVbDtbxnj9g5/81kitYRtS1CUMAy4RbGFZhcAc9vIozQFLk
iehjdh3MBcVmoDNKgs60G3Pv77AmgpqY+XhRNjZTw5ZbokSh+4EIqr+m2B/Y3OT2fJ6m+G/3nQg7
O3i42teggf5gcdonwjMGB6M/ZsvPcqLuUjiLBQVvF8dy6YcsH+gNmvnNZtk78LYxkG512APjVRRM
9l37jC0x8dfQMHRYOc+GMc06DMF5v5W5w7UkxMey2X7IxwBEoj2r1UCmE92QRQpsNVz1Zxz5MM6U
LnuczzY0cy16QCtK5VaH73dkBYZOILGQuLgHL+LTkinP3BFD1bAR1AHomjtsKySSte5aZ0x1SC0M
/3XgY6kLSEuR/mYRCbf5Q6p6pzujAzwGwlt+F2MkWGy/3MSrwnss9tMh/NKYqEq/AmBH3FMR1Nb0
r0v3c4OP1Fq7dvHN45ripdBp40QDbbWTC/ltM8Sdn0z4JO1y+ndf6+IEYlzNKQZksZy0M5xTF+r+
+qY0F72ugdRPOoT2aTAl5CikEfZu03HER5RfWnjt68ccwfFVdBYFiRt9+9rudQdkQy/goYq40OmN
gVHxecJGVN5Ie6g2o52xI4NTpeYHt4QE+62Ud/EqRp4GipwEbBexpb68uEmURkj0Fay2HcF+kiIo
BzCpZltHeXMvNhpuLmy3R9KUsGJ9Dad0+xYEy2UrDUztBJA5fgvCx8i5KaH+XVlgB5+8tk920G8J
0CtUHDXFoVboO/Kw7/a+XjovnWTRlcdNSTklQN9/xxGH+rv8hZmT9Di5EGa07zxOMNzoiGWwGsTJ
52TJP2wsOuiROxxq1kROX0+wtMdl2X7PDDm9M0zsm0YSQiJrK+c5qqkpmv1aukrRvDkH4wEIHo1i
dMApqtBI1QAkq5wtUWbtyVU6mLJnVO1OhAKRsRt3fvXAbOBuY5VVeOKR0joL4wks5cg638fRV7UW
K08Jy8zrIE3/98wGttrgHpDL1Rox9uVz4YMbU5WS7FI3/BZwlNDucSciNQ3fRTexmsfKQG07tkZ0
XrI6e6q+56N9Pr89kzFnh60rYVVW7KuYxXOI4IHl/p/oDNRU+UjP0xEJ4oBGDjB1KxjeCBiQbXf+
pimJv8+zGjVp54bm4vnxNysjCqXl3CzkX4ClaP4JLZ3vaFraNZ/ZMqCEMVJQbsK9z6bvEaWADsW9
3PsetwTk+ytNBrO27RB2Hk8BP0vkThbGijLlzMwB7HRqX0nDUSOWBDau+BaiAkkSu2uh4hrQQjky
KNvvbZ/xtGvgqULe5Bp2+XAATkd+1EkdOM/bH4xIMcAnnE7GUBk4fSanLyxH8lZMGUFnj++8pq5q
7eEtbOsPzkt/ggaBOhCG+ABXVXGcGgSwHX2l2Rp4aq+zMLd+cy6Af4VxI6S90VzxKSL13HCFCIMi
sIZIoxXd3CbRyXu+wFRU0sXZJvi6hpoywDJ2dNrro11XH1hYIL4c9CH3eAC9GFyuaVBBDaDOZz/e
snrtGWjAwZEtpqKB7c99WTzgShuPII4+muFTUnornt+bNbhQw6nmYduSIYShTeVgXiIQEp+zYeLJ
2MgziTinvkWj9WW3Z822/FB6eRUpY+E9BM4n0bbkaqWCbBwr2fNaBt2+tRwG+pHHm769/Shwoo81
IvTmSff1es0TI9bI3PGqhsLvDtcLJ5zEQelRdCb1xb6xZvVJT79r0+wdvaTwogxMprt//2XoW5Jk
j3FBgmSzAzl5Cx5UaNmq6qbT092eQ3tzEoy12poRqjxuzOr9lTRLiwy9r4yGhbL7pNLlstqYyy4p
3ntcQZ5/4dvGaZYyhTaSuhrQte46LAszHLRax0nEGXNkPIiTrYNBWnS2I994TYv0gQnYtpath7qM
A7QFSdfJp/EggbaTP7e8wRE6Xulxl135JkB2Z2cKB1OiJk7MN7clxQ/13Y0Y4scQ8zIPgwH+9ok8
xW9KLzPrrnxgpavNXIaXzKU1gCn07pjsXIV5RPcW7rOUtXga0E7QYLhRB0lmDy59U598xy0u03x1
N40e/o+W64RzwkHhb+7OJnfb9qJ4IJ0fiKS+2yQGmhzaf9ucF5ecqBv0jkk5/PJFXmvbtan/9WuM
4oOkSxjx+NYE8xMOEf4aFEhC+UuA9ZTDw9iO/nRBbvVEEoXkj73DKJir4+vNYBM7DLehAqaDPPdC
rq8sh1pjrW2arlVh4wKMD64+mm/P0WIKcyx9JR+J/sxsHyE72rEu2R4j1JZIgAdjEIwl+eIDuJi2
5fMsozOO7slNBX8DVk9SfP+yXQHcSRTInSbhmOiPkB9ZP+pXKNFVfzS2KAW3BbtXaXIYNNkVJhEB
cLfznCdQ3dt2dGmZaUJ3u12RQUlV7BoOfEN1pIp9yL1T0msWUaXOIJ0Hg9Gaky2k6mDzV6ht2pDF
/R/y+Sh7lz/f+7pDqimcN/gwRCfcwOrhn3nG2m5PPOtsZb6oGdBCbOICj2L2gXHv4r5uf31fajbI
kdns3/oxHM/waClIpVH+ZyXaKOVKML+ltdIsvIq6xtLTAyOP3ZmaB7P/mgfaovB7iKeRnJE59PFN
YzUOHZpOuw0wYyGxFAfNGN6zoP0j9JfE/vbtCgmHWhsq2DG/Lso0v8nyymAPX6kBfjjYmJQOvXsh
ahgqFyZFcbNf5hAVwSOuhaQNl0fwViruMKznPslzIKh7UZewvv4g+xtALDgk5ODpJHQJ98DJUgHI
i7kXZjvWBVOXg73IosGeRLAi/PZ/wZmBkDjbIV7QC913rUvqBebxyIPbn39xJNafQmCQNIxV94b3
FqYB6r43vHsiRwdGki/jF4qDZGSjowFZRJxRqbeiM5BCl+9sC7GVu/3Rl03574Hm5Bq83oHvXcHS
GA2e9OQPJbhTUvH+cQ8zr7N4bkz0hTiiHLkG/eeiZeC3/fASDXx8B65VTyMRUt925JxOpuZ0s1BD
SDNRygyMxzYCY0w75dwETPwpmyk8Rh0P3aPEkUkNeFbdXbDmQ1SQn54g2F45g3BzteJQatnrYRFm
Kd6FtRXNHNYpxZg1Qs2g8x4TmZUA3h4QnIia5Fx7wIuIQ8IYlp4KDrO79a4SZuPxDiypYJMfAiun
43k+kedE9+BQha5Dg+rluccCxAoSM8Ir6Ins5X9ty3iSXuNzEpPJdQ4hLkiT1pLlYrd2aIUf+JWG
mYF8YXOdAAB9TT04mT1NQAnA79I9ZKko7Yl78t/TH69s2azi+VE1WUmQlj7qwVC09GhvRDxCXn8f
Ln34brio3qjU+NFclYjog78zCvdDW+93Ha0jbiEwk+Gnfvw5Hj4/s0UdrWCzhHWl6F2vm++Z51CB
S11Z6hgU21mba2CQqcs1zIFh0y1AslxIuXdDLekG/UD4OY8or9PbGrHB1n9cRZAugNtRNfJ2iBOS
8sBIhcrcftz50zcXGD2N7zDsnn6M1Z1JN4u1TGBEuE5Byl4PgtZd5q42r8CStvy9oMyUOJpu70mU
IXhxU39R9Lu6ne74MJg+86I/ljcOag9tX59zYLFvZmjIujcHcJ8nNLxMqh6GMt4JUWqJ1DwPp97t
1N1Nw1khFbSdm8/cflN2hKWMg9RFc2S3KhsQB31T5TQNk04spXoGPYzYaBU9irOuABfnzHqsvcDm
emd7N1ejIKH7uzDBXG4LJ5sG4t22SqzyVyh6pfLjQQumKdcHtQVbrgxeahqzyEqd17LNA2lV+/sM
W9T+ykmp50F0ksYgAcQMC0vQUdJDwLyby06FAvpCCFOKAR9niLwR5+zGED4Eig0+nbLdvsLu+XX0
S6dMMHnGFhxcBSIbTcE2A8W6NUtYkbeXA/TbwqjQu7QkA52g45Mi6JbRS/BEX6Rx/oulaXky7yi9
rGALxgM8XhekS+yahdsBSwASZlY5gl6Nz1JapSuBh6oMmtNfmtRXPT7CwUOgPPfezVVXXmCjKMZg
T5vD+SktgIxxgPKPfGyT0tU05NHYP04CZPkvD0YRp1r/iu3F+z9ZJpn/z+ABUMztCi7ZtoOF+NBL
Lgj5aP3ztFarEzWOipoC9aKHVAbkWynyTePAtpo5174hNLnVJPkEYnaIgXeAS68QwuW1cs+5Z0I/
lD8vc7hOTp/YJsQhaEb4WtpkD+oOouw4XbfTRxJu/hic/o9Qyy/z59zkb6/2y8T4NTR72oEowXnl
VS4+Ce2RxMCsEvAKqkIH+otSA4W7I9q5KogDyomaxMoCE9tJIAwR69AQ2nCefAHXSakamTQo/bY8
udu+RjtTeXPQngUhE352zzrrXLkr+u2FI/YY5OXpB5Qw5Nvi39ZE9ZoZD25oYmWXZWonFSCd8/s6
/kNQHLeHT5CE+0DKY3hf6g4hO6GLdWC3uE0IspOqO1ucnbEDsRQLOL636FUmVGIp1PbGq/3qmoQ8
+G/cW/wILT4poNlTcxfLm7TD/RDweWWR6PaRv+8Fi0HbBjwwtSi90L9PaHRBPVUqfxk//Yxf9DVr
KPw4Ir0aeX44FF2NaiA87U4Vuf3Kl4ds2rLNgJ190YGrKwsuIP+/KsdX8C6S0w/efrJY2IARgB29
8oRujE/PJnjclHaG/2ACeFOtZliuBzI9g0LfIcZL2oj5JO4DU6Sd2IO1mtW41k7t1+gIh/rG4fal
JudLYtjJHclnQnlvdAySdgDf8bDs5KcAMcbotXjIuSQQL9jBegLqq6nzFmNyivwJbAFzY389c3je
my7N74pmI0eCiJokyiVlmZUZ/vY+uixkNk024PlEmdBPzhhpN/8w1MtYU4kBQpzBp97e0D5Uxp8V
pjMvo1a956iMfiDalvsD5vxLguBurhW32bqGBdMXySvC93/YAKxb1BxX65oQ6VhD4E9ywOH51A7u
9CafZzVzoLPEcJWX3h6+emInPkf7Bhekqaxp3m//VuYpvzSM/kkS/llpuWLSmFy3W1KFIDDlUklG
gvg0qt6KAqFO1GLZsiBuWBVMIXXA7k5aK/s1FJQWVmt/rUKQZXF2Vc0vMX6Ueil5KV46K1yJRX99
bbF8lNvX3bK3TcnV5ruGLQJfzq9ee+vkLFm2HH24czyu6Vs9wCVXu5a33VQbtnuLJ/FN0+mO71dk
NYtHuGZMb9ndchUC/COVo0Q/9ZyWqM+pTsC64U4YTw2HGCvZ2Tx34kvpHmySQT262cBTgfVkcCC/
IvJlbahSbd+O4vtnsV2NIv7nAFs4Hd+OHx6/Aq4HU2a4/lZ8TjqHI/BQbUbiTqwuErjwLeBt3j/r
34wFEaDUCsuelJ9+kh/+1KPS+NVquf3tdgzQL0uvwi9f7OYJBAyY31QJkhNpP0TUMebidxfwIcVG
smGnC0fDVmrNlGKAkwTZNt7diNar22qf43XC2/WmdUh97FbMT0sua8+EZyioP0p9g8ydnCljHNtQ
lntcMynw5VJXxg2e0R2r60IwQFS0dH022Nh4vVAWbcf4xOtFzvGMBeA71MvC+6RrMg+iQL4mdLUM
z3H8TnfMsp5h/gh5LWDPSwNh3CLdYXfbUMsGh/VPlddc0HE2a16NC/k61arAp7O3zF6haXHN4QNm
/oSNiDbHj0Gvx25vifkuCg5sBXZf51iwZ7ZiSDp3nBcAhTh7e2EPJLNRCxo9HLdy6rn/b0+pOEF1
iXCDzU1RJvNqnVmYbISKYWl2/x8c8DkXH8t2UHwCXIFczkdnsbJdwIMQqhHZLrVueRGzl7hIjIvW
y3eyB17zRxIaUQ5DPlhtzM7B28+gNhZMKAvsoS17UZckpshMFspPPHEQAM5LKltTQsDngVNoAaPV
XJHO5U+AEcjrxnd/Qtv6qnamlw6M/k3aJkH+xJAwdbxhHOjNM7q4VrOItmdUBeAztQ39tzuzv6ZH
3OPEjc/O5POQdAYSalndKLH7coY6Z+2/TQMPdT/Y7nsdQ/2Svhug3HdyIkP2QsBQT/wCQWGIR7EC
jGDz70Hsv1XM7aGDZufqTNvKeW0EOYXScXXoRJSo3swFAx8Dd+Cd0xvthluSnOPAFxFLQYo94uvR
tu2Kb5xLBRtFQ5AEvWkXfZ2ToFm9+N67oLacFYCdMPhd+kuKkZwDVHb/mkoGAyAyADMgM+ng/NY7
Li7d1QdKu3Tvt+F8HD+aGtithl+0M8a65BvLZipAC+/4RaGkRUaATwWo2MNcP5Dv48RBFCrsuwRy
YMkI0tlt1OaVmlfz1midYapxW/TQH13y63sBrFJ8Br6yFY9PPzNkyW9vey8dx8uMLsSJg4mm8nWB
XToDL8XiHJcqk+up7xDDo6HSSCdA7nsvXXkABdB+PVGZTq31czXgPFAlmKPog609AVZxK+eQsYid
02M6imGp14KQ4tRl9jrVxXjRecTxH/cQqVSdAD5vZms9F7TwFuzGkquVHRjsbjwq7NtI+OvokgkH
O8tmr8qNU+tRoD/zNMYHkADAhf1ebTmXldxGjuI2Ab4Rl1gDlqH7RdxyHh8/eUxGJBSG4gpHo/99
4boVL9dQg+xFNidqdoYJppu/+3zQgLKEGmt0YtjiUtKs18FHD8wi/2XB3bufbZ9rBHT0Sr5WP+85
aKK2+16s/AQi1nijExZRoUM069Ls/c0MpksqqCMpsH2lvVAbRGhEHpZO3B5FrGS1/hWYylUEDQPV
+WNw0jOssG4GBFYqE7Y+rXV/ZxvERLdf55JFsqU3q27VMAijuQj1+8dqOScK+BjMcd0dONglBY91
hYP4KphfuN/G+QAy+54/qUaCJIwdo1OCjis7d0IsAopa74R3ctv/cIzsHHYju6WMJr7cZ2wzs1Ni
A2w0e6GhTmZwauAeRksF20ILUFmrABAGpu74+ANKN3lysFImHXdLM4Aof5xtxOvKRel9kqxuNSar
s57LgPtvFY+k+ICrgN3vy2zS5rZm0mjkLb8KEZK/kXkKZkADSxdGNf9ZrpfLcE4xNb2VTARG6m4q
PzUplme+FJAvfJP6h6/GGXukef2Tr0s7o/tLh9yHTM2CZuNA6fmUS0Qox1CdFg5vgEVnmiXqL0BQ
wH0W89ALWjymZH9MbNm6A5+ejfQe1AXHoMqryBuhjvQYP/CpeX6DjHx/3jm0GnqT0debF+uPiHNq
wAkFqtPbUTpUvOQI494II6yayJ99VddhBelKW65CowyBHx5tvPCNy2po5S07eeKLuZXqSjPR9y/k
HVg0gAddKU8i3ikge5GgqJC6Iog0yeFT2iUgY8NbWXW5SyNavhKvC8CzL6JKBuI5aeY2MposgtvI
0b7U7euHcFo25BSDTs4zayvjxmgu106olizl/RR04mdq8Cv/Nh2D+6+KJfYxVewyfpIC5zJo14Jv
WpriI50wi5BaanncnBLuC50TrHWnJXSlp8uRC4ZU+VDZffeH5zOIL2WsuZMolHxd+I731LdE8/7w
+wuzwlRSYJUSafDN8/APYVBOHzdlrWy7HzMXqcSIbEvrQ1ddaex86mBqiglusQEsjY1zldThmgGr
aKR0X6mtFWqsB46WotX1sQQveavmhqpLbel7vkJa82UdKZtGcqdchHBQj1uhieI99aCfF+U3/ga4
l+4+V6aPCOlXK1OrZKGkvs/HP/0oauWoWzvMi44l5lCckp3KIgbtHSNArj099vX9ixOWVETK6HWP
gxPV8PFsNGaV7nW/vQIDnGsbwaC9Q328iU+T8xa3iNaAXodjGPJTGHo5g0SQGwqH3p+KwvRpQImC
OTpTZ76eH1tfEzEcruAnXjmHzov7wObDa37XWxqE6tKqEK0gFNaMlZ8oaNu6zvW3fYcStV9jo4jQ
YriHPYeG3RBbo9XgrFbsGGX4dGw5rMDMJI5jzl7DN3b55KUJe5x2XjoI9qq5G4byP21HA/7tYo8z
fmngtM3v30p3EOjwscEPks3kwC9s+XFqX7gGXrnIyUUr6ywV508mZZ5HVjuKyeNgm66e6QT3TTvy
2rr9alaDRx6aJ57Dk4QBRrIA2BkziS6yG6zLN1eZbf5aXkSAtdG1RogqlX/EmSFlfWv8qSD85A6t
NWDogNir9YLqvyjLLSXBNGkPXZ5u2myRaOqfQxs2+x1Q8hGwlMImrIt5oPoBVDlReKR/hPptKS2J
959gAoCBMavoWSMfUnOyIgaA63/XiqTwKouQ7/8/xrtCPjVXePtbElXVGL7ZPHM5pbH4ygYNhawz
o175Q/kB3w9NJbcqKwQqj+qDhKlg7uRZkMDGmIuCNnKNcOMcwQKGunyWIcbjBm0kpOA04kZ9gE+r
xg8dmbCBrKN+/i8c3zEgk5yqZ4E//fKh6SC2i0hl14f7/3p7HYKlmk2zfARjnoWa4rKZkOU+3VjY
Ml+6IGctUjrUSRaXJAP0JpZ2Mrb1Aa0ECXceOlA100r4JvgD5pvxb5+U6ptfO5IQ6IoNHpM51Raf
OHABZTHynnubKkW3meEiVQ3o0WoV9PgyhDM9CI109knIdE4ob4udL6WDrXlXA7hEC3GuLy80Ruxt
W/5zMS6W1q7K+65WbWnxIPH8cuqXZrqKFehEaOfDkQlAoHU82ONaUHqi3Yrs2Pz89vzLN+k3ABMt
OTs7t756O8gN/udgJSDTQJJ02eIcTkNZP+lcIDMVtFTuPmwp47yuLpMEODiiQ9n6opCiSZ7d74qQ
D6kPm/X1TfNqgYkWVJU8MKzkGID6Ngz9kUo4fQA2HQGhnnLw3xzc7z7lBqH2bA/r7eOYHpwxxiCH
2uZqw6ugrl98HWwas2IsCy6iac7JFd76kh9o7xD4QwkDJDCBW98NjQeypLV6+5DtqGFOdPcVvRGI
Y49e0SzItmdveI5xNlOInrUoqs9QGsKgQ/6RddeOJH3DNrrabyd3b22tXVTLenRQalM4k5bngxYk
eClLdPGF+dqVEJNknnTzYim46Fcxg313eg15jO9txjqJsJ3e1jVE5dmcrRAq23vASqMzPYqtZI6H
9u7T2kpRM/tX7wekhxUXZ4VI1u+BGPtVxGqpkWEB8IAATUbovEsnXVYreVlzmob+b9C5GiLfIX8m
I2qnMe9giozEVj4qubs47ing7LFmr6/Z46e9eaCQ/S75fFuKSQ4GvGFqHZkzm5CkHwAjFztZELH0
BHZrt+f8WJDEXiUfvw3h0UYBuy54Vvf4Q7/cqUe4wjtk+uK3PQ8gKQ8lJHx684XpLktXpOy5axgD
zxzJ+JNQTFrlimrTNYKGhcFTiB8dpC/D3bDxn4qrFC+0wILShsUGKZIHdS6eYcEKogvf4Kpp8bHM
2NlMQCOkBMKg9DtcTVlspNYMKPnlnr/7+5DLuSaDzAT37jXr0YRmh+mS6EKynsynBpbDlIjrjP75
vW06JcqNbVGb9SKJbAJRuhJ0NAJV6MSiRcmQj+WnU7ukOYCklm7hf7AKAqr8KSe5A1iI0Ji0Dv3h
kws8CxMRPSjmgIgEpA7Zk9VDnHvYEUnuy3tjyTouSTCuOBTL1gVNLyC2RL1nPTKSk8ZqyEeDjcjJ
Ir/kqJ5DJfUgN+nHB1OPLl5NVC3qnlSHelRYVgIkHXj4kUl9z9YBxqjUoVbahnr2asaM4ec0/oEX
L6zpNrlVD1b6ZN/vyeIAlxzJbOMbjORT+lYLjGPT/1MFzUbqSgyHGnt9hq+lyntF9sO5uuhUNsa9
2jDZSzetMSSMZvjjzucVI3UWYWG0tYtmqq+83iAXMvrFkLfeIvHmKl9SOeJR9tWWzWB3D6l09qxl
BX3PXW6pG4cm3YbkdtxSAZa7nAJNcIT5kl+8aAdfoS9ywPmsM5Jd9XGy0XMXfrAhnmfGuhy1sKsB
6r6Cz4zMFzU16IHxt/JJ0K371yBmFevKYDjpoAEHtVgr8d+1pgeHL4fAe2LRpFkd10tT7TvZCGQ8
KlKOLWOt6SOzMIB3+8flFjMvWj/imi4tWpGQERjFn7B0p4S0IY9EEtoTCfXDsrhck4Ru/8EPAiyv
rZlC9nY0P5bex6C10cty5SuhsOikmmtzhC2WuNXGQf19DgUaI+9Il35ayHPr4Xp26tTOw17sIcT5
Rb2ojKMO++XLGMLL9aq9CPi5lOarAld8wnHUgXhWTZtM6Xrc3jk3u53zds7lCF24pzGj2cl8KBU5
+HlfS1ar6uB8fJKxkNYNhllP85fZHVRmhNO7O8B+bk35ztVoA14VnINYd1GSKFTgOKlgU5nNvbAx
h99a+ja4qJv+y/RAoHDh8SNQvJh0hk+F3xUq9PlLHjReVaNlx++XJra9ckjVZkfCZ7GdrfGjgyof
wUQKBZi/aMKSLDFWt7g6WCivupMi4qN03SDtEXfx1nWiwmDikJeBSCyGSwrO1b7sZ2ipRTyxR1X9
lCdy8lH3y8N2vhdHqSRaJAy8NvPxfIsp4OaCY6x/jj8muPqU9r3R7ltJ45Xg6MtvipKSwltVwCaz
0AyOeRpYCjyXTxPnFktjotgd0b2LKjYWzI6wmkHmZm5qVBJUAVoqQ5un1KHzIWu2fnJZ1f1i0Qqv
WH5qEz2wGCmQlejSjaudnxjLoPCMU/smhceB/OCkwiLLtLR36X/OYWzo6MgY36Kx0GIf8v6wPsQc
PUwZBAmXry6DNAT780dUZZXpM6u769ygDyDYS+Nl5bppuMBt2NdGGvlvjCfvu6iiviP5hx8RucqI
32B1vBbofcxdIAgeddNFqMuO3UWoDQSxDRlLnGW6XcXdCTSPeuLFh5Qjy7qUtQm/KotS00WYI+LA
YRyLHpjn6i4rEe236gWjV/OPJLyvyPCp0OFEk8j9XzlgNiYbUnDvjt77JRE3BsKzb54Xa9TUXdYY
tK8Jt5+EDZO9Bny/10zK7ojA9KNcXBiwZJ0PmyCkn38P+A9OJK2uLiUHsbbfneiM9lXzn9ErOGyo
ZbMpOjey+youC4oyYTqYBM8vBI7KFDM2O9ODbDebXxuTMzvDLSigvaOjloW2xxNJwdolZhh2DzX5
iQttZNugOOGuwljRQoIwE0ANKgnvSVetiiaryHJy3Am6xgqDAKrnuZm3DEbJ7G/ddXf5zdcOgPkx
zqMWmxw/jhrql+0cZZdHmpgylC3Rjl3E9wYAuwdhrpd4c1deIKsMujOlWWMDfwFPo2/C7Yz3v+qr
UCwnEgAYF2Umxhu/Q8rM6a0dIXq+a8CFAnHVYLvnDDDyZcUZoFs/fiVHVPTpIAns04uuCceImhtz
dO+cniDusn56Y8ZTSQnAKDazmWkQERhy4rsKT0VOvmbvf31blfSm5iDuEjnxG9dx6FD2xdpB6lrt
PljcYGEoQYMxU+7BNyEv36/Bkn6LmYxLZEJT7X7/3z3U238IO7nr2vgS2FvzcVqkUb55eQtZqdft
aoFjWDEi6qfSu3OO/YlXthpry0kAnCdFS0Gik1M2yzjHgzVZjkLcEF9tIOvkgX2l3/ZDkz5I0zlu
lr2YjLH6VGmiI2f3vc/fPOeMIplGJsiPdOJr9ZW1ojRC22MnemD7NPztrmtiSQ5w9B75am38t5hP
EEzeVOX8y483S2wop4UtbjaZUVqszMWztMp4kZk+twjdAHlpBwSCIXMC/4eH4RFmPDhKqyU3+bsS
2iSLTqM6esHFVHJT4r+hFqRxAgv0zMRh8RG0wkCrdy3da91zrRz8mPUDgFTxrRSWYxAjSg2h5R9y
J4lOZrW85t5BVrpe529UQyVdaKgcnttxwLZlDa10vKF2HfE+GVsoIaXJJOEZFz9G7XEybQxJaPVL
6kOifuikfCBj4+SHB0KRaGm6aqm4x9paDs34faypZAnZqMQ6yQGeeCIGKmOlMRweRnQ5LYoEPPoS
D3r49DsARMISm6svfTmBLeMGL1lGeKZPE3nj9UFbyuc43kt6Lp150goYpOh2BdafmmWTT9yRostR
2WwSK/yrgtJVYOVpxV/I+Pwd42YAouOUqLEQpFn26uLALrHsXRtNUMjGHt75gxP/dkclx0BRZI7x
dCyHk0THGBI49jxW0QzMbqo2gicYJB29Z0iipPux++OmxU+ZxRCDATeBftG8e00OAjUXpuAGuYrS
sAhqvflL0o/EADquXtW9odAzYxUAfFviYDqzKDGWtP6+nt/4JGkQd0ulN6Pir6qwu3dTWn+EGBaz
DPfb1NnHuXKxBl9kNuVPnykV67vG4vayzFVC69mnOgAPqgMghIIF06dTPK5xBH734k8WsxLiKFp5
emgE2FmfMw2KOU9Yd677pKdMA7Oc6QAozKVQHeeaujOJF7Md3uXKTR57HsbgUTGrxIEf34UkhnkJ
rBJ5t2oJIOkK0xDJ8PYSX+ie4gC/MFInlJXvTR+aBO03WH0rQMm2HpW30SXMWOzu+TGzn5GUaXTq
NuHqqKMgENWi4fMo2TqEa4tfeIropzxu0lusdMYoYHVwMqt4mcXrjVUbmAn4JVz2FEyezIOECj2O
HDp/krhM06LleBh1RfCf6o1J+b9d8YQ5uM6AOvJB5vYlN4hB4HylatI+bX7X6dlKchBaUQV5xe/X
ABZC2s7u3VEZMtqLDzeK0kfLNW5XbJB0I7Yp0PgOOd7+6XyRj4RmppIZPfelmjxnBAK1rMMcmLtg
45X+Fyk9MOvh6+Scqm4nAZdzzCc0SigLnClS8gvxAX1QYX8yX+1wmtx15OmvKhSImeRLJnuSLF8b
RGlthXP0VHqPL8knsfsA7Va+nrfrPTAomqoBTYDSDtSgXUw5kqYlcNlYuSU82rNhMMQoEhDt/nLi
0pf4c0xaJpD26SRYILxxLUXl9UYbHu1b1jYkEsd5jGPhyly2D6kGrlGRZqfP6s8jTWQGCxlCmX0j
R07nF0lyLYkrTu/ZWT/w2yuGEn2y9TTk2UOroJLc1Pi9JNTtcMVriqnkGDnxFvd946/fospmIWq5
WnxRctVmVXUWljpK88kfnsb2fXfpA6NZBMBqHrA7a1LJWtG4A2bPS3RJT5gM5PzuockotGRjjU90
He7Vm8YF10ESLITQpmb6hugH1A7zog2wPHC4hAQnH/bB4r+MqTdlMTiuBi1znqjrGvvRgsrQT0Cs
Ne6JD7tsfZyg3jjWbrQRc38kNyJo7UlNBW17IrGKtmQNZlH0TAAawm18gDeTjsSCZ3661KAGLFpW
mGuLhvdn9JVyDw7goYfioOAtVLB8w2pEUqZ1NVQJdgJE3BGGjB/+s6j2nxPMpCviOw6gPZrO9jSI
j4+vbe9CfHrHFrNm5P/p7qh2pHYcZD8Bce/D5PeQ6Pn6lPqKurePYB5r83lpAyMMii0nAnoqPREJ
HyHrSt6oBLVY4gKDcKCWv4PFi1VgXvesr3pDUsFl6ffBLjJPxt6VHBqZEIsXQMKqHE8gsMLc94Mr
uSP+8Gt3gwhESKnmBGwHWqLKiNZYzErvTqDG6PHD2bKbHe/w3F90jmuTrifIeQfyXB1fMiL8AtDn
K4qoW5GkUL0EeeM7Wj3QlOro/BfmmMGNRV9VtxyhqYxiuTqoXHvYZPE1jZsJjsU+Lbl/EepjOQtp
P1ZnQB1+3zkT3isJutevKfsfj8NB3uw3fZwM2y9/WzrWbPCDE6d3h0xGJEQn+JnFJmRsF49xa0LY
pUQYCLbYcqJ0Hc00+VYQ/4+NVfIzPh8RupwCI9rG6xPVFztKmnMlZnHtsJOyIzqa3rzDmB3PCMjS
N4OAVujIdFgM4umstLXCDCIKmFb3Z4z3TBV3ZGimOg8/lyH4PTYd5qmTaYhSlin3scb3GGnnp9VF
dzCepfFU+f0mCFmb+z1ayjsFpYT5jvniI1HoMBieVRpSdfBTxmSmhetp77+9HleFqmzSly4fsDk+
Me20Dl9iYO1Mkcih0MZqpqmx9YKBahokVQVR7pU5ayXw62UaBgf3f66TgUdSP2tps1i+rxOzDdwv
nRJ66uDU6cHRUZtctN4aareTIAgQF3EZnT3OTkDwgMn79RFtvvclNylRQm188jJg7lmtzCQHMQGt
BVvT2eV6f5g1T35H2uKX4c7anTvaOSEAkD+Bm89HOKSIocBsiLTnKxZpVxvDix56lFFSZClyHQyx
VGjH4IldmVErD7/J2F8V5YZR9d5lbC5cnehaDnBk8w/kNR0Qle9jyXoJtPEzCERZFDaEYoumilxJ
eG13Fw/3Uh/Gd4JH4Pe/GUxgQ2+eInPE6eR8gEllnHjFgsbYQ4XghKagiiPWMLQALCR3OMCXvbPS
N8XQacLxAE+TV/vLPCsCugMCkAJSgy49eR3jlViKumJ0MKtcYGbV2scIAmjhubmIfEpMVaEjB//g
RkRkFndFA9h0Gt1lghIoPDkskKF0GQAIPjp/4arkKtyn795Rv3E7SUHPQOz4tfvu2kouqs85yzDl
hU6RP7ndWrSg02F0LYIhl6q8CmwXu5lH0vCFkbVJRzCDIoBcVqjSTBXwErlcol5PjScpW97ueGyh
VVxEoc8DFWHTW+TjrzmIPZz9uKPY5qbTnLNzr9xf4lKADbb1iLt2tjf78TVPb4XitbZI0PgXdtT8
IUUWhqWTBrDpOq0udaPVeyTB7hY6gvRON1GILer9eC3MeybHjy6ZUNr0wuL2ULDRyECdi58XXPnC
0tstt8Df+UfyyKrL2ejkUyq+GwuFxVA5mRQYEQhZQgb5RKuPtSDkFn7tpCakDk48RKQvDQWUmIP9
MiJQI1Zy9ZDRQO5QGm0M9viyUCyLu11b+hYqTd9EY+Uea3JVhBT29jb9cMcGpByxN20qS1FQfJPl
ru7MwCrSKbUxTTQKso7CCsfiMjPthJ6cbxOHFaPC3IpCwlMI4uzjzi3kkmj5otJjCin1S8XEuYXM
XsFD0xAT2RINglUAFx9VuMjMW2N89MqGwZLd1sdepNl7fee0FDZAOjNk3rjvcy0LrNgfPIRDiC3H
CbPBLdSLKBtZCbkByUj/EHyOEry/k3u2NCWqYrvp9A5NWPUsy+8zXpM/ysN5dZin5xcc50fJaVk3
YOOTCxejP7awFqki8eoFVpHnh5UZPHE9w25QntXO6fX40EuCBjBnocbhHaLkv0X8a33KZSa52jlx
uG2zTzE1zHRk1H6HXI731dM+bc6P/mSCK4QN0GOrz7JyX8J27HcqGEs5UMeO29VklY6uAF6Lo3Qk
lBpbnPk+5nN5XlS8srlzqpVG/7nJ3oiTZ8QITFD0d+ne3I9WptBjoY4OUEsoc/uMim6rPaNbf1sj
syQc9TSrRV9GqN7uv+l8r3EYWNgg2IWCnaI3kbDKN1M0XYG/vCveE6qKMX2j+K0p6R1fHC54466Z
vis5rk0XacqJym/9aMuANWcB5GNOQYaLEHMya7Iv/tSNOmrJPAmD4Cv6tR+QI86s0UZ97MsSEM4q
23FWcG9l3fK0iSQw1jWxlD6nC9YLPik8bSQBKObCg2wp3PGn/7kr3UpZG5qGxJiNLxdKXuToytFg
5nBgdE8HtaJ8dzoTtzWdwRXRtGWzNrhC9TTAPFa5fQFUGZFoJ0C9UwkZDxrnAZHVwV8fzpVmiwxM
41pmL2K4RrQGaf9McA1meCf4M9BXSxB1XnYlLrDNpJU9LwsLDanJWxdN7eS3O+PUoWgQr8Bne1nT
S1bYYkciPzANvfO/7s2dvtW6xdYzL/r0k/gIhpVVsH1SDuHByp45xj4UZ4EXu7skfY3ny0lNbhTa
a1D917U6K9MUW/bnrDz1ha82rfowwBvL7WczZDVy+cSrilYZX3Suw/7g9W8bGngwW58n7wMT0FKT
RSkWI/ylCxRlSBEL/KazzwAe7Q0pzWLOFf79ZyIiHA3kMFi3QNBo0QoR9H1rIwYUlkXOzy6FYQGS
VpdjAtS/sBIzRF9vavLSmErDEltpOxqJbdquDM9WSt/VvmCAwwjk8MRyheIUxSGKCvPnAp85RqjM
cgXp6VDyFQM+lm8XYtq1bgOWlGS6EUsAycrWQzeqf0Zsmx4WOzGaicaKEcMKmO+A7HNOFB9QvoHS
R+9LwHAp1V5fE/+4j0bZdKZlEqdIpxQneO8QOc/KMM4Ll4G8BdlYUbfHGjpqqrQao7qRmueDqHrj
5gjzn2oQHQTPfqX4pnh1V2Hsxstzso0O1IaVK9PfxLMrY6F7dUP9/iaDroeX0R7oTsn7yvKIo6K3
Hqcd/lqys4X0ob5K7mcu6kkiDLaMjmD7oUyULaL5B1GzA38Va8pjiXbe5zRvaZWS2hiOZvZW8BY1
uhWb/0ktubN3dGrVGGW3KejUcEORGjNx7LHPlFfoMxv08wMJ8Gzb9LG54Ct0GN3cIGgFupXJMDoc
+j0prcpqF8ZYfzwoNkR+XIg2sbhnD1rdOyA7MZ5SKc1SGtnXd5jGR4FtudlOY1/zaBr/RHlAVybn
KE+QHQhb3yMbMrv1i6Nw1bOgBt7fxIzwnWIEopzwiE7iojDsDP90sIGkSQljbmUo3Y/7qvkXXNJz
KBqPFm/syjDbrm7getsYn+u5bgTnR2rK9zaWpT93K55JjFxYNimy3VHq5jG2iQ6Jeb1EcyE1ASNK
z8PH2z+IFBsCGU/yShE/eUJK1yhpP4NvLK99Am8q7t9n5fHI2Rr8V9lVUcEuue0I9rRVmIIkvg5q
X3vIDqWYq5xbjb5erAcxAARdoEJpYWHDMyld94ArWyKzaq62G9pyl/6Uzn/cxMIwM6cZ91QEyfka
J9tNNrWy5JaUXR9CvsmmjECsey/oFxrqpKk4y00O0YsVH+BnlZApty7AQeh98jrHHjGiHJ4vzakR
cSmKKQmhZN1+OetEZ6hS5v4TxflsXzaYScMZ0firOtsxdSN2VD4Itg3NVBuq8guZT/NfnsnKRohp
8EQmhTQvt4LrxlM/l0T/3GdTihhXwLHw4l79x9szYwzeaNbPEqarcTb+o8zjs6KHFmukHGOQlwdC
Qxc9k8+A0H8+yNojGaSKunScKWmaG029a1Lc4U80Py8FaOV1JYywztAD+DY6bOOyjCPAz6t3kBuT
JVrRlaPIf2XE5kXutpcvmUGZi3XsiW9UBfmbpceI2U4ZRDBi6+3Ng3gXzw9w+tfZp+p0nbeh1pRz
binS1AEYSTpiHoTdul1xZDvcROZNnUmOtyr/waF4KWjp+rlEOqRV8R7Lw582Ha5fH++TQetfh/vy
x7BNjAUtaFbrCgZm7URg7v0bdBj8zBTh5B1th9ZIP2CLR88X/3oof/fO8F/gJyYrMaAsTRkNf1Rm
4XDds5DZVbAFVQ3b761QNgovnYFsDkJcLvLnMKqb1nO400Dk2NbPHblWh3j2XbhGnoxyILlNU1W+
PeG+jt6w+H0WmGbHDOyEeaUTZjOL6hxanZcsvxkQ2Qdr82feO2Tf0JGsmC36V0gHHBEPhfdBz1JI
Zqpf+d1BNFmQj6nnz+Gx2g8uLz1BK6pqLZjWwgI7gaTEoqdCuvsbBbZpPm8Bt2esUpMRKQJTdA+Z
xlZYAr4W03BVpMQDdNJ5YkbHhGHeFSqqGi6LcJBWyY3YpDH8iCmR37hs117r6SnG6JQ5yB6sNagU
zRwtYy410dvHYrhx86Nf0VpGXA0I4ZkWmplOAw23nrMWWxPDcv5tB+DymYwylbpk8sRt3BZlhXKf
kwujAbi/F6LTG4DOgQvJxv4kWTbiPDJA4TCjzGepjhMCQWUpbHge5p/+5ZuDFHOW5LftcDBKhFJK
X0D2lpJCe+HvAmELqAJJM6bWyFpZEhzOZRZA279VH9pLxFUpEjTXZyILDnFzsGUmRb9puRHBbwok
mNBuwGWza/7t/XnLizH8Dg8jRU+fLtRwCmD2udpwd4ZcX1eJPqYMqGvHlie3gtQfk5OgFBi7Fh6f
ZK89IPBcTChgToxZBvqY3R6pbV5gllOaMlPllkh1H+CfMW9CyIq6+VvEZVjQ5J6FPzsQgLn+S9z6
nVKzU0VAic+Gbhj2sDq5jz+rnx8LJ9JZ1v7cmq5TJZhNtTlBxSfD93GBgbbiUMfyFZXHMVBD5ZDR
5oSKAOg4vPGmyYzOxP2ux47TrIUkQYrWKiXR4+AGEh8IEc+mfEmtnCYbHMRR7PzfwVGH1h/6rQHN
GkLd7XUI9C7mp7NlQM3Z9E6KDlXBI9rx6Dx01qge4xD4jLYjzrtsX+JKTiI/wQRS75bdO5MBBpAr
F7mgcNZN7ZrcdeNJRwXZ3MJIZUWCRvnt9YN++hOqA2JiFwLjMt2/ZZXUaP59PK0rTAIk/Q+moMuG
JVHu7v6LceysV0Bv+hqcSAdGRygiiB0Gx+n+BbfYMm7F1hbTI+960bQk+z9sUs6N7PVcoaeY/7Iv
TusprxOdI6Yg0cm4ZkKfq0c/e3SzRIaR+b86zJctM89e+vSeWCGQ8J9TGN62+UB7r2TtnemxjOhe
gF+FYKVOcFn6ixOw7RRiSarkNrw+n0LVcKOyxgnOPvmcN5wPrfn4FXzoh3jdqy48pEfFWMGJR07O
PAGiOXvoBhTIplHjHaDR00+RV2RtVAqlKwbtF+Z8+ShbPzB1nIYxa9Roi85ew7m7OB5XTGPdCS/7
iZR2wHzxEYfg+Qty2Ngvtl61+ZHlhMjXpzISZzz1BsgzQy5Tr8Smy+fmHiwJFzbj4gWeVOTR0uOE
9HThPxNBe7sFlMqM26MJwUQFU54KNnmNH58Vs9TD4Fli4PiPKLE9LC1+zbNn7yyXKLO43mk8Nk7s
VhACO6AMDP48JVWDku6mAE6WLzKZ+pp1+Ottw5vaXqZpjWeQsb1hKgfTvbn27L8B/oTFzq1oNNs7
DTQAvVEc3/pVteR100nPgSG1JPYPPEGwO2wLmcgu7NABeS+gA+/KrWd3jAblTjprfp24/IfgVGsr
1dz0omcSivO3N0H3N39A9+yXs+qgaazMoavh2u5piJyvS4AKbPFDb5RGBgDpY2Et4m5RvxbGrqNu
DcZVIugASF4nuoCGlcf+RK3k/G6LC92riCGYBLjinvXT82fLx4xOz1eg2Vfh1fVQ4/gDC7e8giSj
l02fa2ll9DiMSVJoWas2KcZvF0+lnm4AuB+8+E+gvNp7gPbMpp5RJdHzTmt6aIJJEGnBofecBMJ5
txicIvzLuIfx/kK4ypUMScj9OwaTuo5+gH/ifwsEWxdK354HcqmLDe54kYlut2gDlws3zuvRERA0
FZyHyBrcBr1Df4wzNysrrcvJygf7ogrU480dosFwDppqefI9P4ntzYuKkgEuTrCfGZG1SY3uCpYv
eMmurPT9PttY/3Z4jy3pc7KDs0yWU8LyyIlJ7kQfiIG70qRgCGc39syEbMvcNfq+m1FKxRKk6zOj
nAr3dj7y9Y41bdZEYzJ38bqIE6eMMCzaUedV5RTPjAcsPSj/zxkcOEno0pCz3zrFfHhznfzj20ha
jJLY1wsYkgpKGvSMt3ti0gQqBvxjJLWTWsM2e0MX24T3tKYC82BxJ/AB9tjXoxFddcTpcOCar322
426brZZbmlrcOozc1cmtu8HkrPwwEnetA2IKHuf1Al4qgp6fXc8VpgM0DCb0cEPb3iJxMbAGh+GH
aPiTsTioH8Q5q2rhRnEe7Tvvoj/jISYtd704iPjAkhWZQYx7BsfmhYSc7uuYlPmaOe9or+PRxd2p
TV2WcnbAoNjAl+vOCmrrqQI8YFOmbSB2vEQdwevfm2quug02pAoe5KFLHwggCH1iqGFxf+u3j1jf
e2paTC9VxYRPYwmC4noxI/NlmHYnU4sSF5vOXSAlz3gEHs8GtCTOdVbVotpmVDWieH13+/JYWx+R
yzyA7dpThlH2PPoJo1MIKfCrhBmdYjBTXlcngEoTyGodrEttdeB8dCE6nZXI+6IDtuzeVPLMhAKR
i3PmyJSs8eZ17/1fsWV3pZu7c08USP8JfZO4t8iY95jOru+1QAMFjbQmRvIA+3y+3xnU/NIaBUWX
mrr/QhW+C5ZvS9+l2s//btAFOrxNl/CgqUbrB1fACB+HKzTfpQka8AwJwHi2YR4Vq3wjpUPxs9hW
9sW9TM7QsUhw9hzKd/1TwbOANW7SJdlkPE2096iRTptGnkOl2OznmCx9BI+EjsNXciZPs6sKRG8Y
7ohbj62BZekR5Wh+rIFQrFV30BFiaayMqc21aku9xmypqek+NlhW3f9oljRi0kxv7zDIayKqGiJi
gEC4Yt2mRaCydBSWBvlMXxLxD0Nhqr1sA5A71UvShP/crosYkFArH+pE8Rs86T5qgvOk0GljFlIc
XDGIRtVH45oIlWjyqTEsYyYEERF6v55pnLCFFacDJFqbyPo4d5A8QCgOm6tbjQ5Z3QT7YbLGPBi6
O3Xamg001rkkHfQB5ch5vFQ059dPDIM1Atr9O8/BQsOX1CUlcZzJ45O4JpW/illXa99V+J3tOmbz
PXB/E4L87ESR9/ae1n5ZHro3SJPnvGEDIhSfynARV+z/B69JMXWTdfMnAXZcgk6rnkUWJdpC7Dm9
+4RKv5Na0ENJohPaD1vRd5pIAX55beqsvBBIP8hxpKqjv0hJ5S/9mDrc2I/2KmjY61oOMgvYb2rO
Kvs7JjYOSJyN5shibrQ4XRr5rIzQDDitMtxZ/aTO3Gtdm73kimQweiPJJ8X7OGOvCk6DR1/WGyIE
MAxHgJC4ccGc8dl9umsmSIZS6xdi+AP/p2N0wDrJ8WMokeTj+Ccp++btHiMvHU4XCd/lhaOWM3a4
eXkSoQigZ2lp1wzDHnhR/MY4YMjsA27nNzFue+eO+ySeoAWrWFazZfO941yUiclWvRVCNCYjT2Zj
CCd/hq9mufrY9HR+m+EGdfVZa8EnhmqP1ACZjIkDrhnQxmEqL3ji3gYoLAMXfUS+6fyaYEvlNNrM
2lXTArJxwVVn3ZeV4dDZu90wV3xxp1sRHhtzlAK5npLCEJmjIjVJIM09199jZlxcBmXIRErzyyGL
7kVjvhCbGbrSTmhdaZd6M7fORgElxsz8AsoaO/1scjaqyl5JXV/psl91ij/nhDjEvl0pqGsuFXDs
bLam3NFgbqXol7TVzuaDRbvpVHF+WF/GKl3vwhSglZFKiW7QITPY5bNqeYaa0jfgSOW6EDSnEG0Y
tSPsF65FuF2OB1h+I1ukMnm6EtiAVA+dcHZQURzB04/hO4s0EUC18VTyZ4KDmbxO9LH3G0GoF3B9
hlILZmCpp3XPL537OwkQ9nayUcD2Yodi2Huf9AbTtHnCSdzm8cC4w7mUuP8ZfeCO9aCsl3V9lRak
qAN2rFGz8I9os1vVNQuwkn0WXlFEtSeb1H6Nvv9g8BudsJ4CzLaeP6kadRIaZ9ob5IwrUy5KGaiZ
fy904THNtC8hxuP1n7iYjVWkmppPz/ZTSXVhLwnQdhyf88h81eD5q6ei09bJOkNrZ9iVBNPTYLLA
BpBjHkizbT2JotRPNnk21TFEXbIXVch1VTVq2suf9VPuT07nsXYybXonEMLhpAORKIzukc0FkB+S
BPyUG2pHwLH6wEaM7wwUdVQXNw5wA+A6j37UAZSYFzYwMIIizzyaeKFnCDSzCosbF6a/GTWnUAlQ
81UB4p0WlHyhqApCkBiNL22cdMwMPW+3jBc2JCDLnH+Noob77zuvkvpkjMfQxUC0xxb4472jcnMy
lYG+CSy/6+YV/55OXro3c/lmHGV4k1gX3dMbyUj3bFQsPhDBFTBhJtr+rBb939irG5l4cSSpBlPC
xow0KppClgAsLnBm7cUXFMIfubTypEzgos1X7jHdFKt5irQKDJbp4scFxrMFu4OqcofKIhNQkpBf
6KhVnGQzFXE1leB4yLdYq7MLp01s7subzfe/y2SPfpK77aHjaJFSwnIueGz/EmUPCZHtcgu0IBLU
2Y73HfCcIVVDQtpD1DdGZnChLbe/cBY92Cs4kVimAgfo1pxhX0B2O3ZWwgzXHyxWVtzSkP4XKDJm
9eZ8TiT41QL0cC9qqZ6Xvu5NToUoWVg7Nb/qOGiRAEVsA3tRYwcX0pcYEForCyOAmqB7YnXpF3+F
JY29l7S4U7wGCQrpbchEz+vL54oge+mHyOwBWNNsjsnkzc/tK9vDpJtq5u1piZxCJqtuZ8GZ6fXO
pNNedtQWiEQcTKvgu9AqmQiqkus6Rp3ue7IKO0pVfQsqY8qS/ipCTWhBQUWqRfif0PdYKrXSQWW8
0zyJASoVTXlELo096yNZQzkAjjx1dr5CYZnqddsKYhIiEVosEyvzNCXp8jTK/6/k8mFtSTyMViX/
zIrifkXqPQhC4ZFMj+ZVJXhwzt1101285TVvxW+YHulMDnkCRZyM3kTNSOiluTdslPtXyBkCxXq1
z39jAbyJwH7gpwwRdVZ5nJuIy4TPWyiJcJyPYzWJs1BUuWXJU69k0aR5wCTXySTCOKQC3j9pv05G
He3ZDR8WN5insWBXH8Ty6DRwodaZsL0SPihlNAcXbOTixzj6QIvqpJLBglHBBiEjcieSZsX6x29y
C/MXYhhkp+sIkLfeTVotgPno0cqbpXkDDTqGX6WFZ5Kut6r/wgKGz3doS9Jo4dcdjokbcVqXtfLN
4S0F7jM9x/llQLcuZR0/KPWk0q8IKXRAuixbMy2k53nfKqDHLsrzO/hvEH2h761cluoVn2byAWnP
2hT60fLTPHDq67RdQ7nYf37ldUuJ+kA6df/amBrKlgWm7oleX4/sS381tWu9p0MbizQe21hmUkxQ
HFONRidAStulSvc57O8OXJQf5amro8KiLH8xrGLENiR+yYkhiWk4tugYM7laZATQPs/jTsWexQQP
Qqsc9XnI/A/xI2DpuYsrL0yYw72cpuOjeByrpkD9Pzveu2itL87d1xwBr6Q/TDrglD9zAIibMI6W
XT2KU22yNcfUWnQcvH5o08GKqoNip7DJCZ+ZXRxBJmoxMJEGwfLp0KAaJjuoAXJljwC8IjXavqK9
WwJvbXd998bUfyPGpRJcAepge7/ozAOf2+054fpJ3CMFgivgNakQmprNNyyzOjKjfPGPPejFWRJ6
Q6Y4ZaMh4LhvTEvbdZriy6AL+2/ofAeyneDFHOz1+D1akgKGV5J9+zAZqXvGsJ3nXWxDOYhu4+Vo
IDhRnAnxKt1qd5Y7bgZaVvFJlzygA+JUwMmvShUviv0CUpMnIgWig4dAVbWf0Lc1jd5ms+KuTBIP
cqcJH1fpVRlg+0k2az8LYRCXoLJMX52rO1BrIbEiXSm7qAyY6nU4N/GBiOph6r/OsEd34abLvvIR
MbsSu3y3zVytV+ogvnmXdL8teRFneO0shKlqI+U4o8ZY5FoeWk9pIXBRci+8/xvOgMpNsACRMPRM
Z6MxMrxVuOvTYsxdN4yzNZCnJysx6OkaSkl//yi4MPjkae+/TACYWu6lIjJgcE8JCfiDOLBBQiNi
cbGtSXY/dSt9FWTQStC2LVup81ezZ93qOjluLCivMMRJuickwHDN9VGDQX9fuJBhjOY8hNDSWS0l
pMr/IfIvEYYKux3B+nWrYrLZVt79jjjjYn1jG487T5NpBDQeEkfOrEsjbz4rZCdm411WTaGKoOTS
1yO2WiJ2scIXMsIg6ArsWXyNnTE8O/h2ZaOWPWfCi/9DIlLdmT1BW/l6PBPAzV4sI7fNEYQSShON
wC5NUH6THwGwwPuFWF/W7YzY7rGmMppnzNmdnR3vLwww2CaaRYzRV/HoVYn09OXUReyGp3yfxppB
FUYKR5EQ53ODpgPvKTshwkFcbqml11mNaNIKRoWvXa1nmpmSX/MRe3YRlNBSQCGtPy2352eFQcA0
DfLiqJ42Gcy57+Yi5O0TYNCABQ3a7HTly178tFXU2Y3dRjvqMDAhM+QUoBCVCUoD9/a4QpPJWJta
HysieimAp+m4tdzcE+aUmpgLT3Yfhpk/YOaby9akfJvChvcbmkdIeXGOMWHMpb/8x7s2QwePHlNu
8+PBwIC3sWw9JxBolQiPpPTONFKtvUa5MTNri4Thh6/fKP3VNEUzoGltMBEZjJGKBfxtcFmhEdkE
tlhY9O+ewp3BHSJmIJjgnbiG5rJeguMRwCOcGIRDJWHuxez9opKSbfAQtUR59JTxjloNqC7FJZUr
qA21/zwQfDKAQGRXHBV/5Hk1OtlOXPWwcjBVKgoZG8hE01aBJLYAXrnRzuRnZ7EjTxvk1qBPNq+9
BTus/Cs2dEQJHIUa8PNmUwLNFKbPOYFdO3Hl4h0XVf9hZKyZE/g40MLD3OKrtaI6N5BVrUeL+tjz
xFNfRGCfsh7ufN4dwAyhXU/3zwftg7KYQxCB6fOz7d54K7bJxzJig7FHXjRq0eE+Be3z+l+69Io6
E3aRmZ5zD5w8C+bZXb09KMNDnzrd1tHIO8CuQ/R9OFMBBj1AsLWe17DR9gZIBZ0HnETVrXog6ONs
2FyTyX5FAwmUy7DnCqmUHAC+otuY7a9TY1mQKrhEOPJAQP34LFviMpiosXgdzLtuWXKzGWFz64/e
VylC2a7I/2VedzwCEtcVec4YHHvNNephIIb6Vh4wwQX+reONnNG4mP887dI3jjcxJF/7XeYSK0ia
BBwgda8MpeGeEWz++M+NIhNXgHLNo8MqOVteweH6km+WWsXaLg9SpCteUTotICUymnnlltiZrCfw
ZGN419IYejQRtH0+Wc/Cnq+UkGOr6jV1UnMafyew9CeNARu91zgfyV34MYTetR5bpUvHIEyOtPqM
WFqWCmXA7afxetwXmhaIKNJ+RHTPMeaGMjHFI312def2nGzmBdBX1YgqbffS/sbRH2OQMVC2dJ9P
zJzi6AKxLINaKSwb2lchnTlKODKiL5AkCJ5UfwR/e1Wzj85CQQk9jRLLQ9xqJ2WJrTz+yFBWOcTO
VM9z4ZNZ5cTvM2nfFpuvxzQpaN3UL1SmwMgfYYLjHfcjz87dPQFRCacQg5v/IE6L5dgf12/dfwaW
woqnL2tw3ayds5gltXqsA+MyRwVZ7ha7zD8vGNdlvOEW9NZVXbTT6VkgCNOL8Rwa8iHroD9ivcW3
t5EMxxkAsVRlp3D+MEP365Q+qyoLlkFFR5VTLYcEwnx64GRyCSAlkW3euG4h72EaZ9SxngQZDS9s
CLlWNmiZ1vTAr2mPOVv8FENwhs6fbWVY3y6xONVypRt9/oHmJj0FAtIYCVmVPGj3L/SnhZHDRD2C
qDZO/rzXrPLZPFBM2yA4qoxdk4yizFOKlyFfwhq6hAZuT93pcZfy2DrooxZpUXmv7RxXkKLCp9y6
e6/9aJD4jmUn3aJeiO/OERkKpRAioQLVumXPTBNCDRzMptGJVqh4sbOCPThj2WVA3zY+qS4FOPGQ
+2WZbm43Yv38ofVF5xaGybQJzBSHdPWmwDIB7kKiLqSejt0SWA0ceGkN7/eBxNLZc6s0tlFF3aGJ
hhjjZWDEpmTdvk2lLsf/r0Tdkm9v6paFx8MhI96duzLuFrlE3TTPEcCa0d8HJ08HGLLQo3hao1eo
IXvHsda3bYOF1/3Z8jwKMEQwuSvpciY87SQA1L+OBz//ZVmGQHLzVehNJWlekQHXMCwRF1xw1lC1
zRZiv+rxVeO8kPWD6L/2WhSVXDQHA9r+1PoVQTqDBmXuBvB0HyEd+XEIy0T4F9xh6J1nIGTRqIQc
g3Z8ufeIPBP1apapvCIK9xb7oHniVAGBastO4LYIboJNvzOL+37ehxu5v/4YjSc/2e/UIkA9N7tc
8c3E3onuHxIiTdc9rogJwpGYFRd/hUzqQjKwS52e1D/SBRPQ0wHI5frOSMuJQGF7+ZTZOAWPqRD1
IH4vsTHxk849KLOgnalJ+uJ0V+Z6t5ldRm0/oVASxWl/JdrpL1f7Myg0Gb9C8OR/ECbTzJbNAVXP
B94sMujtd9uckDYuBI7rpq4Xum29zLpmb9JZvUDhzAOgZWwDLjdNKObzfELZnJLSCb5xtBBH/tO7
ycHbTly8MW5grtRE+/fLQ6sXwF66lI46QTxdPlmwP2kZn9cHf5vwsb0KbUsIaPUct1oHjMEZyXKn
Dt/owPHmdA14IV9nWKpnDUc4ldsNOy1E1XsqGYOdso9hAP3GVOT9xjasUPmt+rrA8fBluuFeISCG
a+obVz/seC8xExiLf9JzmOxUT9sLGib7PUb2iWM8Qqauz/V14t/s28tTaj82tVQDGlGgXCJiSCTR
iyxAopmoYL+HdORSqRlntdMPgKrD341sFIAmAMul7HAMMgAch/oXlNcMQxVGRur5NEYAt09sm9t9
I35FE1MrGYwXcb+ZZZ8XNyiZmHvRKM3WDpQDdf50xnd2E1JmInaPLgHnbY9rM1XQZODCT+wSYUN4
n9UdifJZbBjPQcJZh2CK4TqhEi+5bU5ON+tXGDDCNb9gQCmc1NstvlMC6E9nuNegF15kp5wwlKv4
ulKUIJ4hIoKBFkO67f17ZmB09YZHwho+9KJqFQBcsFEXtweQGqjredHIUXCARQ/lxrO5mknUwzVX
0fkJufkvuV0TEvLSkp8zk1jChhrrICT4cK8CNI/ck6MEZ+sgvpuSTymob9mwI6rh+leoBmGl797f
acU7auJhyqCMJlZ2FyZ9xIRm2O0IKapLmhVh2+GckcwnaL/rKOEAXmq7Ibbs+N3IP6drx2RGcjfu
UtB0FGUuyUd7hgJkqTLXsBXpEmDjnQIUxDaRKxNlVQnZiaItQxYP98KJekVdjB2YG5XGj3TEyo0+
1ExTCOs6dlXGPiZamziUfvGcb37H4RiGPXZDBNnRHRpoSi669wjPF13GqxMwiJv/EqeMrOMLZD6u
rhurdIn0mHDoSJ+rJ0IDoyv9d70wi+Er7iq+d5041TDcGX2zSyTOaV9M1qvEiNxWKwjluc8RYABP
gyF5qqmSPUVOj1Xzx9KxwD2UlQUssQP6YYmykipCpBaBVphHMnyGkymx2j32c0xLilMNL1EOeLtZ
kn58VDoTMg7yq2wXhBVhzl47p3vtLi/S1XFe3C29UrcHEYLeSMLH6SZY8KgKETO5WjjLVThna4rS
Y/uDUhtosZoMW8PLY/R1FzpGNvFYF4xEfCILNNOqStINNrKx4NqCbNc/z9J3/qQ8+WbYfqaXnrIV
D93pEs/DZFNRfDo6pqDnsHCLuILa/2txOxrE7FsudFXf0EyTaDVmVGmMcnJviMiekiMY6Dw8xQCP
/9JKnB+29huAGQpCfBW/wNcp4mI9jQB4HS/Ft8IHw5KZIbIX6LaAeyENFYvPiA722I+05cUl3Vrg
UunegZkTrUVmYxXV6cWmP5NXZog9yTM7/QB32yqDR0CqSqMFk/4ZuTpp+FR3GyFhKraRLaaOi+Ev
g22SAwxRAxPMyrRFI2uK2HlCtSLiNQtU+4KCB0ztu5sucB98Av39xTnOKZQ1306zCfcOwi0zy6rK
x7GBzl8rVeOCwdxGhuOdp9Yzp8MYOTy3FJfzZw9362mZ0/7Np604yaTBqLfTF5deoM6Tr3zblDx4
pjrn63GvaEaLITavbvQxsfNCnaf0C/Qa/AvxFoIcAEyK/Xy+VCLSHa6XUu8u/xQO+DSTHSFDRvI4
QLIoQLbwhUWOU2yUruNBPLcvQETIMQ3aHy53UFDD3K7YrQ/gCkB0e8FibBQTeE8zuJ99Dizocljc
RJgB0j4yXoIHboM5bPYM3RnQGM5NGzTSlfIncjT8q2i4sdF6S4VG+7EQpFV93XC8eZ/C2SBtki/W
WFnDTkUIwp/GeGRbVDbhmDuUqthNacogBeIOH9VmvBmL2H7h7YDAqZR6E/hJvkUgJ/9Seolibo6q
ukP9aZZrAvUUIA5asg+W7CdMEZjE1zO0LyI6MrJv8zAbEjxtYF1mmSn/j63ct1oJlLYRdodj4u17
CW0v5AHenH4qyNXiGiZhzYKHIExL9pV4D0Gxr0sXUOF9lD6fVCd1Ql3uJmN3bqQSOYfQJh9FSVeL
qQ9cSozZSbOEDwsnA46Pw+a6J5nrposTtIGktw5SZhiwH0JnxPe8zMvLbGDnaa48CqcCqUOWqNJy
nJCsO/93j0K1Zwdg/zB9Jjj3tgfsUsmyC0vQz1KtvFzJ34dQP6YT7PCOxj+x+UEwNdsXtgCLwBeW
oIAHTbspXchBZWHZdSRnualPESAjLy2NW2DS7EeLWhoVWylZAuE2Do5TAl2A6dFt5g4mxbWik5az
Jqfi5Q8hP3Xzc840FO4IUHmmDOYwH8SaC1ZGij2vf/P7tb22UFRNwFu1y97/UnEGYVMCU9KZ2L6u
8GyywXvUcio0fbQ7v2/4DgV7FWU3G1v+miDwg6MdOOfnfglDxKx6WK6oMwWEGHlxQEOZUTcYyOMH
oABQAgiICjIkqSsZBbNjNEEEdAUUP6ByoWf5zy9YMhArSn518KdNgdNf7d/9a/L+j78uaM3qkdb3
4vNeQ3N7dTQMbbG2qst+uXa1tFod3EAjSbUp5GiszR8pA/AQOKwT7jb34eqcOI3U5p9O1TGRa9EX
B7nrYZCnPgRRh7Ruj7Nequ50MhTWuUbrTpEtX0XcN1n4cQrtwi/8FUagnpZCcTnhM6izCFXnGrnY
NdK1ZL3N+GGdRl+qmlTtxPpy1GbAdV5dv1nwjWNKK0J8dXZEuL9igP3o1TA/2CGl7fb0DaeoPWRw
WuNF4yDZ3OLc+UxYo8r7moWsV/9W6xPlA9G8oI3KEWgWaeDP8Mk+7xP5pSj5ZmPIcdEZcy2Q2I/b
tIN+fgj/48gALF09KBx/LCjAxtGWQAtYBUMzbUgFoCE1Fknel0TZvlEhZ1jUBPzdtGnNaADbpJ/X
HtSwJyPWAzp5k3/eIoPeqFsal+FIZ/N3uPWDOPmA3i9x4Kzf8M9Qi7a7JLMSmQpEJCX3/Nb3+SC1
J4fnG8SFvKyZLNAmbdT5L7xuHBM9CjYfwHCgBQHzIrOEUVVXqoy1aHZ/Ep5T+q5HyKuJfCQjN7as
D1nGoMDS/efq33FwVQguLfzU2uH+AzBRbxugsGK76kBwJ/GmS/CKMNLSzcixXovQrNakOyEcO3wk
HQR0Kg8h5a3EXFF+HGSmloU7pO7Vx0/P43IdvlxUB0K7Vxacq2noqWycF838JK6t9tPdYrQxMxff
6MZ1OrKfoKE103Qni6sN98lBf6U2qkGnN3bgSYgXh/xPHEUPCyVuJzKnaomW8qTXCe7azsGCn4pu
qPZU6Y+7GKHu59QnAQgLim0+5tsPcoCXGibDUpDIE718vnCzDkswWO2O4ROsKnjC7BlIPRu/Adqx
AJOijj/PZudArB5SxtxsywIYeay+antWMQHE+rCbDAF8GnSL6P7sqZIrG3S128rqKA3f91AUmR8e
G7CrVUpkxillLr56f2/U2Zt40cCsI6b8YCIWasDzXVllu62kXq6MzhuDrgPG08Bgh6fMxgKO9xW2
Kl3n7JqLxomSAkrmotN/TCsLoXAMkcre5eWxLqWIfcU5QiFJU39FjJp1bPG3OH4ftGFLuKk3RoOt
FvWyPiD/zx5uJd59CUbHOql38ExKvLWOuUI8WiriHz592Um9U1w5MDNcwfftdfsoecJ7kj/lwRGA
ef2V9qDDizSd4DSY8e7Yakd0ScOP/goC8fjVZoJgmGzePIFGs2wxg9enOoH5niHTx+5HvGKXqoYZ
co48UzbVvuCUOVxiwo3A0be4cZvIDSC2ccwruL3SKd6lIY9NqNEGa++KT4mFFgR0NgY3AjJkCLtn
Xm5LoQNdz+nMMR/1YNsJG70eYk0P74f6Q1nUivoNhuwF5hbrG+CJLwi6cx5w1T3vZ/VK6CZ4YGPR
rGJkrxZ3NkMKJJ2zKBaO5eyZaarg7CWLhQoB4WV746Y1MqSCkPwUaMrYtHzDrsfcq9qaDO/GI0h6
mR4fNp4nTULu/+Y/WbVeo9e34PLPYRvySYrRFcvfMdDBrZNMIiWQIXXWlkqHJQ+LA4ZcPobTUQDn
/0opnGcbgwBNA48UAZNgX2AZlpbykNIYnZjCaMpRJoN7vcLd4CSFTsaiqORLzeYTJ/R/+Ij51H0N
TFUE/bfcE+124zQnHQSbD7H+phtdH0s/j5yUOBArqYZwd9an8Yjb2ztvqR6AKd0fsGWr7cTVX2v1
ea7cv467GiXg91a2+jC9qK6ODD6KP1tH9KbTFYV7QSUFuUCO7rv+v/pmJAyncWbIBJY3Z816yyif
ZeaAAhQOoernCjqqhnSVTPs5YmENzBegr2wO5r5EGcC/rJl9nZZyZ6W1PDzscghkMJmxwhY6HcSf
BcPm2E+1mOt7LS1/pd4nvovjDIEStIjep7XsPAyWVA8FPWa7mV2sNsWgb5zpkW5/PUa8p3zirgfW
+xfYY6PWwHmu/w03IICzHZmjuJ3jdPFLjiM9avkgYQ7Um/J950WmGesCMWxyhohhSsH6U8kGqMe+
37Z3H/mGFt2by6OVvXJzx2H/ZnBm4BT1xYfxjEpLViTnFAoHMQBTLtTctRlDyXfshF82OtUk0cp/
STRS+ur1CDHzfUa+7jghhAcbJVQBEw3skMjvqYywY9zDgkoWYso1M/sGRv86c7eS1JWd6lxPaAW8
UMKAKLvwcCXJI7daQniS2PS3q4M8CFUXulg7O9RX8SxT9LrpuXxkqNZOBEjzyS8S/7eno41oLuq8
ciBckwylzgrutpitWSko60/dllN+VT9lHk1Wgp0RVUv2jQ90Ae/taYJvjb9WugnYkWK8EYJcoCAN
YrojXlP+P6UO6ANHZ4liQDn5lLiQe9fsrbhZxBO8YLpGiNZGxEURXEUGDHU9H+obFeeXzc/aBwtd
l5/N5rJTPZxnNR+9nG+/VClYksXUvp349Fk+ehKmnLDWy6KiEfOhHB3b3WPK5wPMvFgT2+EOP+XA
COsCR3AyF27cWdWQTld9tJTgZdCHcaZ2kbh9L8J7h/L7tximESW3hY7WcwAlKEn9x6vHYMozBSom
J13mMdTjTDJ2MgQOV26JZmh2ZkrgDszOlWW5WeylIvtNKEaw3iAySAbBMp9TfyFfP2H84Yk0yBrn
QE1w7iKlLfACHzKxalBkPnshOwoS0KjEcIkQOP+Ec7grNXFcp4ZVzFYxlmZKg+j4iPqD4AgjbgFr
HIRVDSpxx8LU7EsInDTtTdWziUOcPSMREDMXxl9LzMQ6A3DM4dBsPsLtR0qT8ddUkp8PGhuso18c
SwwVmOK4Wq1NPnxHzqZdmxvXUlBJ2mGv6Qp1O/iur8W9kUYMUdcnwnGy1+WMICt+V5BpmsQr3L4r
ZAazKKaLdVXlaTix3wSniVXsXsDtbUXOJx+kATYVpeJSUHPblds+E4zNXoK3DAK/UYafYJl+r4Is
hgk2PsYIC8Ka9NuBZm/0YgX6Q9KeDS75zuqVMXxSVGTh80Fa0iEi+K9xxZXjj28/kZ86h8ztNT9r
rIVP9vr0Qaabw//Ffm28hCJeqjszGF6dz7HIAgGo3N1F5hHvRJdNWNklMvn6dp7ZVdanIaU+OD4+
fjkfwq10a1gatTkalAcJ5P3TgNUeTLj2V7CGJ9t9z+nDK/fw9XnDFjLHu/q5gdSo8NemPboe07kD
LkoDTy/jfOne5g+JDl5DBnyVFXBdByXz992HFGDUZDJpeCuDa4ycUemvc1jLHU/wT5cuIGYHw/54
SsVJFzmyKtzo4HfgbQt/ejp/AN5boVnmMfc1DCjRpLyjsphGKSZRZZfem31kG59nUqGq6qWoWCOQ
EmPZmSuw2wP0H6u2yDrOv5rxpzTCeCtKTcDD2QiFYBRSwEkP5Qw0qjfNO/4LZfTNENx293zKyT31
ui8dbxMWEmiy0kbVpIHNxUlz1d4l70Yz62pVu3rJF2lbJZfbQcpuwGLNX9SKmrbbEWljg51RnQvP
35+7KzT1V2iZ6Jaf+Hg3azu2fq0tOXN3zr89KjzZZgWg/jmIEeN+Ri62sIi4NkiRHm4zBOKQELPl
CaihcLrEtlDtH6Sq8+iIMYeXEAQ/cnr8FKc9DrWjBUk9hsu5aa0HJi3UKOqdN779AdZ+5v+UBfVY
BSUr5L+s9QWo/ah/IQTZX3NRit0Iu/LkQAaXPl0n+015/lkMeyZU/9SsY8GqtebkQVXZbmHRoia1
jxbmdVV9A2Zapdy88fp6Du1xvMwXPShKVowkcZ1Oo5JtHvFlh3JocXewGW2zCq+Ub8RVFBeNNn86
omUgHUpGzG56c508vspcRu8kf1JbKpBQ0A60xGgVKWM+MKESzeOKZKC55p3Xw3Z3pUadQ6PO1X9G
9lUktiWNyTGW9MfEnmPLuqfQIRxoeJyRzwe4F5C9WKVMIhdonOsl0y4hCr69vDLhIMekaDEcMNqH
VYp0ikgFF4lv1rk9tHSh5rcv37ffB1Qj4WRJZ4fxkOgB1pLjEDJ6Efm8w4l4SI6AADEV3T0lPpRa
VF73lw1VSqIQnV8QmigD4Zn0d3tJ3RtO/3b3XMxBGrs9qZJzHyBudRatvjLCrp6saM/3wlJmouNU
RQKVuUuMSa1yvjtNOwRQuhUqR8E2KnV+pTQUrfVcYd3Qsd9QxGVqXT7ZkYI11oje4SXs8LPh049K
V++SXiSoFHsLCuB8hJQLBCi4r1aCLsMrurpQS4X8iV7gVXqBWQJtR5MPGpIxXHbAzALuo8AN7inb
STQ+c5vtGhGye1dKrKa14EjGnyvnvTdpmJ4crkM3gNXWtEmKVUod1cq+gRo06OO9x0ZyJpnnELXf
kTTWI6xd0QfB4MrLiZfHyIBpchfEJaEETuGKXZXyMvMzNDwq172h42RZPpFVHox+ufhhFk3rTDwm
FMBLjNtX08vyjsftBbxIo13dbVV67/WYS5HX5CW0PSV9Xd6LpPPJNj0ZbC+tCQ+6Nh86GNd95XK2
AWccd+muInIDdlSMmWHtJ0VV1ey87CzUvR+LjU/Dbnn9dzaOu76OY2E+GEUSm5b+wu/kEmf3v0ws
0WCr2MyVUqEYk4wEBNnTgCfd9yhppxPU6BYhQLqbBbVqR3/PW//bcqGE9zNUpRaTt6t1mW2j9KxF
gwZo9bGQORaZe2wt1qUvtsCncsG85TYCErRJV2ifkcwHFjX+XRBDz9nDQWN6HJ5KXiUP529PKvQ1
gjOQndGfla2W7g7uklhqPy+Gigr03zzj8r3Q9W72kuEnqXf1SagDTUnjG3yi7DfVN0P81U97NBTk
aJjpikCdb/85VVz5X5rGtmTl0H59ye9egtjW5a+EfDpoOS7h8TYiqFf8SJiQrtvFRo8PvWwZsMWf
WRTgUE+qHhzJJQHJiGXguUJ63H90BoGY95tYDw06ADBfJx2tpWjAdzW779ctypRE2xui2dSyUgPJ
7GDK4tLHVd4zl7iL8z87jqdBVBdFVdbrkw0sn6nnQMOi/6fQ3IvUyBvCBW4oOdJL/Leef3uOXGi/
nl5EUEF6rMQZbTQEA7SWAYqa5xBRuL/uZ/Qzuz0TQJRpHKPRs+lFZxRHWM2HJs6himEJhv2hM9ZB
b5KhBt5huww+qu/4zf10jljKtaZxeQ5JBaa2RI6zhctX6P2T0rq3VOkL3fsT+AE8PVds218tUVXO
OUCoQ7kprTU8RBFfnDv+0cu1vvRQz+GthF8/ojLt4TlAA5Vb0LWTB7MwBCQRhHKWeXSFM8zvsyvl
p2ekp28jeOepwh/HRq7RxRI2SJOgkBxeOxWicQS7M1swydfwnGtlaMJH6PPGs63GXvHqBOot0ZqA
hLQ2VwPaJXNZuS/QT6CAnnQToGUWK8ckvdTpY9V/EEs7kzP8XQE7sNnI7LlWYUAhnL5i4ltgPtAQ
kX3cTToLzk2b8bOysjuIiuealatLsUIB0jIbjRJbxO/IzM+wbP/NL5V+F/eIe2PvS9ttMix6OtzF
6M9CCAKLR6L+t47L7xylofApTxPa5pAmRzH9FyfJFoOSIx2EGYfxRcVXJu6XPn54ixqFpencYEDr
EtnL8Ic4Y8o+2Q3gzAPuoidBND6xIiKug59dig+vqZCapNjordTFtXe1O2pK2ekJk8exkJ5lZdPZ
gmsUbJJ3FLtXR6VzOBKU1+BoxNj4xScZsG00nl/ZwEfcfdmJRMOn1Gq2aOKTMFE8XJ0pZTNVH/EI
UEwQkeSNkKALpnS89YTEEeUiDBjzrmZK0V1139GlorymBAMZdHPT8+dZetY18+ON+xbdRwRsKpbU
XgAPXlMyAshFmMZM4CY+yZVZH+S02G8q2e4M7ZE11MPH6h8/ocqHMweGq8UMlqK6Pyrs0cTncGmf
AC286Bm5PIaasUKSlQblbyIUZ/PuhCZ5mdbclJaVZj1MuTEaWuktGxlofl0tWFobypgG8NtfOPks
xX6jV6R3eyg5yEWvoIogI4Q+YpEMa/6EJn+dRlde3puETbzNZVA9+/G492bOoQtG/Pb4dHv2T51z
ewNbJly3/r8mVPvTYcgjM4FoHcKPxk/aOxJTqcMqeyA/5xbFhGgGFFDso8SWf42QAFbdnrXbPpQ9
7126+LvMpwSHTMZnRFWRTIrTbhdqVDLOG1G0cbiYxqKQT3s9kO2ywtrDdTkjvoTOgESDpZ5ZrGyG
iA5mzt94V6M8d4FNP5R4H7d34/tlIDrR4r8XTHdlUQ8o6v9JF+y8ZZdhajyeCxC/dGPPXBAy1oYx
kUUXMAD+DP6XBQMm9fV7CXsUPM+QP+SNjR5HSqOOOcaEH1CguP0hF4Zd/mfOsh3YT+dJ/SrNWI1l
Yxlqkr4Su8JF6rOLDIWmbGZHhsqhAVW12GIP24VbjvPest54vhxajJihrJxqH24Q7iu56cPv2HXM
cM14pwm/YebgJDOwlJkqQ7GulANqy36lNnm/9mTtFh+dDIOVQKKqOSoE1rhuu5/CiwVGztCBgUj8
Py1mTlHhTNYSdRl0z2UMF8M+O5HT3LbgRuD+Lb8i1m/mBRTUxkdDoIFaEY3VzwmBMdpY3gk8pDq6
fH4jXMXEHcSulOmRyIDviYwYYepBZ9i5pH3mm1idjV3c/CzkA0c6OORmw4nBM+rp8x2UTW9eAEiJ
yXBFKOz8LFDSFZvrI/mO503Z/QxTSAnidMEs7rffelE9GDoFyleekQR5P/8ePSRG5TIX50aC35Mf
Rg0uIPD7ZTsomIeEQ6Ad5jKrWb1Z71MfsPoFUQbj8dh/EykbwyVSIuzkBsxHMTH7QGYmCX8xzXQT
poJn0j1KosJFeqTdxGcOndZTcudRUmMurp0XCMbhIjf5ph7V60py9iIjc7siejLc4BJkeD123svm
5UcfOKM1fRbBGDlgEHPNT1L+Xj3G7X6pclHY2ewSFOHOqPHd70jBAfHyyHiLdDPtYa1SGbYzJWDq
2YMuXAZVaqb4x4OfHwcb4PW3H8lGcjrhbkhTuS1zYVDZnJjlvHSkp2qnKABYUB3gpF3A5CIaqtEs
JV3zWcSbGzXugw52wiZBZuDQpoTNvOBxO8UUcHttuBlIIeML0s+DG+XkeSgaH39YYmmAyuHX+yqr
2si4lI552cA0schmMqR7i2dBi91Q3TXu/Wbs8Q93h+i4oIuoOZvW6ooBkNd/Cu563dtL0xaAS5wX
uwFwutzbOAmYV+FpXp183mbRpA5un6azXxJT0+OVU+lpBvv7Wib1c8WXgUrnQ/nX0u+fvM+IuFEx
CerFrTaxwyD/Yh4ynd32pYeD/cqKv6Svm/L9NBhFfiSjC3K3Y/JhaQM7uepbPjPL1cuJ2wyC6ixb
b/VUpbBSaLSWEoL0Uvu0fX6V7aUM89KJYG+oCDj45avkF9gVi89cIJLiRBpSfM+KUTM8IZL/ENRt
926WZChBr/1kfeUDbotzUGJvozofKzqEW1T+ZHMyDf641anqAmaxosE4/DNNGosGLGlgpzF4j426
B9weTnklpkaAgRpLHatjPNpUIuflutcxBTNvKsoOVwUjXoxQpdprhw0JLOmpUJMb/JU5tQOI8qjo
isp8Pe/ppZIvwabRedhkAWrcApS/s0tfNLvJIX3jOUxTWZqL/bNYOwKw/tBvboK1TdKT5ZKXO69J
xgVExvoYbAk5Q57peOwukGThvjhZbi4HwsPM62mvfaHaqSlzvmZO0hRVlJLCw8WMwWxU+o0iR2zt
yk/oOEOu7RNRJjn/SW/+oraTBO580NGAZlWAvvHD7toqKmNPj6n4glYgSAICcSOn76C7DoKSZ72O
88ZF2jYUCNAHvNOzi4sZLKMhqtX9A/Wrcbtq76oVBE0UKUVoZ7+6Ae8h6MEXUq5WRtmpKr3C9nSg
WezvtbEiw9dV5MXGdIgjlNJU+xLrx1z4sd2Y749dO8r+USz9gSPP0P/nAHcB5V6FO5Vj17wtErpV
DzWpa9OLvihOTgKmUiioFgHVOfuGMp2tqBwFkopWb6MK8Ayfo56KbH42W26Qx765IjhSVPtkXs6f
C2IurF87vcb8pTRL5+v7orjBwYtA3U0PWerJ4E0EyAc+ApUcWazlcaiFLetWhAKPZag/ZXfXrsiH
MU6vdc1DqBvfIEav0Mfyj9qVH3P+qoHHqnKJdUkbQofU9f2X9WxlopXA4C5FbM89oX+EXsOPzYgN
YccnzjxBWFQOChaeqmLz9YUqYcrGLZF3ZkXDk5rVa0oZ7PDEyw8FnYGCmcGaiIsdll1WCS9ChqTD
uv1cYsza11h6zkou1Vy9Rj0OCqo2jPLVc7tUwxXQnD+G9IGNztbuRF4W6slp7sFGDXswx/euyS14
FJs77WmJtUfBqhzM2qVxFC8Q1Fa60bf20anBQ21ufY8Ovvpl02GYZOCP+JFQWV70ne6JkqUVeDov
IAqkswAr2vJLDGC8wKBvdx3Ug6lFwL87lTOqfwgC6tkZS6jbjzSEXyY/7yEM8GI7MDjf8l8Jj/Sf
2PD/K5mjrd0ld7ijHrjohhhLND4Cm5fR+Ns7mN7cSKK+5v0M5NOPAZ2ryVJz68LKoTKYNpQNH74Y
trvY5lzIzU6PL3AHlHMLmkP1KX/LVN09Zwh4d4qIMGbx9MoMz2PoyqgM2gagJIvXqhst77qVfnww
Gi4XhqqPC63uZTLpvF9etbDR/S6/rjLzI6RNMwJte1R/ZgeE6V6KYfbbVSKrARybR5LrGutLhCrf
YtYyLruTln4bLjZCfEf4pkm1WsjCUDtr9Kj3JykWW62/p6kZ7b7mbWCOw4Os5h3bty0Zmhu9Q2kl
Gu+01Imzr0bduXKTKMsdFSHCs5vfnn1egxt1skLxKG3rERQlcjxqNqyZxY4JOxgwIyanB98v3o8d
mJFsQJu8Fhv54U8W88faqkSTBpxqNBwfqYtFQ8oBTju0C0SF5RTYk0EfNBrj01n8ibVJEII6SnZE
Ow7dtYujeJOOibVUdMwyHNzhOvMbSQlr2S/UG82sr1mE+q/lpYm/M59ZzgQimm1C2CqF+jimS1xH
3MyJovDMfaPLXxIHXSXZn/kfteVD3wVQw2v1dx6BsfFXVuuxM3TDuJjrQlUcweLspdy8GLjsf+NE
TIzu+fE8jQL4ztjff47rPFJjwZXj4PahgCnmkxlZTgh0KSTHmR+s+4hwMsKi6GypXuNqSBK7Awbd
1wZWFHF3lEXA9Zi/YfNcnTbPXCVx05Cvx3BiU8LHs/mO/JSmLnqDtY+i3PP2w6TseyYdM/ytBzjf
0eCqH7bon6XZoQNq4ORT3g4QJwnzgngseZFAD9vR113/ylPVpFGlmNomGVv3fWn3JLH2o1lOi5Ib
o79JyEvrGpPUnLkF7ZRW1w5+tGpf3elB0kdYZlryK2/TwbtNie9Y19rLPbEfIdJGm8fzh0Rj1Ybl
wLcDNn5YGqqiNhU+EGbKe3X3C+BnUtHz6cWD7U2duqWnKh6cbYDtsebCP6lG0YX6ghGMXWHOKpOs
w/gQfn00dy1cQGSrsFAT+4kd/khonHGXJihuPNRzoF1s9HXGJsgWipHeu4pnDzPndplXPOVayrJJ
p+tbny4qmZunimkYIxFf1l5nlCVGXWKX021Xi7Thk115v2YnYY+E6Lx2tqFm+cI+L+UdBcgymAog
AVdi80OlFWz932jrLc0LrI77684yMhuXspGVT/Qkc+gtZ9Jmm275x3uUaBroY4EXQZIVxJOUPTk5
Rt0TYl4O8R5H3IZT+AgYGBwiEsE/yZBdnhTPBvu4vZioJE7Y5JKooT7rJ60ABgWqNUNl+yX0IPtw
agSDNOyqhQpSPqwv/+5utT9dy8vz+8BBzAxeBgI2qKeGet9kLmKxL1MjD26x42Pu3B2o1fdIizFJ
1Do32e1QETa0zqLIq/psZsOn3fJiWf79UbgfpAJRTayLjGYoigpL0a6XwhioKq/G+4u+QHDflXhG
vwTVFMRpxyDIRe++CCPoUfXTHYpB/knJjhyh3CBd0Gc1/a/PG+g4nqoOXU+OlTeDrg6hcJYCfPDQ
xUWeKv9bAQ6rcGryoaid6gg+x77pkrtLiuvlRMUvCPWb/2yC3ISoj45ipF3vKRvw6EQc0Xy9iKGu
bbFrR5jVoG4/1+VWv6nMG4rPhhnf8ToEjDXGzd51FCfnxHbOc+7zPIM08UT5mvBFGicxYS5L8LHR
QDke7LNLxndYZkj0BtZahCaUJ5bLDpCuH4BzVFzHL0HSDVrJka05IspLvB/SecqqwVH4C+g73bUm
t5Jc3lSzLt/pRnooRtGEZEA0Gpdr/PtFORdhadxXSjKxRw8pXLoBkxi2f2uAfBoGrtqEGUgq1nLk
e6ylhzCDfJBKXO+ANNZnup6MaydNXsg6hYIZVYE+txJ/HJrP+saaz1NA5wSFao7qM9oz3GlZVsUU
dHMxi5SmMhKBFE/ia3VwI2dqQl87dEm+1//LLFLZgHk8YbVR9mNDsC0YMBOpyBvxuEq8m2lZzpkg
cCMAfJLLfcKkw+WdD8kAMEwNDc7qIfTYkpUj8WgC/VunEJywD2Ni2GyI4euzfiBHkvdlIQYJgTdf
F9TdijAVOUeegzQBTB7KBMVZvBZDB4ieYCcPgD4hztlNCHNvowLsjfIHQBxq9QlACIRdY78lR/j4
xquVkgYcPDH8JenrS0IwviP1Tram365LHx+6FVnmWD4IhJJ/zPRSXsi7dXp8/FsBBsqTeDQo3rbI
WDrdWK/3gvy7IQQcVX2J8plbAn84+4Hmw+0KF4g1CQA3nf2tX5Cxx77F68pwtLgfr8esLk8I1qTe
evMUHdpY7ZdXRfrmtPyAVq4zhMiLR+3YXdp4jYzS+DJFsVwkXjivSVYKemh4wwW2zAM9rEuPugOi
oJhmx4rJBN4PVJI6ch085dccDikkaYlhHyIYTVskKTHf7FubC7KYSyvVH5G8QvQi4k+zesNO5YZX
FM1lQjboPdffNXc4brML5ehGCHRtzG5javjd7/tTO5qmTUXqoejlhvfWnbHNrWvUxTqyDVGnv01M
YhiWcC9aO1maqAMCh8/0pf85WxcyLR3khiVwQYc2yoYosafBBAZnCRBUUtGrZWDy78/mECXRK8im
H+IObR8jZ/Hyc4MyyDoIXDsQupY+cSjEoHOuhKOEnJ8XFFG6X4ikKDgEXXdZIqS3oNAr5uBN5ONf
c5/yO6yXgNllTOSrxcQYveCJplNN+SN7uuNkxy5FKc9kv1+RVK+L2mYKURA1YcrwNr7IfpLpRGKH
LD53bq2pukh46HRR5FPDPXGMFg+00HcGHFFyGe+d0+traxEFyEVvJ08qxXNR6d04dkkR5rv7pVP3
Gb03evY0a3r7vxkbpoGhW7CSLxXO98a7+kgbOSxKU0dsiVndb8Ika58ufRPj1u5Q9MplWeGZXMav
hWRCqxef67JcUB0h1ofsLft7FSuk8wWRO3l2izy5V7QXcUnbR4+N2LN257v64xPYAypxj59cjepu
mixMXXkWe8OAwCGFNGSABCeGNpCumWj1cBdG/0ZgFvEQkQxW+PtU1tHVtiBG1oTbxgj1Bl6k3BoR
ebzArRWoWP1UQ3BRkusFhcJ1KLnvR8IQwg9PmuwXU+TD/JsaUUnGExWebRJ9SmfeYebnTrvS6iy2
Os1Jb6LshECIq8mN9niDMMrc7Syh5qfq0A73yQXhM0tDdoUums3vAnSax3YmNHiXDpu1Iajnp1Pu
6DbTMG/ZaCliKzrTJJ6TxMWP0bjzng7oTWCMqaKDpXVYF293byKemOt5+gy2a4ku8Ps/nINb9pU1
iuSMQNUiaEJX/UHf4wtYa4wZBcinDNKLCEreJ3HjY64uxBMp3viEuS6u9uLpJH1ICOzfIx2Rgrkh
YUxIdE5LrZrVDjQRNp/AgJD0WQIdYknEqTHiUx7ltGDWTqh80RbGNTg0fgqrgs5WzzP2S7UZyFjg
ZhbR75GGUZuEWaJkxPZFxUn1IXBqsQumQnjXeMb0gJAHB/l300ubMx5RyDOiW+30KGrRcq01/dqy
lJO7n6Lm2/Dh2+/3O/UuYAkuhz1U8hEpmMzrdSzD8iNYtz0TkocDNPLYoDM7BWH6o7oKAUdLbzWC
ZZk/4Y486DP08+xdAPxdPun1Wnx39TTQaEeVvUhljlM20JNTKosUN/kc9lmf59SEh9dF6F9CeYeM
gpmDnPt17rpFnTIpeYPVwZtJty2+gQcCl9LIyLDButqcyaankgRhROAmcjjAyx124XvcC1E0O6WK
g4nNfSvny34Xk1VbY4RP7oQ6DXASZJTQJ5cu8WGerk3dQQasAmlzkpRdkDoYG6NH9ZDviOK5aHRs
e2kTPAImuATtaXZrlr7jThkqV7NkkqD6zfduH3GHlE3JGLIbXb9zFFG+Y5x0db4Sp80hR9NbXFaJ
KFS3AseUpob1i4+hMSgptVXhaYXmE/kOmImU60mRiPo2t30wNlX/0Dd36TmMIayJnTNCnebx10LF
vTa1q0KamGhpAjUcgNkoDRsA2VV6MPklR2IMd4NUafF18tlScEk9AGC9XI9GIr8H0RKpAZIkOL+3
Cn8RPijaxNhfGiV0hdI/D8fHlLHpl/XM2AFHhle5luR6S5mQYYk9AjWldNbKYfLOWvmwv/ToPWVB
2jRQe81Kmy7KC0plhMj7AxoUAD0zo/jFUjJuRvbsUSWx+616ly00Zs4HlxOBxv/fQVoLkkbnbQIH
v3t0MoQ1KZcwpZpvTwC/h15pVq2xrsHZZ56tH4dvsSIQIhtIFpbq42RYnAzPaSH+gYjaQgbsYlv9
jcMEe9egQmCmLv2KcajMl1bDJ+qP7Gy02UFD4scDfjfTr81a21XdcUoIA8t0brNLa9XRUHMBA/1P
zhLkfeFr446lNX52uock1VneSm/1LcRDBKl1bA/ZzTti46Urz/HqM9AmGybj6svVg09Qqk1J7yKk
FDGuDxQSZt7OUSlZHZ/n4l1m6nseLuqipgHcPQ8Nri7S2D/yfKge1xPj4b1/NDtkjC7H7o0R6T2r
u5NiQyfUxLbZKmXuhjXjs1TOCLaHG+vHgWWqupuotQ51xXx/hnAMVmQBq6eCMZ8JyziR3jxB1svK
Pr75El4ByCZT7avsYbkKZ+/uyzoXGH+++uSxgyN07Y6uZiS0/sIpT2Z3WqhthNMt1RD7T6pmAWFy
3Whx70wRHxAmk0omL7e9PRegRejbtOUvl5J+dYCKybPYCASD07S6NF2YDFR8rC4iFnvfkLY4CDid
Xj+Vsc1MFhz8KDy+t4bPGYhP7NQoCy6LDeXWF/WsZFM9n8c9NHD1WdLdkBJJDgOjmCoFTq7/JYuO
Lda4AOe4UPKp1Aco/MDmyg55AwuJt/Qu4mTNdHgm7C5c+8nmH5NH6cor8NJBtIIvU5SFi6hSQpgD
tGWY9ECt46supZx2AMGMvIuxgxJvs/YaGyt+7mfFfbbijJPSieYB0VandlmpOPHN0KMscshhLAK2
66CNVXfJ2LyNhistmNvIcfEYfrgM3+P7CljN8Fz4CLZrMBlPMVSVemm32ihfEmvs1ynlXpjsKGL9
Ew/usucO0t4suvfr99QMbP3lHcuFQesC3+qxsHrIuL5uN59XevFrqk4jGMNLs1fWQSSuSB5zxzCh
FjG4E39Dj4Ryr7Nur9ZDEr9rVbkf+kXErYBkU/pzSgM9cRm0c4e0hMlckZbVh1b1ihUXdHVpCWRa
HfgSLL8VqA6zHUjDhWSmjYubjHc0/Tx7h2U+aWWm5RMI7O9xYalZj3we05mBw3Qn+fgQ6UN+t3HB
igVTE5eiAYdIitNdSKXBJRhIKqmFz388MmvSwoQ31qqBLcsk7R7F3C3nyORsKaw5W/6gviMT8xHG
j3h8fsuqQCg8KRLQc/XwFk55sojPsQbJq3Wiggy0x/PypU3cG4BdB+zzCM9GAvvLHH6stIKEpztK
Tthzv7o1XB8E4Q7LcCgCfoJtOZj7zPmPpKoSKkOckuQUU0LwPc+xmy/l8Wvl8HLzztmw1BzBMVWc
czW4D5ruAYMrRdV/kzsEAVeL54i1Y4bbK4KToKkVxAh0u2ym4HBhcoK5Lyxxj/vq6ZWaaBKtDWY9
KADL5xMoDOWMaBXum4XStbeY+/20TEIyeMWiLLM3zVUPJjGuloQlxmDZeBKn4qPdKzD4Wk4n41kx
xZGEf7hUsQ/mlT1lvN2Aj/4nQWFujl6G/IVFhr5WbVDGZqUyPL4ihWEE+vq/4S2M+0Ec+XlP2pJc
9MNG6KJ6HQGypJAUD7Mrc83u41NOCEynxVyds0PuXAiJbjOqUj1Hq5NKIQSaw9/48kB0RSkkJn/v
Ut4OXgQsGP/y4bSmNmwmovRx5sJyrKmt/lqfCeIPkQ/Yh2uQ/qySRq6boYbzNV6cnQhZgEJhf+gO
01EecrFvJ0whq0gyiZCRdVtU3Tmi1PkWqccVsEIxjdSPiAPiGdpAq1nOHPO6t/501pWkuQivbnqs
l/dMCqE7JKwtRsVZnNJPZo0N3C/GiKWRe07/I/dpp4woGuhOCK4x8RpvIRY6TyRNxWmdJXQaAzqk
e0PZ7PuMY9TxBHHclwGNWiirOj9PoNreRR+44bJJ1AemPV0psguxVoZa56D5VucytsdYtZHEe33P
N6Pn+QH10z9Lotfct3p6kIFNMQyJrgPplkQEs+4NVMlrdUgLYke5bHn5sNa+ITLbaN6DhO15LMtI
guBhr0PCjhAQ6x1N9XVo0G8q51+Lnh3VEmeNjOJDkCa26Wx/sDMtsf5zMVKtmDj/wp6uywzB6b05
2LK2SSC4KrVDNJovTapHGsS/doRnr1gGQ+/uDg8/u496VDhbVU3ERv4NBNacljC/oi+3a2d46JfZ
8Fn/8gENuFUnfl1k47cXloFPQEAJRL17jIunTmRRqNuWsnoUJC5DGiBOXbDQVbSR89xt9JnhB/0e
HRdRaRw1U2+d5f0Vkf4gydTPgwHFxrZ04rzVaHih36wU8Ti8KaDszuMoowX8rMchEK5aKGa5XWz0
+eFBY8BdY7uHXqpg49kN/Qhakd8fqNvcDYoOZ6jt+n+yQEWfmI6jk0RYRJ9TdM+ILpfP+B+hzqy6
4LtHxkf3Py5O+Ym+9YSK13ugWRUjcUWqkmZBm+rBEDUJpIgY/qW3LMHYdmTPJLHOw9fC8mAsBef4
7/7WwbfkWK+flyL3Qz8JCSvUdqciVOSqXy8rd2R6JFq6MZEQ0lR8uvlLtnQEGElHPyFHtsgMqY0R
Q0YGNqcnUVoSDUuVLHDQ1bYtV2SaKYojPZbOswvrCfu+VCv99L2w8DC05XRPMvEwZtezmWKsdrDF
bZZmJ1RmgxJLlKVwUFw/JEXgL55yQiJIbimsraqUrpN4AbE0AdNOJsSoO8puQtZdhoxhVCHir5n7
WYqL8NYPl84t0kKpLMWtBxrlxReYD7X28avQodGt+tixd4x0ExffALE7qs4gOhzpnUtDPZ+Agtfq
xkBoyzDxDemypxo3Vbl72aFZpfnUtRmfLAt0mDPpxt6M20AkWICXYUCYlwW13uac9IyM2u0Lz+eS
oP8lb+VC2Fza8m+QvnPo7pL1TbfH2Zo8nh/uEds+o72/WyVpFGJYUrx1VUigzqwP43F8Glp7QAM8
vgn+18l4sjJMcLKWf2lEnn3r/l1shpyBK7G6uI+80p/Xbn8ZuHMCPUdzjjkaYBc+N79LY6ZSQJeA
0r+0k8SDOl7GORQnjuNl+EPibDOLRjqw4t18YuaWBFqeoyBBBk30Ggx+gm/vLfg0U3fwxFHEUARc
c+m0/I5fKpvXqxS5j/iRP1MwKV9NEOZOCSJBJBV7Z8nHTpD9igivnonwXJ+w+6+YTk6vh8QRcgUe
xnTPTJ6BIoRq3GEw1886mc2KemqsK2NWG/uMHRUPbI3sh67T6pp/fC6RjOi0DXAiL0aSpsyWsrWu
lRBswq3bnp/CMv7kH/MGqMclVb0OYyGP+bk0lmqu7gzGFxL2sTR+oSiTwG75OtGC4aMc/N6qXuWr
ul7gzSA2kaJS4tKIrrfwhWcpqo16CYBovS5IkS4qMaSlzZRf5Rn982oqxanWbBLb3FiqEZfZtg4o
6enuVu19tlQHkidRgxQQcPumnfmm5eVIZSpOjblyeSAfnaUEl1Zwi1zbT7RqL//maDIKWd7rehl4
AIJmGuHxqxgAuhcrFxlEmB1MD6fv0psvWCCh8tXR4UIAjgBFcXGEoPAYbkuhXWaTanPJ1GdWd6uG
P0ZKNVy63zAHK5RizkbUWjQd4ZuVyPEbb9EvtAlc/5MQD1tiaJ/hP56pw3/+3fXckRV+ZrWBqWHm
obe3NLtuKl8wUzxI4WDYj/Zsm1ZZ/OkGc8vrxMiRKCBOXJsmcW2zSOHN1pcmwkNoOVGtlYhRZsst
gFSWiwGUg+sRCZDnxRS9zN1QEuOHevDxnbWgTLYF3gR6a/5t83BwzlfNt41Z21ztWG0nxABLtjTs
B8Ezqf8GpXjjpYJox8IjDLEweUVaQ4r5O5mYRrHdYM+qnhVcIRxlcnAKts+WeFPOpjSXlybvZoPB
ztv9XTQPjqtjXAM9QreO6ZlKbRUOLSxSnVBFhUXy+l55hZJ2Ld6dpNXtzzbqnfNTMsWdAVzCb+Ot
UxuVOw9IirIDThMqAtYP3acFN8GPOoY0fzYuvF/l6jsAgVK9ifFHsT6N44adNpKar8XhkCya6ren
g6qHRQmmQPVhbWIDwzA4wXMBwRTbLqYYSRuMxj4fNyZI8How3El2cDzK/MiK2KWxANKwDtLEGzQr
A2BfQpnk3LODsGy7uAi/Og4/8SM9CJNE7XOTAYGflwURZtCchnK9XDbcN7/zu2BrqtvHZzwy6VqK
//ssWWic8nNwJPDBwdtD69p79aDmO8gftDXYfl8qNxRQ6UXHaoKbPFhLWlvPcueAeFAoEt6IXCLd
vjwfOdqxlOGLMRjioJPJ1VNGoandVl13gLOUn6eTQ7panvwTe4+aLtg3TcQiKVRrV/Y6WGR0CueT
4GYWSfkWK4AZ0pJjHGNbilO8NqTl8cAcFZ1cmrVVssP/TLsYwnITJEzLqJ8EyUDXIMPjzC4/dBxv
OXQoif6X6I6eJooNShqVpZVcpq3Di0umGdoMUChoCRyhhti1USB13Bl7ZpqnlP0/H7bhTIGppk+A
hY4AMIIJT4TOEhn+AMcKACcYcJsTLuK4iljEw2I2uqHVOL+fcoMMYqviazGeYvT4KAdB5qdfEDu9
R/uiDie5vsixfjcOGNl95wY6VFaRD1Ou78XgJNcXcYt9bhN3XsWAlygI4DS4zhyJU3q0wEfVJ5ms
EJp/eQyW5Cw9TZH7bSfAWvu8Dn8jwXued0Pzu9PZBHZpQedEfjcvNIe5tAM+Uf6QK5RGowV7aQxA
0vxaSlFY43NxSdOMeEwxyLS8w2suT3Milyr+dc2DIwAPgCbofoP5f5hZ8O4kVcIjNEC/bHPNgsft
YHLpCtFzQ6UpPQNL9Uhj3r5bqyDARZc2VS/TJEThNZHR8+pUIyZzJPE4hcxLA+Cn+9isoFk7VySy
GVAnBpij6mtnMSh+PZh7YGA1ZfVxoUCyLF9I/P5hiGl14dZIriBcwK7SdQapZZhgUNA+MUl1ynDn
WvlF50VwXuYqugSJZrUo+F31E2g7Hh5gknLPn+U8+ViK7NWp74vZEntEa05YIVcbREyawJD0S5ph
GwXf8YS2zKdXo9lTVGSLRWoJRO/MgzNdoQZn7C2VZFzWWzvSbydHxeXpma32NF2gufkBgkSYJqaW
VrXyu/Pm/NrEpGRLJhmo2ZDqZ9FkVPxYyj0xcfFiOKjy+kJXvBcghY4SxMm9UB8oS7QzrMH/b7Cc
TsjxNhnKPzFVBTWqYL+LCrZOL/S/BEBO3oHKmS6e0Mdhh43o/Hv5MYcciXtUA9nSjCrGP+uYT+vT
iUnkIakMWkGdLjgYdxA6UWM8egzaR5AoFcVQyv6RQAJ68SQe/zggCahHDnDm2T6hVnFinjqZYNiD
UCJJf5InAxwo3czMle+V7/93zuuellfUvY/YF0fzoAWzr1goJisPVMDV7pQsb97TrbveOrFt22pO
uooituxfneSDFrQ39xr1Zco0qxurSWW+UUdQrykBx5sWh5YhXgJIcwi7bO2ZbIG+kM+eQQljq0yB
TRUjArug37n9JONmQBkR0VKXNbuYogbBb/2iJxMgjJ/pslVb7BisQ0ECuSBxnh7FWZVjRotPAu/8
wMmEYIgrTSNxVFGMA2oArdJVsrZco2q/8dZBr154txjqZS5fAfNicmLoxV5I1s9A40d487WLNDLy
MJypX4CVsbxW1MzZbxUOWfnYnD2hb1dPPZ0SrUzDHD5/tM83TpjvCWzMem6GRa0DCbzoIIKTY2/0
7wrmYQ4WtEzzRsYO2KmbULgvtUPRfF+ZEEQKv4OKkfumZ+bXCWjnDP/vKuHzaL+SyeicaI5aqVYt
o5DE4cZXLUhH3qnEXpNbji57iH1s8qxN29cm6/ltOuQ19FVt4aY+9ypUf/iV4QKbDeofdZK85TXz
Bf69kJUcMz7QVl4JB6nJ7/GxrXjgmpd7vO1HfsdiKuehiY6JEXhpJNFjRz2adLBi+ak59iL1A86d
pZDHvVKxrvVqN0AX4l15Fb3mbgCoGUVEtmY2+1/AYlqIfXUs8a/UjMEb2KqImKy6ojXiHEUTpXUZ
ihELAZtsiD6MHGx74df932X/3EIQGixZx2rWM9Z9Uzzjj2jHOfy9QqnGHu18bCjamam2csMcqq+F
Gm2TOnCWuzr7hELr6pkDmZJGMA5gMzf/3cYFWZP/7Gk6/Q61ShG9ZR5lXZndDBGxtWYXrOOtKo/N
1XiEfULURI3veEW65vrCqidhOhoO3BXKTdQ5Y92tuvgoIHIXjnEhe7mCN26fK7LT3BYTfopsIJdR
f3cgHWDIp8xy76K2QkcoplDoZnNL9DpEMou8KzGoQeVm5W6i8vv78GbNx+F3+bMf78mr7w6cdhgd
1GXOp1dRCkMmWjnJ0kBURX/HxhtR97YbZis3IFCayyJZfMalQ1/JHL5T18vPWXgSayiOY/XVd//F
ULgD+o14jNOB4apsRFKMnxo+jU1+a+omI1An2Ae7M5jEd1Va8Jsi4huMzQPly1sZ79l/v2Au0GrG
r3hV1IflYIxs7edGPh5XNbwRKgYbBYzS2sq45cPjLB08mMPj5vSrcSTfU2yw2QJFBFwxqhl01FKe
6IfLxNX/Cjkq0mSu/iYsPsosJt7G1HvJrOUuow5eXcZTzazdl43Ae1lsMDq/adVPAdAmbw6Tf4E6
tEsUiWncwoRcD5UE3tm4huchrC1004UQux21Fx9QPcDKM2gU11ngSx4WpSCdmMucOpkaDSM6YR8l
aN07us7wI3/FPNxefFDSAiWLxri3tOVHg71pL5ZHbgPltpmVYgOh7q+CV6n7st+IPnwwKFpBEDMC
HvHpjJ+zmhkrEiOL34u1zxkOnRmuFXawmhIWXF1Q6VhPpDbOMLpfEuONH71fozC9dNPEa5T5AO4y
wttsqWODGCw5tJTFur1pYDNIiKVn/yUDaOwzfdQepMZI8G87qCrEOr+mCJJS1w3RJkDmIYC+HQ1J
k2fWSeH7E3m8RLI8tHnwMts1KU69uMKcsrz7dtzn6VfFVGSNqLvkFvGhEGejvn+U42C89n7oLvt4
5lJKWfCqWl+VvjnDr5ht5PvNRZyqQgWs4ho/i1hUhuZDQtZAD9RTxVy8rn6bEPhHxAv3q4Q32Xuf
7zbs9Mw0kerrOLyngKsEmqNPURRN5RPUDazKDv+znNJ5yR+E3Quu0cAAbT3hFYDGXYICjpxrbY4c
FdL7r9ZAYJgVuxKoOGS+6x0SQjmtt6/OwzuJS6EhDasx6DIl18vSyi0NYQMqGulJk6VjRUaTWC6U
cH7WdNit9IkRWmzri8wMQkMCf2UHil4SZuo36yPQjAoQgvIwC4J6bva9b653QwxizAEVeoZ9hS/i
f6644LHDUcomlJq3MTAKsPAsU04/sxP7iIpz3xUjWrKV6zaprvlX48VPjLQz9lJRqQTvpEwnu4MW
H/chQgz7dClqNA2kt61vy41WWjhJsLn6WDi786s+PFIpHB75O2jzc88bRGiO723eWt07KbJQhk/m
zWpNx3a8wZGTxBGMqzIfPZAX3CH/Yrg5WfgQQ7irZrb2BvfiQKGc9TdWJsX0MHY+TrqTWEOZlESz
Ul5fbWqhM9N1HuFMrh/1D/bwfu97/PZwkEBCKzzzZQcLXZ2Ig/yUp55LQ9P2KJWPNY+1AyAILulb
cj+qmLiY3IKAg2L19t8IqOaJ9vbRMZJpfi5pRRiSqxI++0arNr1qaMg2vPH6y2K5+ttf1QoiwC+k
2WgZzXK+Hp9n2cJUDS14RHrwQq+mRQy8NLne2bHH12VOEEg88fKa32+uj00hryCUOFNSzQYX/6hL
n1OIQRIWIaBL69xb6L/Q0a/j8syl47XK1fFjP8MB5N2vfcPTdj5KqRmzjnibRpV1Io1LDmaJURRF
r5SlnJ9uUoE3wa/dkVb2ZBEwJL/WIfGbj1WE+Ol119TwCeRN4liCUkLdDiZ2kItdDeHoSazTNCKc
uTb0izkHOT01p7XbVGKgz9LFbWwfxFQIbvTCJWxmOta+HjiBNIgOg0PUv/Lc/SJodjKjarTY1yrN
qObMx66PqeRSE0maz8xHjsWR2XD/ixHd3U8daU4kTo/9/og46DoUKTz0IwfX39xJ2ynALofetNSO
F0BeH0MzGSGvl+/jVlNYLnkH3DMRO/u0h2Tuq90PlHQCUApS4dNXql8Iat0CfboZj68HkaCE3t/2
fl18zsi5GI+rfCtMuJVDGZEQxFfTl4f7L5wXOtKuoBuc91bMVZiPGEhkCqGOlnTDp+79UqW0aDKn
+cOQBuYFYTuHVWkRNzgGWGA2/V/OwcYqAeUNV6X8czp+08SfqNW7mXIQFdSQKLq/EWORxG9nP70X
OXJn+P1Ik8e8ALD1z6IrXm29XrkeFed9BIGTJP7GllpBsIsOgAbWjQJpGhqJ3qSuBd1YnaePBetc
3dCI7oAAIf6HMfozCpXnTed6cfpsrKxP3tKsIID4N2OpHjHSZXf+DMZ2yS2uPNIE8twrPMKS+UMx
PlNnLtLSHi7xMoTie63ksO3DdYCP5SBJ9/ZvnJJLItiEoncToBohrL1ktjVzZlZawfiyEbKApv/m
B2zfMF3XJpoNX1H2fGt6niUgpIChFfH5+9Ty8ftEGhYclI+lXrCpHfe0eAysg2BljN3D5mhtXE/E
z0B6AAtcbyY418REu/o1iTKOjtDpJ4K5QlHpauaAxu9+/6sEt8cGjW2CNgGZ29N0GBH8/U/1Ky0P
UtJ6uwLLozu/VVAmlzGVtuRMV4wX8MR6KFOl4ZE5gY225hKPKXOzrUq3sDKGQIUNIZWI6O8YHN95
DrBQzkDeopwdLiDaZScmpiu8ZLIpMFFnnnhnm2Q9ILQlH6IjA7VJXkpW1cCyi6/3HTpmUfx7sz83
12zhySemkcd/Qjcc9R6H3P1pWqxlC4OcomloL1FaLERSTpID8i+fDQv+ydj6U70V95GgaF1BqqIZ
emhWPltlxN4lN9lhYD0Bly8iKdLS8rIUJelAxLeEZin0P0MV4OgLWkCqgxiI61tSQz29J4wLb+gz
3xKyegmPwZpWjPlohPbMqLC41lwm3iybRxvRh3GhdDkElCg6Q4QjBXdx/v+3SJIgt/1q7UOGLY1q
jnHK34tKp4TfrtHkT3WCj7ouIxDCo/W8HsXeyVZ1rVme8ZLGkjD9XXDIALIin9MpW10/zwbzuQNs
D6DUX7dbIjNRDF4mbS+/IeNA5/9RR7T2XC2ovbgxK7VoVRvMoFr+kcbTH7nc4VBIkxrE2IrkVEyk
siQL/N7cQAvItUvrRbjtGGgbuQ2niyf/jm3SwEtGrP63MaOOpGCxmqP7wmI5cQmyiu3Ynk+IlzX/
xF4gTFlUYFjfg4PyzZXkZk4apjcLq8mFHbTq2gsbg5wN6FJSXKNQaLkrZL74Va4I5d/Iyy7OCQOE
bK8eMwXhsBg1Z4/yHfQG6iiyIiON40B6TR/2Bym3785Fl/MegCSY76KdS4JiFmDnUcUODEPbGwCl
7OuC1M4fNPEOQ3ahfW1JMF4REmRreUY1wOyN/kpGqQAqGP6p0k3663bc7hraSlpZC5N3uzFYLie1
7Ot7R5vy16wZRw04NsYnK1NflYgrwR6IJeM+4Wowv63pzAGMLRSz03BrVmJSIWq1SH577YZUzKSO
B42VlFmaR00Bh9bVOM5T/YRL3maR/p7QB8B/CUDkeak1+xAfD5IiCdKcZ01iZSLBDgx3whYC6TqH
X/gY4C0dZnS67xsbaPc8PDP6RiiBGk7/2gDyDpiX6E+dUhLIotzQiC2uMWmB4l7ouMmRxw7uR02W
xEQtu0ozk5sFbRA0kWRHbSt9AMaFhV4iKlaijkB3K5vaRpJoGcd6tGxiJx3QdZK1qN4g8BWuzbnW
Q/yduOgSw1qe9ktB4t3J0ycRPxAIrJ0yO0z/jA46kVD4qUX1eqwkukugnjiDj38NYIVRrv6Rx2wP
QH5OY5F+aRfrnAcTV6CAeHMF7QFuIxdz2+iOe8MiV3Ug3EzOcUNQFNivUOR88QZcR0YIRvToVWkz
N65JPK1RZaAmAob/yV6uxGlvQjYQzj5Hz8nUfV0LseD/CqIh6lm8SLbg8eIHKaQTZ68c67a6Pe4A
SdnBKdkviYhx9nywM2A7BCHsEjA9zggj0PVFjmBQZWM/PyvUhdo8YFqtuDYKxZMhDmwbJ1m8Dmk0
mOvhsp/Kx2IHsYVEmh5YWb6MFNIP1G7/9k3Wr6i4INmFIrBEoEFTESBO0S8nALt1/BORPUxZaENv
cFyiY7uQDKyPuGj5N5vSFFbLmtKPAtFfHsIw9K1lRPf+gK/z9suz4+vg7L2MrOSlrliav2mgFcBw
ImhgGyx68v4Q6w9BUxfG3COaIP9wd5vOIZ1/58VoY1EFjArzfGcaugW2kZf2wBFhOQSSICZI5jyW
Tp6y9PPESALVGT5ruEVQspUDGAv2nnswFQ8ftSmZy4ceg26RUKqRqNSFrrjkZPQr5g3Rnwerq2Eq
vORCXBvAjTcsOVsdyl93Vg+wiDfZ3XepR7frN1T7P72Q9NmLieKkfAcFV9MCUYZOPhl+Y17EMWpX
QqSXcgByYZhHOFZhzzgVBoMsGr8uD7dT+Niflg1chIuU/VhLKCeKjPldfymRLOhvOoW8Nrkh5V0C
ZZIXOE7VeGeA0RE8v+nmvFQWPu3d7wfqchjBgdS5nyRgP6s3b51TR3LHIacB5U8XyUIPjUjMVulR
OdWEVEmwTokf+ixGHcE8Mv1S/L4qRgCmS3yXzNJZd0tTnrSlJR2Ddw8ONAp2uGSsJQsvIztbm9zT
ob/PHtNmFJ63JGHHJUtAot0b4w0xwRSy1mOnKJLnT15FUNde/nrvM1JACrUWg0vvMVc8YAljh0hS
urqTzG7BnpLFKCDltsFumNy9kxVG9UmrpcP+k8AOpSPG2Z9bF84QPiHdMmK0Sm+xFvvWC/27p2QS
9lhkvo8gumhevS+9B5rRbyQZ6aIqmya1ivL3vp0OXOxSynvElk2/ZG818gYFnKeUWKDsuYCcg2h+
gwTMrmgpc8nBGdZH4LHQZ/bhpYfBfZXVCNYm8jc57MNj//Jt56VZxIpRe8ev0aTe4whZOqphp4Ho
c7PKiIlLFxgd5rb1GtIv0HXBJX6cc81Fz5h2YdLHEIeO2ZBP+94g4L2dyt3Rh6w7z4YCPn1bbXTh
nreQzbzfO4Bp3KLb8CXmc+oL9gayJ6Q14X9CENKJVs2mwk0wMjLFp6j3drvyIXRCYuLygDxWvTaY
54/OsbiDTCsXsuRo65otNTyWyTZIB/N9eLrPuY2bKBd/fT5o/8bKzIenaNuP0CCO8unRN6qNyLPW
B07BTbUDbvQLiWEq5BTADyp356HzlgwMdnIVm5ZZLvv+Ptb5e94Y86kWqRpsTOS5rnsNBvjLhd2Y
MOBtHXDaryVH4PStMAZHKmnrsHqkpS9NhGIihkNuiF0Rw9j1mdtJoEca/SgE8HCmkzqRKZ0h6U0Q
xTKXQJCKxcO/ioR072BYiSUZp/wSVwW8TSzB+COlDzYJlpjVndh4xWC8PljsK8pHGyL1TYbs3JgI
Eu1njEa1UaW800ma0ZjoQmUL+XCm/pHcCR4XqXIWLnl5bG2lotRWROew9tjkiiVVcxaxy+/DrX6y
9tOusDUzlvvN6aPYGcW0DIFV5upoShJglUiBo0Fs21p0bZqf82YijtvOFrrDMTeGgo+n44jTwvrd
aI6/NfAV3hM97oRu8rqFDL5bP1fkZBGkKXrfYKw+dyJqMxN2Y4xYj4Cj3xwMKRhky0fvqbDsE6Gz
u4sok4ENpv/TKvu7DeACv2uIIUefvBq5F0nYJXFbDSHEtJ4pYPFsxVTzqXLeRDDCnuTa4VXBh8MG
NcX0zb8qD1iDx+GPbv5acbUp2KaJZbPICYceByBi8FEMbBwqtiy5SoZQusf4QoivGklAoHMF0Qk7
OgKDBePXIBp2Omna022pWwP/52l19hEj0++pjOj1aitp0BMD3fd9Cfs3grGMlpaHCAQUdW+gR+Uv
BtG2oOP0zLe/Za6UUqg8OAmlHaGEBcmhxzjAPxGBglcnGmjudkRtD//58wkSvsWWmimRzDpewCrO
gZPdXSsM2MMi8tFVDrtNNzRioTbUFrcKpE+YpVa6a24oQpcCSBv+jly2rgrDGO4SFPWz3JSBhnR/
umPNpJhRrrS6Ehtp4pLhGamnVvZf737JHQIcJNcFWamq5pkr4DGb/sN3Ca4R5MfOt/Ou+/YwqmHu
FWJDI0IzZ7v+TpCjX1YP88qLGgxqrjOQdYQWSRBznv/rCgaAAKdzDLlNqtnUqvGLA3iHtpnDn9uo
u3yiuUULb4u7x2lTDyNIzjtzGtEtBXz1yMRfP+VtXMhY+WilrEWq3mAUyCiwaRyhs9tUjIqRlrSh
tbU0R6oH5jejQUXO5MtK0PV8zh7ThTUpts4e5gOwJUn65h3tAGO5ukEKl3C9ZiNZwkEojDUARnIa
/DRfgTf/ymLSkbgDwgHMb7P2c6w05h0ldYQau8xjGnnD67v+XLclGtUbRzUbLJF2hqcOoB3P6238
eI4yCtPgaKPw3F69S2qR0gE4FuBL/nv493Xj7rgoadV6o0Cv5NlRHKO23hbO+4IfGMw+5GxkQwKG
yuQtWgaMRFBTpDerVQZuZC0iWnV/zAbGBsiHz9YR3udQ6YUL14OkrTNPW+fV/a00qSBBil33Pz+I
uwtDG98D3+3e6bTOOxVkzQWTwu4B9iqQHVdD38Ofvj30lG5IbsfVV0Yx9k43n1kKRIcvtTVQC6Bx
5Ux+RkPUMhsZCD0uVsoIFB7WbUz+DtqaV3xWnI5adzPWPrrHjJj6U6hj8WK0AhaSuQ+Wz4hHtTgg
hPsBHNdrXCYdPHYp3jkFbMPGjE7nrfaNU6KFhfmsq4WWvdA6yDMyrvg7DyxXApV6PWsN5QOGbe/d
wSBR6f4nmLAQo1OQd8F86rDAGDbkzuOkK8uD4N/JDZkUBsxw3dC2Bsjv5Rh/zgeygtab+EK9g+K0
CAYpFP62xFgTuDOU4VsSgAfG9Ok3Yty1KzgsHdoSOfGwo/e12pdYGQHFn9h5o0k1F6cjb3m/IvIA
QSqETZQdjVY5IVOL0EFKlHIegsNSIOeUtFshCI2wVOA6nZA1BChoZnqnlZsVtc9pZPIJxtO5mKV7
QRhzPElkgP7yhGna7spXrUIrnQPo+ATX+820B4P5jZsErsPU5Y3+o2PTojuEFWj0RkEOJvMf77X8
veOGfnhM9lE6wuRxyi6aESPMwwlR+6dpwnzXlzuWD5KkrC2WJKJ7aCaTjG0nj0ME1k0uSg3MiXEd
vbloD4588ZRAs71+jQx6eYFSrDyJwX5WOp7EBCoBkQpmCt0xouSJT8M2f60Kc6hZUGUZ9JmSRVtu
IpsqgsxpWuYkurb6PJmMiNPOSD7M8Kny/tXaGc90eQMZs3swDGbF3emIdGBT06Ig1AbtOr6UemZ5
KqvVBtdUnONgxW789wo5j9ZgGGWIKNZ7rPq2GtFTGN0pLmAcOAoN0H2GinFWm8CB/+QDdL25+tOC
4BL4MyngtTTbKSkgdZjPLYdLXBWHqz0d0/ON+RpsYYEOfjdj8jAq4quG6zxembnZFQwfR7kDASFZ
NE1zxNKiFAAbA+RgtfOhKLXII4ZRliYS7JV7uJVUadZ16w+WddoxWan3plFkkzYPffe+YAQ0haMd
VRueu6tV48DMn6cl91ee6SlCEFXtFJ9uDHraHQlYMCmc0cBsZN3QuvL9V07rinFu4dlkPY+yItXe
ArPTOJ+dGgoZYZl0b4Rv5VdPslPy7tiFQz9ukXPoxerlt8kTGRdrJq2Agvrk56PBvyMpR5FM3PC9
xkJ9ESoKKZcx8deCeYktWUi3eyGExARHS6EN47e1qygQ6CEkOAHILep8uDexfWt6KAA8tW+J7af5
gmc6J2yxpA8QPX1VDtoA5i2t/1Xj7eOSZptsBAe9Aai+83jxOLazeWzi+TBd6jiZJcpp8UoVLZTd
sreepE7QDWgWJjN7zPkgCmpKvnj3gWSSRrdCdJzuMmXDSwuJdSimffwzZ0snWZJltcjCldyNp9n4
BtdaRZIyu7hx3fFjo3R/HKByrpJnTExAU6UP0u+wI7z+kc48U9aSYHXLM+I0qkA27QMm4H1tjfD5
b1jjWHCMVHCrc78fzACPNhLRrU/etvSSQGQ3W3EZuOvcJqgt2wjjYMK7H/LI/Bl/nB1guGFUan3F
nTpKKN7MBFOLSla6XTGcrr6xXhUB/jMU43x0XZEDIDxBGZMXc9b9K+ESerkcICcnWip7JAZYmCBC
vhFqeElTmJjqkJGQV2r2vcuEytb6jSKE2o+jkr5h4W5aFBhzZlM+9xWwyb24T/kJsklg5rzNAu0B
P0IxFa/qJYuF2L18aTXO5H2gAMO6jjQOQXBtkn/c03Gqoej/mj/8blbUTHGMOL81JeKzDFQ1nRiJ
QVQgAfo3cXI9mCPSxEV9dzCzvYmO2nx+aEzjDW491hSA/ddwSOlPojEBU6vUR3e7tygxLaup7sAk
1KkR6Ji+pBBT8UQVB8uptDyA8A+nRkLSPDmjmlOs1jrLBKbZrZP10BXfqUU5NEQPEzyCkDdJJpya
crrI33EabZA+b3DQjikJ2xAmNDzB5J1wwrz6XDTMmNIA2uCA/ZwcuhDoVnp9QpxOUofN2l3EFI5j
K6B2l7KqE4aw3nUBZ0jQTj/ACPevFsWUG1xB2VtPtRl49iswSWxq4ksWNIkIuDqKcFkTmasLXSab
Ydn/To9yPvPdl7vk48e7qCelRsKllIBRdgJF5CsNjrkJh1zXJQexFEQzWSAPKrroQHbrYxgxNeGP
S6QWbOuVNFY+stmyeRkeMBo92+5/wBq6sMmZsGl7iJ/3kBuzMLS6Nvk4aSugdwh3iFlAd5vFV4uf
VVfKnhS+R9fL8q/Lb/P8o5SJCnoit2xwKwbyTIpMxG0AdFFzH/BjUSC/pP0mglu+WOnsE0Q8osv0
aTjDwHfYyaQxHj19oMj+IM9k+0pOPxKlOaDxtsoEjZmnSLruBLZ8BEAvUHRCM6wWLjyvJe1srhOY
xJEXsEZX158oAxGaY8FjXycV5VfpOSxmPdZkXbCH0PxP8QhmcqzrzB5oyl8A9OYDDmV4QHD8sbdp
hqLrBxpyC1z1+kUbpc7HfMr6znkCjxtfWmxa39+APbkSYCtiSrsDncwzA0IDQO2oSZmrGZnPpZpE
al9wyKlwK4Cq5HREYdtyUeFT3qW+0FHngJ3ERF+EO/CErGNxHKbSOQEV0ssm1Fqj88qsGblDcUXc
Fjfv9QI+6FGKUQGQbfp0xJ8gLZniGJy9nFM+iAC69EM1gcwWGbjp5fUoTeqbpWWWGECx7loZ84+r
Asnb4lxrlt36SFiItEpb/WuQknJpSlyjiRya3Rg0VjIhnDvk06WlV8qtjAi0f0TdL7+71ahhr9G6
xosWBiP7ZErvyQcLlv+wUDv9RWNt8nyiqsNszstxI3nVBJOsXYwCPewI4UIwOVFsQQwp7AzvwSPa
qAC6u2nc7lcjilShjDlv2gOdtvLcGigYJB8fJW/irsp5FRGzxUOYH2cuaumT3p3/aGlEWzMItOSf
j1riYtdHplhi/OMMiMb+yCaDOyxrVDktP0jSfONwM4OgfnWYrMQyAhJVymWG7N53ZbTxopvXBQYs
9WUDUVN+HbbBdd0bNIVa8BqL3eiUeoGRkLC0zZYL75RR5XfVg9kH+eFzrCUxtlfK0vIYtxqJWdgV
cwSWhcyDTONlwJtznJ8osxIxhT59BgRvJSvEoXbuk9QeurQzZO/tpOOPrXu8yXCfZbjzoFTIxf26
DzAIW9kpaGui15ADUuacCFVSsCcPajP77K2o8KwrpflUAr5BFDRWBYODYDtokagspPS8FaSMzVjo
tQqaWoQ5coGiGrrIWTg6xmFfv7SoDX4UvzXP7rsyDfrPyZ3bb4M4PjHcAThckVAtDKgQ+vxyooiV
UZJJLrdLTudZcN2cYBNbS1UGoRiRwhoGjsEoRy677W0T6ddXn5+6vF2EGp2wNdLBrPk+3IuK5OXc
cxH15PAFmcSVPAAX1fzTH2o5vRWQ/zJY22R7Oagtfh84qXZswXyI25IHSf7V2h5kOYeOLdxOjpDe
YQih5qvI4budnHq66rX7z3Frt1ekRhJ6eAkziQAex0VZm0DOclZQO1Epr8xuzsoAw4LuNGHukKSq
cv4u2in7vdNFf1+cpxUl2NL/7UdvGLz74P53NAD5ABiGTIwTS/CIfJ08h3v9iGiPVJS8H4IkNGwn
Z6nCqAWIFMMIlL1odGvuEUEyFIt1T6PU6wka8dIpiroChIre3gEQJdG2Zq7GiQ90MrL2hhs33/qb
Q/30/dFFodkeOF+S+Z6+K1FPxNissvmxGJRUilbhdzTfwxs6oemVSQ2mSlupYhkgeBa6a+4v6t9a
RGvfoccc4rWnQb+TWTtrCXYm4zZ9bGNjmxwjQRkyJ1B7khNQ19Ilbs1Vv8/mvt8s1gLk/Ms4j9W9
Ta1HPPsUWr4FMQuVtpKIf6ik0bvdg1brqG0kXXxcK7VD7KYAaezlpeRD/pfuRMgWEMNNuML8VJML
s5JvzcTACP4HfbNIxMP6JOLyorGh1Asm2v4rsXVt/egDeNRbUGf8/MM2LU5tSOyteVRgzrXXaNsV
3hKKgxGUte1BkAQSFYppqR0nFzYn8ZcSoi/TzG5VD1441+7bLe0loeI9Mte1l0hQoaYnZSX7sclb
lfHFWL424DImis8ue3Gs/0lyZ+ZiKV/A2tQ/XPCCehmfgdYPKxn7my6hXOIciiRcV8x76nC+hz4Q
thkvHi4wL75CdxuFfWxBOuHBr3yBRHZyZhtsHYUFmbt3y8AcD69mKzlOFpfkhtWWJUUQeBQzOWGW
jxy/mLE2JRa9Emo8+6D7quZNSDQlTYyGNK9V34uz8h9CRMDqCpDiCIdTNgSJjQFvaLQ6yJV3R99B
m2Q8FgRDItq1uzJfwZNEN5hTM7G8mi+DUPB9qlAw6alWP/zOzjZgQOA3U4iP9BEvJGjYwGnc5Kwp
flh2RS8N0VNGvnyQac8gQLeCegotSJRD1Rv47HEQxtTlFzDdktP2yeIDtgSCTHfwNZ66G1kcFqDT
caxwYVI96hShkLXHNB+FijjaJ0x5IaQ5eh60O0/9Le0fKC5oHSBHMJ3DS1uL+DM5hgjZhCPDAHu3
Qq/ezQ28odxGAicinnQ35RSHakkDq7UU+W10trTrOd1IwyteBXVfSCDkVDuF8dcOqljKJu/vf7K8
KbQ8cxMEZQZKUoWxPB6uQZrkk7tyfy9KNkiO7AzclZWas+IHp//wAZntQ/MPw8TY1JgN1GrkAmDf
GraDXFl3Etua+oKt0x9zH3VeixCdydz0XjYFbmkwWz/nJsJOfheGKYdzGg4QLUoMpYTBb9mQCBss
ptec8naUa6pvKHhwsIJs1+1l2bXt8M+QMUiBlFcdDVVWwdrdTrbS8AesmMvuZ2Lzn7oco3beUZ31
Dx8MZAfa3TY+IVHhC7S/kRaWe4qaUwfg/VK8sHobMggpaFDwhUfJLikzbnpSI3bZPhrweleZJGt7
4tPOcfiXoLp7ZO/aq8NyMWxISBXgUapFNtSbQ1DoONnxNE8ieOoScYulRHymQPTuYIggZ467KpW0
4ZD/13KzBWYRyZoNPT+HGa7cqci9VH5vlKrcyfmaWoMhviI0q890NMisYgFXCQXH92enD6WlnCZ2
ifFa5bCrvJMCyjtyY76B8XkQQnB3S4U5sVRwOkMVvGKntyXuxbpOeA2vCY7fb38evShrM1fHR9Kc
zcxsnCzdfP4mP3GbkLoQlmKcrmefUDo5hkuY40XS3/mlTWlx/boi/d5F0+MAAmqAWRDoivR3/102
QEeKxDfGJqwSlmbu9L1XsqRcWZpzBseLYWpb4qAsDDVFxHXHrLbEriCayrr+XXdJfonG3zFyy2Ea
othykACMVkrhbkNArV1PEvMXZAfp0l8dAYRACFNhA4iWtbPhBU6PeLS3livzQOqOcb+HSGdOThD2
NuaD6HEMJFBTa8QNJxmia3B1932clGY79YUqdHYZQMa11VQFux5pumo1XCb12R8sAkGYgLWQ1EaT
C2IeMAcI+UDanJ9PXm2LSrgTwsNoVHmuOlechmecfULekw6BNEUdUkHsVlSTYw6Hq/n1gI/kVAJd
rSB+7csqPmUMApDrUOVzInhmbZqwiQtskoWFbFCMexnEVkB+beEJSTZhOC84rXzioWICbE2WxxIa
8stOI41ecvX/CMgj+2ZUnFULWQAK7dIaB9A8u23wMcWTcjWwjuP49kJbs/DHzwRGy/I+n90xJlOA
btDcy4ej1X2dQTc5BZ2ew9VbEWxXdpc8lm7sLy6daNc/VyIRxO2aJ7eCNKPiHOqKMzoDEjDjsXmq
bU/hvhQPyJd3v38+Uih/ol6OsImr2tpDQN1mFlnepVIWPF1M7i8QHzQ43qKH8bJlBzLiq1JKPjhu
CbUMelL+ApenqA7UEpk5C4sxnVhonG1q2pCZEDx+IWMR7ov7AMFrgA/Rgi3OJ5vMReNWNuvf6sQC
QaZXf5bewuv9QsrKt8TUs22tWESusuOiOdyePJTuwR/xuWlIJfI3/zRqNPb+3jiJqN+9MmdcpEdm
DtWSkSJLeCKwKNnuRQEAo7pz96svx59GT0A/HE96kPNXRZVfvHJkzsXFCd2XHra8Wel9lW6CH0M/
SLrnHJJkZG5or+MMPHiqhJ7kOo9ETI2tVRuFgEemtoUiBvwVh0vOUKEHXkEkYWsNgDen41Aa1rSG
ORJeEr6ALp/Gpsxqlk9U1e/XSH9OkdsMie73/H3gTr/6fOIbhpt7nrpWh3XxHbyV2GJmhfHRcpll
jjnPJSmNjS6sifxKcN72+reH9x8YpFwMPDd0J4iGhBVZhBejukLOdZ+y1a7b9L6RQ5c9JCPQrCBo
IU8uOPWHUoFeH6jYqRYYNKhRire8HrzNvzO5iH5kjmKcw3j4UlLdUYuUCZM6byMY6cCT08uD7n4Z
JNphFt6OBzV1cAdWFZmemBvbxVwsrcfayM2k6SfF0upeQzuu4qA5InROh8C/+OItfRUZuV3dw8wq
NJoDoFzt4+2tMSKUpwvm49WhOO1mOzuBG0FJt2qYaTxEXuLs/lSRT1fPLHDGLzvEiYe0ZYOiwRfq
BvdqxNVcFAzBgZy2rCetOMvDfdiDnwTHOFRn1fJujJPrTP77gYHJt/NoTBblKYVPT029xdUZkOhN
2doBZg1C0l+xs4dOxgzfDvi5UZsnGmNJRHq1uuwEQvlJZ6fzpJHpx6dN5/hy71pt5OPFAFQG1Gd/
rm/Ttu+Z0p/euqWHIhkhXy2auJqT6ZwVXH+hHnYTEknQ7Xy7SnmIYuFclvYjVsRYRNMcuOtjLUxb
qiPp0M68n+WVxEOLF6Pxij8u3pXuG87y29eRB/V1jr2x8kCJpiPPjvXQvgKQm3rMGzhWXDV3Fa5F
PYbMVxUJH6AMW02B0Q+CdIA3LG/tt6GS2yivNLVNza+ZhSQ6u/UPKV973uUkIiDfuiiQU2ef5rHl
H70urXr3lH5SK+Y/KZoYLOvxz1tmm0EELQPyegB1MPMH6I72QVqmIQepxhTgulXWrAmGodpgKVvT
9l0FMmgmu6zc3ycODNwyrmuGvQ0PeqUhawgwvO5OOjAGQYJqx6TAGJamgo362GrJgEoiduW33yYd
WI9hoBg0DqV8hFsQ7yWyvj1syFqPSOpYDyDTwk2Gy7ll75VnWKgkvRqTQ2LADdHH/yuPZ2JTNiUr
Qww2Q+JdnD0923MUIXwittkVx2h6/Waga8erm9vOq1vW8rPZTpD6jRgz1ERmYpNqxk9tlgnVdugf
vQKsiwsAtcM/r53elcwO9XnW84c41J9W4KDFqkMlj/O03sJJjSxX6kuqWSG82fqb88RqcmofC4jr
F7B0b98hl0TM8K2kDplzX7bJT8vC6CQlt4XoMzjf7ymLsFv6fNzOrqPK8/1Bf1WB0PKBi8BzBAhU
FJi1HKAarqWxZu+fSQQ0YQ3CPbtbGPTQn6ESzuNDAZcpYyBzKnGl+7lx1UlWaigSnJVArsfy6PaL
8JtFPHhj6FNcAjCp+bxp+9/4Wyi/S5sKsODxZj+xr5gkK/xOF9hEItb/SAoM4C84AlODUQ2DdVTm
FYgZDTB56pM0WqyRGClETJgfk3q8W+kN0JAtiOC6jzdM04br9XZefl7FOzSFpv7S1gbPDIM2cTRJ
+KwHAQKdSSa0fdq0BvIaB2Y5tjd9uIdisZZcHeQ/sP7b+Uc2wAlPXn3xatHqr80yHQu0x1Ra3COE
etnsZr+Gqzrh5lbaRsRGlKRT7/ZrRh/lhpNmQsG4ZDtOdCPJo56HXMjVXwANeo1LV6a51xEvuMyc
uuUT9Y4CVjzZIoS9+tqtVAmciikw88WFxHtu/FO5DP0iGytGb9KO/Qx/euB5FA0yrKCFFOHr8cMi
2hGRmNWUce+nZeqSgCod9rToVQsYljPpaJ0wUcNTHaX5/wH+XMIAUZDiM6NxRIsfe5WLMkBoch/s
hRuxQalisG52SGXmnXI6oee9RWBhiIW65R2gvIlS5E5s7Cpjxnp9tmjXPSfWIxWPqsxLwstWhuBZ
GVMw+AG6Pe76ZeYvnAar2nGhr3s43h5ylknqIgof0dUE8zFNyDfUevQ1WFegcD0xy8Hj07r3RZTX
/Cw/nWP0oJ3XIKHmWNJ0MaSUt/j9XSjVX7FMxSQgtipV8HT6xpO/eyNOAA4TD0Z6irOPOfEvaZE2
m4nL43n5oCzuKpC0owA0h5RJfUG60DR7nPVcgDlFud7FadrkTDjat58CJ3BABI3nrdmoEDxKvcKz
aPBD1ILtSJVnzxDaMOeIZzYhN89nro+eFn8k/wlZ9Qk0of7V9ly190E0zTvpA73xPgLhd0FXNWFB
aA9PlQogMl6mi/OWKOyH+BziyWfDSNVKgYlFtkauzZ3wOCFDPC0idTKme+BQ5Pqun6kkEdzUrJmo
3KvSbTSKO+7caoCnTwkdHbHF/GYhxs4W5BIJ14D06SHfb9qiB7GKel/m4kHG6lfRTuLwiRoxirIF
ulZBtzMvDnmlrI2jZwzzPdrjYM1DtuTpUxu4EYTWpNwwqMXiKxJ+bOPvl2KXSM5oTLVWah0lxBWL
ej7Ev43fc9cKWs3uekKTJRf23L6JQ22Amw0pCGGm34ktlC0ujiLZWYigRAfYBqKklfNkDmbMeWFS
LIQuCF13hX5P3tEQ+/PNAzCtK1Ehsn1BSULb/A1NEYLvo56uwUTMLiGbcl5HYClaZLRnxhsHYFAe
GY4POafA6uBvnZeNjWlTI5lCmlIb5Cf7Y5q2YC8FAFDRVw7IWhaWQjZ4wXZy216PyucvGYxS1r+x
VR1rmthTTVOg4JYk+4LDQtLLV8BD/W8uprWpg1ba/QokSPMHS89xXWSNDEeERXCQkojOYtyguve9
W+cekdY6dpF67pa3p8k0dGHlresWyI5CY1Qi9LSJnvO7f6cmI7iSfiXHa56fv00OGSAP5Qdrt33u
8chXKmr6GfIzL0URY5FiIBsH2C2MEuCIPcSge93xzktOiut7yD0KGkW1XVjU5JA4BocMw8/hN5On
5YimX6s9r7Ts3+HjtcbzwzRp8LM6cK5uHstrVKj0XrrYt9XvSGOUFQeT0dwRx79sUxnBtvuQ4gMA
mC5ZVj9Ndt3/aUiZlLgfccffMtWYYnSd2VuqC44W6zRuhNkcnSJFO6+hcOoHwo3hqoK4HWLfrGSm
+xsxqtvFV2MuV176VxsrCed2V5lCR7mcZA9hM16xciVYyn3AEogvWxF/ECYJXBj2JKUyiIOEms6h
1s39gp+OxMzNzPqReaOuD65fn5V0rtgfvcbty+V0rZ7EI831s7rP1iVC7cR9LhWQf7Pa8/FfQrib
lvkGJey7JwYJ03Osp0xCKPKBZj/5fn0qWl1DYDSi0zRv3Opk9ux1G0YctIlz3OY7DTW03O73yFwn
N6at+YH2BpDOtTxKh0eV2bxEZq+IzRKGCLr4b9FTbmk9D1Ufq5UGJXfrc11KiqV8kX/KgJCY7EpH
WWJw6Zowf9UuvMlezeGX8XMSF/Ty58IdPTwLziU+77Kr37zk3lOx+QcQd7gx2bgDCu9itDPrn1dY
viXISFQJxTFPsqWG+5n14uQujIEwjZTwyzINdtoBBufZHA6OwKfjTm3uJ/87RkE/2x3MsjEO5ZtG
d1RJM/y97if0Ypao6R4t1nxykI/yoBr4REoeSXS8g16ojyRLM5z2tQOnql1uyhJ8BmCnnb0elo20
ejZpb6QqJdhMLUhIpB6S9FSSN4xTqmvwtPEAEYY+eUyJvO/HSe15pTHr4REkOOrh5KSLi/u2ATin
cBrOXGf/6h/0Kymdp4a5MGnSHCDZylG6D581NFfMJaRWEZ/IJvwSvgP99eWZyUCMlxI2rJ5XjTXa
amqVzqiPn5QoSwEoKoLgrlaRZT3iYv3YmA90oxjCskfe+yOu9bML8umKDcgmSOwvrlvyfMFhl/62
1e7zXMx+bRkQunLPV3kMZ0+8Ge75INdA/PXSTaAcgpdKKX8SgClvJVshtoFAOoUv/QSiRjsIv+4B
NqGGRsFKBZSiUKRHNatxvq0l9s3urI1yczKv7YpRv6RfPNDnzF8F00VQDFxX24tpHZ7EXWreSDFo
7qYPCGCH9ZEgrP42X+QXOdYZKfkdewyUAV0RwEYoESQ4gFUfARKK5+bKsAfj3IE4Ss75vVK4hCnn
UP93BMLUZPCefJX8qrWNikD13CJ4e2pGm1yddya/80JKqErACtriv+5HukB1Xn+Tf0w/3SR88mzX
4dO/mlsELOYnByOloUL4B0pjFYGuWFbGhp+NljFI77+kdrbTLWC/yYaCs+7AmVNqUeFfdRLCqW7o
gRcbLQSb8+RpRp2a53uKcw3T8bWsGSoDBEdmOYV/XQ6miMDspIf0Ut0MbYaW7S79dS3Lm+lt+GP1
mMJ4tlyTK9b2Eju+Fot653Ebx92Tv1kKwnOYhaoEwR6VksQzVa0Kyt5hi1hFfT9tu9t8n6/dFXjB
scwehBNNmqymUoHK9kRnpKT3QS48rNGV6MJu+UULTVGco4OnrfWhJjpnyAaKMbWuSqDlTjuaxJ58
Lc/O1HJSW8kDMSUZxBoe93Ur9IVNZ+vae+eidXXszpkjXFDVNrDICQgiuBd+dMKACVdprohmDPeP
ylNllNvuAI/qcZC89h3wkZjub27JMMaioPrs5Mdh7inSkUDwCDCn2Qtn9LdJLn2NyNa997b0EGxN
LuONkp91Kr61v/kYoSmGDU5Q6piREH4HOp+dfK2mTmjcHuYk7/nGzTnvMTVTzMKToXmoL6kl5cXg
+M1FcK6d9TISYw6ijyVpNgFTr8dSQlBTic+BhDqvzIIBtCXdEfbAh2AMq1ms0wnIKKX5oHAkJ4sL
W912RN8ZxZ5ZInzaiDCetL71DNufWXt2S+otGcNgwyoGiDWdty9GXIsT2WHwUXdYrJ2AuxEmKrAb
xjYMS3ptJ3aC0CH993WFLqT5nK0Q7Qob7j8iPcy2zPxWnPa/S/ngFnSBLZt4L2nlgzH3MJWAtMCP
GGj2gRHVkf4BXNUHdWdfWTFTaAhxHNHpWUyzNu3Ve1urT6D2d93Dq3fFYKqQzqCR1cb0Ebi9UxQm
nTIz9SZTTLZAf4dX7NYirb61LMVjpp9eKS1pw9Fnp51e8COL3wxmQPfJbnIfzb04+LMXOxoaWRbM
XnGIdSDB2gqnMQjh7jgf1gg2hr2xxf2ogje9oEPwrwHcDWMd58fLIlo35aQCGVA1cK0grB5bVgk1
DqdRqL6pfgif8aWZt/eq2HooGpZe7oKZstzoNRLJG2gsaOXGjJRxdDTGC+3aFgHB3yRUT/2+9rYT
zBt/yPBr0dXjGDRd6LZPTiL5pGj8G8L6Si7YVGOM5Is/tbiX40JuEJpFYU4R6uypJjbcyrpEeNag
SJq2RUXCxYoKnHR4wlR8LFKaGFNEkrjxuZUnqrP/0EaRVDFrKUoMCoS9G/OiGtQonLM3YM9fMAoa
WjiGg75lHEgM1ucNgsHQbelAsO7N01n0LDQW06BJFaQl/przSR6D7NjAfVMAG+ZyAmsD/1ik+Phy
Tggv88zwJnMM0SldjlfRvUeEcprLvowH4J4bKKF1cC6xzaPo1z+AkDBPRNfAz97Yi6DRH4hxMdfg
U9jZ8oQa4EY72JD7g3l328Hm/dRxhqzau4nK1H0qssfN9HadKUrFhYmVzqdxPV1QBVy8I8p9POua
YBkFm8RhhXWowbKO7PQWyp6Pkj/r/hsIOLAsgtXnm1fXxht3BF450Ng+pqClPtsmyO9SiZ3SlxqI
PT4vK1hYaxke0z5SLfsPNeL3z+2SyQ5ml2rKulWWeQRP2Nwf9gOygYAQ8AJBjeLxtZlOTEURUR29
iCAhzpSnKitXwCkpzgze2X8xW2xOmqTLSZpBE0s6g0FvMilV3I3o1CL3RX25WFRZ/eCCUymPWGy7
PeYKjMY/qGObVHH/Okz9Z0MCgP9tOM8DhBPWOMjJTdgBymk6OqaYb28Gx3zIH/gdpjtl0CWosWRm
FRBVJTmMp2bEBeGWEgBxG3c52+FWiO2eoNMvyFIC8opHAAWzVLdwJFvVf7uPRnmWj2vfPdOk1dM1
AHKWlhm13rYiAjc/uGmi8kt8op1kG5DM2cBJnLvQklUe1Tj77BQK7gtzQAmD8UqSr/6IUG+5/PW1
7xXy9jaoAoEFfrkGgrLnlG+7MbBaMNh0HGAUNBVDWUjwOgFvJpGCCnKBdUidwTtN2isThz7YaOtl
K3f2eYdfzqvcU7eIrYYCr83c3PXJmtTKBAyDrn4e7B/IF0Yt8Ef51BmIirzao+Og2+7+msP2HJNr
egCxmoufkS5+8phCVljxqkNZY52uGdgzerrGPcQdNPVZNezh6n8sidDHsesw+2RijPpSviJA2yap
V5trO8zcOGfRwj88d66KPwaPBGnFZoE/ZKSFRfyVVROyPORf8PMDFbLmx17r5MViKfvCrIDWXQSp
tYXuSoFs8H/okT/JbKpWQHsNMkwz4wOKXQ2PYesSq5XZsZwGonpl9Bo9q2T/xopw+M3tB9mnhhnv
QOTPkKsh4gVOrAGFygka4R/pN8uJ2Q02e2/nOYDkkeSFxrC2imGRCztBVYKawuryJwh1QOSaz0+P
sLSB2kMItv9+iopbL28EFudrC15Y/jACEVes0Bz/eJXMrSQHrNbGLXsRdPdLNhSyLRYIn+xRcdVg
+irk0vWUQhoR3KT972nTML8b52e+/ubg86J8o+ExlAl5KGk+J0tj3iVZU/YWCGBThNexjbbabIYQ
SsRF+Tcpf2O+h2Vaau5g97euBVXXkzvQZ6DaybCvh4BbwDOF6nGnuzlgoFf1oBcylx1RnkwJCtM+
nCJzFPyyamFAUwOFDrzys1+8M24RWfSq8USDUJsHZyMtoQhmmFTFfkpUtoBPScSLjl48G8MY1Hrl
dySATCj8+IweZeBjqBn4K0yaDIP6IzatbUphTxRQpNGIiSK00OdTpztgzxHMi54L3xJmtgVlo+i7
G6pCBLdS7OlorH7qoU1UBdLKo+iv1NNBesEhugXVzj5kJpFbv2DGDi1u2TcaBh6G6iDDRxkyCpRE
ZBCE4TSEoss3wnGD0zhXy1EPLUEs3kkKvFNw/wZJURru1yUPwZiXiYOWkJfeid5JSe3cQUO06AIz
U+Wy2tGYDRTRyKzso147rcmH2aF3SGCgX2aAwQu6cZzFy6kKJpWvQkVih559n7f5r1ra6FrPZ/nY
S2RlJnFAzZHvIkLMPCoaoQSCA/v3IDXvFByIc3HupbkxRr4mGNjzhAcvSvq/a2sHZRm/irmrSGMw
wgq4lrY+oCpd+qITCeGPRh6liRZmJr7p/cRtZuZEgEOy3TCMVPEuT7C6jZbtNc3k/UHblgz33a1J
+cHZpT7E/c2MoS5mxbhSlxjAZcgdEEJULGpvJ9SBzKT2YabDaL2srM51Vd4hsLw2h2hNyZ2pEEvT
mLCawpxArX6ZpiibBzBjk+B0Npu2gjzIwbT1hRr2F/sOiEHz/+hDd+0s/LWR2gUkejZ7wLVsMLlH
iBfBRxeXQpegptMSGBidtwHRBTHnEapUvhFwhdjEwylnn5Kc/eQrzaJplJ+Q46xyvOovJjvsAcQm
YLcmjlFJrsDk7CsVOpzyIN8uxj5c4jX1FkvKiXoXBSLYrEZyZnE/l4wBiOBUjni9Gw8EHabqyLw1
6xlUTBvK/2uTtvDxyFG9ky+ct0oj1kV+eHhbeQG2Y8i6TQ9z0HpIgTQ7pB2KOuROuof76nkU94Fc
rnZWYcBg1+Z0u725MSp3BI3yRPcIDfaNI2hNeI9W8cWQq5rDW0q70vaQ89aww+vS8Bee9RNSqlGo
28ViD63GYK5Z6oi59jKJvBq860q8WbFAy8rDYf+xjG5b5pmkcLw8RYzb2p+iff8BHb/AlXz8x9gd
klXlBM/NZh95tiY7RY8Ca07yhBqJAozh8Vr2XjPqiivIrYJIfMB+iVwO7tdFZOm3ILc+qRZ7WxL2
epa9QozKmOSw+h9Yiijbl+wQh/ythMWr37uhNrfXeMl4CTja/0wqoEr0AigceuyYeBcjOAr30vPm
GZvESiRC9O5wo8qRwqA4x6OCAc1t+YasIlDYeeOVuvL8VqNWfub05J+EXprUiuQVl8qgaHYnoaPA
eWPlFZZixRkYw/5s9Xyyn+kUS/eNSPNYhe/zjyy5MMYBqc46zFylgG/Tv7Esc2bP37K10qgVgElj
Ikd9vYds3e5k62qcHmvl7v/68FzX6Gbe+4662UKjjRB6679L4/2MygUcBdkdFWBdd/bWBQte9ChI
yK7LB/iVdMh8OtAmHpfy6wwhbw9+ld0VZPdqN+3BcHqaA1HL/cqyk6J5+qCRacr5XGZRv2kHWERt
Reqc3tnh+QftV4CdZeqIh+sTI9EdZpfE3xZpeV4xoA5tW/a8Gnva2vBTrVPCsVsd3UEYaC7O7GeM
BF1J9x9l5BdmnYZ3hnuZn3cDcvn8JH0jX9Nv59q9PMx4GY6+bbu5NTmppHNgxYWEM7jHsiLGdHep
wG+XiWqm+5J3ranDGCS/ZK8U/pAOzMcaDm+PoYcVPcmiAkMZLIp/niLvHAv95P3gt+YTxuY++ePs
jewlpuVkHKFYuzkeUW6l0rlIc072NB4dDQYFc3o0u+WpH8yst8TopIp+IPuxl6frzo/2oB2iA266
yzAIl6j25sw9S1GUo/byvgO9EHPhn2bRJRMz6oR6cNPLa9DCBaz8/DsnnHIsAV4h6S9mag43RwHY
azQEEmLmouTf6DOjLqbfVFgneGFrFJPTO+gsm+CaxhN7agG6HCDoRisg4/lolTTNS/nvU4OteLBi
H8AejxO49EYwpEj/HCoqf0n9W7z4V47L+nZFXSsFdvzSJ/lPzyHNS12CFnM4expCNxvQ6GmecfyY
ZqBqVg4VfQYru9eLGdgQvLG3Uq9gyQrfHuifHsmG3HVbD139BaT+io1XzKjUt2xzfYJ9Hcf9wqMX
4MObVDTZSADMgpO+owpeRdU+fuMk+Tj1zHkLhuBk297c339gTl4fG59ufhSTI+bPBuDIELeLrsM8
aGUGuQORtrHuwrSR9uatD9o1gfJRVR1ALYEIGZc4uc6D22ztCZgd1q7scCwU8fZD53SkB3dqZ6aL
8kCMEH6f1IFsyuhcuDyUocXnZwu8D+sifROqtyGewaGn4EjCZSEUhQbnkc8wytfeQCoNHSJS0XQN
IdK4k88N04zluWA6sExu/VYstGo41Ds6r/tsP6lNQk4anJBNXps3uJ99ck26gfwGwQnHFdlBTcMY
04KxGgZwN3MKCGoo3ilVq2v/Myr22Cfydc8Uvrw27tEbg1fxLl6Yug+ouZ5Pe6SZMvTf5rtCJiSb
4FHgbI+2Ny1g7cG6QmSPGib/KurGBC4URqGHawbpIeYueJtWU10783O68jqR0vVRcFQZ28OxRQ0v
KYv+C/iD7Z9br70DIplfAmC1+ysDN6UOFzNKsf3/FvGeY53hK7/LOqc/VQOzh8y+hDbo/QME3MbB
RcTQDbvoivTFd9NuOz0AwS2rCjPjePWsGbWL4aOUSExiShUnZB4qP/A8XAE6pAgACAK0jtNxcoNY
K+CKzsxh1HgSjA57C0HmFoLh6fZL9pfum7DfVtG164Ict6BOpx1MCjkkRYKfIWDg/qJ3Zs6tBz1E
bkCqzzdHMgHRUmAs2cIcVINymjGd4+cZyKxgUN1y55T+G++fCGDcE4dVEYcUSQE546g17JP4ZhCx
pE437hKUi7wwhNiSw1mKKmo2N+GJUYV5jDUo5nrnYUG1OHebw047s56K7qDbMFlK+hwYXVsoEGlh
fWM31tBY1qmqGumiXOxqm/tXAb0VV67xZYijFc0YQQHJqv9dPwL9GKdTfqqBs7bd+MBYdqlkkMBO
0ZsYhV8njWRjTR1d/18vTwRq/WihRlXas5J4Qc86TvAmAsPxdXs+lvTKMTR73bLHhCG2wWkrSM5I
6FOLbTVpBetn1AU/xZlmbvG5/TNd34x447nHS3Yvj8K64zutfX+PX85l2XeRY6AvpEdx3D6Rc4On
j52HPrIBXFXpUQxaV+BIeD/HMI6xde7gduWr3R8qNA4iAoComflP91mlFDaNxRksOZXQE4aRUzQz
Pfde2MgyndIVTy+oCFnYd5zpRuNjGKnG2htJcYjAYULU4mzJLGzswLR3IQGyzVdnn9aLoyPyORVn
ywmGMcHmThy9CuMvXFZw1TR7Lu3dbTAt45IahOPKbHBeyiayI6ZIrJ4o3XXz67LiySV9QhIoxadW
BBlli5VuesmNcH48TzIF2IjC7zIeE0q2G3LqJaOoBiD4+Dsik83Ov4FVGcFaAT3Cu2EvJoIn+G/1
zt6Efl5X6LjFxZWrpVzOmw3rcf1ODeiRORwhiOOSB7yqOdeNfM15su5kbONn2vvYKlPiRP+A4Ziw
g3WDOI1EnZQtgaYykbpnDeOQGumOEwWKfEsnGxktjezqra/ymIEI8Ap3nmlu2CXROIGpstQYijZj
JzK+cYEwNvngP5teVbayZgVYaZNd+HFdcDrmMD47Pr3RAEHqC9xFb0FHWAj0dPZ+IGPGyUKhvGh1
VpsOmtAlspeGuwjTBAVXOe8TzHbS6Ig/bx8l1PMgu+ELVWCRsSIFI/j/ZLJIDt2xOqrbii2UEXxd
V0Rq689pETpklEPFCxb407kdWfzfNpOnrlBjbwFElai/LtNC0RmUfQPrCghl7RrzA1Jwmy8uFoFp
tOelIKF3s5U1yUiEYoV4qagXBxqSg+gPf5HrDJioa6tE8Zc5YbRdlUr6hCUDL2zGHc1CelC5wS9u
Zo/hY45m4hRO4kIXuAgzEN1lfUdINIdB85sQFFWvwyp0WPtfoPAduVLW8n6zPTQW9nv9ngiFvFTG
3tFz7Gq6Mls2RC54jNOLQMYLtEB/DbpswlMM6RyGAI5yy/+1SyI661OqBgIJ1oCa1GRCs4I9kWC/
Xzwq3sjK62qPBQvq5rIOhzlSF0a4Tpief3TUSkez/vqRyg9+J5dWEBP+WW0hNi1xIHITdjcu9eQm
NDIrqqsW2JYzdoSS/31LPYotHOqpe4JE3Uq0DK5m2iTX5EVkBsdAuMsrr7cuV3Wn31CGNtT+DSdT
Hstmz8IgfGR4gZkki/WkkVjpiDrEyoJ6IV9huAg8YfoJewwP71zIYhOTViQlvWV4GZ6YQp3eihaE
QvNktPJTluXDGuvdQVP1rIy5EP/x/hCj+raw1ufnKjkjTUohF38G7kpuzBgLQj5i+icm/fOFtj2z
lKZKmql11RfBe2DEPrsL7QmuO2RYw5U4U3fUcMJoWF6H54XG83cUjtbAjLX17BLpdeHEejIUtQf5
iJCt+S+8iMChpQmEvr9AflD6v8lq/ng8Th5Q8xJGExfrxZGn1JeW9gL6ZRNImX1ag6k+9V0LhDJ8
aateuUTsgswUvtCRJLd8nx4KcFoLClr9jRInC9hGkgT352Bh7Ee81QYOiHp2liEs+uOGxvvrGDPN
TR1VOOXcRai/kY9XBbGC3BcpG1pvUjus/IKuSlmQKpjQc11kfhKCZRMnjZgBUSzv40AwSon06AlZ
vRLYz4616ObnyvRxpVc7PfAfjQDNb9NvROqPXliIZBA5QAIQNz5rdVdezzguGmgMx9LYp4172Ymq
c4G0X9Hgdt6q6bBDcoBeR/bNMXV7umAqp8CAdn/dKneyD7cDzQZ6W2OJCO7fvWZjoQza66qX0M4+
96gsGMRig3xd3iAMF/rzGfALQi1qvnNFhaKSfFsIqSUrkPGS07jxiYWXQoCr0OwHFVCZV1hmc2Fy
4f9kfQ2ePz52QXR+IYUULXEQQcqA4h0SN/0ej5DEhOKHZAQLSgovXcnojRxgzPngqvBfoOSKc2pZ
h4E1opzaH6to2rX5UnrEFP2ZZUb2VAn6ScRQJICLX+c6kVCNXustTtU5FMIGWsklGXZAqHCsFQhi
YEy9000usgp42gbsuW4gGHJD3zMhPqJWEFkn6iAcvkBGGdSdJIEVrsOiQLQM/kaEzOBkUPxHbtQm
T1tdvfak5vQLKUAe9pqqiv8feK6bDqAbQMZ80On8kM42IXi7D+5GYpC650wvJXPIuJw9cQ77Lbdn
9XSteMPXiwIX+hUh+/gW7UXZRYhIKRi7CjXvslkFG5ZvQP3cr1yaJZhW+Xs+sys95/OtHRp4ANvA
sWKilsCugyvhOO7guB9//AyAyqfs28asoUKABia7UW2tbY9AuLKbgnCq1dRkJVpvuYaGq85N2ThR
FCnprwMItXIMcTMvxne5zpqhal1fny5tid8tToUP9cVwYl4bl6PX2/82gfW0Nuu3OtIMUynogUDY
TE6+gCbZFqsQn2fjlgNPeHyeJrGdmbMlF97a3CLSP3XEHmGZ/ZwoVkv7YTzDQQU4ymxYXq6rVIHH
COgTPccXMhbLQnksGo1QNsKxtmYk03yFnzMtMpe68O8AzoBz9sqIVWMFG/zTCFnQGE8IRAGr8Uky
pT5Hs7t3yERtcUgVJApHlys4wgOnXOJk614T42lmbXaU8AekDgb2SwVIsSA1hc5lwnJmWD214204
KoX5z+UGaZkbpRQ7GeJKo0eD2zfX8pVofIfpT3+YlN1d+ADNzGO5comP1aBvItJglMg9QfQY5Jcs
Im1mTEZNm72kcmgf65I9yW3UfLg2f4WM7teXB0JWSzDs1JMSsBcq0WX0mK7Wke/wH/Dp7J6jIOJM
dBd3QOSbyYzxruVBJfQmD1OTkrP3MTLNz8ftktksedS6j0BVKYJAzIryIdbFXv42GyhulvoGccmJ
Z1mMm8wuCAFcLVgObkz3NfNsh1lqAzzZk1y7Wxm5iqj2PjTKb5c77eRabMcQySc0OgTXh3gD/5sc
mrL55n/kUpCu0IMsNcM/idQBBPaL+if2zjqAnBBBueMmhBM0In3bHRgjaQcbRGzjtfxuy70yb8xc
dmWXQ+QW31Y5XTfxtR5DK3HZ1qNHjwDTCxk3gpW5omb/5kcztHsVJ/KJT1ytF8bE606+c3ZDm49f
712qXzeyfupoLbYDwCX8bGErXI6anQ3j/QvOZ6N/9RJDIN5fJfdNtP8Rgas57dFQ7O2lBz4P+nMt
B2VUrNkEXGuqyAfxqRWG/ba/UgLJWUnBlY03yavLvLcmmrPDtb2qPYt3/OBXLKY8KAwTLuiQVe7X
cvSLIxgR+YOCHWIjFpnGyA8BSp3OIEAJ0rZH1HDhJPSkYo97vt4zTj8Q3N+qxpNwCR55TaDDdaak
7oK3/JrJOtGrgS4kifSM9EcbQLRTqRpnwQkcKha70MxjzeGvMo64w0zgrlV06vxjWIGF9LTmX4OP
UOvRlro0BjfCPULPzQJ73yXkEvE7elyv4mlOU+sR4SYLxrccqSrEHiojD34t1NXE7LRLVagOAu4T
fTwgz2MBcgSceKFq8KSP+xfSU4VPh4Ne0uBk7g+OOu0q0qbgQB67pQEftYKp8KVkm27mjAC3GIw1
qz8Rv3AxqTXdcFeZigJ3NIdwBX/8glq+jktn1Vfz9fT3mhqdqnaTWdLYymlJi0hNzZYiepa97tLC
V56loP7IgWVFrgcL1OB0MsCeEsi+q7Q2qmlPaQF2tSxtFOGef6DQ2EC6YKecpE9Ph/D1W0IN9fZ3
8K7aMk8uwh7mrkH5nqEs1lqLuFMtQ1ZpuBsSQe81oWe/vRFbOfLkR4Q5nAIZok+RR3vLeUBLbDAc
JOfVBLo2BmqzQyFm1nm82EuP8c1hwLtax4yk9nIXiIPoYHsjiQjiwD/zX2ZqvXIlJmFN1R+vE5XW
wNR9niyyaVAfxg70kQENYSyEO8F2J000y9BIX9/YhdkwNBfHkljTsufWfhjvwuSVGqo8TeLZL4ge
/ZLaFNIPTkTSftFcFpVU6QmZpNsl5BXlEctbQNIo9O7FVVxsZq6BP35VvRKhm5Mley5xQ6G80f4c
yx5Gf1mpujsVv0zqTXn1xid2bUb2La5eaLB/DbFZxJV1xkHlL089gWrAWrSYGm81HmY2AYJfT4Lb
JVMPDGlF2pOndB/jC0XTlNuaFV2RzmfsLfaOI0b3qp+QRvWGRemYlxKdzrXybfmy1Nq7yCheeFwh
dwxgrodmo1weDNJg16JvWG+StZt8Fhkmjbzo+OXxr2obrAHqioIa+D8w939U1LjY/2XofILMKwN3
VvAR5SwEFw7gOKJJF+D3L7xsxGcpwWwnRpSLQBflKg8THMBVECsgxznrUQqqKHQdfZZ/OAjtN2CQ
muCEfMoUTjGJbIPaG/1FcOJiykxAi/dOG/Gpu4m3rrVA0yVxe4GduPv/oExsx2eIfhmdzZZl+3QQ
DcZL09P4EP22SKw722z2IPC+41fFd+dvbIy1dhx0I2GJWQUOb6M6U2n0AO6vHhDIz43XOEz78See
zW6WCknMplm7I0mkuJGcGvX9IqOss1rFAxrkqq/GmbcuVO/BYsqKF7ZdgY6bMESRqz5yULfxWqKa
GUBOtI66tesVbiL6Eh3ldQcBqULHXie9GqHRvDtL5NNiCXJNwfMNo6d8h4qxG1gp06dbObRPAmey
lUk16cBcnzt+pGMzcLg+1oKqmkO/M+8jJM0xv5JqrNrbLIAEv/DbA3NFPhr38ueH3rUd5W9jmdS4
pjHN2GiEA81la67wjZgzb1D6RBE9R62lGUdTW9zQl88ylrk1q64Pfo1q5QBqdbV7vBNDukx3JQLU
J6aW4HU8FA5RsQ==
`protect end_protected

