

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Kv0N+ODrJQAnD45jVEsSEPytnysm3pvAbJ05V2JaqTdEQNJrijqrY29nJXOyqQOIioMFCyAehxdh
SS8dEy2RvQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
wl26nrMFXa6fm7UAkMFkRbwMiWczBO907OqYX8JeRapSfb54ShwQXeaNsbVvqp4GNYQWgD8fiWsc
Rg1ZH/ALNgmzzsXH1hqu9qf40O6LpbgjO9M5gvRZkEo/Tsa2oqZnRuXHxvGdfSUWwgm16QfnXWFD
HONMKYo+TnX1BbyoHuA=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cF9G3LQheZJrMO7arGfYkxyoON6brspPywtxFKpTvNhoNGqsA1QaxZgfesvqKSR6jIrBuWrdpeSm
PoQl517JxEpEF310dys+9f254GuonHdyipWsWNgWjbTCuw6rYLvLG1y7lYwgHlSqKUNrBaGYERTL
bx0Arf8JZijWzxoSQ9FVJxjXj/PfvGzrh6e0n/oHLpafMxMPZcDI+yx5HuAhNXSr705mAXB8bgRf
GS+N50n6SUyWqcyUqw3kHjqQ2U4vJW+j5ZC3mQaQb3xJkZgzHfCaBKMstoXIjqY6XkB5Su6aeqKF
tsdYwq2h1uyBfljsOFo3IsRsUpNIiryBaM1j5w==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fN4hvSzwAQXVTyvBcSPI9qSFGq1b0QWYvne9odu5QkpUwhn44DFKeJSRI90o/blLQLnT5fdJ1IVC
mwqzRlL7DmT25nQgDxB1mM1knf9aPQaDbovHFOWTzAPBPJqGcsU8B7iu5g++kkRlIJA/0D9NUZP/
zdeXDuR/f3RpGDQ9X3WIBcSwde7JdAaZPxu8gycDj+eAg//eJ+Ch+IApwl6KjZF7Lov59CHOoVNR
udrlY4+R4MFUEO48SwDCDlqVGTYZykUVxSqzXifsrNKc0qKvKF4GbqbVHDidoVCoh7f7Jnj0snvM
x3DFGPDnokqNpDBX7xF9L6+GYPELuxQwMV3Yog==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MECPOWJAU4w/UvBGQeSeElgdlWQuUK1on5QTAzUF7zMKC1Dzhpw/yWAmwgERdTOHF4jFwSXDGCYX
dcq7yoSgrYHNe1Z9FD7/4uOTgF7lUDYslV5k/HR/cVW9QWbwl5jLUaoa4U/BsWl+xPk3gCXBhT1o
1qrFxMGkr18FyvER+gYFNuGtJOdwhkp3EWSeT0uUZpww9gD8GQxRUyHQJxyLO7OrJ+p6c8iZL8us
t83ykRj64BZ4A7H8a4gi13wX2JOPHaLBMG6QaY9NxFK4P+cAlJ5tz1UR5CiOSua4Nbo8RZAnEv5U
qSe9Ctk2cb+fZHyT1Jbe89K38c/68dSDrW+q0Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JGQumRp5idVwKA3zzoqht/27epSOGyhvfg4tXP+tPHgo6OfP/FU3H6/X1Nd4Y66ilN9i+iugj0ng
ehLY04ISDe8fLdY/NaZ+qOkmAGDYirT/RxSo79rIeXhylLKnHv9FphaO49Z/wGAPNVJcMj7acDAt
BmSxt3Wb7gOV2zsovZM=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FGXHNsFzSGXjbxp7bvoF47vhF8reHgBm6BrifhO2QcSTwMmIfvC72GA44UQ8v8jHIWHgPlay/nGH
qq6loQoHzagZ/voRdMzWla+HchA2la644cxBm8f8Fq9WGjAfrRKdp+ka7tSEmDbdQiKs1i43XT8z
Q9z55GPf5g5GdS4wXPj3ZM9TkEPcyM6MWas1txHsPj+r/l+N/OJNLRx9g9A23yQcrqoY/ibZoyFW
/7no0S9W9Nh+BPh8OXy4CwqtsvPd0/Zl0/JDLnm5d0hcEAn+3TkTvrZq0NgpjAEEOfrxtp+HqvpD
SE2gPjJVpUBZWou1zkZKYyakXZCQodq+NDtzNw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
F906e8HCnoCpSqD3r+WE7K+s/KYERotG9eJntWqhctwt6TVBq9CoZZVJN9Zfn+3wXVmdnhkBQjMC
uADKRbnudfRGL+nL5+j4oC0KbYfD0q8Ej0UOTWdLzd6Fzv7je3z8yC0NMmoQsg+CJb3HRyTLjtBC
lMwKQzTlR0fwSf+ospe3ALmJ2+kbK72wD8m4KwhJQNbFEwZ6LUJX7F7M1ZylRc29YvbxKBJAmkFN
zoFEbuwEdaoUnr4sO0GsFgDlPg86mV07+1YCTVnWxedGOrN5TaxztIvBjx9nZP57MtNP0Yohrv2h
MoIPiNshx3S2EZfmvwCyMK4MD4KfktUFDrCMGA7QzbZa5OrrXNk4sFdKzdYd+H/xjt2mMqUbqrww
NukumImAH3TQcrnXxCyG1akxvL7Dz1UY5JdivC48nxHVRFTGkXLI9ydMR1ZkPTDcSy7jlEEnU+sH
k1RJxIO/OLv+mGvAKzcU8NFOV9ZHKoQK2HRXzdlga4YHzPcJGrqkbmQAngkm+eEYdmut5bSPH5h4
AyCoBf0b+RwZn1R1Mm3dqPsHh0K0ccA4AhNm5/nX7oZpQ/lE4as7E1SJXn7VEc8Y8wWPnU/9fWi/
KZr5B8ek04yaGYjuIaqZkD+dINMGSeDqeuhYmQIoyHLboREDYUKjPyVDK7QnmyOCpnYWu/U94ZFX
DaC2j3IcUKTrpVXJsMc8Aip5bzh3JSYwgzxbhr5hvSExMPWnrZIvtQoSEteZECmHJWBMG2zi0I72
5x9PDn0RLzLVQLFlFkYXZt/F6Z8yjQlpiirPMsvP4WhNysGpJFAOi8AT7Gy8cSDpWJt9NacNA0q5
HQ2q6N1k7THqYa50kzbkd/wfeiaL78pASOTo2dqZI+eN5IPEHjRhbc40+gLhwlw+qExHvY0juHOT
9CdyJlj3Nt+eIfYYNImgXQBkE3+keAvlEo854f0oaGnccl0fVcaLPwiU+zpBVorKb9TkaUHjFi73
iQjAsHSY51OvU47WAYk4IhmfIwV4/LomL4U797cpFVGiz/7HhQe0m/FqujeuOeG9pPssPjMmf5yh
7Xtc6nRzAkA2xGVoQIcRYHAX0dPAU47UyaaTfp7fZtmBt8FLPQ5jow+O9S03NkuEm6599avBKvDM
fHt3OjONfu99dIaKPin+JIUn/zGlXPS8JBgg3YdCg+rJQrnyTfOQ8N76IAMkVbhDDUvyoYigJWkY
T0sbpubx5GaFagz+oez+YNGRsSoZOTIu+3uX6kekx0AI6k0rxFsQHvTTckIdDP80G3FFna3DZC6g
R3izgFXj6y6Mei1M7c8uDX9bBZQr175z6coEO/foRtCm9goYXQBZJFgFnX+suo1EmQBLnAZ0XsLc
YtLvwzchG50/572Pcz1mGS39Bboq4gP6f7FN1Mr2+ZEZ/uFzOk7bhPT8sxs1xzLhN9T+jrQQMHYz
h0ZGD4otMt8kQcMtrtubdT54Y0u7YbsNO8QupusZgWtLF4F08dj8aTm5tV+mBe5LnwwSBXmDDcm3
67E0psVaTbu31ewxLA7nkmyitlrI+37I2t44gsTIjDKRZWGhA7xGILQXTV/Mc0E/kg/xBFv9OdDt
h0bzywj+nR5Yg9FGLiR4crf/+k2jj9p1RvsnOanem1PWEXg+3u9TFCDR+RPtIvArmQMt/61AVQEd
KHZ1K/kWikJrS20FXCLtwGdP5jA84mPploNs33XlRBYX74Dv/ctjQC46j35UU03d9xK3bm5OstX6
e0Sp2GlHV1yiNWLqRJRHIRV4ayOgxGEsHQOioSBR6Qm+VE5tPQxNAreL+abiGHVxQz2ih1TIQrmr
gSIIo30BUk2Thkv2Z//ksB3pnwH60qI+QA5IDZAD1vEWJM5y+zbiI1yM1Y7OAKWed85q0N4iQ2Wb
vXc4y/wQtKa/x8JMj09XCdtBR75T9bKus0aRbBRpVjdJrRdUeWNFLIQ+nWc+bvHMIs5LVFu9Gfd/
e+EMeFYaThmvxlP72zSrjcr0cUGkXznU9qg5YrH7TrNedPscfcb5H3JjirgxP1Q5lB67qONtnBxu
xrz/lYZgtabdD2n6raOm+ZkNLNDwP859rUMiEIMoAbyG91nbaP43EsQFWOUXfZGkTUNlIcyG3/B4
DuvTlRBusthbnNTUUhBzxDZP+sYNnyxDzJ7IejaqIfrzjbC7t7HrdoTq2ogXzJ+ZZePw/bqbNHsJ
vrH4SpmXtbOgA2k19wkLXgWgmdmxYJ6VQ/OrjBvcJ9yDOfCU7A55rwB+L1XWkyqXc+zEqIH1tVPk
J/1TFTZbySX5iY1G8Rl2gwxqrgCZYGRaYIuFE32uk+Jey6y+DsqphqsT9pC2AZkplxmzYlg/gCGx
o0v2/j/8IkpwNYJcUj6JCX1VWgePEvawhYKuU0iyNcqrxK9T9VcTnsOXhdVchQk7BcXQUt0ulH/3
ggpZl8REdR1hwZ11YyTNYBH6v4RwCIRXs13dd8ST32VGWYcXYfPWQAuHYmFSXs8OLiaUnECRYoFx
SxnMXW5yX5vWUu034Q/Eo+rjUz5sluVI/WOQ/WkSK5o6wMUBucQO0dd8so1Y+GrZka7a2aKT3xod
iFOlNRYIOs59YtnrkVKSQ764HwCPQ1HxLmbvO5QGO8IsyTBR6qiPKarrCri4GzJoaZZriefSQOFQ
ZTn29T6uOOrOSiqF4pkF4TBiaGa1AblH00BG3tzkzNEFkUUShJge+TlNlZ9n/sIN/LaJiGz9OqXU
tPv0+BNN/wmDAwQojGYnTiu0v+bfH/fE8BsLMdqzXaLiqAFRGLjVvF8bGJs69m555RwbrbuphvJI
QGRI8U0ZF5s9UVsHz5bbjE2N7Ib4vj9U1iug+CJ65ormhtro8oUReLMIJmGyhgBa7Ia2TruNQjdD
slDPTU5/8oG8ZV9wrrSR/X6rHuTKutPpm3/tEgANzW7XG7iT9ZPpUFde76vSX1reyEqHZc57yDNp
XuZDr0OhppUG6/e/7I9J2p/5Xv7tFg4RrR9X+/6XuHLRAUkHwgPsXDMRS7JsfvBChOtrr+p3R8YY
IYgee0n1vQMSkGNn4vqpaJeB6ILFOmgKJ2iWqDWx1ZGuaX6/dmdmQmK61SKyKtICmMPUau+JqX8w
l2HKdqa3XrtFzfUkcWddMZgSza5rxeHlo5aDiuPPfr/aeiNQ4/6r3xEmjkrYLM3z55cIEfxIMLlo
550fUex1HkN+3ZLpKDFPZYtwsljqywhsD1MyrcuZSouDeVNjeMwgxHxQiTS8YCArpwaUily2d6T/
hlxtwLfH8XdZp0wNfKhOrzVJxGr28S8ICRJol0a7fi/Fs+NmyIqPSrL0yJwDkjhhgz07sFUOn3fq
eczlJ4qIuuZ886f+OUtWvo0g550I3jXKPXqpLVLJ86khMBWnnmnC1075IQbZH2z0nSdCTBAXX03t
vi6YSUgIw0pw33zcRGgbDDBUVl001ubKu7+33iD/URrKyb7YBc6SnjLuvUn/o3vyNgUuEMDXvAlr
VVXu3ky0MVUfnOvPd7ZzOQSGa4ct/L+WhE/yMZ51csk57E9HbfeZ/VqObLLuCWOISD9EO9erYWMI
J/zX1I9rHazzsCZoCVFOs6+IUF1n7a5/ilgE7SlIbmDV5MQv5fHvSd22QxXfMSfov+Hm9O6I2SnS
ZADAi1tSqp9TOc5cgbPcDQw3ekT9F+60WGxLXZbGQwce2ZAiajEKgrfAxasv84mj1E7m/OKV++5h
WqoWOclPeQQfqk/9dp9zdu9+r1jhnHqSWCJ/Qb/BDGtua2joyNKgVi+yPe94+ctRJIs9h4GfG94l
OQ4zHd6HdvcYdLa45t6OU6ALBw2wVjs8V6AmIbXjedqnryB4vyXTXg9GgQJbZGbS0VPvXlkSL0HK
JYLf6Fw4/OYf8hfaiUv3iQC9IWFJ1LKPBngrxnW4CsqCRFZ/hYthVNJzRx4LVc41f+OYgxp64PPq
TM88kZHjx1qe4Bx3R84S6AVTmYWhQ5E+C0PMAive5ac+LvXX265lEpdjsKzR0UlbkQVwx9NMFOEg
uNllRewFq1oh+7rKirHQ+c5aUZjG0chRRmWMPeJr6Mo2wy6HktR0t4sbmTkAPq0oHmkGLJrhX8xh
+kB2BYOVyB1UtLTT6glVieJxcSzw38+25DKbNAgaXF2HKj1BbmiG5gG8GvJB7eGkGXMeYHCKejcA
hVzmLjkyKQke8L8JXCeArbWz4tdpZYmnF9WUqBQGoScnaI+paRDBUsFjXH739Y2k+QnQaqvALTjp
VAHkWablBheBcQqq0BpwIYEXUpYro8wnrA/a/cihUw2MgIlYwJyKRl+0mp/0/ApvJ5E+5tHQDkTf
dCFZYtTUKOOWc6FGu8vEK1Fk3o6hSYk/MaNnTEQf2euYq43EJuSpoc1SWt5lZwddPTW5aiVq+ZzD
3WNJLNtnEWnDgA0tvpqggyESnJQi2W3Lg37ai8RmdMdUcTodWNxzbpF7qh7LIm3bV2vp8xE7jsFQ
20YloAP/SzhXF+qc0zoR7/ybf8Ofyk/zcbMV5XxWSIoNQbFgSSIyzZ1q6me2uCb1tGbLuGX5chD5
lcpkQO7XL3yh8dlKPJ96Jl2bOIFZLuNVSWJFZRsislgUOUeNZXue0qqcM58Qw7+l18+sFvpeJut4
Kcg3AJm0oIYxqZgluQ/PNYSEDu4IpYms95JZnny1LBnMhTJHuBuDAErMQaDRsBqJj895nZD564+B
Cr+gYYDF68G/DmjRAAbgSoQWgDip8xUGc8FH4YFfH2UumQ/F7EOpE+ZLLRreucD3SIcQlw71NSzg
UWBXMYV8wx/QlxuPwUpciKO+NafWRcMWtYKWqo7icwQsfh8O6s1fsgnGa0nSYHZu/KCp4lc5RQ0s
IYhH0k4zTDVSzl+uV6APpyANmX3Qykw8489lOoM72gVyDqc7HhIJF4MSHcAMcuAaMaQ58kBGaTih
lGAxPMWieOFZFNdTEKZpt4Tnr0wWnYU6WxKbQNFvyOHFzSxb0egCJ/45xig6e0HTH1UFgqOfqu+i
HoeexfKt9UIVTmeKoYKi5TXljXb+BsmJ8C+ChN80S/L8G7+uQ/OG0g+13Dyamg+4AUDrxXRooZPM
Pi9ynCANaW7RL2JcY02wvHSyq73I6d71babdfstHsPADx+Ej601TFKnQZ9/kW/NgpBOlablxvBKQ
enDEcU61cpc9pSvldbvyRu8Mj7Y/kZ1k/b3ili/HC81kc/Fzjuj5USjF3mu8c4vcJ/P+7R7eF71o
9poPiBm6TRfYQL/lVNl9c59SPPLRgZCI83ZoeR4Wy9BrdRBv8f3eZpwuVdAECL/rUVFQ8LYQ1ZxY
A6zxvqaMidJoz8VI9wZScNzFI+MqBWxGRGAgqQoupKD8dqF/is6/aeNvMxUPWH38fg/wNTwglTpp
peydjffN4oxek+RJmZE32yPdnLo/pbopQ05DTcuyhIwWkGS1MVYGM5fj9MivSn/SqHOTzPavwKmu
ZMOAstftUtdxi44LQHGOa8ieVCEEQV5k3W0VQw1Hy5XFh7liNbRI1afqwHjxf9mYh3jwDbYm6OIa
zPjVLNuR7ey+swOc7nHfFeAFsDTlrzR4fVi9bgZ7WM/gGh7Bva1/y6aMEDRgR+r8zkF9LTeP3bHy
fK5945/Zekv+5TkIG4uCVqOTclekfWiUQatSgd8SsCskVLc6RwSNYjoQRhgoJsybfZQB85q9k4Bi
oVGIx/gIF0WJhy9OMMOhn2gom4vL5wWnznrh05JfypqspedttmA42ioGCp7UzmWg8eqND/hdV5t3
5nxfMHlbxBOIx+s3CIhJKlbvCaTQ7W3C8mu61X/dsDz0BCB89nuR4wh6oG1aAbPaBFTfff/s85Ro
lWR5TB62FlSHCizXox8B+xDWxCvGhALymq++JmoyD0H7xgOoR0ZgnDHJ5PrehJzicJzspDBsnMY/
lfekHUFuCUwwnIV5VIl6qO0bepWo85dXfxT2RZ9fYaHdFZb03Q55LI+sk+3sAuSHJMvlW/ffVueq
8Blj53HCrqtv4fn+pK6iC0NiKqgr71u4MpyTXXt+YUDTXCeoVKqkVzckZRger0OYRBWl8+EK0AP3
OCI8BrSIenFvG/sqtQw5QQoDt8DrF9MnMytG0PeSjNWnaBrnqzsYupTHiqz/cHu3a2VPIBhH4LG9
3iR6GDyKz8cxwZzAAbVOlGmVPqQBTdMlOyfrNFmezCOnuHPNDdGnMBWj/U9Kw0vzdp3kf332QZG5
9Wxu1vPq1Phoen1hQXV1ss2FJBG47k2NFzKqorLBKhQOo80dilDb4vAbA67CJax5t7G04cd+6jmZ
Msn6wIEVew1Ywl28KgnCgqzpt9qxQR57pNxCk/NdwBjwIhBrsdfosv9rVLEy7CedjysSyExgmo74
q/FNRR14iksjdRuhlpCDC3ag8Pf0jIrq38eQai0aTQFMcE8bGrF5riIfWVFrorzb4O1CrJ3ljiRK
fVI+HT+Hm6TdRBnvyg1ffqGphcMPuME9UV2CThT1g/XtNZXiPI1BFC34HuZFZQBT4ULTwLP1W7AI
tuPwyo7N4P24JXK7hrYXI6H25GTvt3NW11tyX6IWl/b8IQpLUFEcuJPRLDYabrVE7gGcpx/lTkuE
57liANVpdXn3YMhQbRDl845Yh2Vdgg8G4uN0KXJCAcqjalMPBaL1Q5al/U7PjOqHXyfnsxKWcnF4
vqiuctWku+9pHfMAeMSriIgc9CGNTyhtUszQOBVT6vzIfTc/O0w6girBzErbTRjmblN5nLjT0rB3
TTPXtItmKYmzvHW8334ZJx/6+3VUR9qZ0FRGwNNwVPErehxjNHA87Y0EwsrzWDziaKGMvd/YhWhB
JQvMFCQXL8EZv4bgCRE3xbr+Fkn6hoKfBzWkpRNYGDS9vkVve7bGOhWsXL0xu+3KoDRAtpW5yni+
/Qe7j2frP7JK7v6uBo6VQj4HYc4TYACCxTJ0Ef9dCdaSldCC7GmSaCgUJvb/s6gcFC2hqiWPudus
C5q79gj6kxVCfjx9Ds/k8r2OlJBxy11cgGDrenKck94t18+TqKf3rL/YYIyABFN8T4Bu9+J4JNFA
DPJGqjOtd+q/ILvlJ8a8XG4KVRtGA/jOACpJ7xyq2X0vDQMKpjl+mIGM9P/ylNwoyCSJbaTSzud0
Ma0yiq+L73hKioQy2UBscgiGOwFdixSRXb1Rk3MdxnTOb1DtrxMnspN4tdk29s9FUeNzmmmqETh6
B7bpi/xT5u4tSsejrC2q/yj4kA8/zZ7WCWH5lmkiOcJChDSKvGtVidnbXm2xkrTCjPQKsjBoZLLZ
F61mHydgbWxjUE+ERooqoj5w8XAEiurilcVuetTaLoW9mjULi/Eye1NSeiF/27XxWjKjNgmNBWNM
L3xz+o3vkDHTx07B0l0dC/ni5DZo3/ehZr6L6PgCs8SMHXZh+lo86OklQRvh49WB1IEDisrBoZnt
NvQpGzCu97rUlSAi6Qa7sgBhTUNxpl+XOibUmIR4HdTCadzHKdtX7PGwpMBkSXs4g1Q4KHyQkbCs
zNo8dsayjpr1fCgRMzoFMR1gCzGyD3B67o6+sdB2bSaGWoW7W4fJvMGU4aPta8zYu1wfxwzUDXsA
x/QJPGVt0OqRDIofQEVuHKE0+vJzNjACWCwKXLhdSnimDdo4Iuhor0+xu1m8LsuD/IlvxftlcyL8
4IerMCj9TU1I2OxqGoGIkw1Go9+mG7SpNFDKEFokwJfwtPwa1zPf2gLunwV0lUX3mXcAu/t631go
+qqITgIk3qCB5lB3qKQmjzs8ie135DukNuYYkv27hLJknTBZBryWzddBYVXFP0/s6dzjmI1rtflK
QALFvKrL5Cj1EpQ+kw3CCBX28t1mIWfbqZDd9uwCNC15hQJFgmww6323xt6F52+uja7hHOsf0Vbi
bh9019i4t3R2z4bec/G4V/0uQiyrI7GXsgnMhW5UOaj/ffZ1nzIt4XHL+Lv9yE9Dw/ukpTMVCBca
rzjlcfbzTl/FPMiUHTQSIt/mhN8dEzFT1ueMfBph9xwKCTzMsKroSY4ICwV2h1iDj0Le71D2Xt9s
eNSdAgeAPLkElhI/TLSTbFv15ei5BSzUvgPNbylGUG+XMXUtUAIhKCPlAWCN7lywDE3dZFWkBgb+
Dci8lsbLmxjbBkhVxdF35eUxlaLPOJWWpILrjfdONXcnO3+1jCw5aP+yV8BlvMEIy4hRlS7T3f+v
6mLBMImeV8903WdSxYM7kST+qW+UHy4DSCMC+PSIQ8Qo1HBbdZWNTuo3SBmy9jP9xDjFvbwfL1LD
mVIsVLOyjfmB4BVz1K9nIZ2uNVY4u+bTmFMuwkjO1okS/X2Yx2LaAlkAWSEA/IgEo07iHF9dZOm9
6Fh7l/rxQAA+4Ss2yZBs5FlfiNABXlcW4Bm9n/AdDCuzQS0ehkb9jpqW/3at/G2oJZMyJ2uCyF4m
27C/8Bhakx0SKu9a3cftJ5MDici7ew63eh74wJFaOSB5zhDHUALw7WRTdEVBvCQ+Ekqo3m9pFECq
P2fJNrbk90dttN2YCvDgyqbr56tWVk3XBi/S4RhH6NcF3230v6+RHLO9pRZW6hbnjYaxVpCZH9s7
E9GJcb33ZWSTIy9LTzkYcYm5fxw/Yt1JDYRAx0J+PcX8hP2fMcpUCYjZXdE/fVGH/X6mbvD1uBxp
+JT4j0+wWjN6AxOfZIwh54Ds9HPgLiSEPK8Hd34QvOifYNRweozk3N82BOEH3Wj3K3eefW2Z9eyt
nicAY6pY4up9AcoJimjJgziV4N8TtHrSMuPuPIb4lFTypwEoT7Kg0rR2kfYTydjlbB/Jl1mabY/o
VyCiztQpLu1VFok2SWur5ay1EvjK/JMTJ800EO7ERxGni0xEz5B5ue0uMU8dVmBaz+9Vn4k11pD7
r9XqHpRAc3WoNiJM2W1k17/7uMMigBJH2FTe7T3zg8+2Uus68IVKo55ASsZ5NQzF2iMVOk+JsSvc
ZkiXh+ThjDgHyHLFNDDxdBuW23kEzduaFxJ1bF1mEcuHKv6S3vMS1vuWw0ezCu5y2rXuL0bMiwYm
gmwuTxV8R8zXGY7PKg7qLvMEKnxDxKTEZXrmObCFIZg0RkZnpJvSmiglAbqaWUsSPhs4y5BH0ngr
6pgMqbUKCw00l/oC9GXr4iwAYmD8XnZlIuR4jSrL5Y7ANzfpogLTiPF8xwiiOh4CGyDFRe/utaiz
eT9axjpxVIRKkPGVjhWD9sZTdSPjjOcI+Nujk/8rdK9cr8iEytxc6x2x6WhvfXWsuwu2XcKmy6dJ
0aHIm90/sZW444Ym3QPDRt/01F5UmSioL/u+D9v4rBJho80dQWYRXZhfxqSOIP8/PBEIGeXkGSPM
+t17qmIJdtDFrn1eEkqC5uMxFF+qgX5QSvONKi+h1trSiLLlNPi7+B6+K+T6lMiIFpH22dtXFNKo
xWRlsczT0EzCRfoNWfzwrlzNB4uUZTB/2iZfOCX46pCeOfvMjlQxS0Rue6bbUHswA+I6PIaU57ei
3cgzNCfCyM15+DmYh3kXwX+T9ubiMpFndkLezBZCGcSHLxV6d8NjRo2jKIHIRZN7x6ezDXgKBzi5
dNXKudUhFVzYWJ/8y3gBS/PfdecbD0Wx907nurOFR9gcuIVOQI87JECursydwRSbACEuBCNvTCBE
Go8GTZwVymhdmufI6dpA7mz1rHIJVnUtW/2kkkf26VCi8XVqEiPHg/qP4fKiDmZSNEQziY46K+ZN
BbQem6xQTm5jXLB020pLio/E/DlZDIsB76y0bC/21wqM63PNSoMsR3OqoMkinXldttq5TsCdvzG2
dRjulvNkLizV7Jz8Owg5T2fYOcSjUPzcNQfC09gUGqavHLXXpvGsaAMTJUeGbQmw30T4C6fV7Mhn
dcObLLp371k+8fuUyzn6qQ/txXVAf+i68s6Uth3mUVCXg3KYiouQCIqetifDFG+bzhglhqP3597p
Di/gaccguGcE58y6i6SzFXLDuCjIvwSZLnGHYE4liHMrp4GNz/n6pxBuywEzjWMZtzlQEvYLjVVH
/ZaAKSApWzCtJR3pwaOi0LyT6g3p84lCxooQBNBa3LOoiIKZxLobIgGYvCx7/bZfzOBzRexwxlVb
9Tn1rM7qxsg0f/vM9aPo3vB9juHAWc1Ih+Z/gCFFXmUtm+Yfi3K8bZxfPWogzAi2xO1hn19ccUpw
5UXIBtWIZm3E3GbudYl8x7aElBfy4SUyR/RG2sdysHkf4vj/SfdB4O07zIkVDGm8Y+jvNyGmUgIK
UnTppkq+qfuUxevRWMnH6/MU6V+yq/7p9TCIGCB8RYWcL3g2e/rSZAMnH2Yj8TuFC4xeYL+W/p8F
UYRM40MoHUoLCF5apMs5dO3R7nvqaTPXkU8r2FvY+d/menSYOQ67mHHIbx+BJkQ+SZmKfT5aPmSc
E2WRCgAHtCC4DIlrlJNNGUnnBJ/Q7/hz2mO84gPJrlH73peiawgDmzUZM28A9i613Xt0R6ZNTFKc
tqBpGZMaGzepFWyrPX6TniphIxjK33gCGsebwVMmUt/IetHNZU6eMRUumkTjhk4xPRinoqCpoMPG
9hM4srZdu+qFTMYYHhs9MIjuOi+BaEwTnXogk8lMA1XhXdflwd3B19olpvaF0xOnV+Fmch/cayLN
v/jEJxkJqZQeXtjcc1dpgsOAsSek8F4SxXHXTNXtloxOvl4QxXoOc9MoyiolctiYu53m9daz+YWF
ujBlOZz5qYJlviXrJiHWbhWpGCmP3FsPK67lMWJgT6QoI7GCJqFh8M1sNoQLuSRys5zYH5Z+wUWI
tJeI6B1PRb/Hb++sicqfp0c7XN0rc4LqZnzvEoMKk5QYYUePJKPmV8CBmWfWAYE3VXXHXxVhZPnR
ojZUMi+IcOtVWjv9I1oW1cSfCtEx3NzbM4rnEcZs9klKCqM4XV/+faQr78kh/sQl6m+Mkg9FBs2I
frGrXu/tPf3Ul/zslpt+wnrHOqZFGmSUaSU6cG2gDW7KdFgq7zyg/nvlKI1DNRjW3lF7F5QmwQnS
aMHCEeK/KcvXw3FXgXwjXUYz7cLB8TzppHMshIakDuww0tZjN8ZTtHT5dt0j844ucKyDzqaLA9kD
JQWMg7jC0p5mNrJ3844SOy2njJEzZ6Ii2VGillcUjDfa3TcxJlVWva3f+C/6I7e+LSOziFlvktna
UbRYZW3BjYnBiT6NHJ7URl5Ilpr0eYII8LlSAGu5xSYSPayLADrhJoan3FIQB+kUwIgL99FGWqOK
esZBJlZY4NKC0x4Oj+o0MTHGjwzdbWE+igyOmmGa/A0EYLpnWqxFPc/bZ/6LRxvtg/NP5hipcQlH
VNXn2s9AHNu1yRX/KYqJyBJGZSLR/O43+Qsa8a1+OpbwDwD0dzHOQgnj1VlMGRU5i3MGAuZZ6XXk
ioM5BrTRrfvO5zzVTnr6Prmomvo4uhXpO3b0nUQrWCZdU1H0mn6cBtRvtoRMLN90xfOFP/Ne8CgP
/WNBJagLAxfTdaCr7B0ThTWd1ynAiO37RI0KUMfqSoUg72M4hiuZ/givICZpr/gF+b+2VZo3r0kh
4iACUa18ahX7o5xCoUTcNfJ5jVbpxa3BV+2aeKzuwNaRx837qJFRBVIXoG1N+YJIrRqJNKygSdc2
A9x2MaxSb+nXViMxyiWdUk1iHWH+8Kd8p2O3ZEKEmO4xXxUlOoYOPyH7rlxC3lS+25dAs901Ce+u
fMdrJHB+4Ti8wUXrf9xfaGvudpAljvLM/FMWvC4ahNeH1SshCH0Gj/APwuZsUm+tQULIZXIr9+PF
BXRWGg6ws/+cH1HNo4xRSNwz3q6gQagNABbWhgG3geXPsvGz/PKvYkchvAWqLZy1EUUCBO00FItc
nE+bdVP1PrP94JrUPYhJ7RD9FRgusDHf/niFAzSI4/lbTBX11OrwY5LRjSYhsPvZ8xcrLs9xLa7W
jiXVD9iherbFe4vn1AuJDda5dRnDPB7HnjAqQnI4gBBNtbfybVQgLbplYfZyMM+JW0tH485ajyFd
BD7Vhj7gQrdiGLolTxf9zPO5VdgLKRXnOkIZv63jzExYcxE0ni1i0ksh8J7hUAXctl0KvM2p2Ts4
WWehrP4xkBXj+1jA44iTfiwR16HNnUuduiIxOZy2WE4uVlWwMoDsniVY9xdVrokJrXKJaYa5Bl39
z9IaxqZ/YFReS1/Rj1Diueu0baSmQGW4sO1r8ynE/IQJe0jsgW8s8APSEz1fXoGILG1HGMHiTrRw
CfQS4oS4R5HnXNqnoxgzYw5pe0qRYOj8X1jcYYr/dpStZ6+1wF/xQT8Tw6OVWF+XXW5hGCA7QXCx
ferQTJSwYbXWw7/7Wc3m2ZFXeOZWHk7pf4yodEZw3sNT+xP45+vDTbaYcyU8tyOk3YVLPeqFqko/
dJ4fShDBbngT8gRHJDG2nNQhNHFvTAj+xPvNweNP4wk2uPWaCp4BaUVxdNpBIIP65FevgbiIcwcD
QKDY+zdkWSxKPCkp0JjYnOhU/A27RPbTU4xUFRWX4fCXZxBAJA3ioypbusxRs7XnydBP4pVNXouk
S9ZVWwkmw+rZtMMXE3roH7fmydxTsrenH+1mEMtv6Ce8CglV90wjx38FO0IFTR61rBkFP5a//xVY
59jaAQ/ZkYdkYKY52P/SYXH6DWivLPXns8qts9m4zC6uJdbGQ79uQDZzxoQOi0UWTwgGywR5htBv
qIwwkuKHsMxdxq930lTkPKG3/eSpfjmHq7hQ4HxIulxb6MxFMt1a6zAMIRy2vQzPb1V+1rIG+/a6
Qzc8bcoZDmUjoZ7gIr9BPaofZF+p7satGGG9IdnBmt9Z2SdYodnicETRoaGLV8d6y0MPLinRVrzo
QnK3c4EgbE6PYDxFXpBhllBzodLlnUFpXGenlop8mbSTrxuKq8TxvX0xEaIL2U1BjjC1NdhV89ib
tChKzXtB0c+tqFrxb42r3MFJp275UV4IExWZ7WdgnTE7zt4I/5U5qtWid/KjaDSgKgSkHkI/lirs
j/27D3iIBBY0/x+3qmhaAVa6Y5IDivSKAgkBi/+aS/5FmGVNrSV1w0tWWOv51JaNQcG1Gilhbm24
phak7QJrT/r8vSMsqnuSQu0fBpNy7v72ehDc6D2cLajlicIzQBwCBIFuP5OCM/OgBBsc6hv3FT6M
pPT2nhIHTkRWXvmmV4QGbTFEDgo9cew3sclpUhZoI/EqDrqJsdmrqH3QR9g6UgFvQPgkJityAmh+
zCdyFbcH4ruThsarW4iEVo2C9U4O6F+VFZCAX0kbIZzHDHNJUcPnPmg6jlg/doCVqaiIzi7YK9DS
PKhR2yXaFTJdFrZYsbMh4oUYgh4KFkagp+bAdhl10DP0bdcHZVvRWuHdv50bRCWu8QvRnMfW9V2L
+ne6Lv55eBenoDGZnX4cxdajOXpENP7mUtUNXVYpgU1/aXhvECv82O7lYW0+Y0NOY7i1zuOGWY7w
yV0ORvyYZt1b8f6U79+I6JIrmS7O1R4l+hL06OlllksL5qziDI91t4ddYfzgNPTP0Iouws6kj8b3
jUt6tBxDo4kRX2dnrWeb6lReTNadyRdeQMWo9LDF1ZKrFvRd5plmbm/ZKxQHhDAa1hD1QVqlyiEL
AQFaKmSIoyw/K5SAbGZZlIsl0p4FK36hTeeVyh2Nd5a0BK79yK/eZn5VCDtDd1OIhvzV5+GbyolK
QrnjBYVrAHuFCp7/S7Hn9BpR3AySLmDnllydApm5QHSI15BbX+MGaLTkE9ZRVzxruBP71sp7NfqE
3ohG4Ec0WQ0kdL0H60yViqCp0FOhmja4VuDwW+0ZoWQbys/j+fnwNvac1f1P5YopKmpl70sKpxMk
9BN/ehs26UFTcfVacqeBPEnP1yTT9HDGu+KTT+qzVVWrAMtJd+8x7NT0/yHw79NtcY7UcH2HwV2J
fTFUg+ENshASu/nUy89ivwgHumh1a+qxx8Ix19mje6EdYLeYYSlleFtSqRHbALNv2e9IZQqOkH0U
Iz2ph9AYYxvfc8BpktHXmkNu6IQQsPwnHyrFXP/jNQ1zboKWRzjO2r9TIffQYmdgWlZWlat+hPBy
9i8roWtQeasBE4mtItoeKmxxzgLz6+m7D8YHdwzElaCE/oRPt/+mWPsLyEUKDNVbqRGvhhWftb9T
zoa4j3NeSH4iCC4i09baT3war7/nyfoyw7gpar3LIBwuzIAhXaUfIACuhbUpEVvwVcBjr0hyB67S
bqMZYio2gYpRU71xceuraSB5vYkrLs5/kpns038x7Gs3rjV1Mt9NtA6rj39rsNoAMNvoL04rHpjC
OUMbhu8RnpRxV1hTYSV/+nBufZ7YgL2fdFOxdEt+Jo/3YqDolYWgzF9iHAac7gZlouKrbK+Ul4mi
9tXX2IunfRCECyJP0API0u/63x2fxtkTMJW+jtyxpKVSqOGFizY4IqYlgI8pbnypzACgFAESYTiT
r6YY7h28uKjL2aRJ/8t7lIuP+paiwqmTT2pNyk2bXaihN86foRkSEsJ2StAkQgu8LV+6bhBqX9wE
REw/6fzOENiWz/U3bq6m+UHNz8Xp5OJfM5mtkR5+t2jXACKFc+CK6J3oALfnU2S4H7wSPJvRdDod
kVkhpeWt8MoTHK99ezl6YxK3DNuC3c0zGfM75IKT6ENWH8CpYy91TKdQ1wkhnyM+fOlPLhqo5lwt
voXGU2Pe5Tz0gtg2ZkFCdG+2XCbfm/oV6xI/MJXyDtLvHM/84rjNCYU545sF3OOUBemxVlmRckuj
QkgY4ylKDjTpaKye3KUMQmZmtJeiKcg9mbzlQ4VU6bDfkm0VqPS/h0fb3ayqj+BvLMiKr+f7H50h
7eRyqWFOlARIcQa5IMldDX2+ZoxIzqiiFI5ySG6buT25Qx39v6bYFzZGuwxQGqRphrsbZbFHdfv8
WuIrhS7hTFtUflYq19sn5T8npS7XMLChZi8nCa5fBnBfvtF4TxjmQ2fbXjsqroDVRw0PSquoYZpz
exb4oAQTIloX66P8lL/PzL+jj5Klx1eZC9bnPwVcG7voLbkMTvjm0udNSiIQesNwTHemTz4d+Oco
HCPJLau1cq5jaooyd0tKIE/iljnoEuE0pi6lreIvxgRjjADj94VTmDuSwd1sQX/yH5ppy2BmAryr
EBVD3yNJTaK/BwoPx3MrEqi9EpiIn2gk2UYXd/1uyPf4us0jxSXnw1IlvMkQ/nUXdfBdKWB56zRi
E4Qb5R49KEtiI/fE97aJYG91psShIVFyWgcjtVMCX9HZ8qK5hd1QFC0HB+Im/OJnUO1PB+mEDUKH
aqHsHKY0oCRQlXWE23JdGYU7cxMDFyAatY0HI55mS8IKz5IoU1pm5fg+Uegyq94m2DVRdgPxF06f
oJFazwp2QAeFxwyuTgSBmobwLaeOnr4H9TJT/BJLd+CHEgB/N6iQzji3iHStD35XgyRN3VIm/V8d
0YbfagKMNorSofIFosga7QZ0vum3jLyAhw016iq/lnfteHzvx1znkD4MlS7D8DTsKVafjRPPT9n1
YWJ/8tfZCBhQqsdJ3JsuGe0Y/OlUMYDWQCTI+EN1oD8xUBEsZ9Mx2ZZs44nu09+aznTAd64Q7UpN
MHOhTHy5w7DrE356XoJYdN1VPQWvowZqT5TJm2TEFVEYg7HoV1LZf9e5lDmFIloKIL6jlZ9vZvNx
q+JwJIgZoBqk039IltWvJgGwgjFQvDm0MZLZT7VAiLRIHshMTd4Fb1ziBkY17X+oIkUD/bYBk9Do
s3OVvK0mO1SKkd9QQL3nKaACqqxHMX18lq4dzkmkBXU2nXVkCm8jJkRm+2B2Pjgua8zDPAXmZ4zg
kUr5QhXreasJ0ljM5ybpnJjxZSiK0wFH7mFol/6RE1RXxyPrBQr+e7yg0gCKBuvIv4Sv+cSFJn5l
cJAIkJS4W5R8PqAKV2QcPlinw4kMqWOBnhOgkgwZH06eGzCpTE5AtwgSb8j3WUQMmYqBSBXeAbDp
BqNEMprI1I8rKRUAO7sJHMz61ZCHCdGUZBBDqGGi4OqZakmTlObRmnuOcE48DFPzfpGDjzu2QE1s
894Ti80ffa5vdzy/1tLx/JlTWmUeNHM4jMdcbC8AFL4PwJ/G+6uYXG4bCjMOuI9VXVGtekWepZs8
wy8lEOK6G2A127Y+HdLoyX55TLq+6fuctEYavHTGJlST7xEtg762sg685jPJxjuVSiUAHAPGTJm0
65e+uk31S4TyjUY3tcvrXdScsQ/Wd2JeqtV8k77IQ2Jm8LSoVLUsWF/fmteXnZYjalDRySO9F4Uh
tuBLrxz/3YaEubFG6phUbwSMW6fHd1uqSjuUM78JcLBNaOuSiylR6iD6reMVx8RfudSoERU2CHYt
ntA0A8aIfZArOSR2ZKX/VCJbDYRSmU1epQb5nJmxh8SKLKyHxlnF4rdtSLlO0AjYdV0cC9Sl/NB+
iMG7Fnm0W1+I/AqGOQyq2t1gF/Cgle9P/Tg3KCwqVzjNpUblcHaSgM7QO99p8z3+0D+Npk5OogIa
X9jVRyge6BdmYo/xA4sGL6xrWgpnqVnnD0yU9IbVWMX6oxKxfmnl1Ig278+04jlPo82rfld4FJir
MTAvjJ4RqFHveui5kr0iDWKBYChfEuhig5Nd4YoC7w36PPwwe3v2fBAj1FpZnSlPu2Fxgglj9n26
TqGuhz3j1kZl1Afowl1cxhkUSL6SV7HFH09+mYh6nSohqxIdwn+eiIgY+5VyZtaB2yLj1I2Mkdzn
Xxku5Wih4mSg3TpMrLl4z4M8ehoyVx7knBTeVWPiL/rE2KRMM/WBVruE/QNlBJoXq+UEwiSeoUCA
SJUl5PBdJ++2qcO+vgMJZoysaiDBrKDoNLSZVPaouvGJeuMYIe0kLZIBqbcflSGs3l1j0h29iJHC
a4o00WX1NNKTHcv2WyCBj4cG5mX8b+ruBHaGup3lwBa6zEvz920KISUZcLE0VM+4FUKB/81zZ6R2
pdv7SJeQ6wD/0g+M5JAX32Mq2LjjZHW9v03mMJe+B/BHnkLAju1Wj/5Z3UqhluVTHBGABWmVsYwt
0n8hgfDq14iIpnj5uh0a6qlnAoKgLnJJnkgfaZ/ipuG6THuXb74US+F77qhxaiHvcXUU2sD0pnHm
7tX6u0Y7yW2p3NTUPBth8j4CYDgZ08No+iCsiWzJZX7dKC7lEYRRCfsHjy/N5N/iz8fCDEjvHiUY
gtDFlkHlGuK0x3JF0iQPQTiMuksl3ZPlBUABBjq19hA2cftQHrEsSBtGcWZ27QTODRJ0rP5019/j
Y96wQkwv2fkwcEQ5F7lqUeJJaON+nl5ywuUhOkdbclBvOEyNVVNnwBV3/hqVF52Xu+z+9UghgI0W
uuk/mXaoZczbi300O1/OOb1zMz4wreB6gBBBZMrjyQctzMwbOMzRBgLJZEbOwruEXVhtPNaWyJ6T
WfFf7j1eEjGGv9d4q/1bg+SQfhk3UTjsBClbhKtJGxPIwF/gBJjhkEo+4rMrbEgwcn03s03+6yK9
HD4NBwQwr6uFTBtYI1E5fwEB56S2ZvonugzOd0itL7xVjSl49iWTs9Z4o837za79itjcaUrqQtrf
aWotInghyV6LnHS0leDXLRs+ecdgav8nwmsYto5QAetPa3YUj/yC/syKGYTZPERyBGB98O4nVzdo
59Z/JPt8jF1Xe/davYUq9UfwD2FaJM34SHQZkPTidCgGr7c8bCC6xTK5R0DAYOwDH76aUZZhDdZu
i3rkAqiPdtSMUDltim8/VplhSMX8RDsGGTBxVTVvYo0yKkkoyjYUVNLFk4s8nY8Dw7Xj9ojQkxgS
mjCcZQQu0jmOmvw87AWsojYJv0y4V4CjW5S9nPH17H1d251oo9Fm0CCGgvTUxWJXBizCOR7wxl3G
d+4ttj2Eukf8o5GinOKNgx6Hu86KB+H4Pu1oY/P2YGcjUMgXW1ViHYkVM7yIu5ExWfi399qalfxt
dNng1l2cmucB8V9puVcDz8gt0i1thlcuJqjwdQwhU7R8j/PAslfRmYrj2GMI1V6w1J24mhxGN6TZ
cNtrYX9P78Ihift4SG8VvJqS3OJduc9UobspsFCP+fOUkIr0uZAfNgb/M7XnVpNG3zHAMHwpaLGS
Hjpbl1hgCNQPKQWnRQ5ajuOEvCIjKEJpqB2E3LpJc52kAFVIYHCfmE1mRaH82IJQ+PtNJ1Zp90fc
sTtIjzMsgORFssr7QjscO+9WRQoGnGOi5OpOdeUpZbV7uxVbKcB+eYg+CXYCQGKQgEMrYDXi6FHY
2Ii01bSAsbq5BG8dYmcrWF59ezDvaBS8WFpBaolclRA8G4XHU488Y7AhmanQu+HdgvCkFGNEJPsk
VEjSmuxeuzZLzhEU7iNGunTrnWdi6rQzTinYtapYKi57sx4haN1mxpBFMgVyML6ZJWjIM93fO99S
WhRPdqzpWZHVC0XvwTKPlluY/MdpZSQuoYv0U91Pr8dVFExY7EWEJWJEbUvOXoGAkrDBLw64/8lC
EkJ7WnvB8N+brh/yDVkIH/I/n+ujTTUIAUYKoJMLMn1FRUTZJNb1qM26M/VWEeO6U7vkKnqBRXhz
fdd5oyTvl5/r90/fkmWw6pSJva45dMp05uOugJN37wrDzW7QvwJxKSDI+TLDvP1euYtWrLk2gHvn
gP/3MRxaMFQebqfUspwJrM0E/rBNTIKus8KNh3Jli9V10ZeunV2qGO61Wr58HlnMXK62gRxMRT48
aG3RqiJJ/pD/EMxvEzrvYI0wuW4eBNNeCTVcvxfYXulwIHzndY2c9nBcuER++HNnWUyyDEFO1SZI
NJzXO2uPZaist+w0c2z1Y7OoGFiIsH5k8xaxPHHS+PPSGrueSb9NbR9QweCLoyS1ev+ht3ZGsTJH
dcPeUhTDVSLhozpZjotZGGrIk6P6xKfIkgZxGH70QxnoQUWchZzSG3dDfM21sRwGplM/FhuOVsgg
bx10s5/3sd+3VvOw4hMG004IAJ3NTboN/D+0PKEJ/ZYWZkud/jAxyrwXwMgfbXiyor03yM6i/6aK
NClRykL/HmnoqBzV8g+POJPx0gXGBR8FvSrEx8b68Mg5eFsr2yOy2UJ3JY+yOI70u3BPfKz3z1MA
qgWuNTRVj9q6b6OnMDqGSM95QzAks97KBhXmSfi7whfjxpQ6NT56OYNx12+LpTTAGTR7ZuhLQh3h
LE3cHW+mbn45/Bdy8sy8DJJAgk0e6l/7tVHesYyLKmq0jsmU5od9g3RU2/mI9lXgrvosafIu/ux6
J2rFVzDl+OnlwUgp8esrHAElBYnYAavVrTx47QlsYxg4G6bxdUxuXjMVTUGRZhPKJ8rbzJ0HVpU0
THABeVXzPqOPBSO+X8kxDfGAhJNqe+S2nWqHBKrQz9j04jQfu/k2dnxpwqIuJXZXLb/n2y90kVTo
xlbmVe2y07ve5DE/y7g3hW5HtYXiDDk9+uTTqaex3WbZn6PeHD/2wVYTclHKYZp8MVtG3t/ql0XO
b+3iYiGBHTNKixh6orFWR82RRSD/pjdTIgsMMpZ9a4OVMEwVC+wmHYsNwBco51+/yrrULd6/N/pd
xU7vKkMlHoOFnHQD647+kNvLm56PWryNJJ6Eqc2+DlXtxgpuw0IinlakxPtlI6/Ml5UV8FwFT4fC
1vC5+gDw3KHAGNe7qbFbLzK7KzhOHuKtbNiSJT7PgCu5i+s/MHqQ7H3bjt+ZHFJCY4+lUWC5bECJ
UpP62wDhTX5kJ47PZ6/X39UiXsPOifVD0PK/GCX+iIWXfLCGQ1GEhIAaE40ufK9gzVA3O12Ic8c7
MXluF4DHGz7U3Y5Rj5awcbUHSvJJNLQ+b7o1egiMndumHu1hHGQ+K2ryyIONL3bmbaDavYsthWXE
cFsu+J7swFpAgnxYIhQfhTL1j4x0JDq2Su1VeliB9I9Z5A9kuZDb7sGQOBrqNUAZeKzXdxck3aRh
oY9nv8O38P7qPbucMnpuZFeoc9kbSOBtaCvz2+kdew+8vBaZ8PwNXcpE/JbrVcp6599dQNcpaNzR
7CVDIqzrWKaWn1+vccV3UV9CMXOnVDcZDWbVFTXHPqxy1/xidZaGxyQu1al906CtOUZKXYECDC+f
tf9nBHlFU3Zi3OIfqWm25yRvwykG7BQ8QJpqWbmXAVS4oZirZi9O7YXa90yw7EdAPAsWOgAuqJbs
Lyr8m/Z8238sYHidaXosqR+/TVMd9IG6kSP1ac5K8+94leDet1uhR+wWEmVw8y02s1+9vxnIK8+U
HkGkH/e28JEl2TGSI4k7JqG30tKS2wefoZ6sfV39Fb8mygHpblffddiONd7BO+NpJgYLqKIVxzsm
BhQM4+Mei7VBKeKIFXVz0sSpb7CjkD9KhRTD8wS+DN9riEC5saiBIzplQXLtYatcbPkuhqlk/sax
HJOOc/2lyX3wkhMo1yJscRywZpU5EcbwlL6cYYuaQci1Jxc2vZ7fDaNNK/qaOOXB0y2BIwkVzHJS
DvpFldquzYcx9Umtq+8boZu5sSdc/BnKA4vBoo3kJ9zqfHbmZu61BXfEEuj2Q5wKBNWiNKThVa7Q
Gx626GrGaiP6Q3ZwM13nth62TFYGRXB4jMjqwPZVJdPjTi7f65g9AaJP+5aMa4nLwhOsSDkea//2
YVBIgIgGvXIQkKF7Re7U8yS3/b0EwjppPanzfvelfKlXY8dDQBsp7oy9ojeq1gHh0JdPcc+kcPqq
qVFGdjGPM67TRttfvZgU4ucZDQOgu43y4IQZdPIDv5TUOgUUDIpt+V7MvsJ1yXVsPooLv6WM5Txi
ZP59gaPO1iySeZ5lzN4fRlS2f43VvHxZGsHJgxIZz8kaR5mW2WipG/nhDt3u1mmZhz4KCcuSgPuM
ABoQWSgB6IHzIPyAhZG6z9YtI8lKEJXkI20K+SIJ6TY5/cOX2qvXFLe3FONdFzVoG9oY2LaOLMAS
sraPHyWC8jMZZDGl3qJr1VVUxIuZ+HEXVMD2E/Sgg25HxmEPq1AdKaSDO5xVU0z/ma5I700gMYju
G+VuTdVojQIIXELHdybXm+qcYqpjip7/688ARLz/s1Dq6agGhC6TTSRAc7a1g3abmirHP9q++Mpx
9qjJb6y74Empl5fR9O53PCMZY5QviGSWBEndtWRkw7PxjbQ2mo4rw77+jbyC4G2g4tfi1DDQhMEA
T7Y0IlHCfSW1ZcQCHxRNgfFvUZ6x2Mv7bGzZ/UPMPmliLjHA/u4fPgy9FEIatnBQleUJSEgdfT6T
mNIupKguRuwWY6brCl0S0NVJXZe2XRKx47gBq3jE9SXONugIiC2euRXLttgBHNT05A3a+aPre0NY
2E3FctkK9wOyXCi7OQXxr0ob58F1WSnY4RdcYkN3u8GmuLBNSJJ/RRaCR3VCdytu4lvlYllu3iWs
eF5F4zVJ+M5qGEDRqqhQLySISYnFFI2cSVsTV20QjKKcLHTl8T/7FsJCrTOMSYBtdhLxaSQdLWBO
FI+xnYmgYa9IEKi8aGJ+XxZtEDipAlgHT934cDmWFJkHtQQU24szqoLVoQ9Pqpss+B0J/o4p4a5w
KeiM4WmbAqJMBPsbd2mLFEH+XnBkIWBau6gEJwvz2LFsOchFtUo3AGgDVQJBwVdAY/Xev0rSTRE4
H+5R8mjO8majRi9OXeFnf/xM7AHDwYdGqHeAF3rqMb+XmbThXc9X2Go/ebjpV1FCMS834OXH/CfQ
JWJhDcgcYI3q5Tc0YBFlyVwpZYPdTBaAgn2xiKokUks5if9aaooKXBcb/Ho+YCNgbzEnefu9IjWT
HDN8p4EnYwH1iCHdEAeVM1XrXawzfZTeJmy+5FnsJ6QCkCrwFkNBd9FyQuRdz1e46NeETgK9sJAz
i5Xp7jCr38crejv5K2b0tQi0wKi9rk7+9AZMPWsDpIG2zG3MK41Yzktc3qlFHDdojmFwOGneYqzO
Uf0H8jxDqvtpz87OX4ejOSi5przd1OmJkuibBapRxweJP6RwCVrxC9j19XDv3mwC8RJjnMPr0Plt
L5/xPGmU2/jnPH8/Ew6O4lvsmT2Wpa3rwNehFZATEm5/LwazvjxcEch7kCxQu09EJfb3E9ImnWBa
At3ww13o58xHBAL6RaWfKj796BugKAuzrRzvQ7I4YNRzOJdmHwf4tZ+MIFDeLpmspEnvmk9aBBB8
KVzasec0eCEmNeQI2RsBBiBm6nblswg2I9DYOHIFg5pRNab1x+kiuWh8uIe3Ulw6Q/Upzujx8ss1
8uH7VC7hZkx3OJlRSdroihIzxxVjSsSYZs0L5y0uuK6OcpBgxNkt/TP8ycp3gB+ZqhHWKSBdcXcN
rHgdV8INqDcD/ywGHxjq2NG0WqhyVD08geybh14tcDdMhxHBMBKqbbX1zaEWb5hrhnwXzpMwnaOl
/tqxLsPCRZndE50AzJXao8Y6WjxWekmkICpcw44xevOkNMkYb6JwMgZVSBb/R2Hj7AW3YFl6foKp
eH61HnzNkoZI53PD6fbwYaoSw9ljbxWNVTU7nuP6ZwhyYsPzBQmzp3lc5bR5yDwo9eeCyZSLNr1X
HazjjI8JHywB68WU0JF5awlFYyIHR+ivN2ZzYuOFyCD1NHGRUgIeZFGOe1ZQvF/rsNMUL68bMIbD
mkF0rZEx5vN0WkJnwZ6OUJatebd7rY3QwhNE1GKSn9zSmNQLnEE+c/5Hm+EAB3zdwJzOxcHh2ElL
iiv3w0iNJdME3nQ2PYUGX/u9yahuTKecHKU+MEr4+2Dqz64m9DGqx7kS1Yg6oztJOOtS7FKP3IEO
TIF6FgZXGaS9nqZxMFNYzOgDnfhiXakwkx84syaRbdVMFHGPgaX8moArg0RB2MF1gYEpgUepHjzI
625bd9PDK1VV/PH4jH/pIzVZjaS6sqNRxOoVaQZ8iVMXBXCCQoSlVG9BrPoBAse9bgi2r8ZJx90+
kVGRkqvKPHzKv8ujmnDcIu2+OABnfhrim0D3S5T1VQ8vJDA9U2bbXpiLf1su5kmaP071/xL+UxxN
SSBvsvM6hBfaZ2z9wU/wF+wvOSPGR4znDU+c30Py7PHhsptPD73HCmY2e+hgS4E5lR+Wpfx8h9IZ
jJvBkE/c+wOuNPJGH/by9Xcu6UZ47lNxCr6+l8ltT4HBT8LrTXacMY8RuUqh2QAqqK7hSC/3XWPP
AqDv+ezQC37wlty6ySSS0JpXRBNjB/MtOAb0bNETRtgZfjB5MLCv+oHvG6GaLrb/j8rXM3Huabgr
3Dwfwz0BomzPlTh+aJZ9qwCRGUkYF/MaL0qbw0LhJtZBx2LuHs59InR3SS7OV9FQxyP7+5uEqNpW
6UMWJndorSWtDHWHKQuLgd3ES2KvOJot5CJSiURw/Pg+mpaM/eQOxuJ9f72Z41/6vIQ9/EgLbSY9
z49kQ7ug4DYcst+iuxJm49qDQ7yWl9WphDDsYQClz+y7jHpB53Qcuy/dtoXPkEGOzUYROemusKrG
9higx+2C+fQKEHUSurT0uZUXp4ME5+b8mzqRmL/fpdCuR5hfVy7FP3IlTdhORTnyP0fIhXvKZoSz
2r7/ZmXhoxbWSxJ1z71kpSyYgRGCeaKUIJX9X+WXAUmYRPQFXncOaY/Z6LzAL279hBdAqCfA/tZO
19mD8stmm9RkFy50HOPcd2u/Zk2aJNQ7DwZlECBVFVcBxsM2Yx62uZXN1evORetCbAb4DfmkpwRY
jv+67bz0RX/o0aLATwOE54VUB0lDNDKQGVD7FaL8iF+X6EQap5IBVt2rwGCIRTHVKmsFAzSSuTOW
KQRPRMKmV+65O59cGBL3uXCEdJ+bfSMe2I5LC5+GxQUVIT8oHd7Yyp4UZhDcSEpr/AATMLpQc3ew
HpFxfqf4Po9RfJunPpp0b0/RU9L5yYyHkQms4uPxb+942gPvGo+B9qNqqcKcWQNoqdn23kLw03d9
zkag1O3o/a9H6aMXzhfR8aMwtOixkbGT1GcS6RH0Vi5sD2pebh69N7vo+OUQAcA0UBapvp1FZ35Q
12X5YfXnB+Wh45INCHDHrYbNO8Li2lJutGdjCGmxbadKa5g4hy+H6JEHVOngCcylwXDOtMVsgZdp
cSSGp8p7plmvbJowi/1aOGun7cnnpH0wUKsLqeejfwAG+PcHSwc3clWsgBM+GMfl2LrtPPr+5TWe
OHpOFyyt/hgVfl4PADXpzs34H+a7T/gUcUJ2oxoF+y5VLO8lCIMWKVCFvJrGT2bALddz8nWcoNKu
YniJiKc2Y54bmLpijV3qKgirfDtWJaUaz1eJLMEs0R6eDESrf6J0ZaoioRVc8kiyv79sD+shPI+J
YN/2+TmezTKCltcBa2GW4LHprLHAXNi1ZaVCLgg6Xn/gyKBaILnmP1S+R26bsLYSxr/5PzZPcmuo
8v9MtICCjeR7XIhoyiYK/9spSr80BGozs0Vw9osUMaHAwAuIY0pJFEHy3uEVUmdu9QSdBIJk47WX
hIMmCxVmNhZS5g18+R/s/22BOBguIH9ocDdaFZSiihyO0l3mmg4Iyr8lgBe+z4xXNtlET4hLVgr8
85+Ckdyff6WCz/oZtpWoTvdjLhLRUosUez65peAJMufnITaHe/U57wCv2gpr3s809qIMoVP+Lv+F
8P5Jd/Yr32saWu6A/pvP4QwWE7TZPV5xsTlfBJWDjxKd4EWNxuk56cRIFvIeLivE7IV6drZ+00Z/
o64OWEfSrtaVfh7TjQxy6AZjDyxWwL/GH8o6VmIxpvJBBxmszW7I5CxNgeWj6XeT+sVS+GoNn2qt
V+STyAcVOfyOgyxj0bJ/+4CpiJyUzHTmmesgsa0dIILkCUEV4XiLCPVFiyIYQyHzgVzz+Df5BRLw
sJc4hQ6F2fT0QMY0IIu3wsjIWS5sT9CGAe0+cHzmVRZs17PJJsLICIAOfHJnop4bPAbmgV/KKE9l
d9VC6xObVUGBfksOnBP5dlDY/4HFQ9vNSW5u7PcT+YLZ4qKCOfYokQuoGE0eqnUtfzRJxVNrmGHD
cX70342d2fVVkXh+w6btCoAqytwRWRj3Eh0QALXD1ga8sfWolpdLPKWXUlzam9Ob7nsnOZuvARMV
Y2/LmE88ABkL4ag3B36VzrrYRrCR1NtfS1TXV1Auz0yEYWKtOldvRibo2xEo8m9P2LmLmZyQShw1
7i0V8Pm9il1Ytq4N2POtJ5ZGY4AfdorVDtEcjZPzkYd48aQL4nZkCSAHRpgzE4WlFtV6xkkUv3ws
/0PJbw0aMlHcY+H+f2uXRxD4GKlsd18b5OapwC+K3s/pwvO6PsdWTJ4hsl1kADMWlC8sq1QyfdZa
RNkb6T2v4YwUyw5bWu3aUKcNFdimWT3ETJrFyubrrzMBem+au0hhHtpl4MFki/zr2dWIpwS7kzq5
laAB6aKxae5EXn2GNDKmSSdLtfhFrbPStQLV9Drps1UPRwqk6KN+sK5mtGtGB7cf1toMVW3usr1e
MvIZMWrm4IiIO/Wgbkup1+4ikcGEfpErnfbFLhasdaQrdD+TJfzWlektD1RQIYxzjV0EhBHW+oA0
iwpnijAnx56qAGlNfe30Oat0NdHBERuWWGY95kFOf5Kdbjtw1O5rr8ZsL2se8s7rH5St/eZZ9kvO
QCRPIYUgIlGaUCKvJrnQS2AY4Ly0fw7ivOMGVqwyKSjsetHt0XP3nOHdMrlYZAq/FFk+/qwK1gtB
W/T9a5zaJnFDrBRVOgAbG9uB90QgHAr78jjZZyISxFuukzRTyXqd6DVd0hLeAL/8Ons5QezOWPMq
WpGVeh/juxZoAqKK1E4RAHDDE5zzBgivb3/lUsqF/uCvEceeXiYVsLYVWwG2E8PLAU7+cDwsPu4x
oCIb0rqws0YqXh9uysn3QLys24COZ6H2t13DV9veGbDDXKHyj2JsSS35eD0nPOw82yc3+Wq69kIO
NnYMi2TvcPhM8IxyC/QjRsbBWbtZpJtja7Yw6Kazmvb3OL6dDUyIY7i6d5HG8txMeIW6L1++pLFe
kvzzJuzLFD0P/SmQH0Ky2C68Se1BR3/FhHqb8/S3YF35HB15cMtlGljiJfDTRrgTgD8KZJI3D91F
8PykUMu4jF6T3TMpC4pKmDUFu+Xsb148FYRl1GqJeK67iGYfxQ1QP/hun35Pr6cgmY8e2n9B5tXu
v55r3fMUUphMXYrUFXt0BM/u/QnkFvT/W8PGXTfyc33iygLQvTz5hXv36V6EOYOvh4TCg2dyFXHf
ghEcTQl53R9feUl5HOwoQX46rKsE8IwxnJlksXdxQdUkaDxH6VkBDvCE/EU0t4vk2eYkL5xDO6M7
zA204tQQC1uihjak5cOIxraMluzNJLm1byMwO6bjQXiWZIDA7/Vf88ohum42amxqHg3n0yOI+lsA
9ImfoyoY/aFU3B3B07pbHopoXJycxoEdrvNr/xin1DVQVkPjLxytGTfqdYyjh9OdtDUIF7/bs5mC
1Vv2WUkirsEaMLbQd2aXFWgSbbyskm63RnuZPSy79deBqMyCAMu5sH0rKH+L9kC/QPHGfLezWZx3
YSYHXkaCDSTdmEwQPbmPvNsx2C0Pf0quuoaNKEE/MnQDT09K54rfMoF7aqF/xtGXi2XmJ4/eA9JU
rvRBbZy4GDuhPzhiCo9f1vm/J1PDp6gXJJCiECJwfDLL2aODD5FfJUXo9wUGms47+F2IXRC4MEIE
eJquhQR31eD5N+va2jYQgCwgZ+V+/8C1gloppPIuO/eQzFrhGT+PjI1wFDxknVOb1toYgojxsWxy
5JAFkzvRYGKc5u1lOUTXshRgawhDD1ez9SjGWFmsGQjS9XoTeoCm/JKSo+PO13Mt6syG4IMjVeCn
OfiSQJG3vW9RxrJU3EQ59AtvdjOkdKvl4EX4+KgUVAldMBbQhmMtWRxRSYDV7Cmo7k0x1q4J5N8R
xv5HpOPXow==
`protect end_protected

