

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GWT/RJdN/UcIKTAhVxs3scTnM63xEPkso8NeqXOmx+sudHjUMJ/qSt5GFjdXAqexLlRND8lEfssX
Q8fYY8TuyA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J+phMqmkYiPgvjvEjlpcdWdxzP+34SmYIPyc3dLXEqt+h9EhMcqfQg7r/svpEBV24DU6CyKyCXke
3gZaY85pXANGRT/lW2K8drptf9l9vYajWMSy/HjvETFYNanQN5XDicKd40/UNr4NV+8K3+zJSD2+
6HJJVC0iWa6RgWieT3M=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZrkwjC6jJHChQhf/EDIYzNRopX0ckXH4NL9s7GZmKhZ5Xuu3xV3LqvLjlAq2T+/3AXtko4HEVfJk
jD8rEKHAwLnqMbikHpL2pup+LY4/a45y7duxNC07dpJvYX19IW6mqYLKEJTs330XVwBLE1KOyaGV
xhWwwqThGo1V39JpBwMcpzmL4YnxHaTlERiq7vaoQpYAMkwdoBVpG9MMAn3CbeZJI8pLk/zNkztm
rMeS9pshqNVtzdUse3pl3EDxWMB2hg/4/G9fk9okekAXBV0rv5NMqf0xPrBsTvRJGO21aW42nO++
dC8am+sI7nAhoG4w6z/WxE1BGkRuZGX4CGhIDg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iexpjlh7M7dlTcv5seskQPlqyHreGwsr94b5YKwilWQsfXW7U1V2aK3O1/+pXS09S+pTH0rKoHNi
ofASVdK1RB4/i9AYD0Ihai7zYaqt6eRX7azypmOnO0M/ZZIrM+63BHWcDodlNlh86PWfwaKQSqJW
hLVuOmY14GXZev020lRZWg+2UhI/Cl3c8nww44erkAvCrpxmrhaZg0s2YPKI/KBqZbZHwn0ufJSY
5EPF28uCCS1urKeejeaSBUmimEDyf29zU/xFd0fvevSdWXaFhwjT2mOL7DranIxEzj0yQrN0jiKy
Towa0uazE4xB+gMrElDuwpcw6ZUMyEBsaW08mA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DVPBxTgKjw13z3lZMl+QMKXV/uHfXNCgMoWbgQb15TKXtTCmkLiaCYkk+UNjnupib1FZuwkbZs4q
pFuDW3Z3x3poQoD+4+Z7IIYAmkcV2VNFgSXWGO5qpHWhRfkulPfZcRStTLiN9EUcwXJUsLi1Rwk0
oFaVSUr3p4Mr6zjC18beDCFomH1w+aZiTDmIDtnqdWVtxtresAhXiT6k51hdPESOpe/yPCGrgQj7
cckAkNk0Y7ums+FtMhs5xsfKLV6GQGr8vql+qoCmnMNbYofWKIq3pY2FrW6f7ZGbFhW+vgaVatOo
wR1vGhSucCD4x9efRbKZpd3HOhDW/vOAo1pd2Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uIb1xi/b1sGS9N5+ge4ctTMaXcuHePw5wBb1FVa9aecf3hzk8F8+/rWvK4DX9IjVKEx0PLXI6xjb
IH/rGtJXdtbDJdBaXxCtQZnZ3bb8a74BAJHYm3BEextG398AX1ZCOiiun/unyz5EkREGrSg9f1qp
tvP1wCaUgYbP8iAi+ak=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qK9lK7oKxV9h/658uwPcMAAwYeLmnKNpsdduH0hJUA8HIiT0JfF3YHf9Z/+4sugCSI1ARr9LlbO/
o+J2NPNqOXlyDgJW0FGjeX+G4wdX5LlxdfSIcRGs2vzyXQiAWVbMq15jqJGV+qheK6QIsLI/qwOR
naZ46kfkwSE8kQXhF7WZE2kD7kLSTF5QPnmYFPP1wrSHpjD9hfcjmg2768Oxg74FqPuAHl6cX4Bj
Enf4+hzQMQ+IcGssYzesFwyeHIqJFbufwMH9hDnmz2bOveVtLUI33QRmIvvIjsEuvmQwCu/AC3gG
UyfxcM7HSiPQe9MbxhcS0KjoubQbTx7z04URRQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 504864)
`protect data_block
YKRMUPT1vhDJoaGZHFRdELN4vlY8Ng0BcX+iD3LwL3oPcUYTH3/JHjbtM/jeh7JgPJNY1Otl9nEe
LSGvA1B5/RRv83qVu3BSxEm3Zi8ztDz0pg1MJc/ocWlz+hrrMGjaknjTP0m+CslD82QQNXp3oDFc
L2uzZLjERGallDkXCS/Vhyr+60X6nSgKRjK3fh5kw8WJaGM3CSy+5p08ZhcL+HyPABwY3F9t4SgU
8D210M4XmynMyCactwIMYz2z61PPILI70SZ7q9e9h/rGLBnlpJVzduIgwTP0fmqDH+g3xOnpqkB6
0ggWyngepUylcNzZd74s6kbulY2J42S39G3H/OBq+IcYBLay/lllTlD3Q/J7ukyPmpduJHHGQRty
ra3m4bxj4ntkKDPnOawibq7fhrr5LTbBq2PJ/obH8ZvlnsjPp+zav2lZwReIPobfv9te7a2LFk8v
f4E6K9Fwd/hxd7EKWyNcrhacBdUs2CDYQyBpR6gr4jfLTj5LvlRET/miPnXHvYzvObc6RxqRYP2Y
84NZw8uaIK49m/wLw0CJWzR6bvys5gHBiKKBUZptwOoQxZ8BgDP94HtkZBps7vB5zutrDnDZYdem
5jlM7vSC/yROwt6cF70riwSagzPjydybjNpworwZPPJyFDt1ToEYLZVenwTNx2MXhirgtF308iZf
5sMKqIfUnqvU7ufkE76n8f1DRTNfxqrKiWmwVH/EwbFNtKT3uFJ/PmDizM+F277iiEQ74ZIpLEbx
g+n59m4eqX0DJJDNe820mFOGteWiEjJJhYbvSI7qOBzhegco5b9sBHL3skhYOSP7auNfQMGnwJx/
2Vj/TEvkv4CQXTkBVonVfiPP1wSfhQYSuscpj+K/81NsUP1f7GNquI079vhBV0qO8jSTvF+5Ogtu
Nnf0r0qTLpG8XxK93qT8MSrsNYn+eh8+HGpPNwSqmIqj0k7FpwlwlFDNKGSYZZdxOyt3i1ta75tf
FyZfhM3rFu3LhY5m9rTi24lga+sVMkKOf5YUvGTSzDOJSI8aR6ANa5jrZSaooLn56cX1o2JIiTML
CFVNkQSohpyzdIQ7QrQTUVJkUUJgenTI3VUcj/SJdAGu5Lb7wzGy4fNr5QL7nbmA4LYVjF0yqiLi
F3j+9eYBRQlw8Xd9+u68jcfTW9ZaupXpdgY7bNMembOYjAPaio4TCo6bNJ+Ip3wdefTe20xF0lYG
gN3+61cgCbtBkJROZKu/i7wOoVkiYcw0gbKc+j9m3DMo34CBNgRSbilWpCsA5OUwsH6aFYLZH9pj
LgCt8sFR/YuUEAhWaiOZ2UPNakmKlPnjPwN2oMqazt/6VXizf8waQ+ukJ+o8yQzzOh+KlNMK8G0z
Y5WoCu0Gnm7L3CXvrEN8SWjKAoQAwir796aeMY3av6Kzwkwqg3SjomEgQm8H+PdsibHXz0Ysgmbw
zBXrfNo9VosA1z6gwZUQsXo2Qwy67R5HfL29quTuHdZvrU0dum2EEP7BatKOAUHvx1Hydvu9ulIx
5y7OCmwQLoYp1M9Sy+SnFaPCQZnmseMAxRdsQXDvvXw1luaP0dQqcEjuYU2v1H+ZiH/P+GGzPNqu
Z7kQUAi3IHt7/LxYBi9OZPulJAU/h8q4Pm7PNcBWb/LdMzoCSYzXAO/m/QxJb1ciZooPnXemwV1F
EWCJ0B+lCrpHyRhFoGqJeJMqxpyKcwRYlmOtNsQEVUOHYaqNq6tcNxU3LXe5OXDKe7e5JXNjEXzg
4jUiRBkvRrbRL/XjrWu5CYSxsjKUkgtpfmwZHJbpU8c6Ci5iF6o09FxfBEP1n6ny+s6XgHn/Ohqw
4xQhiD0z1HN5IEr3zg4vB1vkjq86cvDpBndATowWeuzbMo09tWDuF8atawhgT6yAghmRbKmCzmL0
PcyL56DXRqMcpJ8e6PH7qMgOZWpP/gpRPJkk2/WHJ4q2Tc5IG4kUZUZ0VKpATQdnu2PPQqPmJoKP
4aYreTS15TD4IWt84VpNuD45XfA2MPKLTKzVgl4YEkr04IpQ4xRu7dNec92lP6luN26LpaSVNQ4S
LBPNJmIQXsR/WqS7WHRWW9CciHIQhy428tcp+G64kXjLI9xYgEPtF72l+OYAcDv1jKHMrgmAenhX
6l1JEpYg2e+VbJbpVKnnMzsPsDr4mBcPHON3eqj48xskCmPX2IQc8beELSr6ClMC8oAetj7q6RYe
tr2YqwN6VA9iQoOShoBnZzoPjIMlb4Rqgp06s5d3dUOS737//LJHEkJmD8u/Z767UwQOeY87HsAl
M68YF19O+LXur0NEs6KRm/05oQnPQ1DQ27LNEHKwr/4vviDF2jcE2RXoXSOHvqa9oeITyo0viFYK
1LAgW+Ic+oOqkqiPlUIhN6QXUnuL3P1dfpodwHNuPojNPS6AZlWLIca1loMQkXKBiE8euoksMQvS
2hFGu7LWpreZDHpGKJQLccF3pH/uLD6LtuLXNOb+Ylk0txCj9NtSqSNAMGxMWCM5Xi9TORpV2HPz
GaJnfujahy+EyqWWnLwl/9KyOEXMyPRb0jyKPjgqXs65a4OUzfZaTWj301p01eX48OcsoLURrJ6r
WwGu5qH/mxFEIZMkSxy9PwYV06iQCOkrkooh9rt1DyGTFga+gvFHrUeZGhfw5nGLbJ7PTuvAxZTi
QMB/bhiELyCTX4qNnnpkdu77rUN/j3KOm8MWZYzRv6Gzi260UW8s5eXLSJGdX9BP7CI3819ERVGM
enfyql7PzRpNGgiKcOAfUBm1uw2GFw4tZKfc1JBKUii/aEMaaPVKBu5dRxuDsepg95Yo4U9W+diE
IkMMVKAu18zGwqj2IfILKRMS+Jkg5eG0zyUZX/4EmNIaf36VATuxVfdpr/4YfbaxjgE699/bIQ6H
Nx0OPhvTAnBU+1cIvxL31ly/znH12GdRaC/jBpYNmiOSf1T1yY6jSDRm42oaRW1knI31aLtPWeb6
PWpvYDqALIoNyqBVrPs+Dq2K3+i/Dv0zKfJfUx34SY4V2OT732ShhBjxhrC0cfy51FYiv3YvWEGu
Ly9HPNlkp4LKt0D79CFwFGcfc+xAPnvIOQX+vPwNDL5Jj5KaF27z+POxvLBOTPxbmXW1VheRFceY
hL2NYB8IJ+LHAmO/orbeHXnFYVOrNHGfv/QFv8llnT4TVbqkquZnPbHlDdSOdXofJ2gThMal5tJL
Zv3MHty2iHQiiSo1UkFK99aux94j1jQ7XaioRTixlBt1Mq7Xz0rRCSHTu1dNjm/qljyA8rnqNFRw
bn0SJXFZsxI2GzFTFTk3rCv2HLEB86/6uJoUcNIwAyPqW9e+OSvzI33Rsc5UTE8crv777zTY8vKK
uti4P0iqTflRYRsHexVlxtjnd8Ea0qxWtn5fWZwvvR8gvZ1tT3Et7uV0YEj2uAXuejJO5iEjBVbW
4pZFY6nAQiAXuOnYMZniOxA9accEoV0m25xsJJ6eX5Z1nwPXAcolq/t5hNUydZR/9T3VxajyYSzz
KLguUxRYSMcTNYHjwu7TTo3yBnWw51/RGkZ1OUnW/3RA5ph2Rvr7jnQHsnG1bVUjM72U1z7r1N1a
T7OEcGsU21l4LRRwbl6pUq0s92003+oZ7dp7qDNf/nEK6N++xRW/dgPp6pEGWYtDmSvk+iJsoyZX
oARv7w1+M/dttQzYYP+U89sdEjd8K7h0zsFUwWat3k4S5L6S8FqzxBL2fBuOWskXb2KR5tPKEE2m
M7oj8oA44SRWdeD3fasefAgrfkIjKQ2f8kygg4BJDCLhd+xa4URcwb9XDWsWFQxClENJLGcOqfLG
fgyjzRfFhwLlStBsZAOpkPWElx4uVsJ554RtQaJd6ItapNmzFLRoOvZehSO9L2N1sHq6r5Ah1yuJ
TnjPKpj1stPQ9bjMCcav7iOJ494pzbhvmHAcTs4fvCnpQ4F34bzMVcAlNxQN4uyZa7gepooHJPMG
KTVGGhE6ydOOk5xD4Cc0vk5BvZDuylhIPUM69AEr/5SwEBnSXbfyqG3AtxGRvTt9fbbgzdSoL6bq
NAWBT6Ch7sdRd/5qhlzE58+BtiYloSGl83DKQbBUNIc1pT5VxaumZN2tNYIZnkiSg2Ezd9YdPWzn
9lAj8G5PpBAcsEmI2EtofxY/wscSSEpkf1vVHJTS4/UCJcnaks92mRTLu4QiNPt9BhxjF0mWvHqy
AbtcOaNE6TrrJxO3cDd/Gwn2/IgHjP8/ZfpIXDYw7AH2YDbb6TuSoSnbajQ7pKbSiWoLtelm4Csu
p1N2ekxXMCdetaNRVf3xCZAhz/NN2gcJXW/n/O6j0IoYbgfWCrMoztHsbKfYqmPXe07Su4hA/NfF
0+4tK9e8JJQigMsKXY1LtyOnVE8ZAnyph/nwLbDt9qbLWAVOmHSHhdJbTGeqbKQXIpqBGSjkVZwo
CeZv1ErTQRGQEzERPaq3KlxXlKO1pWcg1Uab3JZvm6fOVmWZ5AKShlZU+jREDGxXvLbu82ZvlTe3
nvZTS5keA18XSbWQ9m6CYWnnaRH03TlS0Qxzn9KjR7lfFQvBVmgvfmDb7xyXEgI21ADROzvsIQL8
v5MJvfPi31fZ21kCLpta5ioH5rryJuU8w/VQN+Xsxd82LTzx1XVZ2+JodDB7360HP1p/38o1QEQg
5k27BsuBu/RUmtdT+goS4wGdHCtbnhpN+GJYjLnjZB45XY4dKuTrQwUvET1H3XQR9Yz7wLcbM82L
zNyu0WacnFEDK/qbD/u+kFI6O3bV8UQ3AN37Naud1IFLfDAFuxsDXqUU/OtE9S/aAXMsgoSYC2ek
t9GgJGAo1kOYIjLgnHPjBQKnvvxqGTH6xsfiil7GuZnX7SOKhpq7nKN8iKOetYNRkTEngQs4XCLH
ul9Y14Gm6tsLrNe8R9Li0IlbPUiH+N6ttby0DaPsmrDvFYOj4IogK9wRMWXOcNKx/wlGuJanLoq1
d35Mg8a2N96npoNbU1BH/4RkdewiMCp+D/MQSvEdexp33bhh8Fp+kPJQxFh0qJ8q/HyjsDVd7wu7
n3rIns7mHlgeVTi7/eCKqcTpoYQ10pjR3d/Nhh2Nr963s1ehhDut5b9mBxsGJ/wg9iH1DvUSDtCI
7gKQKMI21vIhsWd0A8qOhFJ89VtabdG3wkqfBpGKYFal62fiC/8YfRogGcfkZtkdRTtq8HCQHkog
+4lVyiU8pSn4pOJL2YwtHbR/QVrVP9b7xdRh21DWywxCahk6A7wujKrJ2G7rgD+g8sW/cXEhApja
EJ2z6Obvyw5Av0jXeGv5qtWWMk/CMyEqQvpntn1Lk/MQbd8/luKk29JF5DWOgusk6hZHGY3sYN0b
6FKSRM6X3wLjfmTWJI4pMLXEmAGzFE4pGthlMTjYPIe9qe2soST5u3cLMRQ1mHbcz9Y3LEsL8OER
+ccZgDZtlMOAOL/Fw2/zBZj0cExQ/wDQ8MdJoINJCd5Yx67YdWIDfUBVRVxjNUuvKewrK3oL4vqb
oSLd4vGDjAwgamonebEMumXV8KMrdQkNDfjk5eQx2/imS0KCfvdmL2Yo+FrTCmly0c2u25AunrLv
MpJuBWgH89a88W4E72IdjyUMbsgjEUQDJQbBauG5DAMaDOAaISGBkwJHeuyWaFP/9ykzep5/sMH5
uRhn0ngjftH0mLH7jKvWPpSs1OXlpKxgVHGPlVtAv5RHuy/HEEsUVdJtPBrtIz9kERut5Lrmzrf7
e8Gy2QQLtSgguZm8nJ3LjoI9mE5gAysRYDveHUvzHKgcqKx54SUe02qucWt35t8qXjwaR7LT4tEm
fFZhjFGFQnQt+nHOoAHt/vTX7nSpNMgvZAwi4Yg1ZtxO1snWMen18PKBz2k8heHh1/qDtLNn/C/Y
qUkWQZsog+VnJtU+6kQ8GRxcxH6T33Se9yEh8MLvqZQWPAe4tBi6lnC8DO3D4sQ2uSgAvmHUEK9D
NfQz4nVZUvrSoPl2VDzwks9ARa5zyPZhNetDoRpSjTfApq8lRIrqWAOhZIZfs6oMAsHO47Rn3rtu
CWIoRSzjAvTzDDHX8CChd6GMBJi7PglZChBCx/tCJgmmz9B0uBkibxABGqPwA81lm+7U+2C8N/lJ
JbrtpW5K+2fjdpfnRrhgK3TR5t2fh1JrvmUrC1WIBDdzflEh/LwVjIBOfjfKyUkJBw1c1QfJIfzW
BpJQ/hpsnzGCQCZ2b/cT1X9VTXnRRw6nVjIndhDD0Pv5RLzLOKXNvyGAvYbuMOMOu4kFQmlYLmZP
xFQspr5XK+Wzp4hvGk0fzymmjEv0ep/XHiSJ1ByuPxFR6DZ0JovEGfA9aIb2kV1C9Ad0BIxhMvEg
GZq/msS4DnPNvH7tJI87BUcbSWJsv6jr19Xzz+5/XZEOA1RNs07MqRjY3KHn/EKEEs5c7LroCiA4
vM7ovtWeXrr5BPYeOtXpD0y9XMlrCi67cGMY7bBXUXnQPBeO7VgTovWMWsqZqNb079ivztJ5p7XR
xXb2FtlVGofRm8CSkvVq5PPJtVYtVO1P4FDb14u0RaPhYDXEXZ6tQj/YbUJNtbv9NTEN1qNiT8+F
0KPJ8wQfC/SWvlQjEKJrpRGtQf/+F6X7SZJPghLgu0c8DAVqPz3cEkQew3FAvgfpZI8O9PBB7Bw0
1CUow7fJiJ5QW0ylSIQLprZz9Hak9Q0h1JtZCGtYW0pa0StJi6RsurYb1GIyorGRELe4xYQJmvCj
y/Cfivw8loYVxaRzOULCjoUR4MFT3B55ltS84Rjb1ZMdvh+QNrlNklD+Dn0neYaNtQp9GvmTgWL3
r7Amsqbjcg7mGDFuoxZajDQZg9teFuIze9gUYh9SENhrb6rGJXz1l5AtirFoSL1tYc+vEHY+542t
ZND+2v78JqSQyYM6n79KW9RDwL5Vxg4lg48FLDY3xASIyConS5QvDAU46MUdUBByNXfYu83S2hTn
CXArS/Ueyb7Jrm6IY1SnLQU1/Bzibo5VvRwoLKChAom41QqOXkFh2S0JKJH8Mi1FqrQALEwKBuqD
A9Px3ZEVwt1C00WEkr8LtNLF6j2Xjur+qJI1kiZgY8oEkzsL6RKbKp+pU+hSzWqizd70fealSt9+
GuxHF507RmaiJS7qLLHv0dCZNcP9hnjKb40uUEYgJPJ0IYys1MgnM5OvOkLmqd5K9I0yygnhaftc
xXCUDVtH4F4+U3EpRHwFeTtq2IvIJTtaBbLVk32Gm1jFBr7bPZVrm6ROGlNOlXW6yYiXJwbiXzy8
4GyISLpJJu7rE2LGIOoGUnk51RUKdQ0roBO9WtOMCDgjAuacVbO5l4cSovmvGm0YqU2tELTPDvNJ
ETHfmNBxYBKkoluxvjQIXs5G8L16vKGNCXde3fCeuGwLgIMw2c8m03u1wNT/R48vBKNakM4GL59H
62nstr23gn2Uzse0VyY5DrO75D1iE/p+jaqRQgK9bxn1Rfp46wpQyJcRc3KB06DL7PdnimcEc8+D
Y+wxPtov0jLP1gpx7+NBUXmcdqYHkohVE1mVK3z/0mAMDP6gdimuLdO1uuHl6si/gfyjuOC9xlvL
o/Ceiy99FI699GebpRxqBu4l+7V4tnQ49RtwQkzLh4vN1vUD0f1w4eCnB9/N/WzSK5UBpQRX7/Ai
MZytqPZfkd/x3dw07oFKCxslL84FOk30sOeaiTHLSt+M3FA3cz1USBsqwlAXykvDlM8E0yANd2T2
eHNpeEIoNuaqEWmYNB+PIt98F3NujCgUp+T2c0g2NW/vW1EIaEGMvZXgQIWaicVYPO/UWe8g3UnT
pzgmb7zg5jQfua9e69hOIsK6yDC6V5vrO9lCedJcRXvPX56Cz1XEcz/L6ycK29mNPzmLCptTLp11
wltO97EY7f/5XjWfJ+WyiZRDTW/QPQAHwhLhHQMNZqvRmvCmhzHhJvbuJMWwDND6z7lpPo9kakth
R8qggXpmAgAAz/iRZn98xnjBawGxtCKppkmoZ1xXMAQp3i+EeTorD/XRiRgfU7Yvn8YC74nLVewp
tE8ylL85f81r7WQHx4XA3ZFRJsX+HBX8cJ6YfrLHYm+GbLcT4i/oDya+mSYGzpmR2vVDxCxc3FJn
9OkpbVCKL+lRz8XodkKDQxjnAtyoxzG6d82tI/o7G/91OCUQMpXOYBsBXe+O1hU3imP+0UeoF26U
w9/O3v5gEAoeAXkMAJ/8fG4spm/NB16TBkRTzrxpD51k/ZrpW2YDLNkRt98qvdzT5HCzMfMPN8mL
dI6dCUcAC4LbD8xcJ12oGBa37zzFBSUShWBqjkrBfhIzns7eeuf1t3R9zQOGtXgqSNveG/wANm83
g6SGSeCVQg23j+3xHaR3QhNVkiGJeo4R2A3k5xUXfUjJO4wU7xtn+r51ddaFepfZ8xYEGcGjQTSz
0e4qlYdxrOcycUVVkZj7Q8Idf3Ir8BOACGMaaSoRGUftzGx5GvrYfm/TQqeXas8CWnmS2u1WUkJM
OGZKcsfoTL9ObcoKPzFmiQVUfqw0d8PLL2Dg29e+hOoyYaWACgb4pwJqeLOftlYix0caufGTLdvW
YHEIJgX6bRGQYx2tY7I4dzs+k576cJYl98uAYmRF9r9F4e6kwK9+/GvmqGaQ+5h8Lsi4FDed87FA
q6ZBdwv8yqtqnalPVLuzZDLIXmYJmZEJY9dO/Sryk22AWPMn7msuHlRiyx2yAZpW+vWatWbobrto
P3Ezd15JujcBOU6fLa2hYdktj864OO6lEZxRa9Zxp1eHHYYKS82c/VQ3rLsl875y0Hppemsas9RJ
qVDYT+V8I8cpaHGAI1EaewJ4wMRwfdkJ9frEW6jfOpE9X4Cx8zjZ7n0GAKTkcsUg2M4Z4cgDKtEh
RAsy5r9n0E/FLwLg9aQjtsQntFzY0NWFoJQTNJncMg0ptoX5fogsoGnrGV6XTDpG/xTCCH8W2Og1
gfbC3CX2To0vukkBI7NUS9bjw7uYdY3JgJT1LqwJWZwECWXralfs/9QadFHKFarHHeU1Cy8ZeTrk
99mEkWwdQVK/A7C8LhRZfiio2gCA4MllZhjqMwkhXD8vjcG0s7Fw6VoBoPydg6WrUQ4CX7dHCz9k
D+Fiok/sMStsZr0E3aSoq3X/hJvBwU0SzRN8ls17Lff/Yrbf+LRkAH6M6yFnfeIjSrltLazNEdpw
Enh0WhZgMKQ6qqNy85oRfD+5AS+pLQfFnDFOLq/q8UC7isDWapvbXEIzN3+hNs1jkClCXV3kRHy8
y7bd6cALHCpyamjvd/YbWeyVyIgc2MsyZB8ZrMps5T+aj06CA3yaMLw0xkYj8D45z3oimIFib/GW
+pUUF2nEeRfIh6cto6U3921HrqrDmp15LJCtmOopsDX6Av3oxjvvY5xdevgO2q7V8dpWqIpqgziM
lC4t3x56Rc0MBlWrif0HfihhwBza29au2bGJwJuAVoXDq/DA4wF8dovTD6B+VGmLFJNlCYOZo1Ab
JnPInuN4EXQY1jyYL7FTIpY5FkhhzJG7+oEgsaaRiquexe7NXlt4N+qVpdXI3S60apYSVpuzAik6
dvgDz+4aDHBuJJsKf50g6a2dwNaAUpJvR6c89KQoBcubrhAYpJWF2rKqsYS2DJ7IwFOqRncRzYH8
lE+7TTK+PBApdeMQXEUqlhLzWdrHiulJUaNPpGhXYmSbPXV7j/v6hfq4sfnr9UxekojCG7n+0aO7
suf3xVjnKhoGHIIeu/PUN0WaysCKFntBsGxD9UXEhD54PNZbgPIOZNuxsbl+c5B1nunfhIgXkxFN
04sa8DDsB4wb9zv/54gtO+fO8y2QFT9N3n+QtxBOkuzYPcFm/TSDNEU8ovL+oK7cmZLE+xEMkCcS
JZGHf0ppqpkAuX654XsE3XNlTX+eR2PLWPCPXp4/NSiykkegMeP31/XV5HEFXATaP2hn5+wZtMIJ
tV1uaFTpHy6zgA+UcomNXKuKknwTvZgs4AQAw53iujF0dSldx7C776lkTEsN2k8f0n4k4yabpuEX
Q2+L2gB93ecKDxjmZJOy8Kw1eqr3J1lY5DFbqJigf6t5RuRRv8Od83zSnbxxBTP0w15QnC80YEUI
Kep0x/sOQrnTaUUT1H0fUTUtEeDqtTov0npnKYVk/kQ67ta6iyhAFC0Rjbh7o3Py7L+6AWRrEY9o
xi9XieGaFFiD1cs2+1DYBevyW+RHQ3hMsbNZkwdXvf1zGAiO04RLAoiyTqDSgDbDhXOyRUiMEb5+
cbkih0Vjd9dDcn/R4iOh9DGpb38Mm3vd++2+xNt0aTB0oXmIBA78sWX53EhyvKpi23srlP5gLEI2
+NJ85hTm7daJpJXKaweapZoTka19L3VOBPZwckCMBoL9Z/ZmbnyHD6GgSPHGLCCwdJ9rlHs6qA+r
be/zWU5uw+B85I+Qxd6/SIoi9rImy4euTAo6SxjPcYWcL5CdHzVdV9VWm9PKjXHbJ5VtQUSyjncP
CyUbFwStWTKC/RlTUbt1Z9Gg/LMr9wVRx8R8pmgcZH+4YASA/R/5uXih574/dflRt6xvEK8iex9I
pfti4XgrglilR9l8XgLXuRWcs2r58ERQsRgyNsdlolKBkPEe5vRM/jCGFpTJZ5qSJME8xGTbQVdo
khuQ9BbflzaibBlPXRb7LrCkyRrzdePCa99ZDjOnVgdbtNveKmPxRkSL8SCqBWV550sHN6jMOQoN
k5qxRWHzOpBb1rZTduoWfnZYP3R3O9zkNyIQ3p+Qp34eD5dzFyvVdDk57G3kWbQe9GV2sH3He7lU
UTtiJdGp0Yd7EA4PV2DXmIk6G33YjmgaLckdBq+qYdIzcCoiQUxXd9hJAmaLsgVsolARNMR8NuOo
yVZqIuSWBDeYulDv1+xPYhrQdaXOScfrt0EC5mCYUtVtBz6m/lPw0C8NZ4l8vR33KQurbGN6JqbO
EhlM5887D35camgpkn1RHbw7PB6A7BUG5Y4++y0AJ5UiSNU6HEvB/fLVuE1eI1I7f8AT8tE85CW+
qT4lFOXYTj9vQNPldgrgF9OGocajeE73Nd45z24z13qH7jtWR5Ua3Px9R5VpVQkN644QeIb+s+Ps
1rta5lXIDgVcSXC9OqKqhCgPnB7uk/1U9Pr+Nh9hqxNwPSVgsegxAk4dkECaIDAtZKAlcLDxqO2D
7x7Tv/VLx2qRldyzREWzhTtAjdYsIFuNwbz75Sq5hcV7UQI1eoG83gvgLrkiZXRCo4EbuCfroRIt
AEDnSidM3NP8UUbiHTaD9J083T9GUQDFY2QyhcecPMemrHLojWMM9a3swjgGgyLG0/N/guYPwtFZ
x7eJZ4NAXLBIlTxALOirFd79Q+4E9UgBmnDtQXIZSgiJN0qdb4vV1mg8H1WebRM5j3fhHg+PAUo3
oGZLxgBvrgKLUeoEzETdq2x4JOkhS1PRNxzHOGlqv2PrXiqwwtwCM1b3pbekKbRsnHp/JdCFL/Rm
BTWB9UQegfdstUL2cM/WTzzL95raCED/5NH8WYuHAIZclk3DRWya/X/3l+C3MoP9URnCHFitN557
Rdsrp85txLrILV/4iMupVuGkBlqwzFbvRSAwwLrdArRS1stt2MzhxYpa7JlWpJpfjWLqLj99bPmG
is01DFb3f8cZSSINIRSw1mPsD97/+/KwKdj6wzWKyzNnyJSJgB7YMP7Y1FfOwIAHW+U48V2sSu7R
Ru9Zq+UBKwDWJqS71yXUZMHDxpVK9W0YHp+EFAhyWRmVNCmMfucc3DwgJVxERUREeuRSegeA+e9Q
h5DaVSplfS8J53Ecu7sFXOkj+3aMruAXvQ5lWwcKLJWSzTv4HRaXq1AGiKeumiS+IEFpTX6MYxgk
x0O6KDUOMVeYv8pi0yBzYA3gYae0XMIHTyjAkGm1FEfqdxCJAYmCq8A5EdUKrS96KyGddMjG5qGh
BriV8IkOdB73sbw/YV/XH36ZsMLYR+ZGe9PV3yNb0siU6ukZyD8afpuGJMVwAnsKnz8LT9+8q+Rr
Ldn5Du5JG3lUR3LobmTaDmarc/8zvn4YxtsLfXTBKLmPlof5AHKKebQgDSJEow8PnZ0FJdqG/gMs
Q0kDkY6UWh5z48pGG07V5C7tRCC+zCap4uzDTQhldYi4Y6cagJij7RCoesEWIxZvJqa+24h/9Isx
+7nlGlXcwJYdygY+3iTcgc5CVjdxxB3KfTpZoRt7QFqgVK11t6nqKtK2Kwg0CvielV6lNa9bXp8J
yI+9q4GmELQnkWNn13Sezgl1RORQCMHx/RtcGyijyKXe/ttZhKOFwFYeZRCrz02g4IaBMstLjOXQ
GrIX+KkVZqvUqyHsJ7rcNIPzmxfJ2kzuVOOy6ExJPTPlRfHzEYWZRbwGVd3KUQRw9G1w+TiG8JV9
cuLwx1o2hQuCp0yxtcMnSvEN4BRgGCvf+lFPMHI+TI7edKL82cH5P4uO9NbRezAHr0v2oWz2/3S2
zt8Yswt3ne8zqvRjRc4sI92I23/fjd/VYcRm4h++gfTRfL5urvby+vv/bBXhCcgJ9rYByxH9DfFf
t5oUrUUzp7Ob5whR/cWbNwvq2nEaH7dLmVXK7V/is0/pgkCVWgyg0V3Y7WY4bpPiw3oMTqMSfSjP
OHoEfl5tNvjls9D3alFwQ9Nlzni3PnKI6iA7wGwiGrrPvWxI3L0vh/tucOluGD/UpC2r//GUtqLO
NK/1aJiOMIO9F2/7YvEDInQbyLB4J0cJ5Hlq02MIcn4UvOIuzysDmczyMDILfwJRc1UM06m088VH
FKOhiIRyw/xkE+StDOyoABj2sOfcGHwn2Eks2QcWZPmcZP8voOOjn6i6hPgwkqLNimCK3Us/wNhB
Aeh9WvQXSa8RXUV0xYPQK5a8KUhVGTXSUYGuEvH+wrkfWFSmYSNC6OKAHzmQnfy95Ht1wp10bCp8
T4yjPtcx94zpwAmbniAMr9vNnp6MZRCiHih0Uqddh81SNRk2rIvVOEwYD2vTj7fzKoJux+rEVNxR
g+24wv8Jy529/rarv81m+tk9OBbM1qQGtKc969JILsqFnKt8a9Eb2a+Y8YmWN4+hxkR8Au4lJ6xZ
W2lsdUgLXnflqK+nwQsDXZkKYi8Z6Bv0FjuXHg6LtFFEzxW+bRghI+d3DVgglaYfR+BU/+LT3nLp
k0jo4aNlrsufPh1rHIEjToo14hnvYDz3Wu8JxAF/CCGsagWwlfLcSl/Ip3qXQWk7pWM9sBAsULKe
kxRBxzAL7j8msuglY1dGRzwiRDu8LzdTslq9ARoeaXQMGCJ8MYb00Xtvq2o09GtrQrzClLHnT9Tt
yG+T1filb0iucpd39rXfY1+j7Gq8+CgltR/ehmh7Y1cmLjuzcwMrNjho9EUeWn0pTtrveCpj/Avd
pWe/NW4TqsQAYIYupJ3Fyk4uyv3CdLy0AG3n1nfCIaZvX+Qqxd9YFv6R1CWhL+geP4ilYPWpPorG
hMJ75Qz07nsms+fLcPN52YcUkpnXOpveoseQ79DCkyZR0J4mdWNrUcfShFkV0Dzsuv9oC4zLgfGs
atJmuC2wMFgn7j6xpn1HAsLcJC0jRWrbntm6eZVI0cFZVlWIcr8we+f1Dk6pGpQECk51JETS/Koz
OVhywscALcUp0VQtI2Ieghnoy5GNmPenx7WuVS7AkuPlB/wUULe8UAXL5oqkZJiRw9xZcnHQL/nD
bsKN82DMDZwYZl0R8m44iSPsHPe8cSLF5mGEU0W8bwhLGHv6mcXKIg6SIPrGl6IrKg04nrMKmEUt
IDXbIafOW/6f7+FI4DKh4yWbVDe5tzlijbK3/VoLA/2sHefkAg9CUv03raryaalUZYcYtQkuY1+s
sb2qab4Lxl+xIqbQvu6LOcP55PTTkni+IEyxTAeI5PgzK8s5derLrQuJbdb7MJrzwK1v0rvRe/DX
vFa3WFScYItVm3UegcPdyfImR4uxWZPx01fwQwlWwt8Hi+MQI/iZhqqPVNvY0R6ODnPbifElAW67
sP7DJokoyrXDiYTTnMqHlRQ1aHxI75xusyjy+KiZBX0jyyqzsXWssSDbeZOQasR324bzNRPu8PFH
lMYXXRnGsD3Y1pZ8B9RboE13uQkQ6Qb04az47yZmt2hZL5QaONl3nXaMLaJ2FsvJ7rlKP8EQg3+Z
oth3ZTTJW4jZlLb/DfW2wZcROdHqh98Z5Six2rL+2/qvtVgt2K290x1RQpziRvHwJqZEV30mJHe0
ql9t0Ryj714Xe8qAWVAkyxBFzgHPa/C/KVw5dnOswHS4u7O+CQVxUBirDSFpvmJZQH3K0bl/Xw9t
lAf3CkXCG2gqCfSpUU3ibilvOWOCtnNS9H+jXEXshpqrOXqoB9V3PKm+lJwmfH0HBv++ZMfO5Chw
AXubVsQ3GxTCyP/LtgZa2D/YSfI8Aq5WHCpgqH168YiILVtC5bVWEtGhvqnZrRZA6puFv3QnCfg/
QtZqPspvD/1GhATfEMeRmVeb67pSXkJwpaEP9L9VoZSdWXS2YJD7p5ZV3F91DUlrqGk88EIKwd1K
3KtPUmB6vJuYmPiTR3ETTRAts5oP5XWN2DXLSH2NFHqLtbg8Ck5F4XTwvGEuhauPuIDLTRl52HbR
AbYfJF0tRG+G0Z2H4wJOoa6J/V/mvCfWxeD6nWnKGYnwC6UPzeAtFmXW71re1obdYtpPVNHG6QuQ
ZbVWnrU+7n46qBkeGYpNecBzC3y63RiBAQiBHz8F4aBy7QYxqtWZpJ1ZDXahoWBjWoCfNbbOjLXL
tbyDFH3ETRABmQDEZcd2bP7LyDdvATU6SMsF/USyzfoe6tXUaPWd8SXTOjV7XJf17Hfh7R52wiqa
JOrxdsRLw0NViQAdRkv1WDo4lk2SstVkrOaJ/eQjRN68O2ZZMF4rKREsP5bgDGmM7aiFgKgJ9ifD
/SCgQGBVgNOSFBNEcYz5J2aWCWbae44BVakB64K2tSQNLY0zghXgbevc5UvcKl5q5Jwzh8sLopoZ
fdIM2Po5lTEfnh3I5ecW5xsGSj9zZ+Lmd5p3dv6UIvo3r+iypR6JzHY2ObW80xDYzlmSyEz5bmAN
v25FhzkBeU05r6+8YugU9T2USNKD8G/BOpZRWuga5zjOvPd2ifGdKir6CFtQfVxtFvbCeXeT9CFw
FEauu9x2eEzmu79QEhUzmlqQ0YygJ8h9ZFUlOZukDaEGzmc5184xPn7tmk1zTH1V4C4BI9SKmS2D
M3Wv9CARHV8U/ErMLj0zTFknGiPtepymUeXZ5tsyBoGNLKDiuOJrEKw3uC5PNHUlwaK5wZkRW60k
KGxcj5SE07eE8xZna8n3hCF+dOcBze/r1SohCqABebDHtBvRZ3/qTsJMRrjnvHVmvZOBNkXtLEgA
6czdDlSRkAPQOZrBmGUCn6288JIX4QFpnPMPXx1E+S/u3HxT5QpaB9IYjfLz6fgD2YRNO7ofefGt
hKn84CV419vTDaJnNDWHNoeNRXNiq+6sVYVHwcPXXRS4DaEhea5+ElHj9NZMdUDdkVO6AQUedZll
RuE9t94Nb+PTlu0RGqRC7p1XWNS3vevhevY3vdChuEKAIBuF0ldxMtegEgidkJld5pUwjNWhDbmv
W03jOCwpWcBv2hIUMUq50mo7Kq9CrgA2Z+JglWfgMCsCWiz1u4vNVsoGHFLC/VuHBuB2OC0Yj+FJ
qzrqVwAOW4UMW8xsY5VUdkMsAd2yL8+Zjsm+WTVeNISZUQjz3jfQeyGUfa6YIEnwpS6dzLr4xCeO
FAbEmBsbGFG+nEWka0IHGmSy8okgXD8A0q2M88J7nUnzaWhtI3fbeDqY5NR0q8wEkiySC2ewkn3g
AeBHSE2geoTvfcAUU7VTyqVRfA6saN1WafrKFBBDIQdjUqW9Rtbtm5daaLfI26dWa0aGWdGyQgJw
imswV+zcTB5huu67Q+MyKs9tPpTVPOB/Fb4rPEw8VXQogNdkrAn7tHbRhBiF8Zj/RUKEyjDql53b
BzDhbdw++M2pG0KYlwjbYm86Exek7ZDr7XSKYArDU/gbwPODGXgHzxABlS1JZuMAt/NR0g1WhXhm
uMtzDBG1F20XHh+iaYvnUvIUgT4XBWVj6YeADpTastNEudCspHKGo3RtNYnHfq7o1Clr6ZNZRS6d
1XJ8dHbStsJehu1Iy6RPeJo/Lh7CKN25EFCp78dPt07V/bFVdWU7+pDFg89YWlwhzvTsZ15oniIg
vpAt5jHahtagDKfbcGeXqn3K/dlQm9wTg3nPNT6qpJBP9lS5AF/+refMSti96zERaDSZizbItzhO
JkdiD26CecxqT8qdGQQXpm9kF6kPzru8TaOIWXO3OZgsndZcejWoJLh83i3VBnHZPH4q746Dai2Y
h6Vw9rpz/8OjU2baBVMNrpiReit1BpAUPDS0tD1zZXf/qL5+6eeu0i/YRvesjZCyg9UOU9PpHmzq
+ANqm2G8Smf0sYJMBI5XYn+NwCHKPZ1VI3iO1KWw5HMGGeWNJfkapEsRCQfg4E9C4k9uTsOlIGLC
iiHYBKxyNpy5CNq7FeeYPs+TH4fDOktcA5Ne2WOdQ1ygs9WekKsTU1c1LGCZVDHaXG/Dyv9gaaDu
jI4ym8s73QkxPMpmyBCn+7cu0pChKvjPt0b2osU9wuC0VJ+JxBFSigRLymZKB1/4AUjWLaUl4d20
vHIbQZyHMPF9/T61r/WigfytKSNfxgLKg4Wc79nbbwfDFPrOkcH4RkEDTZouABDhvAxyNRUl9+ch
tMJdFDZj+6wNpFlZ7XFJIvRBqJOktPhppZnw1ASVIkfcYErfNvIBdFYlf3adjUgAg30Kcbkvul4J
WEetGo+YXvxP0/4Fumb1wShZll3lC5/1QHSlCyHlLDxQVxnMOLeioxc9CR/2GYN1suKsRdaudX4m
hRz2+t0s7i7GAaq4Zdq1SerTD69bRmhwmotuQbkjLfCGYBy5T8pNacXJhm6EFuL2Ia5vhvaOjSIE
htMFCofSDHhEkSXW+Q413lrO2jzgbPMGH8UfimbTVdpOz9eXkEYqJ2WIuZNZZssmD7IIdBBcz3Md
hIzBTt9zd0LMnEk1AStkfi9CqWXK6vFstOuXNstgqEumUeb2GS8NJoCDIGO/Xc8hzSmlBksu3Q3n
sz8lWtfmsI979QN3jO/ampUVVitGhsRIvoNQa2rELJp6k6/VVhYuyIsSx5ezl3Tz8Z8fPDGkl7f8
cRbhjmlQBIjxZKYVg67hMaFHd7xnFsv9KOWaGKAi0ZQLmmwJst3zffeEQA89q3g0xZFX2/qFVOTv
EqSYPbKXieEUsDyI3E7tInhRlC0cOQvr3k5KfPkrlgvyl0hJVrh3lmiyohN2NsSl5kKXV1YvFrui
d5v5wgmxrHR5HtZOc6HNYVsEJ/6Ijlbu7Bs85TgO+ypxGXU1Rjzo7r9HwYK4/Mjs0YsMFxFohbwY
6rMxNBdAkoyFKbeWDDDqEn/akCyzbNIyJ3wI/gjyNLhAfFf9NJpUEQF3QYVdU4nfmg2Nc/S09h94
VIMGiNHAEoEDw32rDyK4SAbfuI/rhf2Lmy4cGJnxSuqqApG9bXyEfcLTwbHkKqpUYazlRTJKyeGG
kNJN2T9zGdh/he3HKvz7xE54rQT5tyz0RnPAYaOEY9MAb79vBMgy/1ZnsY58uGc/wJy4HLlLncZq
+IeJ6tLDdLIiJlhAOGnoE2B6TbNsZVFhUqS8svsSJgZDACk30vL9WdHCvh6W+gevbwC2I6qz+8LR
ybjDjWl7cAhbUB3bOdRRmL19VMmpKyEPwRKH/cz+Sm7q25h9sHVt6DETkeK2Mu7xmlNtAvk+00OI
ANkgpvj4WKlRcN6WV1L2rMVYquIKTUOQ9iTxG4I1ExlP1oNM+EswHBIonV4Jvgy61UFVtxZwP4BW
EXvUBJN0dDrZhXitMDnYnsT4o9AIC1QQLwFAi4BGSqIJyKEXq9oZLffJ/nmCb+6RnXtAtoGfvbjy
fbH/abYCBZUXoj+2puNOSQsK2DLMjOlSuffLuJns61fcIKISjqEow9w07DmIRKpC8t4VjxzxRFXD
xsjWFF8+ehlhJPuK7sxFeMF6WQ88Yqh3p0k5TZZdDKrUIcdBuKmQ7ZZG5cPSMkQTlSK0EN5dXc3b
P8IYwiOJhy1/LHEDh/uksoMVMgkNmOhQgB+GnnMUU3D/LHgU2RK8cx+UoswpY5QIo+3iUNB7JfA1
dtYCIRfrMLvgLDQhVQK7ucpIzFS1T9CKnkp3doYTxrSm3r8f3Slbw+sKfJ0kIts6o7M4PKFbhnit
gEDaCON4MAi6/3kwqY6B4K+zfZqXkZPf70JfItP3pl4WBzIEBU34QobGMi3KUgQ1AG/69okLd/oy
4rdNZXB/BOXxf0okNhEx2NJB2Q7KaXMCzDF51cl49OOtMWBZMIvzWxwjHdlCUg1JnZaARON845wp
QNuQSgasputW+SqqGOxYd3nuDDhLn7YR4Wrwkp7nvPS85SLfbiIAl+D+UXIfm0AhihrIYrm3cfzO
AwgeKRWzycAp5OZFMU69KE7XgwMyCtaeEBzPO3plDvPf+75iLYcbjY32s0mnCA0KduzFIHsPDxZK
2PYVrx4ouFxuB23qPfqUzN5Vyz2dqLvxBAgMu7/SLDP2zey8Nn8fe1yUMbPmoqitOGJxLUZoVKqs
I7o2tVpD3gfbCUuMQX/5aXfQ5/xq5UWWmiGuPOhPf8h6bdayIUSxazGIaxrVOhxsb1kXpGa6DLgo
4WwHKx04Tgg0C0BeIdm9OadjhUgVgrDou/qV/aBKuawitgoLW8PhE5/49xfR95+yssI6sQ0C3oD/
xaTprnToRSClB08OnJxdcu+crRRVNSk3lshLMVaFZRaCWnY4BkDHXl6hebpn5shuQwp9D0IL89Ls
J4nkqgxiZ3qDlNV5jvVZcgDKidrHhgNxAGhh5T18oQdtr8dbWoLFTV5rmZiprJp+s3iOA+X/GbXS
JfzRS5qKhtW4CGAwIvywesCdsOCgZoOn0FXYaBM9uJU+Hwbm4eUB8te3Pr5VAZ5SmArsVhpFWVDc
OKoRRAWRfKo6H2xwftsautYz0e5pdsp21CvCo3oaS5kwQ70WQDDyeeTpMjdH1M61IF4YKJU6/kKk
7BYzs98UJ17UaQWlq0xncqAOnGfLtlBFDa/TxKpNVfIWQMPoCQ82EbtoNomiQEI1jcqWrSjbduIS
xWS5T9IGyuDRwwRH4czEdAL7RwXuBaPaTwU2NcB163sXwaNbmmUHXnsj/R++KRo3rDxrE5X5Vvy5
penP6/P4o9/MZL0UiTQUsnYUCkEObctiefayJIO8GvnXAo+BBn5oYiF704kyYuX67H+ElccX8zTy
3gMGnaCz4WkggbyXDBdMwBSNjSzXksNNcATYQlVkXzx3QvDAJBK0daCKZQ6bgjUl2JeZQeAgkf3P
oZwPpnMOHWx8UI8L9a4ztFOoDE1aNFwAP5yutdejkWV9YSryFscf5evzRzpWNH+IZLcTTms8o4B2
xOgSvwQ1q1eT6HAggjUflUazO3+X6quz5WxZcB+9O7lkfnIJlzENRiT7Yh1c7lzUDy8iaAbrvhUa
XiQCaEv8aDSmYpEj5XFYCWW1zoOVlT/K0vE+vNJv19Pt1RUTdYqQAFvI8gq5nzSD/av07Eu9VZxC
O4mGlE99oBUYNPsjNRUN+451zX6OM6QxdELddrOm2viE3cgPlI++nXRhGXtvJQw3h4z/W+B9POhL
9ijErBkXI+yH/hdwvT6lPhveHp3qWDp2V99ANu1YuBAIiWpmQOrbnCGmsIGihSVXo1XEZ7d24SXb
LaaxwaydelL4NjBUpcikaHnM6ZF3BF0gdtG5sGib9T2WSC//YksnKHZ2bNX1pUBHWPrQnfdnBnqv
mObpjx/ZoiIGjZOO0/kCRm/J0N/532HX/EIYGh8CNngHtChSuP0ULZwntM6JaRxjq0fgS/LW5w+N
5PlFkDfCLPnXEtzzFYfG6G9O/2fRAyxPdOftl4cGKVSWRWSmAYl0LG2I33lFAeNUyFlAqyPraU06
POAHmsDYbYJ2FlTGLaK9ezaheuJGqSOZjehoB3FFBG5+ksigPMUoIFH7EBrzw4pvvLkfakwhMMSb
YsQaI7i8cOSJLyXHsCr1ZBTM0VK40LMqZOf5TxRs6FRUMS0Pkn1qSGeznGh0z5o5p3NZ5iTZucb6
jUZfVK+5Ae3ab6ZWNMLRb610Je2nvnvUF4wTKb6FWBeJEMrWibyD7CO7Bkv+3PQLh1bBakVBnJc3
XPOaYaUiZwe4evoeN6++JojBk8L5SMhcZvDNW+5+gzWmWJfg/6mI99uDQYvp+mX73mVcQLSGlQDt
+9Lln/FClOpOFSZr9dK7FNlqUJq/KNCKOGDjs9GPcjNgWZUucH5tLEClhbhEBrahPFXLAtUlfPfB
WNECi2xWqdWNlwnQ9xIBRkN+/f+mif5wHqLdTaRjy6fsTZUnYxFkkYIwUbusVhUI5pFSn0FxMTLe
6dpUCZk6BeeCOMyCXKUNJ03/VBlUTi8hlCrDwqVIxzIC9CvaeejBJbPRz8+dx9BKZ9E2OeKrIBt+
JNS2sIAUOnzNYJMLeisCoQDLTbdNP4x9nqdO6FVoWHoAKSnw9Rfrs2e50n5q0NynBwJsJIRzoNlJ
AjIK8X++FhxWLFWQGblBxEz5kb5aRTwOUmhneG40Xwfe2pfYqlnksstLoEHUoZlcb26Gu/1nlqZP
QoUYrT/7vOIkOT0M0vmKv2GfGEjG00uyeGEGnEQAdYQHnzvtnqzDJRTKK6u1n//szIOyLXzyuAu9
H9nX+8KKtsDboPZHU3eoDLpHhUNCCkw/CBKOzvMuYLVuNN0R7i13eAhQPIiuiYqLCqeuBg2ymq4P
ld8foFGL7JOgnDsX3+b/LIDkLoCBNrMFB5FSxf6b+nCxqVQrhxdBg2ACoLTX6erBq19G77QcXbDA
Bv/UQAQV5o0cAy0shAs/uJ96fTe5foa1tt2cUcv4n56JRQGRO0HFQ78byLAo5OAtCfvpLp3+Vszv
Wl6EEm2xyHIUfLujK686o+jIBbLl2oEh+KJcbuzIKHf9Ifn1GxM1LM5Wss+nQOdLjCZ3vBVeJ+iY
pKmIrRVxEhhj2BzbuZ0gCCeHocoLKBSR1yGgwrEgwegn+UHekuwCHsDn7RV/mC4ljE1xULOFulbX
d1YV/Y4fqi9S6+oZiSBvo6sQR89Xm147vkWTXWcwxTFR5M1Yej0cUDlg4MsuuX62Xn+rjFUt0bUF
DAyUtLyNpHy++2oU56vudeTn6JTOjlLKwwaz2/ksCli6DxSbOtB/R0p0HdGxvmNnJbc1UWEfJ7Qq
6j+O7YWZoVIEH87VnblfYTIBLc4fZDryvIVVQx/Hh/xlcON4kNNdFAssDeXV0n7byABj9Wy/FdMd
pmE946P4jxaSReY4fpMh4u0Vx5IMfs83a0O+ik3ZC6rUqmSR1GGrbwFnBxENPMxf0rJ7X7c6hGLh
CUbGpDoJge4EpJzDwV16fsvHuaS+zdTsDbkBR1WP4yVb7LRKxS8y8sy+eTxQCpIT8qzC2TVSXAr1
3Cuh6X/iKEvRZbrcpkm4m/qPKCXkqkMwttPbj+8oqVO0BWqtHDUVtcaRTea2iI/yydQu1cf0EyQ2
4HVhTwGupK51FkrSUYnnpBXNzDUs44uUd2m9L7LiAW2fjFsDXEjFk/IOEYgM3Lopg+ycL7bof5DM
Ulg6Tq25iq5FCMKsPiIifiyDj5orVSr3hxKFUEg2R8BrBn57SzyZI0R+mD+aFncbCjIqOoHPN34o
w6voNl3RM/tgaT+UxDKwPvFOXrLSFHEU63Xz63R99pCwCfcKAeAh94WyPq67IZxqtcGYFcRdXMFx
anTkssJpD1bzCKjzohafCfPQBmbhzWAO4cgpYa1rnAb/QHwJdkBNHJ7LVcrCUg6hhSWtuOOhus5p
JFPHsrem7nZDBG2rPBpJtw/GZ4Sg9VIaaCZmoLl9zG8og4mUg6i59PeKZw43mmr1zdfErjTZInMj
4HrgSecsYfRZFtvamqo2WpudJkKk7vdPFvjQlchRjhpFVxw/Tfv+UOdNXWu8eEwT9BBa0lQsdEFz
LManCPwDZwMN5ty3Ox+CjeB0flydLEFXeVq6nPhmFbo8C0I3TQMpabtL3fxRlR0Z5YvTnJ4F6Db2
qamnKuv0NxudT7Y2XOxOjr/ye4vlPg+eMQ4nQLkQK91uw25mz1YWZTjyarnCtrd9cX7KXuDXesnh
RSk9SO8M5k5cySFf0+HYeSgOqIeWgSkUS7ofT/qI/OfUlnY9rpHvkaUSFfSxSBklFqDbdHrvGwmn
z6tL3G+e9qvgBHJiUi2AHNmqEEdofXYH20TOwEhXJF71PNgHi5zp8876lGfmowUlTdDbYpun4cXe
YoqtQ20XS1XVgxCEAOsUN42tKsrfkPfU73npXd/riy0Qf6CX82OGhkdMtFvqLMdNsPeNW8MCVYI5
GcZ1l6TOeuPr2tWgRHxKFfj1TPghVjYPlf+j12+wXsBvQYx5P6HeB7aWF9gBmG0fnK5NIEc1vTon
25hasjLR7pTB9dEDa+BPRMgzxzElNH/OvpR4yzpuZNKgejPcGENqZ39ZpqhvEsqT9nWT3SULowOB
O1+CeB4L3IWY8dnlsKYsfNhpmHttSp1WCjNYH8X1zfefgAfTvT5pX5LXbd/GX+4NuIo4WfgMSTIn
4SGJT5YxKc+x0G6TSbMGPGe6s+s2NeYiW0sHADJGdUPUz9Q18cW0G+AR7bgTr6e4HQkNjS9pYCYh
/QrieyGX0CNpUKqq8vmsvfW+w5+pvJcZWLZYwqk9HlA3UdakmNMeFBuV1mQeqlOYX0q/qPi9gF+v
lkRi8msvfnusykrRIB6WUVq6ud5P/w0ARn56huF5/vvsaUIYwVlSPXLd+fllNPQx0P7eB9yDejld
Zb2zyBfc4+zoge0b0j7euQwc3HK7Or5ohUkMZte8ZZIKuD1Qk7YO/XwOx8aaQodORzJeFm2D72nQ
umWZbL7RmhHpdyOMtCugvHbK75Ku6/hW98HMF0D6aqsWMERkjBFuD+OiLcQBFiHLi6dAWqfEDUNL
1m/P6UJmQBNguQmYR2y5Vh/TbqPRTp4KjJbvktBIqecrekl8QLqbWpws5CgdnekBioA8zeqo0Us1
rjc/ZZS9WdPFjMfYDZlhZia40jw6FPoUfnupNWMBM2RpAeAzKbhFg8zR0eq0LMXb6LSptGSRpF2V
H8jf8HpF3t1/kIEWlh0SybMjxkwqcyWruonlQ1h+SS+gyr3P3psJ4zDkJdfSYQ5RkGT0uKY2kfnW
RbCaRG6v+cP7o3+46/EKojvsQk3YgQp8cWIFeYQhoo+oAe8xThh+zotxmIAzilVdgzNW94YIBSY0
HPYyCLaswF8jBgexYPlJ8p/ABfI3duvaPZivtapd080kV3uwEokUcjJtDKiLmEhALW8+r4hh3fq5
Uo+3AGy0Ba5jScA6mtc1V4IzRA/GhCpRmKeiT8ap8fZRuu9pQTUsIeT8lWfxzTYFK9Yz/FxnaaKW
3QjoFUCDMPgYDfxwetVGDNKQMT985IKZ33Qnt4Nxp4CEy+D/Ta1/PH2k3CA0gSWBPnoNe8ueMiga
PkEG5Ku6WpmtfeyHS4QJZQcK0lbvYOxBkgK92ELZxlfwiCTAwm0kUP2by5M9UHFcVaawXzyYtIdA
l7SsAR9Fb1SMeeAmU66zASz0qEIYvLcZh/VOLOuJDZEMSzphYpqhvy9jEy0W70t0vaoBT6wrAu/g
IK0soPxQiuNgNxgeX34gHzsWUT1gQvQQkeNERymLK+lA9BcmmBpWugMpiy+DG9cNL6Y/vcsdqkov
AIzjJhQrPLKvYDCAGE1xkYt2qpwuFtnGwAV7Sz/fIAnMl4+mZx7q4JNGlYzA/dhtx13nxsHhpKpq
zxc1T1t81Sqvvb7wu4P/+Sh9XwzpsCfjO9hDXcIPQl/lYYzPCQLC263KavdEZd4VskP12DBzCxfW
fYZ6NBPJ9WlZf//b3oKN5/ey7K1KcFcZb3eUquXwndl4idls805leyeKJF0240/ZkRnEhOhn/Wmp
Cgwq4ibsukOJYRLU67e2znt+8m0PqCWYy4zafSExlJy60DizIzkBQ7p4CdaIDgw6Kd461eCeFFXi
BSPg3yu9hL+afn9Wh6QedcGSUiRByx4nBwQeExxLd5qjSrsTYLcxItM4eagyGHd72UOB7hzZdiJt
SGXND8eeMxvFFijaAuYJs0zEiY4SMTbLjfrJpRZI+p/sAIWZtqoFzkBR2FCy9YwpJXguUqvIbPjL
Tr3y3WS7ynb8ILBVIAAsQ/I1DSahwlUP/BqP4ZxUFT4sFgtBs83a20UAG2Nj4Lh5Va6LakOtQHsL
cMGmpmbJt4J/KfX2p81IyPgjocYTAutmtyaQte+vPCjZB3YLR8zsgeuy4jyREyMGxlz6OvqE885O
sIOne5acv9VUNoy6iyUtz1vrLbkYYX9vm4F0uZFQT+QA2wmOhybdIhkPI/Ep5KKSJYjqoDUU3ToT
StkOX2op4woTLFk+Th0uh5AefeD5KmBu6zAWlQb6+8bOV+XwS4Hg9SjybAP+wJMXRg42ge+I+QtT
VOmMBP2Tv/orEVuvg5ltNsIsKcso+5vvBTbzu8RUIurJjClZ+2af5VhjqOXmlczs8zQ5sq4JFuop
hoqipk2VZf+Y4cMM9DHlkCK2k1sxCRlX6tz5Z27xuF3yI1OzgYbkyXUqbASr+B0YRxirAOIHVqce
6uFADhipcpQYUb90nDrhhi9Cn1pO3yG6FEILA18ep80ngak18NryKLT3b6Eq4yb0UqqR14wegd+g
/xHoXjsWUtfInSqjBDnzO9zoSw228E1OttYUlkIVNXTFezNihdPDsBn6lXMP/mcZSRtXDlYl7om/
+82pqoOCQSLlg2jPaVnL57Om21s2nUeYjPIaSed3iKr3COQRXQ/s1YFnz8vCW0s0axgLFsz2oPZh
QnFypyvseVBr6tTFwFPEoEzaFsQxvv6YXtSNI817OvxeU0bgII7vtA6zHtdrMUM8G/YP0O1/Lt2i
QWkpqKv+JpXgQoRMTOZctj4FmuTxNI/hAbZtO4EjU2OyLxA+Ajy5aVksIPou0N3R3DxIihpn70xl
NReErXlLlhda/CYIJpn6Ezzd6T6xDNI8U1apUcRBr7Zn0ziAYWr97Zkjumt00BXiWQMDr67cdla+
zgg0YwfWkWh+nDvfYt7Hq568l0pUBHjkVy+jhy2ZWvYMn2ZbydIvD0EPwTi2LksPULfZErby82V2
RKcmw/8HJbvwiTAq7J0f22gQ0WG0y30/ZDdoOCtBzJRFXnYgwRznj38XQ8e0EvnIdKAtDNFsPmEp
1K9VnjH/tTWAiMWFWQqgAUXuhMnho83olcXr+sJVym1adoUoNqevAt9TZelLcih1auVRBux4x+WY
E563hmJTF32gmV/mkrev19LlCH7/QeEOxHynO/Wu9FwtyB8saTpLK/Mmj2Nwa+f8JdI/6/h1+yDL
eeam8YGfwyQlhAhrBq8CMkiFZWxSEY8Rs9Z8fRZCB3fgZS48Ioq4+Pj2b4P/AF5V1B9pPBCF0pwG
2cw0H4XfI2wlRks+cG54EHi3YfwfA1tvoEpcSnM2S/0Gp/jc0qHjWojjVUJQR3dYrhByOVO3wFxP
0wpJHxo4lWxwC7SDUZGgjkwA/d4CTz6eDC3dG5o0C+KrCvGRp/qpXT0Ecd9pyIlUR2XyQ9QqlaBa
is7GSB+FBY6YSLlxONlXgHfySWjC7oSNwR0t6E8c+OoVMMrx2sSl/NBz2YW3GWWA8VZv/TL+SHRb
oXyieZyRTYKBgWp9TDzlysi/isCEbiTRD8K3jlyGjMrzQTypGknMa7LuwjYKHuK+EhgZrBNLN3Ve
5Eze6S//R8b1GBCvqY3/i3GhA8RvxCY9d2Q7D02PfncPJDIuLY/0B4qqAIcyKsbHWqu+gP4rYBLz
Rn+vcP2NoZJK3fRN8AZPam3Jr61J8Na2l02DeP6g7pa/8HChdZVbPOsV7XAAfUnhJGbvbZ9/cQeL
n0ZzyyP0x3D73aUEiol4+JGBYEJ/zMlfJAAq8w4UWGjRbZ31fJIHyep7uh5AXSgNCpWRKfXP59ox
9BkRrOGRjDoMcnHi3GjWjdbTxUaEL24aPlknivfTOxpm0BkOS5OcobPGOmEDUzIElIVKhtsn11kl
ih54Gry4ygwEfwJ/gBRPg2RTLgYOXYCUsDJnnXvKU0iqgeqOLKxIs50BdPNAfnSwo/u2vIM9K6cX
1oM2qBkj/H8FDw9YJS7YkVw+0mG74s6l7zvNitUh+aJshsxy5mQ/Je5IRygu5DAuMoFDQfVPSwkv
2kWidmPoGUqAfWUphZIz+K2sL3kZucVk+g9Uyg8aG/Xd6uZAP/ja7HX+zTtvAQXTIUDR0hZddQHx
j91Y7DyqcxFJWv3jgAwP1sAPseTK+zezir/EsdsW7hPCQWl6ItLqCrDP/8teT8ojy9zdGNJied99
MDYPfDDnZaVzATumAm4QDZ+EepRXovGyVcM9M3Uot+f7pnmSA/w4fTgqKW2Z0YWxOU/Rf8Kxr0vR
K8WJe3Wq0Rd+GV2RgCOBlcg0p3Xw6g51AYVc25gNpsUKsi7auoYPjpmlZuTu/oSSgTvNVZtUXgUt
xCpTShtOzaHs/mKpNM6COSg6rEh7czwLuwmHNt8GGqFXPHsaBRQCfUlEffH0UGnnDjKuKQA48dq0
P6OQCKpp4wDE2bROTmZOFrFxnWe0862DdFzWO43hAlEN5fOTQM7IXcDVroE5QfykkUqwXeIp0lXQ
zLAHzG/qd6YYTQEK/I7UqNrpTk7by0GJZ9g30ks9lrtB0kslX27tnQf6msxPSmyBwudnkSXuuZhF
LC9f9JKoKG9qFOmPoQ1LDAQT2mK8JxgxNaLvI/FeYmlFtJ1Zgvqpe0o4DunkaGIMyKx1fVe62pLd
yXiXNkj/Dt3WpCjhagOrtljnib1EMRl1NZNhPabPqT8vIXi2seb5dw4RJz7HhchY+cx7Kmavv30V
72vpq3Hy5YD0niErwBemXA9NyW/zOf6fjOXQc+hOj+GcG3tTp094vZW2WJJ46m7G8SpkH0jX0sgQ
JyehJkNtvAEyw2217vBh6ko6ZlbbzLCt7NWDk97+yf0sgWVEfA/A7lMqphaNX2DuF4y7NyA4T85O
LrwtZaH4dVqOr0c/cjVrkmPBBVZ6LAlwf8ey17xC5QJadw+DRSdtosHZY3W1DOMb9ed8C+/BpYir
IstCsO9qZiA69eYaplQf7Pj/SrzMnuigvTgVGG0y6zh7QEWIy6+quISAFuc2KumK+wDDrQrHvOlg
o7wq42C2q7w/ODbclWpwjbVohynx/p+JbWlSThtWFSA7PLMSI69TmTjmJXlWh+y95ZSmUMctKfya
SgR9WLbQfhND9RuFqJs2ngZdvFIa8ug6+qEPirNR0sNggg+dwlkSfPIsFxEkZhm+FTc/1RdgzltL
l0WmoihcAGyz68OctTn2uzOhsjfLGg3q5U6zAMcG+sm+UzIouu0YFFctDm2Vw6eXgxKowrI43RnZ
3qyTWIJVBqTLVRlKwz2ss0d4ZGRrOPvyrSxwKskg74UV4SV7av9CpTOorye7L1WgTodSu6IfN8np
xoxG8j/VB5z4yh0Wi6njEE2mpREhT4L+77aHe1MQZpQ5+gw3D8FRuZhxg++4DwjPODpixvVUF1vp
pjUjQn3fVSrvKsKOIQVeqk7GCXPuq0KESUCGgrZSRsABdsqU4SyczLm/8NAvEOMhZUqRLNKKOgwT
KFTfvd8uy1LzkgPcWVpCp8eRIx2R3yaa0Hqc3e3PWQuCP+c+FtKCx11adxnRO9lWcncdN7WjuuHx
QzvJM8Tag+sDSiX24I3bvlZzK9TWigiRglWgiGBHBNa1yVtR2CIcM0DgJAcwmjhTUZEqCxjrIbnY
oJyYsZPTWGZkMODTsy7BWAIVFtSWaSA5PG7DVuGDmQdwt/Hb21Go8epTgwnVUZ2ptMZpAmheddHZ
CZd0pSlC5tK2n4E+uHImN5tZFz5S2YPdSdIjC7dFIUr9ZA0dy/g4rq/bgwG0Kfjt3eeaNbZ96xMH
OG4ZQV0B6nA6LtAyi481GGbTjt7FNLpDwEBHg/ZKLRHm74orSnMzVbrchZaJArjWA7NuVamN/o44
eQer+bq+3TEG3aw8PGeo+preX0VpWHGljAI9jOB0RgqcKmXnWDr2kILW+qIXC4jZptQkJ5Y5ENy9
ACbXuAux4F/yobotZdFrop/CBATIEosMX6EES0sJTw742LnwPZfJK+NcUI337bSoPDlt4AyEKc7f
V+ctlHrn/T3fhKmZyPf7sAxdy0Qzj+ch504Wa2BuxFYTQ+176VhEmzWklH65Sw5ilmy8edSF+3P/
JPN2S495lookLqnqlBiZrnLaFMyh/KydLtOq3rc3wI/s01K25M5g9zerkQY3IbEXmAgBWBdOfEGT
I8HQpLyfrAsOnGDdZ932kLQBg/5UnLVr+oss/Vam1OrZYcf7GoJXAMJxKP+aOMu6mHeJWYDs5pAL
P0IN5TyF5z8ysO0vDrn75jNAotUe2IqA8S8Rh4m4aPrknTiwF4we3nrhO5DjG0UtOhRsmyzcPJ1B
K8VAL1ah6iZFl25Z3MW+xNOBegoTqaGh+Ebggl/RLbUKvhoDXOCtBNmU6RPBe8ry3o3J+RCDuYta
U8UBy7+KlTBCoTdBxneig/e3M81N05yDrAxHmih8lFSd1RdYfF6O2UcMmCQQn5WtxqUs1rRcLnT/
Fp7dRl8f2TAbAW6rMJfxZTZ2T0NslRUWtiz0oQ/w9gD6Kv5Thvv5gBVmBEcE9Tuj5OHX5gKRU86S
zs1TzXoqgi3fCmaLxlUqnLOCupUWZi7RbZbE8F+kWQIljZrO+THXPHwnrE2re1wDmNA/M+E6fLNJ
w+0lT1b0RoiAKqfo/LH8OnpepaKrQWp4jnAlzFWBI7zyIU3cD4IEktyDWGWb26wlgGv/q3f/3/BX
pJPgxC6FvZa4ozAmx4nur/evPcsRdf00f2YPXDhmdHmpuWSWshg9gvBBIMZl+BPT8A7ccW0cbwyC
AryXiZAmOBqAb5FABsaMhxil2paPXli0LLgA2ZMEZwZZzh3oHdIwzUXzgRaKtdem5+Xz/nuPJBP8
kFk3n1x30A/hke308OlJnAB7luYOoa1Ii2htJVRneVHTz3WM3CRHYMaVtJAxINx1cM3ban+eC2Rt
Pr6Ep/NihRZBjF17ANERrjmH7/UdSWFrETPnBFyqh336u/2Dq09FYtY6HCx+QL6w6R+4PaNzEQj4
wKizEbfiAvHHUC84kMscIPwyo/sO5RxzrjkNUh/mk5FHPvAYD1iRiYyZKP3cK0D7z25ljhQaWuQ1
J+8ZqJ5c8ciHPcRHgX4JoPxCcB/+b2nGDK4BlnJ+gD8b+4D16l3V+9/HAZxqGQd7oZmS23DIbLnd
yttxemwF4+s39UcHOEIeRfXThBFu+xFPGhFmEj5Hp5pMG9K+umF92YPxQZuGILotyhEXODVe7q3k
qdzMVqRBd9HH5hJcebeZXRKb27WctxPRu1epS3cq9o6/RsL1Mx226n+fZaYebexrS/zXM+9/Abgb
I4cpN/dyRD7D5o6kbmScBXarUlrVlAJttLCozgzGpMRWhUnznZfbLd1T7xRNojEDvl6Peou+SdEQ
pp4S0s7i/f3hVSUYXDmMJELfMdsoqy4niE8+9u7Q4BJc4I/ZscCIwRmmI4/OXRnUhLH/Z6b89/K9
x57Ft0fBLxJqll6Eh7SZUtVMR8GpPaWsOg9Hzqv305CM6K3Ks4bGqQfx3miCiHSAEd8HfCpmlc7A
uHX44jSblgKLuv/YciDRRirjorjlZcZPuQX+EFTR2GZjGcSUVzWpDja8q+q23NVPMcPxBMFF9qcS
2vdTsF/YNcsT/pB9KxKKg4Y2fQE8u49hjacPfb7PvBVdKSTCwakpwQK4P4VxSG8NP/pTNVG7hKiG
P5RF8t8N8a7Sq0FQ9IaTvfwhrg3O7IFys/zvDW5s6YZ7UhVxwOgLCE8X2BtaB1WS5ipmzio+rS42
31RQ6qT6Qb68qG4ofNtb1N0JIZ13cPtYNKV/0nBA8+0JgmzRQpfrqNoaISXdqyIudP/VgeoBoavb
iJMXU1xh7lzDVgFMvC+QcWmfZ6PWDaaD6pdBJ8FBbRLu+K+l2Y9wm5Nmg6KSFLkWT8+RriZBYIgz
Spd9vLH1Jo+c7B49rnX9WYhngezeXd9wOxqlqKDFHUVqnDA+WMcwghqkqhVoz0lZseZdTgURvwfP
IvbwYzfPcYz3bOIV1IoNVewXxCVmIbT1blqFgaJP+QI0ReoBIo6jx5KzgJOYXxHWVIhi3qNHIJdw
npSvz6q8Y4lawyxCXmG0/4XspIEo2oKZCfI4zao2lA4wTBwxPAqIFVNjyJvFy0l/MZk3frwieTBv
mocGlaPDwrC0RxFwOFoG++OR2dX4WjUq7UUpDW03gyJsNZx0bzYTL8rxa2vaPIoaANChqZBTwrBf
U5kGR2SpvHIZQMlnW8n/LKQF7V7qyaRrVI6Vp3CynscdMUopq4b6tuS2xwWbx7FrEOxRv4kivEGK
9sYqQ+ShbHxVn1wL2vzVU6pzPzfZaaZtJJsWNyU7W/3mC8GFLSF9JnloFlrWAsOb6d0kLNDBNtsx
a7AwqFSfgzYBBudn3aKrqcCdSOlwaVSk4Y164SO4X4F/Itu2YvR2jnHAv5UpPWVWiFXvJm4Jy/qF
HOkWhcdwepFT/if6MDkzEIb0qO12dmf3LtVuY4svyEzHCDNLku/ozEX/HDRFgde571nq8oIIO6N/
9miQqirnyyB7wZROu7Y4mBxJUFOv4DleCOCypZRf4GrjZsHMMlozYuLXiqe+YL3ZAcC6PIpJxy2V
QmQYMnxgqJYZt2l2QDrzW5n1YEarTWjk6abPkvqRFdI+0OW4Z8inmihljIJ5R8SNARJ6dW1T7YXr
xmi4TXvT/EBaMxOOMsS2PDFYaXhlB+U0CUXLuvsiISanDayjf+aVsZKDG+UanRYg5ofZAkng7O85
KaJ77/tFCWGyBXDoRPvkdTtbF7PzUv+FSVTthEEwxOiTeSCzvFjHUfO+sfbTs/J8HTWeG+nlm/7M
9CwUG3XrfOSIPvlA2VUSpo43o46CWUClX0s4sXFQaOLvSgJ/7YuMp0bWs8CYZsnjKth+GDscKOTV
NUwRvzZVuZ4IFeBjBdskh+kvwyCu0fLLR4ER6QjgLvbPYCr17euBQgdUYhKhgFcXdti29Ne4LYpt
vd3ko1lV3kz83Rnfm+DW8uR8Nb1CxX6btBs/9VAqVcaJREaLE4IYJT44IMz3dv4ZJzfRIQgzF4Q6
3gxBuH0yblUBJhD6TnMTIm4RBUQtN6hcw5SSo277Zwbfg9E+Gc2ccEXKboHyXXEd+/HsD14Q5CXj
1akGieOp7gAKQ3dI0yvF8JwRnkQvCsrxSb61OcvIWyg+stmsTquGmd2m8LpG5L2McQzqavnyvgwv
6iBDbKJW94K9panxPkBsurlYfzjkxYdXBNIdMj96sW/e8rcI0WMqbQjvN29KiFSepS7ykNKSAEka
hEj3XVMPIbQu6TbfyE55c1aT9WlKNpJEZrFBcvMrnY7onoY3LT3EhbNV5SCFXlbv9yd8kO6YRyLb
6/vgvA6LRTyBRHQAuRl+BFS0Yg+GqEosG7FNOhy57RbDhT69YI+j/zWCCUXCkVFg7o0hM6dTZ/Ze
VIbVYPkzdETrUTpBY9qzvlHOh92nSN7aIADYOwZYI0aYU6jXR0IW2hrq6zYheqBzcdT8rWr9Io9D
uLx1HhKWxza0NbTTE4HlKKOQqd0A3XHg5ntN0Thk5A7oZOrSbPpGRH/V/7j+ZuShKs3BfAK5V1QP
aCuydnRkrmAOC+s2Rwe08UcSiWIGNxmqiYk73sa394WRMFh4fJd3sCUSdn8kxbRBM5V/wjfodvgG
UvNH+m/LkqaFP6LkjmSkMHqZWI8FOkaDSTh8HzFGuzXz0T6yb0tHiUwIH51ZbLU+dkYsTGFNImaB
cnNjc+nkfMbZONhCt4W23r6SN0bgxY1h46yKujCcXXsaBmI11e44V5eYAFFaPYfA/uswqft0vV8g
W5vrXf5w+If1h+GLfn6VYeMl1S5dYIZvmzYXitxLyat5wONNqk70tKYWBYMg5qVE3HImk0ag9F/f
PXOW0O0ycLtOlFVVlQLKlxbqDJ34m6SlrbtVLY2YcaDOY1wDYgXof5kP/OD/vkKePb0Cx0HWIW/F
WrOqaa80vTrvhV1x3nKQyVvL+QzL6Sp84Ptr+PpFgej1ZRQAYyf0Qb575elITEFvpuGjEVwBS6aP
C7l9pQn9TWoiBkv6+4Y6d/yf2eUUZK7rqIhTURO91n2+k/o69Wu6ciJvGxdk0DJOdfH4lcmGO9bu
RMFFWjXkB2WaTgtU8fXxD88PgkI2m3OHcMAPoZs+GK4MNEJ6psMedTCfdritHjePmbwyVMMOcb0u
/IHAhy505dxgK+xGNBVMYgJmyYfsN/foBs0xoYpTiaLtpqT1GNOOwWA/vV4g68hmNhTBpVrMA/qL
AyPxD7NXNErXyfXsnzSerLbBOpOdhdeA/i36bFyQ9AK0FnnrNR9tDKrX+37FzqBe0+sluLpuZjhg
/6BfuwRjUcQK+wDDTof61wBNu6yetN/y6UBdnPSTE9JArSu4mN6V1OUuRXRGkwLWdMRpbI61WGAh
ceudO0Wm3lPIdKIu9o13yFfvwS3JRHQILYb5kYyQ140jDJ6vORntCWglnJ4aIsEa/iw6FiWVjfWd
pWjG+n3Zs8VoPhjgbYtvWtZauSZFff4mPk0MZ5kZ0qBpXMjxeeLZU189W10wyHiDvI3C8HDxTW3t
Yrk5DDc3jIJ/sV2yHcsdLqWS8O8u2SU1h9A59hjPJpMuQXU6Squ75tckeNZ2eNDdBn13a3Ht8Xbz
Xj7WwFGh85CRWo62fpkcbiXIYucGoKMvnGLshgEUNCnsjqetn0xW9vguorVBiPikfwetZPrGcNZU
xFEvoj1qS5Ad6rbdELoeY/7f9TXyJw+Q+KUqBbwgrUVclgbsxWJ5pP83X9rPRwIxNUF6mHccmj0f
IAdfsEuLn+fm451h4tz9aJB5cu1n8oseR9GAVmOrHY+GMmknU4ZaIDGMzxAAD6wXqmkCw/wSxwb/
U6uUMmIlWGWYHUsysnCHZBbGJjMDFgGeMSMT9oj9qcesghyXtZKEjgymZxPF2ycB2u/OwNecaylf
r3ynyqNI+c3D9wJ2/dRuRkayd22YzbBCV0TV7BwQj7Iqw9EbwuUu1I3VjAX8b2PiFZYBB1Mqctj1
pmYU8R0ER3dYxZFAPL1REjPdF6pGFk6sBWFCnn4HzTyIxWT22QFjJ9/lJ3iGobK4PmfByeWy1JAY
+blB+PEeLmqGQxg0UI0Cr/vzhKFqz4othDl29aZXyGexIvcXsqsxTU+AYyzmL6UcUjOaD7xmDtBu
7dEiV4eFYk1ByXWgoazzH0SePp7/zYiCADnwGThnwMqSdBjZcLq03vmQh8E+e233pjsxeyVtJ8Cb
W5j9+qLEPixs1h+9b1RGGcKV5Bf1eeC4CYsvFoTrceFkSSQ0SDRKCCk/do/Ipste+oCzc1cI0Xop
FYx0B6Iq5korSiNtfxLlB1GiGLH9Gjsx7Ey0yLagvpKvtWrvp9cDVEApuY27lBRM8SFhMs1zHJcd
PdwYXLjg88+4YdnwajePFYEkPN7XgnsxcbqACvrwqOQw7BWlzCRAE0l39ierhCn9dwd3JBBYicvE
QW+sdtBbjJiSvzcjWmJLwDi3hsf9a2PXDDRAvNqDBzfyHaAAeLXnpuBjMPq6ccLQrye2tiLqQaSV
xI8erpt3fHUXzkAZOw92/M5137qhmULnghDyQ5zum6ZGbgb4mxSOdAHdehRNDEzw3rhlX/T7ueTj
Um48HBFwAzdk/HRJuui2JHU5iVY0oE0kIjtY0czl3Q1YuiZWmjQLOdubsKOaF+kj6uZE+dWI/RE7
7YW598/lww7lVEVDDN0JdPaoaJ6yuE2sgBHP2gIoucdBOOL47SfB2RpLWCj0FgWcnG/jUzhrW1ZG
grNwgrdWRrECNAStDFs5DN0sBUrjeDGgrCPDvrd7P8neBOe91k5UmKfu+s5FnIF5io1EAtaTTEfK
zwVkb5QQyw3TQYCXOifFr5w0xQ90psFHR4xQT/jgzZ8euCluJ/G7o16ct3N5x5kNLsJYxRo//8VA
QEbQKWqJuLEAu0Vwz+pVbX40NaenLJ4QqMhTobNf3RQqXd9/q39BHqqbFuAQ/UkXoNeOFRocIKDi
0dOITgGdOvSGIk2jB4E0TEeZ6THy9baOC9FkZBLnZET1UsN0RJddjH6KfhfFcjfD3A5Nu6JwmDHY
vYbazBBVV+BOf4Vv/v+U8EOysjqE7HZN6l6RI9HUxYYAvGiGL9aVhn2FQ+8LqrdopiLMvYKAJc59
uDFtZkBPxcsQeUBkiudXqy7VkEh01I4dzKfHnTA9HTxbjb9tuuh98+PxcNa7tX9qxJCP9thnDyeT
irttg9vtG4otpM1cYyMKwHJ7jXt6JtPvloFEsx675e6ZIgJjFWod9gLY4gLr7tV4u5fFNeU/iCPf
RrFOUrs7k2+59HQ9bfj+y5+6k17vvQ+dlp6s5NUCECiWZBRtXq0r++SKZhDZ4r+S7QNAFMzlExoD
1ZTu0IJDOgRGr9aLHHi5jj27kLitvWiBCcA4Bf12HxNVHMp7ZVsln6Egt4TotgcQOgIA6REth0PX
27uWUq4wwtJU3DhTiZUyFyfXUJDx++4ZsRmXjnwH9gxcEz3+EBxtANeULwZKWWRBp9o1dDD3kxJs
WyMqCjhXkpFBBZD/ScErxiesV7ZEdRkiOFttOH1s/V2UKJVTcEziggbvmcANRw4irHklkE5WiKD4
Wi7QIBnWt8fLf8nmYwNH/rve4ipN299FPKW+OrDQ1kANk2haA0W5KcWsZWzKiKsAsvkmhjBuNr1/
tg84xDN+Am2XJddvpqk7x+1gCIZj6ZsdhZP2DbSqZvtL5oyh9yWPnLJLq0JNxJM0QZpeyoUQP+B7
XSVn4oFtLzCf2G8R64hdBPGjq577KxYMKzjdOmNxtxAwvCRC2EY1DNSD2p1wR/NOyqAN4p0F2Vmq
N0nyEs2zlS5OnoSKSw3r0MRq1C0berVmfCjINGpOnNz3B3t2PX7raHKML4jNvO4LbK8ZL5Qsdd7h
AzDj7j3GfZfDzA+aQSpWh4bgF8oRU4mriK/H6qKDUbCjkJHgFPla9mZMD6bSErPnml5O3uTN6hhW
xG+yco0HrEwkDKdszu9gghxSPd/Y2xZ484eUXlCPsIrL7L1WHczdN+9194shlBKA2eyr3FoVwmvu
5XpxrakXN1qOdUON03Trhrmk7Yc4MfzKtzweXwJUgLfnLL+Y54EX7J+5pTK+iaWv4kpjgggp2BqD
HGE2lg+7JB9Ftq3YE1QIXYRLZgS0TZXazgjpEDi5KsAUF4X3gViavn9/RQ3/Ava0t5E8NFpLK1CR
cLZ5GdRfOk2NkTnn3F+7LfCHS5y2mAtPUJquODuFpuJtdY9hHCKIlt0sVgHHc8rfUZnJM0iIY3rd
IXHn0C6P2OgOCYjYc+e4Sq6+YDlvTOb1+VtidYyNdBt/zhmauiJLAcBroO7Yu81Dv15+606tIzfJ
i8b7WLRi7IRoGoNJxqDnVKw8QuduWYzF/pQ3RByosWCKkoZuMJykyDzisTcyV3uki0nYXAFFcUCy
KdWVZGl780vnPCCC/MPbt+pizGO8Ff5Eofj9Z3A0EqFmcru1xq+YAR4kMZT8iScRBCvSbANlDFCw
MRUb3BbyBRf1MYeaz78rfcGZ5JkYLleKzc8dWsHP8/p70/wrlnLblmZ8FzPRRKOMVnV9W//93QE0
aXzyQFFicf01QtbkVkZhoK0XlGiH/G18BYkpLoujUfAl4NyJp5OA/oWlY99+XHVc/2OdEkr26FIl
6nPaTQ+YXaQgKPhPYqAtLeJzr5Tv9ZVVrrx/yxMru6jQBxpuovGiFckRShGbowo+BlsAa1PkQp1A
gUTxbqd3csz6EyCGUdI9V78ddUcHT6fS4P7pN5p5rO/jfs5LjDHJWfzVHH21YKKXNiAMbqMQ457t
1BlwlBrW+t1cUWcxxpUnK2Cru1OVp9DvyckLR13hoxxeIvtytZ33EpLRfGMQ3lDCnyQnjgthLsGI
pON7wzmSlHE7vXS2+QY3E/AaQTTfGD/eakYmf991XU4kHfX41zFUGS25A4GreIl89SG9vbiBPINj
lI0aiI8mZqM/g8xRfy2wnzj2RV+2ZB/GPmlVHyRThQaVvcaOKIgfmjGxBAH8Z1c445L+s5sFDnc6
W2zUNnUADUQMWTpj5Ssq/xVy8WkFVGVPT0BsixTTvrti1LWeAc7Sngit1ERunuDfjsy86dyfY/xf
oEdyK4HBWXQQhSUGGe3G5Q0Fuv0Idf/i+8FO9eI6bj3zd0lRgRoum4hLUCLZL1amIf0Rk44We2TU
HiUoIiBYSekOggR0lVhtUKdC9YVPhjYFmD5HO3170TC7e73ereyNwzYVoMOsaIrHgHyOz92rELVX
s6NjmE60jqfAwMgNAcKy2o8Q+xjyEr//Kajl/ZVhi3gJ6KhaOK4FyQXpMWDK6l44YaOFbPLUqIXX
fT/u3xcRRLd1VNBqG7euD0Bo1d3BGWSO/OAawnhvD7FRrlXf8jBA8Xe5o2D6vAQf8vVxJ/nrued4
7EE3zxSJ6EqnS6nsCn0X1eC4fpE3JfM7K2rZwEeRcfZs5OE8p7XRzv7pUlhwArrZyxWVEZ7nAqWp
qGps5TBT9BKUMAwYaJhcZ50u0C4XO6XN505G8jmRjrChCVAmA0gx8YpEEK0yacaT5rO+zC5f8GcI
knL6KEAB9KXEXvUswc2JHFV5UUmh2IwpFe/o/zUbxkFCAMFg/vqFnoXRI1kzvLBUuhp1/NihLxLN
WsavLpc02ExX/r3Ac2SwZT6a4DYGAbad1dhAUgIlMW8pMkoC24wkVvXojV5/iRaEZ3vPtLjB8Us2
R7FmPZXL+FIfNlCMQtU5H3oDw4KzlnL5U1QrzpzdfarCs3Sx1JqZMYdrzHuuofmiRk4Wmn7fhlop
6QtXHyePNXW7FzR8yzNVdgef7zIId9wJqyEcsOiPPA9uliwu6oOzuSrG4xcGSYEoNPwuaObCNac6
zUaSO1Z2HTSyZWDsOO2ZOShcUhwziQ+ADXC4dzxMEMMNO6xgxTIFztHMLSWBw/4xY+e0YnJDnTrY
uxBmWtT3Ceg+CyoZMfrlvNQWjoII6+Imb/+l25jhNInmQbVNbbIy2sFpb2H9CvHlgFpV2wYiZ5mQ
DC9DLRTmdBIKdjO4kQIZg85yxcT+s/opcJpp6KMWC9YJdjkZVQge/V5lPYh8+v4Nxylj1NCgYGgM
YpPzoOC+63kFwZg3RvikBc+k9rDoXGh9XXwcoZLg/rwBxQEfqfeM/PRx7trECZKhokpEfIE4321q
mRkforOaATv4aJmQbfqNaSgq5Oekw/ZswW6Yd0av6Olcg4eQBEqGef8unbsAibVVBKsTdHrwSo2k
vZTgXQcff3y2fOW9old00C8TKpbCGgnQu0D9Fyu+OOCTofS1UuSRKETpsG8F8XAbgIQFzFkMkbOt
HEFIFhMDZCrcUeov8Ke8hUQZnbSZ2ADA+r+9NwJE6qhznBCgtkjzDs+QsSjg4meE6fqm+BF1+t8Y
n/xsTU3ZIZhLuTlniPe3tJE9YynNsEickG2Rqs5bz9Ys3D3h5IG64kEwuXkVoQBGN6cmZ1V6WGGD
qWzdJvpiJxtX3omu+0aAA2DiLmBAlnxEiPhV1An1/a+Tl6pvUArQnuL7Kjx0u/lEWFk/H5SfYxy4
hEsGjMvsSKwPbsPrpCfAHKsuVqNuiuK3Ei5zJqTnPUlj6oU5HRf+f11DsvCrZCm7Po92WTaQEZI4
UNfawZq1Bh2iIt+oqL7zntpUIlGwdGC7TsjqmyrPTLDWdh0RAL2dCV6yjbz1CThabKuX8I0rW1wc
bOMDvju2yXAP56FneLV2hi9lbx6137Af7p8PhtZC3CdOCU8+pKemMlo3/5yVw4FSkMsD+39hfVC2
ZtsM0loWuv2hsKMSMBf/qFnme8s9X+ghHD+ESmcwkwyuh7LjqgBVW08OKICKXQ6fjHW4+y6oG57I
uP3mo/2nR+1UnH9Prgqvyvz8Pyglc3RpHYyg5k/O2Uq5DBnDwAqcJv6DV7O7sAACAo9+XT+WG+Xh
htRMp6PrZzf5iVqbQdDj0HQEjZPZ+IR78RgetX5UqbCta734gJDYGr/Fzq5fxWziP8Trky3qNBy6
U2SPjX/vwL4cXGQaqUslO5AlroAtos7LwjvQzu9JCGJ2yCSELh//GuXRg18ePYTJKRzdiQQHrNlu
Q5D/RbZ/qCW3U5RmTBG1/Qgop1KF/AUbQf4uYKk/pKT8ORHWJ02tLx4GzfnPD9zfEC27YIn/zY76
onfo175J55l8IGcNelreeGBOoz7ICrobcgq/HK/wRuqA4rwqrUiYoBGaSC39Czv4stZbPJEt6X9n
YoiVkDcxU2M0riIz7UAVfE3vHDaLlNqgCv7PZd8GxA1IqBlFca5MxdbrJ/Rj/X1lgdoWG+cJZp2S
elQYcMrJc5AJ9J3kfkvD67weZmsOkRzfayYyru5ITZEHjCXwIyouiaxq4euiLdgQzR8I4lGy7g60
ZO13whwPdVU+dTXALwt3R2YE1KQ7YZxjLFXNG2Q5dgNdVZQgmX6b2HNCZ4SirVEI4XeHhB4eYJpI
Z+nujeLTOQx+VYL6bXWUBO9Z9tNzJO7mPnkQvFNT6taTb9fHEiBWmG5zdFsLJ8VrEXciLid4/07p
T08nKTQlQWEZPLgwtuhe9neAdFIDSy5VDCD7GMbQf2N/Fah/JJZgT5pimTnUHtSkRy7RioEsBJsX
KQRMEnKF6RILTj2O5c8rfDRxdGb9JFKASFlUxzP/zzoCKXUVOJIpzLkj0QUTBX2K2ELc8coUrG2T
jAWdUMzS5avFd1ND2H8HKV+IwYJeo4960JNqb0y0kHfMPKGSc2+i4A0g2b24gXfMwKhqGMpcpo+p
pLeViZXyouShyp2DGtCDqPECQl3BfLQy/H/GhCIZCmdCTh6G/i4vMmsHjYIp08ewbOyA0gGrmQmh
rAW0Dfeym5CfDcGJL8KTRf/RjmF2K2qNPzFAzP6WwrKS6TMotkmmH26korQfPlmRHwpXf7na4bx4
0uc8s4kIZVpWWQlCm/9oF5ub762j/LVU2kuxTR8RXh8q5Kr586xfmk+Lf6vXnh3TsXqOcKm3YWht
aHbr0FgUxE8m+NiKNk0Vbs3SkNtV40SrKKRVQAIZAKgAV+EshwAx2Bi1u9wLqxzMBInSNXq7LwIj
wCtL4x9XeNaj5IhOMyKIs79Vs6PT4BsHj4m8I/9l1cwpLM2kdHqOHVmOW0EKOf7EW+q/CSrC/2C6
XN4U0ErFL6E6iJj8Lky9BT3Jzjh/QcZbAUEjTcmYX53bNrFgUjD1ZR9q7TkneVGNn+mXpSHPHYeA
ush5cR1sYdHhUEuAyt7EIZkGT0ubU7h1/HmEgIDKUSaoE+uVRDeRztZ56VspCD3/XG38dcd9+afD
VmGU3L3KlSJysAWxPnLY0yvKb1TSqCY7eqzxMnnBwRdAumo2SOGZUSLWyYIyWuO5bwTa3LuuFkoa
WEW6jswcibTHaQGFPriT6lMC0ia2JcSLFaUlrudQZBp1T6eNlpbDc9HFKQnw4vgvcUZPsLZs75J+
grAb2YU4VCz5yN7jnwcMaa9Zv5AA2n/121yC5OmY6CYIsCb5fRCuJ1Tb3cQXxffq9X7REt/nEAFg
ATns1bTyCMC8jo0+rqTkXcfSOJOAULz5HfbOUIppXdWAVlxgLTh7vaNjPWf6ljlorvLtPGO2PB43
exWLIqM+Hr3An3QJuHdRNIpyQ/N6ihV1ITqAT/kFXZSl1q+O/r3Xa9P3zFRSTMf+osX4lJUsoIWg
g6mOXilVl+e5m7BOhJ+r4AND4PppEeQ/XJv4Nkzw7m/7Q1ZyloV9LFMo2y8x5mQ208gjmBIVPFe1
2xC6ZDwTBx9Q/ukUK7YHnscls/6uHoLSjgY50wQCAA9dWQspEva10ujr+mzpquGa1i4MPy0lulpH
HFlyLiq2WUCXIf5p5pwTuMEr+HOqq5V0HpIU80/PzukmEN9nvUBnJZsW8Hhuthzn5rEVcshtJDQ3
GOb/ph/Sp3PRJLzjjUknvGxe5SrON3o9+KBQ6BTsEhUwPqdtTjPt/i7MZ96Z6QGeg5vz8uEKs18X
eiPSV+3RsHoiP/hwgK0ek6koBxGcOUDyTY5uxx9SmIiJvj0hff7zcS+W5xGm3yk6luLVO+RbM5Ax
fJXIlYboH2ERoVW6sSnHXSvthb2O2/zZCCmzQOuSZm4ilvhr1Xr9nK1633x2u9I+77aAE5z1hcCN
AuFBE4h6shwLs6RHjAovuCRzmGCH05xfoYZM5eraKr10gUekuO3f1Nklf8T1+zmd9OclYgd+0aA8
hNfIKStnm19sJD0e4auojouWWZJm94WXiVQY2n9U6Fh7UA0kWLLx8ZlNeJu8ecknpE7GZIC2IkiJ
bnBe+6PBfb6zAbn6q8rsIh3W/46RThpaahn4UHTGDEWOHZdyI2P/aotoSP6+kDUEFwLHgEtBEWhY
lSmWZNonYo8Y+Zjv/EYvlxDOZNDbWvCY1WdP5kTEeUv0lyh6F8MYeredjdLKlihjHzD/oeTIqytk
VoxtIplWuTQvJhC781a6XM7bqd67PzuJl//soRTPMaPeXMYbnkF6wRkGR62NOpKnCpyXc2is8Gt7
VCbughS54/BJ/RdU54VsfnWpYsxGtDGOWPK/Rpw3eNHtRPJ47vso1Fq833DnoFqyssYdm/hoorJy
MxGPzYSxdXKSuS3IUTLO0iz6BtyTBy4eJ11ONoNS/P+BNkHe8hszDGtfqrB2FPjvfOYtLUQFDilv
GAIFvt/Da+7Bo2gCFgiclLQ8N0Mb2s6iqcyaF5Tqhy1a9sQhUm3xV7syvrRCKwBwZf76kIYnCXjd
mQgxgxsWnU9d468pnBSJ88qQzWCfesImt22eHysU8AwaB8DaV9Yg2YA2JMVa25+fCkKj/hIkwNO8
FY3iADpL1yGJ/AuWc56oms66CRrPTX4uRcpI5OFY8xoJ7k3Zkw8KH2UkkEJkzTk6JmgkiNAdEI5B
4MOqRUNXfpWb5EK0EhO8W433D/k5BwlvMQZWHqtkiufnCyRbkncY/6krXlZuB4FpBdP32IHVB4r/
97YCz/jNsg4gWBV2aqKlWMEOAIIu5DQaxqbS8Ftb7/d4CcuJTp7EE6gxDKy1DgJFY80yNGQor7oN
rUU2TlRyDiHe0/2da8a1kZJCkXfXlaWTszmO1kOiP0yVkEuAvDUiSymJcrFvvihVLweUxMzIXKsC
609jbNNAF3nybWDJmtiTD0QXlyU/1wJZIYlvHTtNRmOFTiPVaGan2ggZHaXGt9xjJWVySIK1HIeb
T5KDN9nvfGShPfQdk1eldOMpw0C9d1jxEVZ5Aj5B1922l5lf1BR/yXAunBPkWtRQ71xWy1S6sThD
XETkivp5iqC9mtpZ3mut94HrJXHSb2mwdWjlZdPTK3PBAMeCyJTccOk5P1kC4SJ9/c2T7hlaYJu+
WYSVUYRjb1Jxn52+MwbJizqZPV6lvyZJHAO8Q2pYAnCySQ9p2wQf2wvGVq67tuBb/6EfyQhuojxe
ktfgAU2n+llUWj/AF0ze34t7O3cEoux/TgMH/Mac4OmlotlCwQPxIdKAZNh/9Vg+gBNCU9AHVbgo
Ich76NqYQTqzfPKTBEZ1DTlnzTfLEEr5JeN/sqq4H63vDY0xMrLDHKRgFdIu09SawWfw/+BkfmKM
k3xVRGAlhY87Fe9PlOKKKzcsBXijYlSAIhH162d35LKgKY6oYHPo/UL/bWgsxVOYFH40OH7YALRY
dZ/uHPzpRkT8MfPUTj3tXFw22OqjCqWwle5sCnTRwFyOY6lb00bQbxW76w/XSFIOOV3a7KTcYmx+
yMdY1vsJAMawHdOPa/u/WJGwMReFgeRyOm6iwflikZQsURPZ00IXrs7olhbdRg0NsbdGyJHnX0oJ
+q/dQT5ShsWYNI5uGDYREdtSOeR5irlqblpW4MGybaZpdXLZP2ZHd5ujlNs0WdPP7Bn1fDzqzLwL
u5UlTQI6M7COPj3VThSzWmr6BDXw7j34BIEcfq8E18H70iphruSe3oLIYojpq6iNvOc7Ogjd80eR
rs23BPLN+FWnbf4WVId41DphKXkf14GTovbFPaeg/odpNbOxSvYGMTkvgY0DbyVtsRbqD0gE1p0d
GyNYYs9clnaCO+dueknuFDSKUHPQvdFDZWzIKAjTcBGXBvzXlKc7OKlRGAhHuduvKebeCOM00ork
AUQ2Jn7dktpeytxuE1saqGPRagPFhfUp8iVBLAcEkrS7wWJKv+vseXkdK8qH72Vi5lr6wLwYER+g
MVjoMqbpnx9pJXHQ635Nu1CuvStV87PA/gxiAkOG+nPnJQEaw9kIWtV+MBFcKjQs0hFV96Okx4GI
O1U7PMqu6rN4oAf4ie07t1XWaAZGnJ3sWwuHPNBNKRtz+xilpCubzC0Bw3WRXDoTMHEmsoUF/FhP
TxU90ym3CQJYq7QuvDxt4JU7LcKFeLyEZvmnZlKGVhjNkNX86JrkECE3QsVNLqTVP8qafUP80CvW
K5iaJxLLMFEkNxhUa0xBCi4Q74wp8x7EHnzk2897Iiwz5/TrJZBpuprqyp1rUaFNpRbNM8l71LLl
iSZoLMwcTeuiOfeQET2kBvGT4/Gwqw/cfM8okFMsUApKTImL65hZmxh8QfQ2TsYakU+38NA4xyZC
Cxnf+otLlfNzCPmqyvhVsy34lKxzJsE+kcEnUOKrrtmgN0bHrDiTPy6uQb0ztWd25nguE1TaOj21
mbFDECqaYhNkC4YftFwAATLn0jKDmO98fvXE03hnwbR+2olVYC7BH3J9F6tvOBAzsfrhz+XRLqgV
MVCmSzOLRXq6LtwxmPc9U39LjqJZtllsdU8tlzU44Z4E+YplCtdRoUgdM/TjL8K4AsTOHB2wdGYM
xuRYs72JpRY2iXU111rbBVC+Etgkig9ji70lKDZGsvvVtdfbp1sQpc96v0FXUcWWvU485jzwsbqX
mmY10iERHtZsTZghgusnH8oigNkqHpT35zHhPrAfR8kcs9S7I5ddP4VuRQFRfioft5aeb6vTCCK7
Eb9hmccb/uwunlpM36JvxcvP13onbg5ybLKyCct8YPoP+fmFsYB6gxgNyJGBlBxWgWmprIGMtt8B
F+VJloAwxXEilLIlHfga+Rw4USMSPGIHfE7qsJ/CwPaVI21H3IaZErFm5SoQfbR5OAQweVY/6sIP
jBCSuhw58EGneqLqdJSTl0Gdr5hCMXTHMDkEa69gJNJ4xKXI3g9STulrUCoY0qTyAr4YS5pEmAMy
gNrlP2csbJNIId6FPe+NxnJgeoL2+bfeT0ygr+DsMVntorjkb4LOsmy7vxR4GtQq0Rg39yEnH/Wg
v+aRfsVn7fWrOT6iQ2lYxStWQvMFgNEh1NZZEaQGqVUc0Fi2+rs7r2Mooul9kNghtMQ7ZHynymsF
zLT5liNRW6ivmpLUAZ5cS2NHN6wD6ckrsMpSSqCY4r+l7BbQ1UmDnFbKILCoq7ImoZDu3Z122+CB
r6fi0Vdz1IbHnD8tAv62Gjubt7GwSd41oE+qsHNp9uRPFkcXAC/UVT5lu/fW5U4+sWWIDsm4CMLM
kpv5UpHhLAVKndhtqrxlIObme2NFYY/d4Ewqe+5SsIFydJ+gDojKek7KaE4jbZyMuXjs6KEoKKu8
mzYNg9xcJO9gt/u+3+1AdFJ3oJfJ7yZwoGNfOOaImy6EZkae/+qdadDfS8JeLDTI9ULG70KmfCq+
5ddOfq9MVywRa1+2SJp8dxiUVbEf+gtWsC1k0253fIOyRWy+P8PKZzIE/y1G3+2Fb9bcHiOAwruC
na+ossm/+gEYRymSZyeYdWHyOmb9mWL++lU6pT3ME3sdh7VHyTKBWCpAmbR6+plcFS3tOaNgxQ/W
zVMPBUi/v8MMyTjgf75GtC5mY0Bd4PYnveYXVnhOvm1mE2DLZwIhj3s8qsN6eQxakIK9dCq0pR/w
wNq31GeCyOtETZvWRUGhfRQxSchQYJVW80K1dwXuv1J8Dlykg/2ns0O5Q6wWlOFzftLXXoDU27+0
fmaPrQWS07/YYwbal1ysvmAQUSo3nbdzSIeeqT/UVwaarfKcCcYh4yg6pKgYugGbOcTzWCraKN6B
HnJ23LEEuNa4EElVjU4LgCPeAI3mILDypTaqdiFSN817GgR08/EOjtHPL4s8XgVcNmVnzKlWNpax
bttbV3vbGZyrtiiLfFQ2Rmks+jDcNONI/wZxdPP5Z9MbQx0pgz926YzeL29CnoOFksL1pSGlfP2/
ygr1g/tDwgzYhI0t+JgO7B7ZiE5ab1EapxLnwlYGY/ujwZB7qrmzBnwcR6cMRSWnXeDMswukxAUk
3Zbu+3fPZiDROBPRzJtD+tlKRAqx4o+e5r0DhjELgM9oGr75KbxdAu81JLbzZ78tXp6oPgpxD3c+
m+zgVOmk7s7IAkVnoAdtw6h8ERFsXvvP7CfztnHfXmp35SCu9sTT1sLNYeLxJTyd5chp1KzqtO7I
ryV+bRgZY9rIjKG+HgIrHhUuYHRpj4aGIttLdIrQYP0DMELqsWpUz1FQRp4fSjVjSGKkYwSzXB2g
pIjdpkdJl/QiuuY1C4p/925gi98tH28Sh6RqVdFoF3NXn+dMGp23U4vG4i5B2cFBz+OFO1gOIFds
GygybljcxZvfO5oDx3wYNfJFXBLqQ8YdnUl/6JnF6DBs7aFiv5HOCDqKQStl0APjg8KmzGaFn7dv
S31NpUwX6fdFDfOzID26yFXfrvZAZxO0WqrRCEkBA4G0EtvXIBvsMFsOf8OZ98JIZilq5ck0UdBJ
QPDAY42VUoRNkDWeLRClOr9Hq/OtFmqvAS48MdL9PRSOygP/yK/DqfYNK5TKYxRTsRaOtJ2DrHPS
thjoK+6wMeCbNGT/ozOg7+/HGD8zRp5/Axv+YkEdK3odSDUe6XDz3z9UO6pVIkxwFE+lcXXvSirv
YVMDBDFH+tla+c7OuiLu/6MCVeei69kq1rFQP/PTxkRvwgG110w1OLct3OcNse2NNo5v+WnD8Hnp
u5NTCxDXJwO6IQ5N9I9Ue/306SzXbQce5Qb/8k+RLhK4mJ6rlMgT4QbMFiBbCIRiJ+FOPS95g9vM
IBbidPIjmqw8HLxHfV1r5gqQ0ZoserAFvoJn030l/SeVlybVojJKKyP+wkzey62ZkIBAjDyGwDvt
nFtslp0r+KC6ND6yUh3/hOo8TOpSmZQiMK2J0RfjGRBHyNz5WbdXPG02ZZ7nlwvyTgTVtp7cwGNk
XU3wrwplZKCRpaWNtzJXv2e2P4/4PXv+Sjrf4IZIW1zXUQS2OHLeG4pWzOw2eiVB9ontf1UKivvI
khPyJVsq23qwJGFeGHkcEfiJSal8XBM15jVJjkfsPxBYe7qT/Khh1Eh54/7LsDvz96uLYjjt+UJV
llFz996YEhkpyI0fjSr99yJW2OObAuZPTweIrh39yBhmMVAvg8eRxkQRtqKJ8RdBfX14y0Tu6G6y
VThbUQk5gxs3/AuT9RaVET6B7jv5KzY/o88X7OI3P4yZUvDgUbnnIfejmWMEwvAh5LyXa0lb/b85
nYcK68cBYmV16+iPnovtqJr5MyVYLBFpvPyRngc3g4/zdmpow9E5wMOQ1k/TZ8uPebwpfxmfJxl1
oemXmj6XPZ1PFQCpjpM4EI9/gjzd+qr289tAiXtWg3uIs5iCFoRND5HEpupGUdclguKIYut0XX5m
ekWLpSseit+zsERaXAgFINV1ukTLoIIdyDnbsH9iGRwIo7wBWqnJ160wvgUZXs2BjeskeGlSFBA7
jAsxo4E+0t3ZDW3bZOkI6Du223HoW5ieEnFso3gPp85+Rjo+jgI4YwIq7/7s4D3eycC1jgO6qG67
DWYrtE2XaTkX6Asb0g9QOuQX8kzNMJJLsUYAnvV7oEF6PO6BZVawz7Fx5q4o4HuX7F9ITEag8hk1
/ARFWZM+DwEzYpNDyeWL5p6NeiTSaEnJfacx7TXGxTn7kA9P3MPdM5j/cVpOHFQko9vDGKYys2k8
BgKD3Ve9uYxBR5RbhRQpahxPbC8YVErQ1ZHvB7zppki0m3xX/rcWviw87RzkDTwQYu6qos6VhT7M
dO3ZJ2DHRYMJqgE5Uo2KfX7eRjgGMlz/NRpb/g2/Ejn4GyuzDLxF3UrRRtwSO5E1XgaVhYLxU7fC
3WfQeQ7/gQaex2QhikIwqTonbEkYmi0AdCZg9IKBlLKK0FpNY3XP4gEuOJiAQP3uxs+BNAthFxI3
EY+icQHjKxWWsvm3d7oCGZkD2iYqfGOuf62R72Yjk2rYr5QBy6ES1APy3OZHAhqE3iQV/Osocdjj
A60MXNTdl7KWWfMOgRmHT5Ux0szbtHZXFeCC45y3rhi18lN3wcnwPfhvfy0uvKtPMY78PnhaA78n
hO6ocX6VuUXYLQEkZ5iG5Yq7dtfU4/LeyBcJ2nRwsv4ReBuumLHpXC2DDpyXsvwhV1oH401eYrZv
NcGMQM4WpBfGhVUtWONEBUWKBuu39HzN0p5ufsIVt4bgq8hOLweR9qtj68EaJ4x0Ppc4RFWZVAMF
BFPMVPIigGB5u60kHVHllXzxDqTZ31vR7zGgfLUZAixpW/ghfBzKhN0W+FpKACOe5gMcCh487JTS
yem/Nz2CAae1aYGPfV4Ar311DKHwzhFL1LbeV1gua23cKiQELyamqVgQUCUcoOrOQOvtfPRx9wLQ
uDkPa+gxjv6n+2ZhNKf2ttUuSJ/jnhbocoe/Vn3r2qa61L4zGWuj85mRTOQe9tve1JmnNebSUTr+
GfUHwJWWTV97kEvsuUxihFs4F2/iP6Cs71Hrg2MZiQZhMhQP6WJqulDRW2Xtdkhr8Zh6m5qZhgCl
1tbR3hrkSgr46ghh8Pv3qNaglXMX+Wghl46XXrM3Yapbqqlp/tLlhrutvJwyQeaYKw+aKCCBusgj
g0j8pEYi8GZZTiBny954lLSE0alYUJnNpsRTAVfbKx1v5M/23zaen4jHzEvKjPTvLbtQHJs5at9i
3Un1ssT5U7LfT6aAG5xqFZ6ccGFbc+BXtVNAK8vQjd4KsPBjORiBpWRQ6ke+/fCbq1FEcOTskTzl
C3zAgRQFQVe1rAj3e1aYKk8MogFZCRjH5kYlT/MpP1rBex9IVEytSRPfDCWKeHQ6KcQfHgm/sKhs
4NU0zyvX8pB5rsqDmEfiuYJGuvT+QdwSjg1go0oHxQ09XDYr4jdy1ULR+VR8iGU4cwMdNUrg1DQK
kj8FfYS629qi2shfHiTDEGleKKQT1m6PwkobMLO9oboSgmN61WO+nNCAaBZenq6z0NWHVAFksrt5
k43IPrZ0Ue17esp1D4J/LXv9mULTlZxn8dvK+QFGER0w2UkWH7JYj/8Nlo3WvFAiaydncYEa2rj9
ZaaMHLD8duCnaDAIw46rHVtxEi2ofcAtjQTt33PDl5NSRhvhJetxx6qBX3Qr4FY1T/tCqOkMLke2
dFQD6mLcMnDuHceOFzlLIfVErhUaayNCJ3DCH19XqI2TY3XPe6dCyuZC8d4GeTmwCe46rs86sEeH
RXEbvkGw9AFXgA2z9SDIDHZT8hBHqXVv0IjmjaApRToV4uWIInjGZj7K43dazYMGG48DxWM9Zo85
vFJm1plxaQMkCl3WiBuQY0xVBDbeKOQokczAToWWdnEPuW09ePAFRIjQkUqckqwUY0rfNRYaBq7y
O08HzMsHf7TN6FEcNiOW6O6+bUx6yhJXvQ+c6HmQEBJ7KjnBcfSGTytCt/GqALn/A+cvQWTR/JGJ
whcI2Cz1XpwDz5o5UxTLgVSTkpqhZvPMGLiI21vV6x5tBzvJITSNhNJvAsn0OiituMy+6sWZwkYB
fyWhtv4SqsixhA5uNV4AovwshLr1D8oEBLzwjWPWobyvUWXvfBoMtQOa5SaXWQFSPkMLzamKsipy
xUxYBsYnTj3EKmGhuieevXFp39Co90KlAwthI3CJ3oLQandRyXWGO+yEuyR3eRPRWNELC2K9uoWO
jM/eQkSz1D/t66Omg3EJ5r+raje195+76fNpmuwkEZxvRrnrRxwRnlC9vsXUv7DQp+HEQwt4EAUu
2iGhRVeiEGzlmS3gMrj91Y3e80cXEcXFN31P8pldhbBQPnDSZY2FJ4O4bpBVcqZhP+kk6iZ3w6L3
da/IsGuFSfgPpL4zknL+lyQG1hcS6CtwGLCFwqsjkGm9htkWjZFb04zQDjiClxetAtAVsyQxnUdN
gHANStA9jNTtp8GK8ziCQdF4nh+y1IVGkkpZiLFGY/MU5hF+J4NgZkzvTawadyMOzk6ZPREvLciL
Tw3OTV/Lkpfu0YFaKgxlDs/OSFuTRVlHTvp2sVQsgIOSfCqjisTZ9XPfDKyRZ+2R77G3zfGHFxQS
DKlza0VArqi9LJilnguY0GGx9Z63rYMOWAsSXgjlgIadQ2W3xH3RYDlB3czoCKRKJaK7DJIzwRsS
yphsIWtVCW9OGK+H0tnQSy8z8seBak+fETcsncbUbuoGxEz322EX5gkfFL8JfHqkifDSKZRoEuSm
oFq+vPxLMf67vLnFG+sdDFiuNcdeweTzuNyVOmZ04oPapc9er96ujeC/FYyYlvv5ijFBVsRoGPhM
zgPDCSFGyMaaGo9/5wkxlpewAB96NyXJ8Lvpf0sESZYvjnl15jVA1yFbp/ZWaFDtd85rDnIySO95
BbFe31jDFwFZhRNmyfxqnROC2KOtGvGJK6f0kwYKMAQULTc4GOuX5rYlV38hkUciEyJnoeuUQRYP
Ay0zS54WPRE6+JCmSSqWaoC7vAblzpMrnZdatDdELrPQry1uk3akwNwpUtvGb4XO11wrJ4rJ2QPV
1BTrhUWDkkYHTsS/qmcn/Aov8HRYR4vdUatIuD5yfJ4K9RTDfUvk3YCP7gv9WurIPtzHrmPG4tS3
CnIxG+FW5qQK9D/NhWwxVPkeUHj5vqFi1B6YmjtuJANivyiOw3HJ4CJLFSzL0hUyGmG5HQ6SqJHS
LtYdrHbAb57VXJf98DdYZF88ZgD8Kgc91eyUbRz4qKbamC8NYuaRKHPHszYUzXd2aOJS/dIubM4I
aQAurfpV1y5Gtb+035AX2nQjLPJg0ZtgZGbfn0wFuHMC84YMvHfSZl8u8Tt3g2pxFhwjyi0Br1ZH
KqrzO4l/CD+sbu3AxwgaIPL+sr/2lDD3n8WxKmfTEkSbQAt/spb0OljPvgw33Z8N8Y9DdJ2gizkX
zni3tAym0cyqoSr1IwcCs1q3MS+sJtWz6JOeEKFcWGQgjBTFX6d8s1n1+8qgPj7gL+5wpYVEeGVG
rynRdzoO4SSwDdYHM/UBA5pFlhlTaQgouQW6G/ots7QLd5QHoUMJ46DBuJGDVuR1iZr6L7/P4tLa
59hnOsYvk0seo2fXe9xJdgec0lTEMc1ACaUUx7EiVNiEXzwR0SoM/TGG+ABS/c1ZxdamcCCSYfph
cwzZLw67tZ/XI07lf4nqiKl4xhHC7S8ArXN5tatYYgiRie3bF7yv/N4EloyBlTP8T4LW6ftPC4Kh
7gHzP37OWDZoIadElhpv/VQjxxJLZjzmxa8sJ4Ym+HlMAEVbwWvmRtJiVKeLaJoUmmiHzKR7XSr2
iizKEbBAh4RXKwIbHL9wtstagKK6BNUs9SGcgZ65Q3X5ahTDEQmaRnPMW+ALn3EGr3gLCZ0Wopl8
cLS7ho+++6vc5FW+A4ddgJxxQPyHThjYJHFQkKzGNv0elJXm4X/CWhdC3c347/HaUw6IYM832Mj8
Y9YS+RWv04fhspcuovPOWK7vAIIHYvGPCK5aEx7xT5ukFf1bRYrfNXtXOrFjglz1ERUj4WIbzXMC
0mXeZrpox+Undg4jWXmq1EFU3TdS4c857lQaai2LIlBDiy7hob8B4KpzV8RoH2yKTP3uqrIY9e7q
C4kQ0WgbzhTfiz8mS8yVPakseIjhq9CTllQz5xMhnOOalPIvraYzNwEH8XitcTtdMHUKIpGlSH/O
GHMAv5BXewnVtprI9QDjQCRLzEkfgNKR4VwY6+jKmJ67NnQNP97Tb9vt39I9xKr/iGaxySpGmdBx
JbNQssAST63vQUbmNUlZCvnzBnYxgmto24EPn51fsp0WHVjZwvZXq0Sn3ZAlp3H/Mut7w1c6IH73
SybomhWY/VT3d7uey/2tqZUutnK90JISJwBB+95m4Vg1kozLmzU25FLju0c/2zlOcVn9u15crea5
eDZbXkpQMUHmADtL+bDxYv/W7OGkJLnjfxksXRgVQQ992aqWV8vNSW51w+2vTxsAU1ehElwfs1ax
WGdDt/pcX5cvooJJ4LpV9mFvqW3BAtFwu1REAJZS1RB57ZNz+hvm78AG3BMpJ5mJTwkAfurMQEEo
NzXFcu0qzYx9nYkpZENviZ+hdX+8invH+Yo+x9AypsCjAhfn9C/AICLpJnRJOEFD3LTZe7jg14AD
rcJFxSmEtFmqBtCXDBU+iDd53ihp306CAaqr+qC114yoPza/DT5bIYknXVqanB+geR82Fhs/K0ek
REyIj98rqriwdpf05FFpCAsHqP1Qd3tMnxwdEwGm5pSVAuOUHPPzkcErE6s/uqaDACkBND/tTs5D
N7Dh1Hk91targHW7USKHZ1XhUx3PyIRxbgzpL10W/hihJIFnaKxDGrnSlcJroyoXxumaeVn8oAze
shiuHrR9SmhwK+ngJNsODleyNkFPyVCNKNK68/iLMNg7Q28wkbCY2o2yJeTAFP6MLzsPxZb8Mbbn
w9pk1jrMcYpN2COAIxqHclPu33QNZ5ZyD4W2RNiXvvsrXqX7AIdWuLL7awIMDqBoG5VrYAE+vDvw
SGKX4ak535ZsrwHTk29aPHrbkVHE5VK6IUNDdmLOVdaPzFQZpslU2B1gMyDaQmged+fhKvgEJoCO
FoQvkpWaA+Spn4XdqPcdpthNSnOwQHwfBqMR6Sm+S2xjkQP2QhQXFSDmpWvdvIXFSRWEwY794Ekj
OWz6oac1zQeK8/oE8hAkZmgivuC0DyaXB94jZmRJEW+Q+CO0ym81YFO/q76V1OxCAJ40mCFH+Lta
HIdrct5DbAu3QU2G7J9LUc+uv+RBIawJ1T4fs1ZGuKD1LXMNe/8JNWKTsli4ZVoOGXBYrw9xtNyz
nuwlxLOPr0F8sfvZioiu+0bQ0eqEb6XKyXwAQSubtDl6DLgVtoORctLSfVf65kKWRlxguY3Nwta1
q9e2iFZ8pYV5O0/CJzleicLHi5YA5+sxmUcKfpLXFxy/sshsVlNBDAsxxiP4vlkBAq+fXdrMrb5D
hAxvnBe4PFqwEQyxdD0nycRnyZOyqaqL2lRs07eSfppdFZOKqpmjufZpeDZieAF2ER6c5CDKhJEN
bZT+b6JbYlIvjjr3gBi0vqZTRCKUXu3Q3ncWCvb03oYUU9LaMEFPmX91iZTCOcC5T19/d0gsjQmV
zbp2mFMIPMiUNgeWqKHADfGrkmB7DpQZ+QMdWWT80mGqdSM+0GQDH0RBZT97v95M60naUgFl7ime
AzFG6frVlc78CU5BUqPAhmeq8DS42Z1apneRsH9CW7hv0HOwJoPw3zGWUrt0MvrrCptJOP5+i5LL
PlaG3c9f2BNDxpGQ9kCFff1Knx5kCM1Z2r1TGw/1+CutYDU0u6HvBelOzYPdomMqh9ERgSJ2gkce
6FZvObuPnY91uCo1Pjb5vw0FTGsFvlD75T5e5JmYTguZI1jHIxIQzwMxSiueNBwTDcVuzSQMUEzW
T9FIDNtEX8OisuLrrtha8kCOGoxaJuOp9IHy9iTNd05fF0NhifsoLpuJBnOAqagsRWaKeHXTBOvr
rbOr73knkB3/zCky+Yld0CtpgvDn7HEoWkR4h0IZOMTihBI+uekUFoeoUhXsGFTPmcvvK4V6x2lA
qohBRkHXktSq7nqC7/vCFh8hSybBbYAVHpDd+OMY36W1VmCTn/coVWhUtmwkW9YFTZUJp1U521ox
Y0KKzrYhmp3WfM6slmjE81JoMqXWY8hwX/jDtrfsFUEjdZU/y+CwwQh4uETVOWT5QcKtAjywQ9c4
vioE0fVNvgWIRWOmF8bd7l4nq/xv+FwCEnPYu7xevqpAT50cpX/lyx9/2a3K0QwXmVSGpxDx8b4E
ZcXPnJdoqq1RJLUwQ4VRGuJ5wz5tdrDkn+aD8nyfJQmQBeyf1JOpjmpXIQOdRKxJZKn1YGHZ/WIn
SB4a7zOKsWbRzHbGfo+wJjudoJVAFGCSWodJcpvqjo6u72B5yREtI2IT3i+yJxVlY9xN3n3nxoXV
9GbzwlkfqCFluAnBfLfXbmeX13gmV5XOWNsbxMjehn+0w1H7t02V69ULuGaLwNN3SQiIJJ25VfSC
fjex/mGL0LZkUNFaQQ/VtyPqpo6pfyk69/UQy0POnBEM1P9Am+bcCb0rJckk/MB6hG4rDhqseYOf
Jkj35xQhFJcs93fa6JeOs1602PSWcd73pr612kjuNqkZMIcyuyXpoMtRE6d9ywyivzUgnUQ/SVPO
XKy9FCMAth+i+yy9YE8+QJHIlPiiL6amqUTy8KeJSzwKM2FFKR3LU9wWfB3NtS/3vUk1Bpr7h6Y4
mN0MSwrub+IezCp65HDLSdDrYQ4OA9v9l1uN2rEVzpaXKkfMf7SxCcad4VK0jMlUoVroJHsqoVvF
dJsr0+LPNXOGRFZyWVb8T3KNaezJjrky6zKDdH8U0NHCFZudoHGwxL86GkfYAM1SSvufImMiwlsS
eAxEpUFCnzPMHvrq0ZhvmHb42VnwbfM/rHl5wltLLTzMPts69Y+gasg7KXjN8nMHa+QX30oic+Vk
n0na1uCXmeUtLJslZRwtu+N4KVLh9djFXG22YhZ61KciPUJ857WO14nE8iIDdp/Pw+HnAePpVJSj
JdXWFeuyAeqRtQq5KQ0wynnykuLsJSquKaZuniKE9SNKhV6uVLirXMYyODgwtSH3en1b4Z0nQuHD
24LTL0vANTdVEhrvfUVUvh4Rj1sJVyG/NXJIu0oWbZ0wLzlPr5u3PQlcrUjhjttjr4LjtgQGavH2
yfql/kyVpv16KMJmoYj4o7ZBuv0Jx38U13Y22Dn//tBd+C+u7oQM7JcNjrdtdq+6Il9aMzZKjbCv
HFryI+VKebU/p4pZWhqgo+l2fBtZsNzqoCjkUbBpoua1BB0XhSj/FJv6pdj1EwUOeQuvvPXokobV
xI2Zny4c+0MtGEbvBRpn0mxc2yahLxkKN+4eRuvK/ABZZNPMmQlKvPj1LuRKUFI3+h/Iq7NHEAQp
C0IEhpp0ZUrj3ewUgJJrYdN0RuqJp98Ppj0z1s8zuoBrz5KFVc/VngW5Cr7zf+i+CQXczmAgZz5f
CLXaH7U2m+paOTj7+ZRMCh0lTT+Xyehrnzij87EVSo384/MI2u7bCFB5qpdhsDZ+c40q72tHEgs7
GOSw8NbiQKj+fyhEF9pCLeyUS/dV+WWYPDNSnhElIQf9fpxEsuEhQjMdNCxY5/oMqRBYakK4V4xV
c7ZiUZ9jL4ibEISHAMyVb3mNuuUdihhQdVNkBd9T7QbS1Hp/aWkeHSh1bKwj3ZGVbliuhLaz9ls5
3c4Bj2A3QuLJ04Z8C5Opwsx0LJeEhgQ4Zwj20Tsv542BXxNFEj7G4lTsqg5K71QHZM2yMSgYntLM
DRbiIXIk7KNTLVvTQn8f0NgtN0csWiA5Ri1ImGWU/0/H26RpjRepcvOJImx/yt1W7iTHWtdB5jLc
W+/pmZyavYA9RQdO4VvET7JzfOZmqDa9b6wE9C53vRqFRlTa2iy0npWsrPQwyZ0BuZVofftMJEVS
RR3pYsukxyRs/7JMyBlyt4+7bMru+pGy+BbuSYFcAHzAV5t/yBIiuw0WuZUfGg4uOJmDkyh+oNHD
tOoxB5OFmctl090DWFiHfpKbLF/PPMFHPCh3M1b7FVzDxdkgz537qqrZX2uPBRigprAdQS/mhnsk
b/MVwPTqYZbuMrV0WFIC0FzYTX3qBzXr5kt/D2dAImHbCV4fze2bM2s1/VdXTWUMDMkq+uWO2OhM
uKfd6KSxmLQcWrzIKrUhPHoEa+whz57scaKAVL5O85msUufw5cWzDObqnsRYq0bTfUzH8z7KlDuD
hpwFtbCH9JCVwC+OB9sGBGj1MGDRvgXeseVkBYgkxxQt2QtdSx1Q85PAiKRzLg45WrbYENKJswsK
xeBj1HwEHmBx7bReDZDq0yI58yZNbc3r792EpjMN4PiITG9hdvxW0S+InDcMlirQNjTYhyI2lpN7
dRsGn68BrNIgiwNEtCtd3bNrAZYVK2hw6nQjDr7KvwnSwzy3WCs6Cj5BEJKcdMoO7FW0ztlWcroK
1pptmKnD1TV5Ld0rGIsP7e1L6A4W6M9YQmDVck8WrEbQoKLKVA+noXSqEMLSR25/LAdV1bMIx6fU
UaAR1IQt6HBOTU3BdP4l0LF/4ziKsjEFSHYVad6cA6H9WP3f8FHfrX4O+IueSJktLU2Xp39a8n0Y
vd6Dj7vO+KQUNnHRFcb4t2OL0+7co4mKWYIl/MibqeUBLJ/0oE7gbpZu1RrBDOO71cRVD2rmM6mW
8/1nYGR/DnBAVOzzYLY3NG2TxDbw0hFhQuUiYSfEIQETAQ0tGnBBwIGSFS4td5fHgTaOaNr4TbJe
L5htdDSES17OefytbltG3b7CIr6qjBfOkOc4gNh0vXry+Rx+t6gnFExe2q3CXfzVCeCOph5cT/Mi
nsZYl0eNij9BgLuVY555L3SgKITE3sMr2DWe9WptcKAyhKu83N1FQcj5jZuaLgaDPo4hNHnGWOkI
c+0B6W/MhANtsJowNgzYxl+oZwDc01iWxCPxWwswZ1j1QeZ2v1lxf7NRQJ1eEfBpWGGqNosjQTlG
PuASesw2im/BSe+/Tz7Xv32bm8Dh/mbNcz53sivQFjhkD8WMJpA5+DInZ2JXrRXpQaixbiUNsXdU
/dLkzfH4sU0POaBFqkoAE8xNLx9MqhuSaDkiE/WX89UNbKtxq8DFfwM4TKVnCrRIv67kDpmmPuz5
YWQEVf74mRgbcqQGUAf/Lem8cUVYa+F+ajDNL+HyzyeqctbdLkC8BSwUT9TreIr7hJz4B+a42pqb
3ua1EhZJqOJFdCzBaXzSM6rmfaXxlsYLu2sOweg8b1ExpPDt0AwUxRi89+mEbM+5VZcs8gh/5HMK
mRsOfn0YSh1bzWuCiH4wc7kaZ3MFjdZCHDtjasHzVAPf2PhyPxNXW2KEQ4WWozZmF7/uG1qGLYwS
RAhmsG5dOpHsPv5MegvibC17ocR4ty6yu2fHRCGAtmuS3hdtOkq9Z42nKgbrlEF4IyQGr8z1udLC
8QVjJKUqXV8RQqIpoBExI1NnOK+NrejvOyml4UUOa7N5l3ywri2awaPrCz+w+wMd553+Z2cGB8y9
T06vjYddzvi21oQ3lJGcDX5pDrHsqVDlqLArY/MDax7BmGYjTKBnNndtmz0H7V9+gJ8EUUelmRFB
2Ah+nT6bJUuqAaT2yF6NEtrLtOoCvfE1+5h9NynuIA+GfMCT+6+dSzDnlONiZQ1zEaldiE7pVEQv
L1G6sL9nFfy3pTTZ/qRNb9paDrnrXN2NLb0wswZPij33G0aslokQkIzQp80GSQ3t6QKzvzKGGqPO
zFhPxk/le8rwGIJPdtxFclUs9ody2sh5UYwGQDY55hAXNEHNYFwwvfR9xquHKHGfblOGyC2JEO6Q
2R0V81NBpSjZmrbA2bmhC/PLJEvTvga3bhSC/+eRNBvw7LY+4rQuebtsPc3+SCPkIheRMWpgP53X
sEe4aBg6gnTX8JrAxj+c2UFmJVpt0L/PUDrd7JjbyD3m/znCNZG6E7bks2njUR0ltozCtn6L+OrS
WmPFAz3KDZQgDO7DTp1Rop+0sftma03hdgYsJQ8exLmu4C8NtsAj8SwxJxXFeje1tXK0mSrV9xQ4
gIOlj/pHfiqUvzBFykH6aD0P6zjvRgiZYgavOur+WpMekuIJyNgN4HtgTEe+YRMm5o8SKmReb51E
vUAW5zHmDkm7XfDvKgMkpVMeuZjnrBEC7tXoUjvYNo41dsjophm6FR32XYtAcjn+IXkTEzf3LVn5
436GhYujau/nBcXHaDok9wRTwkdP5KqPLwSyZx7naU5Nj448PpCdaS28DxIo3lsuVYiwuDIK4rsE
wsf+WOe+UW3qlGerpf6MSXpfYvFyFwlyCnYUuGpbeVDpsQLrsXeRFt9wVh2oY8EmEa0a7mJcvavc
/7jL0JxMYTITpFS64HZ0wZ0hCCQp8uua0XjwBhS0NWBaGNsAPPFBdWp2tixJA692DZ8RSNoat1YL
Mgz2GQYpDmQbE33QXQHFOwwf7B/weE8NeCUYgFsqM411QKp60H+1h9WxnPEyJJZlsX0lY+sy4ccB
vWMfIpVZmiDQWEjYKv7P5sthuVzwZJEjYvjwTkj1pqkiDvUgxodV1PB+uAQtp2fbDp4awG1nU2sv
9DA8vZ/H0U8AOwz8k42jMinB5ccnWJblTRDKO1mf0JshHHQ9VO6jzp/T4a6pv3KReyJCKQzQSGiy
pY7tX1YWC5U/ZfeUdfd9Nc53/QccrBODDEqwfrYd3VHLIILckZNku3Dcpkc+nTpBWL7PbUysjY7i
NQ7QESKGWGSh72xdCCit6xXGwZDANyuT4uszDRP7WlS1jvuL8aZlE8KCSXPU5XssWKX3r/3pROiy
67XptynD0oehX8v0pnrq8WvpCFrFxS6vO7b876Ap6nlvZspTHWiYaM02HlDYjoVApld1wZv79D4p
6bOo8bFrnPxpTVZHvl+gE312MLe9c1d9gRVQTL/wE9o0+5U5/upC79LVpUI8vr4BVh7JwOaRMJ6q
NlwCH03PvU9tiAMNie+CaqgvTcwulvas9HzyLWr/WwsyfSBaIR2o+l8cGwsxQfOHnHIunbJStGmg
MbZdgW3zNNCzQGsDyvO4LtxI200eOOm9YHtyhAurrest7gV6BnjnBjTP1pTQGeozaVPxQIg75K7c
IKGB+PEISF8NKf8aR8fi4MPl7moX9qnl5RHUwvxsjT8WNoD6ZYqFvfw3Qi4ENthzbLWHojTPIojO
fWhz1iyNzvhw60diVkO0etVs4tlfCZZeLld0Zw9rxvktyMC6IUhCpESikWI89BLZXtZnYl/2+NjY
OZDfE+9i28tukkLufQt/C8JPKUFwxr/j0DAfPl4VS6z5+gcvt4c6Q8cWFktzXq/jabM/nYCz6d7R
DfFXC4n/Wk94q9WL3eHn+xzr0fBg9GMPYDNFWkVPzUvXgueTaXTbkudvhiuEhaTwh7+twuKTo2UP
sOMd2jvKBjfVn1+rABwbAhlRk8fxo3acziT6gPly1yriL3KhoN4fut/ZscqH2a7tVf/PI+fxJHBC
WBlKnce/+JDfrLn/iZEIWCXrZ3CdUXsXSA9/5S+c3jJ4IA4Z9EAA3OnGrbHwMw75oWUywtGz0Ob8
RzYlnJX+vNoZG2GpxEiY7ymyqh5Pbs2xMSh61X4o+i8iGsbQtPrWe4t1x9EqWCebXdH0e2XF6mFE
+OYn8gGpLhH4karlfdl1yRXnkPUoBEaF6ot3WV1YvQaH19bHCW44quhVgk1RtNwS5bGTwl+HT7kl
e00LqygJZx5v/4NrMg/hXek89hz/d9s9WOtMyBDr+dEXVD8MzkaHStwrywQXs4XsT/pnQ5o+QlbJ
YbXnJxxDJg+mdqY1vi2qQ51KsqngcmGw+H4shmQ8gwWmzKexcC8udAh9pB2xicbUfxO1Vybtb7h0
Vdk3WtAsdyLorTPUglc/JgtulxafNSptLUA9JszA9wE9ua1QlSC+f+JS2+buCzOC16CUiedAk9oc
yvIZfT2G//kWz2eB/aHltf7jNCFZCd8o4NdrSZiLWs6eFvKUijPW6zJzn9XV/+qobtaJ+WrTwCPU
2JxDGXHAMtzdrUSuWYF+XGYnORayWCtIjVni7v+M5T8CL+b1zgY2fGJEYojc/JPk/PH5EQqiG9YX
EyQvK5l0ojSiITYHp107PkdqTYZL8FREb6Ch/o+kICdjtL3RNc07Owp/HHRqCgYiEg9JlOe4nAgg
YD7Ge/Ws/Bc/MdkGxBReBMlKY2PCdigFPpjmucwm5aZTqjyuhklDJY78w1kUg+UZtjy/bv82DkJW
cYEvh29Rx1B+PFdFoo1hSEU/gqi/OiUJNk3xj7ktkiDEK0Q7t57rCR5Ykeev//XhDH4n4YgRvLrR
0XUao+F4UGSUlECeoU3mbMEciL53pyf9EuHfBW6TlPy6aMB0okSJdGi2jbpzGvVKNc/JTgY2I+Wo
9Pf380ulCKMGyo7SABY6nK4dRA3Rv3ioWMWsA8g+ep/xQ70JmJHFzQhQ540PDyDv2kCUZUumUeYO
KUKaUfkRBRAiVBDdcRJXzvSVqtorlmRMm8kZtF+j5dIknncEtCqA7XJdwGy6qGXAhITQLC+VzE6u
ETJzNhGEQWyOvZZAuie/wz/HQi51IWzRrV1kG7Mb3UsFO4Gba1HwAL02HHSC2pEa7EIzBy96iqxn
HvikPJpVBBDmx9aD8P9ZqJXOsMhxE+pJA9qV9IUcbF59h2hNv+zwJhXTLmKr8TgWQ7CG0KxDseeF
g7v5QSQU5b1kFPvsoFnCmht//nh0gHErwTaqLAoYJ64pt09eEWy2m3iKDTu/quaViw1Yu93axO/u
8tyPpNJdJBNVInI6RWI4hGThT45A/UlVEp3d5xxXEYrsZlClXhHk9D0f1sNq8tOPV4/uVdjpXLmH
jUiunx6BLvQeby+w3S+KBuJMcvBzjaCzbkXBZpX6rWpsdkBDOVpHDG+oLu/NFqP/8iItyMLr7yOC
n+aCMNJxxCTxnJV/7jacRumbkDtzpMy4EJF4qBLXzZ3m4zqHyk9Ezum7qndGq96DPWVLR6oRvEJU
ZcT+j2kyEeAbyzfTAxq03rGvskpXga3bOT+cBIGYQpAXLdRCNKCcbYisHPKBPves5MS/D43VQFDu
phGkKVSQlefUCNRtf9RkcgxNTcu3d6MqoBugiO99bZe0pFkRNQUzinGlq/B1gh0vXMUY2n7+VQqn
so/m20+G2SsfniM9UqeJrth6vbACZDyqait+8Eazc7MW2YNzAdBfdTb8XA/f9pAG5iSXNFvJfrjm
JYwBXd8r4kx5T+DKbe/EkZ5kZyMHQYKusLv7Pbvbr/7nxuFjsCGnNuxGbJosGO2ISqfI/30CveLh
Xt+uoY27y+yhOTPlQ8FPB9Hd4T50HNdqJqI7n+wav2aHPVprRfF4Cl2lGt7bay3AHlmLKXwBpyji
5x4+4IzvBXrD2gbar34WxFOHK9K6cxBhfk70sJsWa1/6QcvH7a0lz1v3YLsXPtB8GYKgGRdeLUkX
7PqF7GycZf70TGZXv7eACWSK7FXPrbB240EpxS+/nUeN5tt2qYj/A4Dp0sVzUZ9lmetHN/xCEy3k
W6Arhc0PYtXXLteWXQN4M6AKzxP0OecikDcxdO3B+N431J41iOg7DgbOKenQYC1NBJmw6vb1NS1Z
CXoNzL8e19iVnuuNrBas6+x2AGFWchNVtv5BZS96m6C/0XZTgXCXVg5TXKtdnF0Z/JeOXdmod3LE
XKA+4gx9JhJI7OaeJebfG5e0KWxXl7f+sRcAQtuE75mLA+re/HixOHEbbd9HApnSATEiukrJQmyR
fxPiXUGNypkHU73sSQB9wtxNY9uxn8wfOofvy3UsMfFyEuGL/UKuP5zA0PSPmHxpczMHoxcIB693
puK1IZe2djYK7AVvMbkgw6WZhNn8hqkt4EIWRcpETSBZSlBFJKE1QBhWt5bOoVSk10JlppMd4JUH
qlH49/pGn8yC95fZNDZ+AAhGjdK1rPhqZOU97fHTih8uqJjbvOjVMfU1MAOlEKgasUMfFyKUpMQQ
duKBjJMnJ4NyJyyXsLNybSSaIOTy8e/mcDR+KN6L+DrSOTkFfdGHbkYF5TytznNAypjmNxWXkjd6
NYH/N8QeStr2wSmXu+MhtwzcdIqM/aSoAr1kVzqC9sAjms/7VwRblUvrO5f6PY9+P2hiIJQxjiSN
1MNysUj5o+q3fIXTGM5BT/nYAfoynSWbLyfUWRqDPn/TgbnzxvRgjBf5qxrJuKint5GO3J2ftDUP
MzAbxef7JjkYwQsrCVA+2wIbCNCPOlnIuZ+M2Ym9CpAdUjMO6gRJKgBB1hWB3n4NvJhVx6JR3t5P
d9BzDzQZ4U7+GItxnY1ReXO9YWBGg/1aSUTFeo7F3I6ycjK6CHlj45SXsEbir4MR8L5c8T8Oe6sD
EuRR/jf55itE7EitzjOxO7a26PjLeN72oO11jmL5c0UrR8521VS+mAWJaHJvDfGR8JiWpQRGnTIi
yWGGLdhjA3EVlwyluV3e4wjQMELqT3NEVEntxFBq8Gc5cL5D7EMlI+ox5W4dXRTh7DE5vaXpwVX6
L2iMKGBn6XS6MXNBUtnOM1+w+qR/Hdqvm5kmMvQWrN7daK5P1tER5UQf/K2Vb8tIFYuIsUElv4TT
ntjSK2CGuidwPbm9VSySjGO8MPNo3x//gjQcdCIL7/Zeuv2N21KtKXuzIIPS/AHbBDSQPGSwrTDW
gKgddU5+U9eShB7/ZmBDCO43GCa5hufLFszwKxFozNuxwJ889uSzVcLFrXuOurEb7E3Ohc8D++7M
ZxxpFBMyTHRmLM1zELz8ETxDNvmgOOY2HavnyuKwvP7/Rx/KCekg8Q+t9fiLc/foBAw/DBH7N9QM
WD7uyF1lhSk+GF0drHG2B0zdm/OxhwCOtCSbTMUJMICFvdveA/ono68rmwGmjsrk0dWM9txUeG7D
EUFcD/l4MRRJf+k5twbzdxl+itovotDEuSmBD52nSkmOZ2m95TMon/CjbdEv4/fNAO7CrIdnzxoM
7Pp387mhZET/2K8YWKnQ+HDFSsDVsebexacE+CZ18ikTJMhZPEkCrfl3iuZg6AqEKVM6TezMIL3y
7QcV4aHuJ5v//p7uO2jssZT/os9hhq8ksfpv8qtRGdggN7nYdiR8XJN9amb2C6rW84z0LyJ/BfBU
7TTrvWAYMAtyXClT9wK58kFyrEdvFL1Uw8gdBkdYwSZv/Xzw2kPBTtUTeMFzxfRgdMzPwRRY/O2Z
6LVfAAdayDCbg4cWkJ0pWq3CZnTWwwXhKbpYH3dssOzSevPbh+EhCz1IYTSQhl4MUdManvdFzrJ3
vozScmUyTNwQpkX/WV04eKMv3Pp7pa2lBUG2ubMkELsYc+8eEJmKsyPOBFfnZBjV480VflhTXI3W
v7XfE+pao6tau1nW1+mCFkdH3bCt5mOofyqrFJbHuLj+ocHjYB1z7HKXf1haoRAMi9c1DfWQy0Bd
ryRJYMpDSnambSB8Cyn8oobLNa0VJ4SYcWIv7Jei6hqHuFCQZttG4L0Y75Bw4KC8GC/5lrF9HOrr
I+N1QSMe2Swar1phFIdT+WRPA4R9bZ4uomwD4oQeEQ32/T1b0vCN6WMFWQsrI2V0rF71MzrB0M00
m1r3ZF0K2n7MHaGSIFK3ZvfjaGKFQgInlBYUqLAkg4JcMzW2ceRsi5Fu7JvLZoMLFHRjFp9e0qho
mtSOCtBc72mdK0J2KT5LWHSqOWMPW7NVTm2xE8/u8olqHXHd3gRL9OOjCXSOoEZkhQumlSNzDxTP
AD1lQmHNlxzrFVT1qKgGl9pJF/ECJpgB7SGdd9ZHt4NgU4TKHouSJn11l5CnDZ7OdqCcRjSVwija
GFczMur9zuaOQX3+PWhJ+rVanDUCxXLO6dRc+5pA/punVEbhDDs8Hap+g1J+0MqoB7RA5zr6Ku0L
YzARIopJ7cSbuWYju+dj3mcyXy0oA+jxaOp5TAHtcCDLSzQBouydGvj1+S087IIYtCMitLKQRFYo
+NrjjiCoR9/7T19Ni04akRb+lPQOXo8k7ZFDr5Ge7M6A9YkH8fHJe5k8fLYGZylQ81A89HNGKaWf
1o+WVhfv3N2C0hKPw+hYnFOWL8V0JMrg3u6v1T3lxXqtD5g1gChBeY3RCqdjWi5t40SFsK74ZluW
tSmnUdYE6ut758NxvEOCjqDIPUcEtYm8a1Pyh4iU2sC6uOCi5tIXVIX45Zh1fSwwewXcq38x7swn
D89NL3G31bnz1jwnVIf+beDlDhHc6IzA7MECSJEcRVjLrt8fe1Zsxhmaalh+AUHj2OAXApflnY7o
yReTxv4bLbNmTTaJXMFiv/BVBTGeovy91OzohNPP0j1qnzM3nxPOKZerKvk4+Nmma7wGKPceafJJ
sk8PDmx40gZ8lWl0mWFs05dChQaOxD1ERZpwdxfkxqPod5vs6YAYHuP5yC+Mq70SZOw4GBd7iLUh
eMAGBvdfVLbDBNhb8BoiF8JeqCTjNRMFKeXh1kIyxt8eTdSFj5edg5Vz2ISKSaucGvii4it7hp2a
6PQ6hTrBzRs0Mv5i6x4O0Lc+D3ZtycCAvKcBLBStTAcHe4nzJEAZ1X+LOC5JF7bMQLVnmat0Nlu9
YJG4j3v7zdARfn3f3SKYtaFHgwV9M0rO/UTtJLfxVaS+2atxYrRB1hyZNDP7QuvSKOJOQGoav1TB
XJMX8OIFHWDiihodKTP87nKb+d3rhCW9NVuP0lA94KIF73QxjQKc1lmb1RrkzsFBaaBFN+r3NxQM
4KO4siisjEglY5gI+8XpqvpM+mz5z+PNja1kFMetogYSd/Wthbstp/G+e7gIrO8UVpNk8YkpDur/
OvcrGtqhqfb8svvOTJw53dKnKCrEJxVpYcp2jBIDrVPFu99DswLSbA9OjvX4gjOoCTrhK6pWwX5X
/Dp3MdcOrzTEoj7g3EDSFfih4UspjjpZ0kdVLVngS3zoXM+TLhMavm4PdBVkBfycTwK+zNxJlXid
jtQVBdsRSlR8xoKsYt8uerE3LHzAxGICEI6IJK0QZluTitzmCDa323ppsGgnt95NcKXUm46EnbhK
VaRu0vfwI3HCylEdGDyZNzP9XSi0xmH8dHodCKyNmN8vaV6ChQ001boZz3ngrKWOAV7P7jKrgDee
fkThXyGPMTtgd8dduVByaZFNP9+Ih1VfaG66n62+sY4C4va79N3A9Ij/9elPhi19QJo/X2WKDNRI
ap/vJkJudqsrtOLT85Z6n98tZEaLRUHBEEALMY42nYP4t9nkZ7Griva+dLNjoRo9xcf/h4PlhmO7
f5qyrkO1mi/AJjFdu+szQ7PiZhVkdmoOdVgKJHMAoW3Sgha3Woxn2STlORrlsC/hLXEz5V4ucHml
OlHleKMlX3tbUBSD9nq5BK22U0QKbEVbgYl4Z61SYIlg6MfWVFH6dDlroOGdwkZIcF2D7flg2cAx
IsdQyU/0bKktKl8OKeUHxKuYYpYFhPy45CcxOeL4i63jR17juKbjOJ1PUx4bdzHW/CgGVVnIVFeP
1hdw1oPaIVlq922a3XWzap5riKBpyV4Lc8Euy/nOWA31w2bXF+KpD1gvg6MqMVcpPhmkCkyTuiqe
knyzpE+ZO7M2rstECS11zokcVUN5aqDuQMiwSmaEy1e+nbEVJmSfYqaDebYcUi2vssfer4OaVkVZ
8uV5rxt9eZzdT39+i2al5iURCtd3j5Z0aRcTbsbRZpSflX3Mh7mAtA3QzcQcMCpEZktrM+Xo83SV
nTDuTH8C+5gF4ls7FEyG7xQsGM1950o2TXjdDq3s4FRBgVL59hF6926vOY1Bcbtrfadb+QN3M63E
Bqk8kLtifen2YctAPNak6BfQdj24aONY7oHKmgkOoGXyEjVG2jUY8kH6kLN16FzYuyDM2oOofEY+
mKapMEuXb58nD2HovlnMM4hNAvRnKhXLCAduI2kQN6bhe42HCc4uomxlrOkMMycdfw2nO9OWQk4L
+oMmvA6Ao99vCgmCyYciF08RujdRh9vjGDelnUd3GZITU5ldWD+aeq3da2Zs7jsP76kegE75ka/3
MteXt57lGerPYcqX/yaj0Nfk4QUX9ZA7hnDlwNKsRmjKLYCE9GeQKfnfLbyyDfOdHXbzEBq49z70
JUXfwUO0cXbqQyoYicWb3KPnLPNm8NGlD+6JOFdB80vQVq6EGvUpSiTUwmCzQZADS8OovBcQtogi
P26J9B58wdgLjJVCv+rmLfSi791xJLe6LmjaU345DbNhUMFPwN35XgbVwD6GIFLfqxjHdxQ3yjha
X7zLVDo5WiTdfeer4VOB1Gc2OUduNQvmS1vL5+FHUlnup0PIaQmzLpMwzrvA8yMx4ShzIsRv0+b9
dOMhBrF+I+nTnrFc5ijAcI2JVO8uIbDB1ERY9PuKkJMEC4Ec036RR/Mx6I8CIvjF2BqTvdOShvsQ
ST0P792WfH79vIixGv3jsmLEio5VRYqQNE540fqNUWo55gX2qhGVYQdayEzquQt4TAAU9qsLuaMn
Kbdvf31YRcWv9TnEfh3ploklipCWRKbUblDBZOemppxpfpgFHJtayRTFzt3Ft3pPpmtZCsy5MfKv
/bZte2ITdKnpiCu5iHZhWeDeh9rhqD9nurf45wbazJmJxAjyw8XD3+3nzaAiB92MriyrzpM13kYo
Ohhj65x5egp9QL856C78HIR5ex3rExnxZrJj0Z1g7ajbvtxRfM+t19vE+mywx9fgk+wVq/7/JDcL
SNrYBh8f3d10l5r8hUR5OP6fY332/WZbVwRGaa0OyP+kctqEpZURulXGe95Z8s6po1bHQ2eD/JQo
ZqGXiKx1eq3TWjAOqCN37yhjapbh0X7cYAZj9Xz/f7pLwsPPcOkZxmrgaQfPOpdPr6ZvR7tPMK0b
5LrE9yTxP+Gh1RH2g3kYe0AgpF8j6E4Rx4EibbWnQvExzWt4ITRJun+hISUAZ1hNeeKOWXKjZ1wa
EXW2KsPLPl5/LZPmO2UP+pplQeecyPy5te6dQvOjzVADLRRmBFu++LhZlj8GP6MRVz60OijHQPu8
HZ7k0UmRVS7Dtxz0xUWDOXvQ4ohN7IzYNjsrTdmDN5Eq8f7M+5XmV40F8JmDmHSD3A5V5Fa+Pu6y
7ZNShf2krkJ0vhr29eCxPNSitoL90UL91EBn7+6UY+uNr2Im0h7VkCv9ZUuvmek9CltM+2+hn6x7
XV9VwPyum4DAUmCh3gB4/Ng25kE3zGnsnpuzgM23esMiVDX+KJc01Ez/QsmI7TneX3EeZrRWhwd+
zwdQpx6k6RuJoo47jtifI9jZMtW2KgW/boJjmWpnjR6yjC0yqEen6q+mmZufhPMRyNzk/thsft0f
941B6x8w8bwF4weyAxor1drLvJi1Wqv2BTZ1XT7df/8pzvbA0faJ1yQEFv41N6vnooz0xdI0ZFcf
dcPwQk+Rf89iuxaBOPJl3Dfj57flj39NXvukcC8LOIXbYUea4n+A5f3EtD8BbHf07FyspP/AOVsg
FkGNf9aGKB4VQyLwBWv9DdwkoXLDVyRKDejpciq4zrvodnICevz2IxwPdGv32uXvn5yBCmPfwIdN
xEkvTEMNzFXTOsuE914yyYpMjFVp3Xf2xyjANHUwC4N/1F01UzFcBYvXH77ldoWKcUPCcT0cKf3Y
fQs+p63XsIaYxMNPThL+KByOQkux7eFgufnN8nNLQ66EAcUK17u61uKyAftIPeNwrPSU7Vx8cZ6G
I2Vr94+X9+ZfJJ0j4lQyLL2oh3kPRoR7v10UP2J2ujuwDYjSzgyZrXBICynFDp6TngcU+UKkVT8Z
9ncO0QeNRqZ8i9K1tgVa3K0tvk21w/j3wIbQ5qGUhLX9WBpu5BWaeJhU/ZgbzhfP4DT8XP0naPL9
9AwTT6FPjsMhLFH7gxsdaN9c27JbeCAPVIvxcpQ/4nzo6QaPHRR4efeXDu8clca5mcjOL5eZArj4
xhdRNdyZy3ieLbFq6iwlsiZAmJU9iSBaGw/4mKolhfH9VXj2McuNsMk+Or2vv7bG3Q9myO4wLBQm
D4sYBK/o9cBrQod/GOuS0X8gMJYgfKLa5ROf3va1bMOdul130AZRRjuFy7qNcm8xuQnPZyr85tZz
dtlCogOXDWk0lriPT7FqjuaPRkZO585Q6+0Wde5pQIDC3z609a7gtZAyuJ3qRv1RlefcFAFbFh+Y
WXTG0Bth1cKOzawlEn4aAHbZYjxWATfjM2baP/ETX4q4pyGjHOpdBiLCajArqNVKT2giPucPeNtW
dwSEE4bqutPAWNQB7Ji5W2DZB0WDWUFYq6oKfM1JwipdChTevCBDoO8SKBTxYATJUchAy3EXawcA
4xxH7eeYmEZJmIGOBz1TUYD8F2WIxBBOknhwi/podR3u65HNcfBoCXCPfM+MRib8iuC/pT228e/N
aeuIrfPawdDulTE4nHNzZUA9AvCwHD0qd5t09ZXiz3E3P2inXsSW+c+nVW5VnFPVjSSJ7By7zm4M
DL3oiccOtKGezggeHJ/qHiY0hEmcOSywIBVVHe9IYsDVk3vYB6C8BbgB7qkvX2mUjRNoUCYnMZaj
CaW/YUaABud5DWHC0fIHhK1NvpT5zMCzNfAzXLHDK//LK4abqjeX5codPy6jTKxAWUZvCr+YPbyh
v7reNptuBLt9oG2VJPcDiNMA4YJxbFveEwBFkarZk7zoRb72kGVunEM2CMBfwRKcHo3vtmfOsIo9
NulDvYoVfpkR3RrnPPyOPtpE/2XwJRyIMLHZttIDD6k30jTwnA6a8a5H9NIg5asHu98XRz3Rng8b
hnIJXwZLWzYnlrP+51q33q/MR7Gvn5WBP63+22xwXxSfYj9X0MQS3iQ96SRHsbQtZAYg/jjuqfNS
y52Vl2PxOMifAiwMGvB+D/+lyBCxOgog9azC4qQcbg+gNpJCLMzvnaq7WQSOD7lNdNkzNe0vgxbZ
8ACP43SBhPmYxk4HwKirJU6kNOFs2kA79Q00hLwfNUoIO3kNxh4oSomfxRaAh34t91Xn9VDdVCaB
l+cG7hrjGwXIcjg2H4DZwAcG3xkx7mPksNZ8UWrsszlxzepCZrkKzqBn5OvhYIJ1kfYzUIvBHevM
BFPJUmvDKsWJHUQtpzin4qVpC54gQQQ05o0qFl29JkZWdN8c9HUkwSmgq0/0feGjAjeZpuGIiB93
PCdC7l4++AcZXYilwdy0zgZffQobjVUqOTUK88GDohASL0us28I5KPL0zfj+XAbzkEc1BhwQHEUV
Ss6o6ikrhoRZJDs7ZCGGjWdhVf/zZAkirxRqcF2zfqc7m01QrFa16ZUhcZtwS6sOpsWvubh1LvsA
5O5li6sXHL1ExtXglE9l+lCUlVW87mfAJ0VKf+X9Xoptx5ctb95HdJv+FjdzI4xSHqDLkiJqP/tH
lHC6nhehnG5YgX1YFEkiTFh0WMPT40pjRCtypvCB0oO3xp3Bz5Ogtopj5n9169sYoN1DDUvcqYv9
x/I4F/6M4Z3r7XA8AcGnNDNywGZFCUURmrwHarpzkgw7A0dOBbBtJIsgqNqMhfQB+CrunABGPvLt
gBOXwZ4/edMosUhGTcSloUkhrFqndDotatxrzwpGIGKMRM0aAfRnJzaG+7YtZ2b8DIFMbwyQzJll
wqLkK9uv5rMYZwqi8Vh6xNCFTyCKHEc0dXUufoXSGtclNJmYjZZ2cVCQx4BFxWOo/Uo/xTHEB/vt
dnZnOEfHX3lWejb626O4QpfCvn0AyErglZWAHzDojslTsqUYcwlqZwgzR6vIqqv0mfFsnlfeEAAm
CCpsUTH4iLQzVx85UT+SjyyJAVXXiDDDYjhHfsm8CBQmlQLC6XsuDj4Afq0xjVmPpPN0o/k4ddR1
HFBeGu3VdhyRKCi+QwqvZrMwoPp+ANen+9a3lqwkol0Pt5Ll59K8WIKHsbtUcTvl+jvtHbwSQtdZ
MrJdfPA4bYX4nUJ5Hn45rAini2d8NfwP38HM4+r9+OTmbXpPdV1awiOu6HIw6wHfCVfcJI4oBujR
6NUIIO6df9+FEQTL/yO3b81x4UQDyL47Wlw1geAwQyUls2Fdb2qgOax6ifyJX8Lxmi4k5SdDya71
YYPnLK2YJbskHpY46tVNwLFx9TyGdJHiapzUi8wcpWv8KL4QkeYVXOVF2ZQQD7KBopcagMA79X8z
LBxCrpV0x5x+Tr/qMEaqPzmRvPDE0T+kPZuhsHDmoxOPmsaX2CCq8065XOQqsIVBu7UNqWCNyQfO
k2hkaFKldpSi7gF9vmREWxCcARGq90XfEXmDOhLk5rMqz+BQaqFstugI29goI2h65ZVGpR7eZPiD
j2syO5opoCCNuofrV6DUV/fnuHZKRcjkKrHQFPpZVQQhzgJSKml5OQw0LdyZxnWT57n2JghEV3m8
+dS3rzU0pUzeKB7lXEoSO1+7HYc5TVP1rH1Prb5zHJBJyok0m+u7ywSodiEWjVqnCk3mt/8Y2/ZN
NRYq4r8mIJwW3E6L+hlxJ8wyRfOT+4K5HP8Hex7LLkh4bI4qaFUprncrjiJnffI/V1fh3fTgUA2p
AgBE+j9XfNKWNdzbfzTWOnExJsougMQAHS8P0IArx3bGSiq6MyiGx0Dvg96Hxy66RmgNahEI4tIV
VpKbGokkrHxR/f38Ovy471rsukgjj+7B635HOMAWmQhgXdgpyC4Yt148xZUlVYibQA3OGx0S6VOT
jtTtHkoMj3BZ72/hdHtwOt0ZT1rLJd/h/a3QR+Jja6rYBfvft0b0F5w2dKGRSkFBnEjA/l+jMo+C
nsoyJi8VtPE6t/g7NONPxDhUXnMuCPBJsFl8ipSrqMA/nC2io1ghoieICBhsAG2ItSsx8l2UjBst
NOn4TruSj563PYAm3r5ZM/NR5ypKiS5zekuXPgRxSDmBWYk2UgmkGtK0yDFSyFK9CrRU4ta+ydFG
WNYo3q5upZ8N4RWTvqy8zxwOkbJNeEn5aQCphDJLlQ6KbSvCWwQfqujRVC9bezY8SP0+TBXjb8jQ
pke+coCdrxGGkUhQFf6+LDlT/I/EkN3yOZjmYi9dJYx1zL2uu63NPd8lki5TpT3YVzBOB2uOXCv3
vXhWbnzaOzm+ies8AiBm9yZjHsLbR/XM44rzDZLsvCZaJWxLZnuN7j2DHWaBd9nk58BM8xE5Pd1/
LSYkLKA0+F+6h3vbR+fulgfnC+fJGG9GiGmSJrGjc02WGNcf+4C6sIU+6WXePtyh0ag3xVsGnPr/
k3v0EmnkHDAAvqWXoaJJyRjQhBojk5QJgXCbaDZacD6JZlZ547lkObLDU4609/Ae4+wQZIQOQC1E
K1TJnmdDbAUuy53QPtw6kvRYYh5Vz/21gKBi20znoXMKiLgbojHcNeaEUycRy2lkmguZojZ1VwLD
HLemCKdeA5x3rn+LZblKkhXhC8Lk53xhh8FniW0p2dbAd9u0oSMZFY0k+RS1IpZTQ/i9qwtMccN5
0uADbH5r1ZtrbJgDPwoyyOgkburPFhOidiw98UL4fU58reDP3fBZkPxzA2WCy9vt+ySg/YFsEeyG
7WMpB+f8cWf9/heHC2XjY2yIQWcevXUOkz9bWI+Kvk26VpGcr91Y6TVqRARfHQ2pazNr3wvAJCZ4
noQGmAK/vLGeU6pBYuqdVqIwv6jMpk6vTWC6YzVlFd6j18S5lKj0qlbTrWMqop4H4LMb1GJWniVr
G7Y+Eps6oOsv6la/Orcgf/XUKnUzK7c0+I3d7IkCw7KDpBYhrMq40P4VxPDlxLDnOscvpVuzh2BL
/z1kAShSpkjJ3kH1nBrIoFq0WFHOYjdJXuhbK6+Y7P9z06fuECGcgFJtHXdI75/ljuLS0Cc6AdtA
7XEMcCzsx7IYLkDmtAlPs2P1J//fjS1rtbFGEZoysFBJfsPXAvS0m3AFuT+vPC252AYj32i6KxVc
SZR0rgkaDg26jDSdvbAsGO0UBld+iVUKILwPiGNvRAoFdUkB1ha+bj2Dzze3Qob2epKdjO6mIe1c
IAaoxYokv15HcWG3xx1eXZKUaTCMYHUdlJPcElXP5GnGH8vdEzk9r/qFbdf/sLIOJHueQ6jc9DdB
T5ucSbTQXPOKhLwJV313rcMs4peZNJDEBqDu5NIraFOO0oGfZ8UxFh+2GozkyiIIlX1GCgTONkXe
Q6LYfHCUOf84LsbV7vGZGe803VVElQb8zpt9ByzJwdazwB0RAgEwD9e+eSCzf+oLSuFmqxIQ5hTD
5Tm12MQYBlYNEgHHWI9HL21pcyFFGXZ1x8g3jV3HM52Oh7k0JP7s8SHfRKYorxydUyeI8NWpyV+j
ApNyhDFsz+zTnRXrZHRTz/8og47FDg14tZYVMwbJUK01+tqGTjb8Oc7TAJfdGKNDPM1MuCb7zcFz
Ma7A12HQp5sXq94vE9YDWMh6FY636d5t8AHHJz02kEPbAAlaPvtFsD+9T7SmJ8hD2yYFb0WnCWXe
mV/khbMdlmiXvK2wIF53JUzwWBoU8s+g6+nRlpNJelCG5fY0+FhRHwB8jSABgZWgECHV3U7+4me0
pSi/uRyegeY4pOCKCUT55s9XAoCqgbRh6dDkE11k9JW5Qgb3emFdQ2Pa2wvq2noWYgaVagSmuaZd
f6O7TfnA07Afn+Uh4TQvOHbGin6hsmQamLWX0CPvWN63fw8KfQ61kSDycqlueWL+k0Pzq52ELvr8
hmHxRZpi4LBgeE1xQg4fYfnWMGRsr/FcpTDS0z/L+psIBd7uhFiP45VAgR6ipjg7zkzIH1YpU4+/
Xp/8T8h+uR3L5oE3DFEmtbgxNmiJiGZmHHw749oGSYvvsUOzW1MKZfbSaqN1T1ze234jIrF9jZKL
hrzS1KMSM30PG8I+4lfMLaYrTamQp/wlOWnincdX6o7dzTQARFdL8d1rggJTOFwvCFBTLSFoqL9p
X76By3j57bAsIWHTsdtFUrSa7+PNMOLFE82nilvR6pIXS9z1egzSlK+JocUszPzMK0XT2LYZFJ9Z
8S0G8vl5ncjWSa22Ev7rwG8mYho2rB68YvVTBvkTcr3qzVXby3GttBnqLTUzuv67d16dYHA2qhB4
YtpQzF55Fctpl65Xr35R6jr3aVhDt/L8wCBtKsoXVcDmJWtLZ5fAABReymh6WP3zC7sigt+T2oQN
xYgptY32UKFnN9PbsI5VxXH1X3p+YNQ0DlGbHdnAAmPP9pSSbodfPvbiOMfifa5SzyTTYpcCo+YF
0u2swSehlQsckb/DngJ7Y9dUC/qXLFo14e1Lc19KgBTCNG2sF5ymyaDnlFREoyK4DdJIggVcgNWZ
BkJKyqvO6N3QpB7QwGEN9OD+LBP8qMdwN5UBQiIreTcXJ7XkJgoz7HBrPJVQKC/btiAq2NMTnKhc
/Gy+YiqkfLyjNMGKeWWXqAcdCKUdGu0SXuj7Zx2wEvrwTOJqT1J6UOSJt59b6Dapi0AJvfxTywC4
o12M50CrI+xmCzT/jIF61Nyxp2ZZdf40vQnahnbWWFxN0Hnt0a15ugaDLiMtNj6KVRXaLgfxJoA4
uHcgPY3EmVHAaXfIf8kH0+2GUqnpp3K0RoKmh/3z43c2isnVkah1b1TbR8EAy421u9GuOdb1mVqR
Kt9EKOeMa4urMOkjIQXs7lJc4Wamjd8+7U5clsHijLMbdOqua4eBKPO7XYgb0/ECrv4azziwsXtR
CfkEE3RcSPD0FJwald13UK4CPuRyacarfY0K2OrRd4faQgKW538dmDHXQNCwwhqJlgTD66Tn398h
yysZw1dMYXPhYU/xB7JegeCk8IJ7dN1n7BRRFTSMtpYPCsWEtCIVf3SyJcM1x0XkOhAf/84Qd+k6
xu56FrVGYgs0NI660xLKqa+acERA/kTyf9OdajlLYO2uLYOLiBYCB4kZqTqqlYpT4/o98BD07/Ay
vfFwHxDyTaPSOnFxPsAH3cnzpBLen7/12fmwrYsJRLk+JNW5/O1Fn7lvyHmuapJ94lDv+BD5KIK2
xz0hy5Q2Er4qmVAscXZ6LwmeixNfLIUF1CO0+NeeJDM+CFyftvAnoDNYVuaNRJR5iRsGMsnAOqUK
LqrgFSDK6plYl1kOv5LQISt1CXy/p0kETyn+hF7MpRFiS5+NiYZpwLuGFZp/WeILP12+PgcL1UJd
7opr50TLhXTUGq/mtCMK9C48tWB+u+69e9pyYyYNYNsEkwZEJZqJM8P+MmayVn99vZfmsrPr0u3y
7UXyAddz1y215b6H2PiLA7C8mLOqYI98IA9pCKi0qZPMgM606370icxWhdLMIE4QZKo7tVDxgQw/
7ifOceCL7uGK7SvxdX0gkqJrFOuLis7UvDB9Wug2xcXRr0o7kMEnZY5h3xc9XIpUB6rWLxhPgUed
0EJqSCHq32SrMRb4qWOvZY279Vi+kqM7H+rFBnqSC7+Q5QjRUONFstfkuGFUDMIWKCmA7jwldECF
o0X7/hAPrtg9iGWkzcziCMOGQhL0g9cX91q69ua0T3Za0vO1wCTuieBUu9zDyJ6lsZJux5gPTIrP
/cBDOhUKi2kOUYcXbobmNiExCtyPjvGA2DBxgHsvABUDdwXP3YprVVggk/nSEb6M/rJq9T5Krlej
WdQ2dBrh/bMRWea5D4M0NQ3q++lG13X6xwuHC8YSDk3Y+Vsdh/zI0kLzxUHQznCVNPbY00GnBqdx
LWwU4Hhbw7UehGLjAVEksrlMd+Ar0lMJyQIOrPDzSIsYIKsIElnDSWtX+awd6F3KGu8t4dYN8Zr/
b2NGsT8zkO2owqFAJ/sYddea9rjHGcfZJ81ZFmHVtnBm3vh9HrCJRISzPIxvSLAQ5G2IzWwpj671
Z4Jei1vlzlbsXTn0acJN7mne1IKfAfJxx0xakNTFBa4SK/7DYT/MsfW0mtodiBHQIwC72umqTrzX
xVDYSgpHjaLzh7wkxRLbugS+5KT44BcKZYb9SWhVstvF9E2cvaRhCxE5VsqMUByaw9gjoxziso2A
aXzhAlRIaVbhj19Z0y93a9Hw+HbgA6De1G3kmlAra+mEA4ZSU77gKSeAHPe5iMknZpjn6M2iAye9
b8KVEeABBXMeEhAbtq8P+60smQxevxVqCTeN9qZ8iEjGgT8zkt5e/eWjsOc7uzWlIXW1YLRDu7CK
hdJfuolO84sjjUFXaWm4DWKQIE7E+WiDHZDPBC/VJbokBCP7qk/HqbjUz+L9lfpFCacXqIa3qzOM
2gdWWpnLHYwSQ0vfTMrKVVIQgXMBQ7spuHT5KaumN0bhm/hCrmK+XsWgzOl13fzSa4mAXqwPvo+z
ZLqe/PgRyHYZxzIh08mE2KGtOurLLYHEPijbfbG/68vFE4PasAhmw/UT/exIw9H2NiErDjepNZV9
11GYPJoJvxn/S82oeYFd8oOF8J8kCX337+f61nHXgBouP6x+WCKaKglqiExZbfaHmd5VuRS0hCSg
BiBVXFBjI9MHIAmTiFUOfJ+JUkecHL5NQdF4xQRQLUMZoSaaaN7mKwlvh2rUCz3muDzhZoV5CC6f
00eDwHMeAGRitZM90TW6YbFcElxpAPGorYS/btgOXiEshgJ0nZABzZQtc1KzAMnUTiv/xcVBRCuh
iFuXLw7o7OaFfl8Pf4EU5i3XGJ0W/3jooK+P7CgVt3k+WWcvoTUhhtnlhGq8/cylfn5x898+kAAi
VwfNrfSvPbThTZRjZiIQd3J8dtk1N0HrDDoRofpKoaCH02AmARYngpfdw3vAeNd8vvxBZ37+uVAj
wXpN/4dByhc8tRl8O+7tqNr9eHU6TMf++HMgnd4Wpc8/WD9gl4TWPn+7AvYNtuImChqzG75QwJE8
ZRPR6eCH3kDKHH+ZWI93oXiZjxBggmCujwddqirctMqXTG768U+yYLOmSVYt65KvgGAhVD4ZiJLL
EyzKM36a/FuvuyFfJwNn6b7Yv/ZwApWVxfBT0xTDGLa3kc25UNpI+WuWP6TOL8tQ71E2VxzBUYp7
jJPAxOgaKUZ7YwBvjMP+m3vRYgIIQRG+R2TB6xYYWyfVsJUNw9q4II7sazXLe03U3tkAYxlpAYGY
YGxNwRUC7GnBiAbF2sZ+7iaA6UV5Ydrf6wxpJpPWfs8kfhFSgawR4Ien0Sip8FdpPIXw4TZrQwQn
9QiSEOC+PGw4hTdibHgqLTRvliaHn/bzne4guV3J53/ZMw+nFNEoj0Gq1OUK5akQtWpqgpQSpJy1
/mQ3HIM/cTk//t2egzTzq013iSDH9/bn+B5XCkeKV8l7UVfHEcmoHUv0EC9dtzNwMSGDluEVPnjp
3+p+25pzTFXNG58JubdCwtCEJWrs5POKweX5TsThmWmPBmuuGGrtOEhihWZ4oRzyG1WBBTkL4eDE
W9eiq1PMtVytu3Rqj795M2BSvQyDtE+vOfad6y1QzPEylb8YKK+vfgHUd4Ve9nMF0WbGwTaBtdB8
Sjbz1xdCfmLnPSiA6t83dqptQdvP8XWYSKSetXqEHkwue0OwKbPWYJhJyGHaf46uXBUvcGkFB5ko
z4XwU4QAw4jr/nIfCddCxeuK9HdGmtYclOCGBhr9czTaJeLiH/JcM6cv0Gf79M2fcGiNpT+oVvnv
sh/96NIiZA/o1Mi4rERdl8WxnR+5wJveh74vFuexeYGfeAjzzxaxPLWYLwanzElUGqlDjHXhkG0a
LCB4EcKuoopLwZNVBIaLhc5EExcUMx7B3VHQBeglO4lki/zU4nD/DxPUsm3lYmqAiXZhMWnpZ3lK
8nzmIeuTgQY56R8iZ9Yl6BFHKiC7kH9/VeNi3EEUVWJsJ3ayLNSWYgnA6Va0OBCYOfthAf4gBCov
CC7x+GVnHtMOJg706JjcEcbgJDXqs7umo/8AOoPwtHzI0Fq/DRy2eQkeyby/8G5KIbkhuuAChNxC
j/GEgc49kfiS6bi7Tuz4ChTUbyuPRMg8aLHnEGbSeJs78VOM47fJO/f+BBGWd3teOP/5+LP6FWCS
H5UXtX6m8+Tu7HbBTLoKZN8kEylN+eD3vqvSH7RQsYUKvcLoHeONBHpSq1mVTKhqy7CyhsdkZqqa
jCriWtQUYNEcnnXgVzKfHy5rEMQIf9l8Ms1DSzxmlohg5Olt/NckHZg4w+HIkKrLFrwf8hWRp6SN
+JsU9a1lRhgkB9gWJaFwEfWvdJAu7j+lk9sdk8w1HTYnwtwKY9YCXuvp4xmtW7RfvwX7QCcvZMqZ
5IFv9Xci/DuuCzRMev879j3sONGGMv5hNx5J7BWkOld4e3tWG2fPgvDu5xxrI2zYJbTA371dliR0
BFlhHWeMgCjb3a6mVSpE9/qnl07Nb+k9AvkUp6MaM7PloL5YQOguK4GI0rK/Iek6Zy6vCpn2oTLQ
hO6mcyn6fDdVs7QOTe9O5isKc+6a3ykWFbNW49jw7ISGfxlFKT7V2qSmaNgGyDyJDC4VbIxqtsDh
pFlWhC6rRZijmV+4VZOf/08Ip/XiVLM7wVjh+iUJMRaLftFZlVXN6n/vAeRWI+nYuXYni5DmKwkq
0FGsUyIJ+SkCRkZ40inZd2JqYazJY0TubVm8k026pYAihDRpqh2q8euTijK43RfzqsCWQWL8Wote
wekLSVhAOe9ZZhRwf3v9PoTyeMfQd+Xe41+QAZuyPaE8znHe3Wp693uZz2i52sZdEBG4VQO1Chf2
VqfQYmVtXhvJ8x0sZ72bbxJz/vG5eL+b/FfY8EaMd+rZOf/ftOk1Fp0gcYc7tIS4U5URoVx8fhHj
FcN/Xt54sonHNaqW0w8Kl1rjBgmvdbiFvf5hCtpxt095+Txdq1cJFZ02/FoPXWRD1KebRBZ6KMYJ
u/qX+pz/Ud26eefXO29waAwzG0x/hy5rwBu8pvRO4yw3LeKdrpAPj6rM2HyYbNtZF1hbtAVNmkyB
KAeOnIrt3LrMTQMJruG0XU+IqpUH9MVWAvoSj09WcuKdQWC7xA64eChVBMJW1ajfrcK8zt/yIo2W
0N+ECtnxH/ZkwyBqsDUVmYPQ7uQDNuxiVV8XJUbuaUi8rzg9zFaV2bWqsatMXd4uT8Y2f+WDotdI
ejPURw6gbL2h7fveHLVXe0cWTP0Y3XgPknmpjW9i9Z7ut1DoXhW3wnADUqKF69He8QJYOK5imY/z
6IfjPXyXQcJNiw+/ibPdlMaKv+H7nat0bdlH5dEmaZfEobhrrKF+xY+zVF4Z+Tt/pMD9cvrJpxkx
Zeh+IHOgxTw54udTJ5j4np78gpeiZUO38NZoxbQQ/XtdpVgekdNlcL7qAIvb7Vk114tGwAjLEUMj
1rurTQn1RMAoizFwouuzextuh1Gg4w423fqr0kEzQWa0iCq1EZLoHygw/Lpzm/x3rRWqSQ0Wpif3
cpajx7mKedcQbwupInMqJ9tAJCbOWH3h+lGSQHucquVYLn+wS0Wgr78CTgrtPTEKN/syCREZyGEl
WhWDsrzdkNAEIzkOtHcEqxi3NWWzFfuUGBj+BiWsl27UXs7RMlTJxWUF4dGmikl9ADVAHiSjOutS
29KRfj1pPy+YAcIYn95ZTHgmV3OicXwQlgkDz4z5a8oUtGknkaVXjL10EZM/TfKaQphwRlBsuZsF
v9TP9K3IsdB1lND1fh+SHgCAbVHKjkyOviePYawMPoJPg/FMcFH3HDojMSYly21L8/9oO5/39ueI
12OGtznW6DJpWzo/ifPncL2sj4Gu4yEOtCfVxIHLM6dehpfdln/QZrw8QU+mygUpUT0fnETAgKmi
yjXuLCwAeCXCGWmBizJ0O4bCPJCOj7gym70bWb2a+BpZoPt8B6yTJ93dnCzuqVr1LwUqndDJWWj4
n1FVYwB8BaA9ZRqVeDEnC8gmOxuONUpnXMyXVK29E0cmwjmF7Fa/dcwEg3ZNOTV2TioWeTo8NmaK
mKBGr28p+6cGvQ4+mf+CgK1mLCA02/XzC3wOVPZEPCXZjxiGENdFDdLnrEbcq5n/k9BvuGQNACb3
ouuS1JdGxijHSCzpFv5vjXgLvw3P74LWp5OuxVVwqi1/lCxtxe8mlYBeLOcra44AKT+hn4S4E7Zt
9vQH3OhghU7Dy5DOYmqxzMgqRqwv78XwwQBomBxdUh5WSD6JJAn3jS4JWUZITuktxl9AU++N7WuS
cKm61xnt5+83WDzTy1vFRlwaJx438UmFDbj1zmh8lIbH8K2xSVTIi5ILwHAzfJ1VqXcRumdug6XD
eyRL9AlasGJdlzvh0DIKP/my3zTMmyxqTWB44pISRTuA9pK6rIOVJydyC14THNeOC1GhSknplS19
CjB4DHpDLthoyPtY3oUN67/Y8F+a0/YwwIXWkXkg8G2qoqWcoFcd8t1JkuOR5bK5n3hrzrGZuuqa
7tCawd3gnGxqlhCA2hr5HQ0/OsT8yfIc59CeoeGHYHkzy1Ge7zSFo9gfOn6SwQeBy5OrAsFvn3ZC
TpkJNBzhkx9iJJ+JUOCz+Rirg1qK7jdD79B0OAKEUKD1vEca9g6rc3TzDzVFLXlB73PMBLs3fNN4
k8lR7Rny49aPDOcpTuybp7Qqxyt16O/pZpNEXgbSZYz/G1pGqE3pP9RXYro/IhKuydUUPjyRBvF6
rDYu23T0SGx/xl/cN3jWPvIQmk3utwXFVdmqmlc3bBtMBTjIgEdojS4dkPc/e/U89nZ9OLYYppLm
NWH8v5SyBy6oH4PQrE4h2NQjlskxWa6DPnWNadV3CATQrZN99z/5MjJcmPdYJL+ot7fLWXH6QCoI
hemOYBw7kHsDfvGN8hiSFqQkVRsh3aqVFIfJNth3U1TPgoChMWaJLrwAYACgfDLoIduGs6Ra3U7p
K9rmc+FP9vbdAKeGwYVYZZGGq8ZVy+y0wXdYYMQFz1PEO28wvoE9gyzURwktHnHXHRAWP2v437gp
NDqtpgAVsQohrTJEF9J6LXrTHi2AryIYI5m3lICufLQuJ64uPcGQkG7iC5hqd6FtzlE2nb7Y5gZF
4/Qr5VNZLveLHXOuBf1hSG9wTKBlD8KdfG2prl2dkML/mkF/nurf7FSQAQM/xrw6cwFAM/LLqUqC
09ZyHjoil/vgR64limBBJDCbdvrx0VCzz0ZV9ACQUvxoahKDi5uIN1pBQyQy4NAWg0v0FNxLKj1a
cDklOxNgoCAz4QmVquh60KxXEznQ7844HhArnmIt/aV72UAHiRl9CeU0IxlY4QDXCxxkDXiT0IZZ
mdJwIpPBYdCU3jCKAWk6YSl1PoJTdSY3+J6SrvjmlUmS7KVGm8g4iUqEHy9KrsctF00yG8mPeolw
+D4Uh6n8ZuoC5K6hsL7VOSbRX7pVw/U/0s7dlkUMPi01PyyACF5EeDTAhjzJZxf+pHSfgTyN/nQF
O6coxKEmHJLJXeVTatWNT5SdiUnNCvTDKC/YNcY8ANMwGaHXkdiPD0a6PY1QoTmyYdcyZhKbx2Bz
zdANES6BDL0t/8V8dOX3tb5a8w4y5DzUuL085D220sIIiIapy0ADXwBS0zdEpnyU/D67z/MIWl0a
kUh5rentCBktIXQMLmZuCAXhPbyiut/vD9niS4dKZcNII5qu+hEYcra2FPE9xnzb1EOgeXle5dGe
qjgYIzKAu5nlROAXB14CpMV5GWSpDNOeU53jV4TWr7gwFVId+anT38O7/NUGSRy1+l5OejYHxYm6
xmbFjqp5tWrA6PYdDko8ENovsoeFfnsOvNaRwxTIVuMsQ3W+C6zduSwyStSLkqSkaPqYpyA7UP3B
ZtY0nipYbmgt7s2zoT09kIFyW4rqW64g8UAy923/tCR6Fexqh5ZR6M44P8pTU8xqa+GVyRPUilil
wMtKBtRkBNYzLveRzjJ/Y30muzHXTUxC8zYKrCWxHACpD1R1FhiycQJcDG5e0LNJZlh8oQZLhiMU
xPMWyTM+K2VOHumOmnlRBy8VSJeCdtgNlIuVjdkLSpG9eP2znvVwXQzVlITeA88eLI/D+p8pPMON
60zKfNqZ+eJSRU+E9IcZsZKHoIZ1UTZGK/IU1eo9tiev1Z0PClg17SBSeqf8r1TvxQ47+t2ZIsTS
xeDH6mZtbRB0NsEP2IGDL7bA+zZkiVUlqXRxPJwUep6IDPoxLfe1rf+Y2Nt7ECq+PaNEuxTgV3/2
Bkyd7tfxUlMGo8J/fWIcWyoSNf+rqpRGLiXIGCj+t5VeSAzfvIwcmvgNOfVFLOhcu8ygKUjZatuf
1sq1gta2rHKxOSBPxW00stsrFKF2loVLuRYZ/Uz+Z+Wx/ZtfxKeS5MXP3MJ/HEUqwWFT5yMhw2/0
84UYcr/vUeraER7VzCBhY+gKSzXEYcMbvSs9e5kMky0nGNGfm0tUdgoIRSd7tWBnw7MJ2/sjeLw7
VJiQIdBuo9bGQOlhs1NUdxKNpUNXkKNbhFtp9XuuDM4eL/k7XwvX6NxnAX03Zlf2dOscrCZLRgY0
OwuC4HD6RvDN58lFBRYoJyrRMaQh3B7Dd5TYbjE7a603kBnpUvhDhBYerrYp7U3wf/VGZEei31bA
0iiPfV3hs/YOEa+U+JN9ojzfQrihnlA1gUqtu9vFIXnL2NKoEkgE+tmFfnCyqyrW9qyZKVvzbX3j
00ovejEE78Q/N5uH34Od1GnIHpOh2PaQjd1kIYvwbVyV40jdTf9D8uur5g2dBGjsh31l5k4ZsfaM
x1vRyawTg4zm0gyy+J24NVDibRVzWfWW4/WwR6Y/MuTqZBZ4g7QKOo5uX6KE5kDKjdsDACQbz3kN
TPkro/DEkz3YlvDRIOn4OmVCygxHQyI5KBrOmAaAwlMKxHYisuvMKbLT5C7Bby9SJouXfEctJubI
cJuO/Sz3isoktVeJeqixmvMqgUm/74WPZf7jc6cs1Ves1avRkvg0u5Zlfoi/9rvXAp+jd51TOGh8
g/zLyVHPSvgRAMPW+DXs7sEtykINa+DYB24oFEsiIiuNFM0bAtcQ/fHsOgE59Vk25Zr1WugIb46x
D1Lx2Pr9ko9u9fQsOXKz5R2KhNWmHUc9QhmiJPFfjOx2TGpRfjQFH6mzaivDMyS51sywnAD/mvL+
SzQAFMyHzR4au3xLNixTfRl/QlbmdMWIrhE5+DUlTIqoOiyM2wtvQMYzqNj2qxpiuXtOkQOUlEzX
BkJDEitDT1ZVuFWaVq9YSEr5TRivgIOcUeduIsW9UJfdA3g1Vmd8ny6gCNqh6850lk1iwB2JYc5u
HWjGUwnPEZ3TK0UJujn+FEojy7KQ+Qj+9Jfl2d/sN3x6pzCXiY/oljxc2znb/9H+1b3t2SGOGI8b
bM4kSK2p+Rks92PQC79TeYLnwpRfJ5ltQ3q4uLDKzPz9uhB3CvkQQC04AremGukOIZk1OwR59nmC
x3flnOgIcW/WPD67TYdM/c04SYyt2lWmc4hEoJbr8vQdVfv/YhNqqa/B5E74bCkTaFSNSP8S/X8P
DXHUesVm13g0buCz4vH/ZsvJdAx2OxULhUqXVT3SPZmGXpZY7GpePFW//w/AAkpG6nI3IYLpFNks
W/JXJ616IwcEEUSmZbPShrVgupGuV+HeYmTe9X6lPrz8Zi0YuYPdUBqdoGRMP8j/VpMo1nO20z/v
OItPpdbX6b9R/U0gtDvKvGYP8yPOTv/wNJCIsRCQS7EkOxvU2yjtmuKYVlPVPZiccV0cJZh5fTTh
NowcCfRmDi8IKMnUXKu98XFfTCzwKujOTz9f+SWU69WHK1SOhTKQZ1B3Jme1Rq4zN0Cq2kmxBhAl
2PWuzfnjqMDgknL5rrNY370QzzEsETYv8xCHSlBRi4FiSZN0+Jr9su4iTpTAVwn6Fzg8VPVdQzCu
fvCMprAGU1Ikbr+btNXo28ZpsQYGcfaeDe7mJtWa5s95taQeuXKk39keIrjJRS2ZgWkVCwbLtwag
1ttF8ZQrm4XaHTWKOYNmu6U2+2DSyLQ2JxM5pPaO4Yj0Slx2ZERhtfGu6LlZSS3kNKHgdizkDucL
P6mDl7u4/xgp1YlkxsQ3P/Pudodr0SLjsV1y/UchTyVBYNcG3lhSSa2JFULXlGnAV+L4hHqBuUOi
EUQQyTpNI7/YCtwgpOUbhZaaJ3u6ag9bf7OY8m6eGMz/Wt3Uy/ebuRyvRADe/8sGvYD4YfD/+NDf
MWlnyyf6E11kDIuNkifuu4k0SFmGXxgROpPqCzlwFMOy9z/8HZb0r0Pna7NMqz+va1bZgCXdnFTD
BQROKN4Y6Zqa3pPHCJapCEtWnOTUQ2ULjHeng6CtiPBgAMzxGqVbW9QMi8JCLPKYojASsad63om7
aoaWrAH1nK7JlelFP3yKBxwU5VWNqQhoyKg7NKs7xqQ9UqmzEqE46Ek1WOUS/ANG13GYxqwglrvX
uAGMDiztRXxWzDehjAx6v4CkjrNRFZy4B0UjnXL8iqZp4g0TevfmFA8HK0OazIMJFBKHNpJZLt8v
vEL1yQH5qQanQjKaHgsRWVOaY5/NL47b9XntVRWfxKjg2cndgXQ1aABhK2IHEVRlD5vp3grQIljB
zX6Q5niwxPnbLrlOtM+iZF4PvBYKkTSQYM1AecD1vHy5Vhvbvh3j/o8Trix4IMyFHOsNDHNrbRvs
v2jlHbx85BdVc7dIrI3AvWxtZV1aXhTVBhAT0Isrp6xazF3PSwrrP5nUW6rtvU9FaCYeuu41jOMu
B9hA5xmGlsES2qDkeYIy2K8Wo2gCcPx5a9GwkzulwnMZbYFKg9hY2ULLEUShbD0Oakbh6KWjDQKF
kPeuli2AVGQqzVtPqXu/mGP5ESsiS15nsO13d7TwTY5NT9uIxlZRA7MpJalVuRJbb9jf2gcNhQC1
VBFg18/IQTiWDc0bd4lflB8qoYi51us7RkntPzJAJGJLhtTmEhHEO2iSBkHtMfQt72TVKHYnOx8c
FdfiZoHnp/wNwe30RzWABJgxFtkW0c1zilVqhbzTLdvHDwVzG1cs1b5RuhL3qrachGmmt+u+qud5
EZbk+tktV9QvCpTB2KQJkD1wCDVGIHWcPx0KTw+Bvz+pZue4kvwKErVhwVjQ3/dDgz0yX8w+xWC8
HvpzO+lRtmHs0tFuSyBfqP2u7xYmvHvbkHhuR//8jXkinoMldxmXq9ns3WLEhp6mI2iB+On90Wzu
hZRCNTKosv8la7du5JGBdVl/5wl0m/PgCv3+nxlUr1CUuB/r0X0L1PAP6858dNYMiooDoPTQiA3I
c5i+iyhvBeuqY7p3ImSKFTxoWc8sxo+phHv8dawuam0zgCtp88U3LsbHh8Cl93v+XYFsO5Ltp2Oe
ESsD8CP8zLgcB6Y3VwYh4TwLViMDWqT3pKQ/KGUunjyJBV0bmqhVmdpxNYGttgL3vU7Q8IzoYF/v
LEFCyNf/MxiF4lRcKvqkBiI2dOFXIQQMDXHejWtQhhP4DN4iQVyqwYYX/g3DLYwbTFzFcfj7x4Kw
OfdrESqIP4YV7+Z/rqWW0zsoHEkW1cxJa60GDd31If/xVOf7bmylUmk8DlsG2j2yEOoy7lwfHa8K
MYHBX8E0FXSyElR4oG4UHcGFBcRaJ2NbMxnd01l7IUk364PghYYSXRtM3H84POn2zPJnM5j7bIah
cHq037V7Ef5mE9CnIBCZIdsxGwNwG7COj+7XWzm/GEAdKyi7YP652nqsSr/q8Dynvtw4TFSPN1Wu
X69NZseY+lSsO+O1QZyZ7lxea8g+Fnf0Hchp2jRIKUs3wYMfcMhbr4rqxaRlCJHEz4VPp5rJl6A/
vJRHKiiiEpDge3krHB+U/czGwI/+JYG16fyVXqgghS0c9Q6KILtJoJ/0nTyKHHXp5ZLRnvUxY7gS
049Fsdx1RsydjBvLBwXw94gdQwmEJIl1ybBKYnr6D1xftMULP+D1DNJNM8xTGylLs1Q44xHxiINP
PpF3wVri4AAQ6tC4OhOPHXlfBSrDKfIotq4Hg8GLQB4GOOGoAf0VSJZaOTtwumXlN7nqUw6OBm4w
1SNsckvXP7rhJeH1+e1p5CP4oDXTn7EN3rhoYERan5hfHGKyo8KsJ1uZ1WMuIaWnU/Z6rUiGXG7h
XKDUS5e/Trpn4J2gtJLCWPjjXW95F7IQhPiKUjKaTcXtHsmhuhDrZ7fG0Oe+nflHH2rBNedEfZcX
TeFWQu37G4XhQzkkC/kOcG6QRpX4rpLdr15oVwpA5zuetVnqt1cCh7XycGpLEausj0OKW9587ROV
B1mx9RC7+E14Q1+2ZAr0XFTFQKhMwhu8BTmxT+t7jVnOzh3P7Li7B8UpprruAI1JcfyjvbPOApFm
MoViuUpUCo0RLbPHCccJwvnI1XuXelBfpNkI/lPShhITprMNlTJbF4szFpzi4En0mYWETABB01yt
BG6ZBMVAi+Ndvuk4OWyxO2U3MnbTBpMd4ZkZQORakwl0WzF1DjDssplOuxLCzl9GTLTaiRXln7GY
TelBbnpGYJ1z+vJHORVD6NYcDkt5bU1G14+/aQCY4T/hVZ7TUlypTreMuABsY9lUXSRk3cstCil+
dl/7s38HUSC484RU4HR2pX9EdTkUxuOqd5mZp4OCoCOdcTYmSo5XFEwo1i4u2L2h+j4E692Iej5I
GotuOdalD6rZFFm8QwdzXWKn6UW5aqcJrOnqGiNPQByUC2Fv9cecAKjLJMIXlE/1ajpM52Ptacjg
0znGHin87sjhrMOeUSa8lb2HqUK9NQltg0jyrk9AWOypBVnQUr/i961dzp4g27CZ2AKCPyix2Nez
eqFh24MzQyBXHaFr2qAJdrdFaUuoxhnp6XbsWEAK8Yo4HvhBHLSqmQZMiRgHX2PBL362i1lyID1O
+MwG5dRAsdlqL99/Wqy7KD3WvJSM/kBE7d0AoNxL8tqPrcWsK+xdwisGNak5oJ8xcmYWstnuVwrU
S4a6Gh9/M610GnZ3Z73QMyLkyJsl9u1wCO4xZPE0fyh0sUhzuLC6VstoBHu+8iKspipHyb4dAcv7
pMc5C4zLOhE+z1BaSd/7+MAsfElUUPpjgTGYrG1lq97U5RaIgLWT5kb5K12IUN+e7vX94IxQzUCB
DJrBAhX/dRpNO35dp/RcLDr844xvf/16ePjsKZ/fKudDr+SeroEuuXzEVuquqZWbeiv0jy2ifmMk
/S+mja5pG7btnTq3Li8BgimiiGx76gzN2nJdUH7Ev6UReNlQwVVbuo5n9fdfS1E5vU3eZ1dm0sIG
Io4ULxMjhRSrAx+YEBlUYPG5chGFlLlCoxIj655w++tklGDvI7jiUu/2FIBcShPWoPEDojk2Od+r
kR1Hi0DGQAzUuOkx2xyEwIqS2fJOFdwnt1+WA2fbqRPHF1rMu6RTiJ41FBcyGYhPK5YbkaxRI9E6
pAvcpNcrc9epHk5dj13i1mL8zZm+pMtWeEEw2Ai8SIXjHvwgD0HkQMoXGkXDfx4YOXRbMVoSP8aP
KmIgDCCowzQ3jAe16MX3p2m6fQ/n2e/WvLpM2jJ3MScvqqRNbWy4ynyyyggDT5u/MUZ+kZBIpIHE
fNVu3DqhYs1MFrtt+JWKvHpyf7GQOkDYsln1ExmN/eNB+fZVV1vkX5mllvk/hxALwrlRhpcqm4H4
eYmdfaearmIchqeTLNx8CYd9HBES0tNbCe9oRImh82Cb6Pziy8UdlhwhBhC9xBS0nfg/r1vdSinb
FIP/DmTI2ngL1+Rtr3G2BlwhOOSNZVkRQlHCxN+FdTJAUbMXgvdFx/80SdNVmduJy+Q3n7FK6IpB
lixryOfXaLVWRgbpcZLQN3q4RT9suJfGCRGUbko8/dfbdE/GcKaykDTX8SAmyA2i+ws9VBjzJ2iw
7dhejGJoda0pPdkvAV2ypnQgquczSxdR2Ss7bVCw7BW+/+JDPiJkLfeJPMWuygIWGKhGpkYhfbfd
ll67/PQ0k/314+ToekDK5m4pcJ0AztKIYjqBNYSKLvdersVG+j02MlMo6QOPLoshEy7uJSPT4sSG
btO40dMEALU54SkxrRxiDsR7rj5SMRV8mhfGGYbvVlVeq76Jc93OW04tl6oPsTaMc/+wjfkjp4kh
sDBnPHMx8Qmkl47jQINUwSrjcK+rKhHt2IKmw+zXdTNjFDvjM2bCaNTeB4IonbDivA+4koNTVFQc
k93tb/pjMH1e1w9hLsOfWYzuh58rwGMNgyN0ITajKEjfGO34DgUm9nOZ8lNID3r7sfcAcA1Pv1OM
+DZ6su9KpMnChailP2WG0TU7IKVGdcBMQ1o6jwv7ujtGxzxTKdswEpsUcY7MgEqBN6ntxbKkqUAm
gPOd8xFAhCma6SKTjVRrfh+E+h+t7o3JokP53Ig0Cjwj39OzjnatI9lfwzQCWEMm1CTnfabVEXzR
PEXffLz8biS84r0cUeEB52YwSm0owPf1YIozojz10upCTYaoQ+Ogi5ErPHcugV+FtGfR+l4YEWun
H7pxfhBvDLu+4hQIGCISo9k7YkT+zKzZwL/QLfudAmVdQB3YTAva65p8JoM5CLmhkbh8fv7BPgAH
ik7WgbCui1GE5zjRbDjfZn4bNoj1ojznq7+lOiipJA0X1MwiiOjOOHxQDkws+xZsCXWTc0bK9sMc
awMd0xPX2mbnRRFq9w29disJLNj03WxvFCPFnbTMZytGyjVTd/EdhztFGm6Eo+TXG4O3NP71st1I
G4OqIUxEXXakvvV6ftTV3eJSYbZ3EbcdmHNqF0fctxuXG73uMSn+hTl3mofM3c97irKahyBQd/Ul
7KdvrSCmcpNuliFd4fd5aRyf43nLzKrR6K3HyCOL8WMCAf+puL6KNWDVhAlZ3x4Xth0gXOSWgxRL
nuIEA9TM1NiH/GWwpucFYuEM/LpINdnSaBP8THXQmme+bxj/i7xuT3nIUD7BZRPPIonyimWn2QNI
6wyW246g+fqmarbh8BeYbaz3qfHKpKQr4/09m8YS9r/XzBYVMWLUNQlQ7MtJC1ZeMgvBBS3bpfZp
RlK+/20bzLdcVseoKz1wxcRE4+eK5VJFdIMg5BXh4afceagKw7fEmJN14mIR5/nZn80J86wkHfUh
yw7HwH7/TiEDuWcXoOHqTO075JDPmArTn5mgpsIkPmb4iPzA0QaMVAIQb7eX/TdXIHC/69uasqja
T4eVvf49CPZV8K9hr+VMQR6AayAoFcokz7Fi5PcnNUaNJTsrCrBc6VqcZQ31GETiM/vyXh5ZwN0c
aT9T/4nXrJ/n76IN6EqJXe+rTzJSbxftAM3QK4Ino847Cvsifb13t8loPuctei2Fhqa4n8Znr824
b+o5l9MJlzmY1RNLmlP7XB656mCuVFr9QbWHM1U7cmimZ170TQ0e28AmNpyhhO9w3ZBZ+immT4bb
UXgyRELm6hn4V8vLDtU4Wy1/rr+xD+LmPkkWLNKrTclTol2CrjdckZYrNPkhSSi44GC7+OO78TlF
tE/8wsE6xxsM9jfH8MYacaLCFUfzUkWqA2y5/X9F2F2Sv0PcYLADedJtZEiJp29MS+kfZqyJUmcH
LzsHE7J+97qehzx5l0/fGdgPrsen9oYkYRh/mEULFCLsdsl3RVV2S4gYcJB8eqvyCgLesU3K8deJ
lHvaw3lgOJCMSJgXQ6M6T3NMWVgKtw9ah5qXF907SzQpi2qoXAJAB2MSrJ7krU6UjJeY99NeqBHI
rhIafq0r3kObnw8fgETK8QYL0oUr3e6uAs0A+PAAfzWbmKPUNdi5OT+/8tdoCKj+fMr0WerST8ig
jr53PCft8RRwWutQIK8+xv5N4TDHoRDD7mVasIeVPokUYi9if8WSwnr2fAoGlvMXMZSQ5fAnKoQZ
88zrqBbNwLPdbBAfqwtTCCP8WwF4nFaIAP4OS65vhCp/nECaKgYrHwgsSbCF28D0vC3FfABwwlVV
/BoUIG5Q6TmWlHiPB5gQsiZnw+G8slwJePuRtwNJaoUAZ3E5yJeRjOrRaRTAoziaht3moyRT5Na2
fY/+ucp+Hd/+XQTgDWdIvD7oZ7ER3BllrO39mJs0x5xrktOH6yrBQ6qIXvy1VkAQ5evOyR8sBd8i
8fKjEAHCb6On8FQGlJpND8tZjgU3VhhZxX35FOffMnL8zuOqzuw3H75paDhWJhkJA1AaLNq33ekR
xJZ3AEwz6tVweMFIe8ICR3WkB2MwTXVqbfbgAefoDJY1GMNwTjYw/pnSCdzviGtyBfrYmktVA3db
9SjL7tQ7Kr7a5sIGe5mjbVoqp4Qter0e1vvfHOQKUOOjO6HwYjfmTm52wQ/6LC56eJTpbU2rewzm
ao6uI6Lbb1c5jENo9DnxkeRcjbTdEI8/lR+gPQAZ1rmMkpRp6tpLeYpQY4zi3ywSBE1qJfJSw9IP
OpdPsEMNoFJvNLZgH8x6Zl64xr5OZev9RYGDAfnwVw+leCgdT9PqxXxDy9aAJ2RiYo9m2YAu3WGs
0YOaGaDUcDd4cq3WmC5JJXCNWV0dry0fTWEV7UuUQqZyRdo6GACEWCWh0Jb1eU3lMx2Fn96I2dUa
ovSRtePLpE6TlDFEYtqqoWgBGmAsy0w96JzCdn2aKV82jEcEBnMnOvO7JY0aagOh6aXDne0VSL4P
pJkvYLFwzefVol7jAo6DJjTK5jq+BQIU3ZPFLZ1G2IduU3nL2Gbz9NguUtwRnINm4zL9VjUbSgtp
BBZXaS/OD/YzukKBks9SRB+/CJpKCtHElKfnZAazfKMGh9mpJNXQqHfA8W7Em/HmtYmNndlEgfHR
Cxtw76rhXJO7lDNd/5oQKPSwcFAvVm7ESa9X5L0zVAPS2QzmJwcmAC7pLVTsjuNTjtM+F7rwLyUd
oIaRCTdZMIoNsxGzf7WIgxk3m83rxU/FWgCmAJjcJUrFLDIjxl7HtrWnhe5H7glSGkG8jT4M3CSD
Hr+64kv/8khUQkIA9IycDfWuV9X4SBmcs//SpLwGkqEesPHIZBR6JKPN1lTsA2lYoH91HHwvw+Dn
ggTugP/hjEQQ9AqRTe/BThHHoq4Ntc4Qe04bWXjOYg6X080D/KP20RSbqeMVHq9IQ5TYpJSkSi3f
ThnITWY/4Ayw6c1Y1ENJFtmA0ZuLVmcMl/WZGVuT16/+7153OUebAK1z0umst4Ozk/lq2HG9k8Is
vM7Jb41ALtBnz+OvsVNceTEl8dtJjJmg0syY4oDM8Uu2JrNBe1YQ2Brj5z/cGaHwYbK0TjG2b2b+
w6jhexNa6/p4OS5Apo2/8S1gCUg0iGXvW7a+MS4+63l/9ssJErSrOT3kGycOV3inON3uLVw7rJdw
taGO3t5wE78x4sgbIj0apr4rqljDMOML1qgunwD2hPXViXGvg1+De+kJ6ytXe3TDYH2IJLvpdWZD
ygfa/Xg/n0hGmb0iKvqmWq0aekNbmPs53Ow1f7VlJCr7w7HPLD4DsiJ/+gyhMFRc5fIEJdjKpND/
aQ0CHbQ10jciehR9qhg6/yPA6sCULCcfOsSjZxKr1cRP4kjq+Wgi+WjpfG84nfrLOJzF2vxsAKFg
Q8rOml9I1dm/TvhPpA2C7D4mAYQpMelSg9EHQ2+n3XNimuLStCmPO1w86k3lXGYgEhGTQY/XpiM4
9cTjvO1CsFWTM6tx4nrwvrLmaBRBL+iRSpTeovjvP4ncSn/BL+sLzfGjOE+TWb+h5bN5ZAcHdVTk
17EGvYaYX+dqFuOXCz5fZK7MjxGMLg5LbbmGMNmDsDZ/zpb0SnhYpY2jJqahMta38SuXyj+3WR4C
J7YU2XlV032xPrzOK+hzwaI9iSnsMAZbKzzvzqo1FKTxBHjR/qN3ASIVnMQBeISBkLF/a1PYMODc
aXJW+03AeYio8ld+TKh+aVJggSRs1wRcrLpKEJA7VVGSmoxiecU8W7Ziu9YcK2HgclW6/gxOkxGQ
P8res4QI0tU+5lpILfOH+I7fm+eE1Ha2vvjzaBT2MPmb7DXQ5QBcR2mi02p28dBOLlRP8er4xTjT
qBb7Ix7J/wWYJxY7/yvLheGC/ikl1RHik4DUHChv7YwF6+HGzU+zDhwT7tTY62wGr/JwGjbqsKzR
O6m0mX8tByCuY6V1HFdY6EjIdubwgMQmFvDSndRcR26lNcpDWa8iz+BFCcdzQYnnSirp8oJs9Ef2
LvN4a2NAn3ev+R4aE+Rj6+rXLvyNKyBSbTpSj03R0SII6NxG2LD/kwt2n55+4/Uf3am0Nf/XqyXt
70eDrv+Cizdiw0UN4bluTKtMwMXNvGAWkIphzeds009kl7tT0p+o8qHMBlHZCAmd+uR3Y4cBXZKp
+OixCzUCt3EHJTmTMILvGo5KzMoxY9HcDR9D85iqV+RycrXltEtJM2Yp1WjpymNq5VoefMlyzG3a
Hu/u9OsP5pqX2zbeJppNtTx9dZKi2qixRKWNfv9KvR7vjCA7ZKWeKJsAECrIYHFsKHIbqNfSuDYY
dMpwRYrFexVmisvxrgrF/j8atdPJ2/yGIyCCF7tK8KU3hGfYEdubbtOwYDSFxM47ErAK0WWm1mcL
qaCi7A/U/ca4r4PIPj2Gr+DWGc+4HmWv5mo+V9xFAJRnonL5NWILQFQzf4XBKBT8wcJ/WC0Z7fdl
JhTYX1W7FzMNFM4XPL6la3Qcna0MUxyKhKjkPas7uVtcKOzL/+AFLrWBENGdHFS1rfwvurBib4AH
YfgcAjSBHmFjfsyrPiB/0hftg/QTYkyYLENJX0wFowmHy+11jhQQi5Am+mXqO+Fo1ln+gAfM0fbs
09/ZBeXO87Gf/+uLjfIU86Fan5BWslfQpPSkLbGcpVse67ruWvzU2VM27PWN3WfhmvTTkIVzOwPt
VR2jS8aN0nbkG+gVVZzG0IOxCgwj5jRCudozdWE925OiHNUF4dwrQz3o7j9gGQgoAzbYRr9zqJao
IJl7loditPHWReQNBXjzjmNF+CLuiQzh+UMvtUBspjWYpdUepdIDUoXiGMqYD47ZWQJGfKeo1VTn
yyW1xmC4GsEu7WzsLXQGIujQxNSLAZAXdYPqOCq4D7yolHvMcFrYlyLShCWCY7rwYpCO4H7XevNA
4plAoJSaivSE0znsSnN8azki+jK90MCO5ToM2KVvwaubxhSV+EZ9qJoKeNOvDVSGF+k5MA0IP9VH
BRHcKDCQ5MrhSEaYveDZOUTtM9v5tVXGEmVX28SdyTPoZfWu3jhK557Y89IBAW1zA6V8h4+Iw2Jj
XpJbhHAiPyUI1VAqvfXwxcMOWzrlSKUDgu9AWNL/a3fGWO2AjfZD+ZWnbv+sehH3aDxEBmfyrijZ
Vz10kFMYHNihc1A/nlqNO6Sob6TpO2/g8myfp9ZCo93jrCDUDob62r+h3t5MiKUC0xPtcai5fOjy
MP9l4MQBRXvS8OgjsV3B07mmBCV18t7qxdvJ9uX+z7RpkJ/TJ5Bo/eEAYXLqB8TeLy21jH1oSHJ7
2kB6ZSg8CVpodmTilr/O5Ly6T+WczZjdfLOBe3g2gwHtN8SENltpnnP4Twa36QGSdMlyi6OcVm9L
M6Q7TC9yuPu7MODgw7yt7SKhg3oHXv2s6LHTjHPxgS35Xu60OB0RM4nwoWiCZ+LKo3Ux8XVghzOj
vmkeL+uytuoc9mg2vXTLthi0V8T6UD8fefokaVey0UNf1AYMn5kHII3PymPbtg3LAsfCRNd1HgTg
7O+fktssVxVHgL9ljLHPoQI6DV8HksIXOk8GEA/LRj6aW0ixwIKcDmYACxTJ1sOPg3AuNjN3O963
fYN/cUYu1FJdVAT1Ah+QXTAa9QH9dwm5v/jHv9hA1O6JkOROYw4vQ/mCxzJbMCxlEJDzK03jsQiX
b8Pa8aLPKXSFpEZEbdUK+eyBjKMxD1W0epmpS2IzCWpB7+0wLWtYNFIIMR/CcbhwSIEOhA5IhidE
EHJ4J9/HPi6JBAuxhutNEP5J+/KXDjnZ1xsY5LINmVecukXywO3QyI7KA2Ps5fpLxgOI/wt+Mz0M
A8LO5kpcNydxxOCWEdIKfQ+P59wFnVXSRjR142IDzfpfASffbTKzh0kZa9+iHscE/doidRszDeDf
hcwHd7MzRazDuIg/Lb5N6qQSproKjCofst2BELypeBU/rC0oitH5X46DY/mArcQIpJ2eKGTbCtyT
nA7qlcFLmmRGeS0FypFvr6zPMvpiLXq2v1pKOcPEZub7+6ndi1Y7XA1k9V26yWLaNIqB6MtUKPeT
tXNzDOpfryJDSoRbSowr4tYkVj8mC2xQpFb68InXe+0CeR9DkBjBz1h0wEQ3x4mGmPUx+9nMm5JR
G4uXJ7I5PrjVoSKHlDS2NPBawdoR5/hd9B2vMGuu2TjMuEF/3E2Z0LxhHR49f7PUu5UJQMwuN+O4
UhARhWWY01iyGqxOWYR4dCVsSuQYd9YkG3fMuxnG+pFo6q3AycquoEHFc1sVRPzqpFAgASUhdncC
IeQybju86+XB7ZucN9vMITH3alPxbxuaiXWA07wOsZthp+4pxYqT4KwTWl4x2zWxrzIvWmbTmJTe
hYZWXBetoYzWXo8OLOOn4I5TSw+LEvhVdMFdbv1CWIObmEb9D2kCI2Ht235uZMz8ZUWTbY7MMpZP
b1lxaNyzyrHUD2nRtHWvFGXopvavFErps51URcCdVy5g9SO2bdqjtVtlxO1zEz1UHVcVeS1Lbb71
wehI95FZPnh5VvJCK1soz4rwycifxYaa2Om9y8KGpPjk16oqrGD/nd69fS6O0Hm9oPxx8jtZKLbD
/4CGL3XtLNW9LDqbiKHsJLyQpJnoWf5NdAq85aetKLLzbS8g7WAVbdNY6EI02dSfx499xPVBn65Y
ZZZtHXf2qhsZCcw6rv9kyP5JKonW72FhSwgc459PN+Sx8qtWh4VCPqCvnXix4vp3eWe7Jt+C81I3
tpmAdmMETnd+8fsm9wrUzVj0LjOcN8cuyI5dmEVDHHGKkKy2oQymWfuKl4JhNheNY6txEmEm8h/x
rQziO7KgZ+Ldh6tStKy4vjtInu3l4Ws0rEW2yRGzJlOdANVE9epdpool6uhLJedHEcd7cOBE5YaT
tPBFy3tvHOR0PzQDqOt+0Q9xRsXdrYTmq6esFpH4VshzHBFngs31ooNLPnGtiuyxsJWxdLJgH9au
UXf27gTwivLGcKAd+a4xQrY6hddAyC9Rpr9fykcGqKiHJZv41x3knDV9NTyFBMGUMt+1UUVtvXRy
n/6CN3NReRZoIUIpXgkbkADZFqhYZ1k//e4iubdrh8rCd4OEuMMH9JUFstPeLbPxCaALmvSKvPXF
eSR32USeVGqh2KYPlhDYCtIhR6Q9f/tLk1XUXjLK6XolAE8om+XqHnTbXrr9mzFJRaJ88dCn1fiH
W2O32oVT6LA2stbVHZMCn9B0TxraI20L/7P3U7EtO6Kz+A6eW/O+3XU/C/xWzjv41+1/tn/xIXfF
mA8ea88ZtsVwa7LESjpnsllnGuao6ERQTPcp5p3BBUENKIDKFwvAhrUOo0+H2F6SooYv7JRl9g8Q
kIhfc4iB9KS7pJ0R03oj/hwUEOWyAYma65gieCjmT9TGkHmo4pRCFja4nry7L2I4otnj9LVVD9zZ
Mcoq7nqAysY5KybX3AIfq00qjgBxn6/zOsusGZPrHcea4xBG8KLR8EW8vStqy5k2ox/osPIuXUiA
yVMXX1T91dwdCKDp0LeqlCPaMWYWjL30DGXeNxv/W4doWOrDjuusiWZTDQsjvnPobik5BxgzDf0p
U+qYwlrsRJnl8CiPnGBqyQ0Kr7RdPIqyd4M4Wx1OXa8StD1q18IqumX7vaWiiwvqksqhNwV53Gg2
3cyGFW19AlLqBm8uZrHawG4NaAYUq6iY2SOFAVd+OAjbvmuCgcF/NM+NKJGbwu89JD7wYWOhm1q2
3uwgfeOvwPRabAvEbUsuq68/Jm+5H2/YHKCL7HrhSV9t25fJdb004rx6WklnApUKqzWg6Low/lmY
aX0lCSfngYwflYxphSWdL7Cv3kiFrcXTNCozodjTY+tBEPve468jK5KfBcrOutBiDhBwm3Z0XLgB
jlDqg01LZecn0PvDnpewc+A2JLBgdkPNVB6AAuhGw/w0k2Ci2rnDOL2v7aBUF+Z7CF8LxHUULb1+
sAB1V/kDhMWbEi9l+mLaw3NzWVxiIZL/7u3L4SltFudN3/vFAt3mQzTthe0fiScx8Pvw4wkq1ax/
lQ3Sj7x5OOBCGq9spHSRolDcpMxP9yT4tVwa86A8J0h9LgGNarp9/s557j1notg4QK1yt1Uv6nOO
wMWAF8LGmNx156jlcZaaHAgAY1+zx9wG66p+9cBOv6oupVj28Ch6Acpnq2zAAhEyxc+Zl/ye8tYX
dedoySJjSTjQ8IsW2ONHjLfayQ33KX9eVpqvfs5/YwThR6D/eY5xkzMZPzQQEyMHqIA0lemAu0Wm
VeEZXlHpJgLSfW8Mym+N40NFgKzFM5WvByCsj/i4e1L+bzcdy2iTCPJGd0GxGCNK97OALQ86XzgH
oe3Qitx829sT1kWTFyXxyc2g53gD3YocCzWUcSS2vu+pb4C61sECezq6k6tVzSAacHFIwv0+Hry4
250ZmW4YLRUZSgDvQ4tS9UjeRI+CSy1vaGjmUyUutohtV7Q99WgtrHLj+wse9gQGcWF4zeHJRm4K
nTMK0e7s0ZNopT9gamrrFaLZJApL2wYON3ED+6/TE9zv1lVNowDujBW17QlOVI7pE0V82YjUMIiX
oV7lt7OZ9ZTNwgpUFbof3GCrrtdPIHLR1PNrfQKjtHgASh9Bs25gIrxCYceRBui+DOvhI10zZYgW
hg1yCpnIO9Yy/tm5icZiF2pCNLZ535wKAMKaFJ90/kDLxzYdNJLrFOCR2ekQLOYLWo5S3fYJkcD1
T/LZpnnV5Plmc6u3zGEtC8TYpgL0W+J3q+s6kBGc7E9u2uXkb1/ksGmUpgbzI48UnGG7DgmtfmkS
9rnb6zh7VmeV3+KIDs9iizhs1gI07ZNSRwnc1Ogb0amxVS8LvT3HRNjlmPTuvWBz9QOhN4vAVdei
9HY9L+Tv+PRx0gIuIQTHwP5o8kBKX36Pos2YKnpZaFw5froLaijm+/OB+hybxQ8uhY3uFyJG+qC4
X3jOHi9SQju97lsfBENiSD13WrXqM7qW4fsnSebQCFEP+3xhMaoFWWIRCpbNz3zD1tHyN54/dzPh
dNM2Upz5CZ3YrjRzIIEhw758tfBhgMYCE35asEaWULdNDFnHwfPEjf14SBLS8/hU/NUYZ/5Ipt8X
9AkS0Ft43AT++cp+dCewRWjo7U9N49WuVPuBGFY53bQyPmboGJxH7kOsojRGQd+bfH49PhyZIL8/
y7cwF/c6Dk5NUTGlVa83aiY7ipdG1vu/iuecnTquEWCFEF4u2DPkXthK/NJkp+CQCg6sJkebY4WA
ZMTqOJw9uQoyOav3MqvpbghB16ZBhPLrK4EkDxJT+0xKPZyjTjvy/n/sa4DrKajqpgnLXYsKxCHf
0cx0XHlsn6FVCFS5y+xbYPMw5X8jFY4vaqhCE4J3d3n336s3xxOQ5ovhFMeieeJUeLGsVyBpwbcz
2bta4PUOgGOPjGx5trAkOCicu12IyoO76dJJYSc6kb3CxUyWXmZFPozWhujZ0ukzOtSqf9YIzNfT
7mXfUxtA5CojYSVAjrY4JacDDc79UdeyUOX1MDmXmxxLNMwXEw6eSBVceasnsC+3PK7N2vh5ge+N
87ffEjLwkeHWP7bpHXS/JYmjW6r4VYoSne2Pbj8odMwkPY5aq9ICaAk3zR3SnJBaA2nn2LqIE80g
hUydfGpKb/y3Vx1jRYJtZXUx5MmIl94Kce2sdq9GU1c9OExI/1EppVhkpkw2OZxXWzZghdTuEF38
PKCubLS4oDJzHajvXQiL74J+ZHd0zk8V3kZYOs3hetEAihiort2eUUdOUwZoLC/QQTv7NWOzBbLU
fep2rXS88F47p9S1q8KL4/Njn0wapbRT+TGJvpXSHsn+LIYoYo+yyAUb1rB2pDpnwVKt3f7SB6ib
/OhECcc6AxVWTssNg+2BclR+8BxlrUtiH8q+uYiWZH4BLiDpBRUV0f2cJui2ZQeuV1q9sTyRtvAe
GwSQe3ggPqXW4PRsk68R4pqaiA4CGj2qt2vPP7DFgi8AnCokoaGTzj9T+iJ9/NgT1OHvrgbAAs7D
ZyZrgQ0CZqv1/1fnFCeCcIFM1fPYpEZ1I2eIx3/2Xk+SKKcceBaPBbgfoVmm9W8E8ojx5zTWbs3D
s5YvIKw5zV4lilTLJTxZaYQn8gn//W6Flk7F+MInk6Ch3aXz4/2UiTtUa58CSKIFwtLxqaWrF9vb
NfKTUDfT+aIYBTtg1eWSIAw2QrRfKWMYQCOqGRejMhgoReP8R+JR+4DriQjC0s5UcFbcY6f1LnL4
JCHQNSAYqiU8bELnAgnjBc/8aiaC6BPVaZ0A0mZOPE/RPzw4SlrUJAr0aZc/g9JYrOh5PrQtrAeY
muKihTBQtLErDsPRk+VF/Rhe6ly275jQnlI7v2nNijWWxMDpOXyNjZDfNfOu6CxAK3jrV+BLNyby
/fxNw05DYi/M1pvnNfM4B2a7/OV/yFveVd+T85SnisAMPUDSxeYjsNpua7BbnaLHMcRh92IMCiLr
lvNnTw1R+CUkb5NrAoNy+MxZ649NnrfemBxZ3BXOjJk7Rqb3RkHk6McgNmM3kBcLFyjYnHDPzFVU
W3eUfqmUinOzbTjHLEoSMLFpgX+eOEeSMTSRJGGNMUXwQoSDAF9TJh/GM7N9+JAfXq+w5DTCDH3g
HMbLNJtbBduaPYD/laAhbES4QI9+v7WsKqahRAnR4HqYaQLpWl/iiGEyCKHhoqCTHLBo6kayvsW8
dRjgNphgmObhGegvQm8APjqag3V7+4UWg7yjWng4CJhksjuG0vmEqgjpTo8jDg9qnmwxdNRB+q34
+d1XtCvwJu1FU9UoNTv2K5UTVWIGLl3BRHDCyqv9fJixis0FKOWIrLo5D8+mkem252Tjl2P6IYVI
RzMGiFsNLhXk2ShAhkigM9SdCl4JAEXvma/rXjbMuhUWwrZOH2fs+F/eRn0yNL6Un7qqy7T3MxO2
ljYyt4a24F1YnUGY5Tv70j7wAAm4LFOTXYO2M7AfpFgco3U5NdKa5UL7s0VnvYmAyTZtqnTNJobU
bX0tRh0VAtz9/z1wQ8CsrRTGxOa9bhPE/cFMqzRUD8ohrk7eFzMZKBMPLsJT6PAEuFrGNn4v8AZ9
nTChVTzg7DQj/NLbk34jrxBDH449QOYeUjhP9OIU8X1eMtD3VB/1/6dFWdmE78SQx12VFwrtX8e0
uqLzgMYujoD4VDlXtT6L+xdprnTfRBi+W6DayHiLqMc9KUeSWOcv5fkSUDv7WcSs+Dy6rQ94m1du
iKwOIWWWakZr/8YHCLuCFvKrgWUfXlyoddwok73q3t1UZIVhZWZKmT8oo5p4wpuVNsN8AN1W3CQ+
TOlYCK9BW80ibr9yWQwAWNxbUvFEsk3mhv1YA+1sIiYechSWQPPgN8FOrE2T4kMz5MXyMjzxWl3X
YZGXhYKG8UTxa1OoXCdp+Hjs1an823uXAKSdFJgNTxFm1doZhrHFcfzMWbw3JZPe8MY613dphBfJ
pahC8KwOoW5WXkhWBx0MiIcOElTH9surz5Xb3uDAvjxiYj3DKyigxeGN71HG8nd60C8FvqDDVig2
o4BiZ+AtR+0/w0sYi+8iO8B5WAgzUprSEpXMVQYB5AMfDSOtkC76RxVu4AR0St/GMFIzxbGmeUNn
5uCEuZ8igBTwOpdVTulA1CaQVYxKH76wZKbADZW4RSHlFRJ1VhyFVsqlHbSKwgwD+V+30vWNHIB8
Fzd8LcP8WSAoGT1XknvciPFRTn0WNsRBJs04ZZ69XIyWl78rOIjfCxiAMYR8EvaPnhGZ3F3j+mvj
f0sLuRURD2Xfa50qNx51jEfzQejrAQaBVUmndvCsU94uoKkPyk29lZqDO+lNsq/r89Fx6lXrI3Fg
QXJr7SYeC9GsBen6iXTYuI4P3l6A/n6rDyftw5qdb2p4DQgpGMR+olljQmKlvY5vP1aeXbbbbDrl
CAI2osv62oxm42Sha4Net+5zKJnFZvuHzEiGSWDg06P2h1xUJDqIji04YQtqqSGB/LERhCsanEkY
sr1ba4BsQTQspFVc8DLeuSa8gmpAxNEecAchDXmkSbrziWW5/+kYfxSPHEs0kNhfb3HoKBepKMJM
0kDnzRfC2NG2EvyNtbS/kiwXN+wCfA62PSLjrq5ohWMpIrh/7K6Uh30fw/2WsoD8DMmxHze8jRAA
itwTiAZV1s6jULs2cG9PmUa3nQs2lfC2mVTf2QMGSGXe3UMGftQYug+iHIpBp4HHwKGa1WoOZc0U
Iz94UJ+aD/6Rdbvjd4tyxXKLgtAzjrXh5srjal/x+zLW9CQJWAqq3/SOv41SW57dTWqYfzD5kQZy
3u8RefDTOyFdpiX1bG8TBhhtjZGjAoZUZAWkmo+OZUpHpVjUkKePQOJhUG9L4NrAWihxTRtzZKB6
5JiC1YEh5H9l1HJJZvKJRK6jFmKF4odGpBUROZ5Znp2/77ZZ+zCsUh36vufYOLQ8Q3WPJ8I5cKXW
DvzKKN6ILw97fl1WXVS7mcI0GT7horUYS4CItX40vGBMKIXI+eGfO+jPwVy8Y/iDeOsc4RThU/ja
SjbBy88SILzKdrpV+H9bMpc9Sp0+59XlkiNx6WkZt1cXwA7WYQIb+PUIKFKIVSosSx8vd533w+Fj
CPsDXqp8eaXt23qr+mAcS/QKyaT/OEEl1H62j881jBadyPQwMAcjXwru/JtuNQmAILBtuWQyhXqL
4bTqJbtWqc13l68Mf+ZQSjPRT/3KzLQiE+ZLAuVr5epF2eExKZvEVzzeAe8/AjctOW3k1lTqljML
kRe4YFt9VQsHTglwtf+dxIzFAmlpjqkRFyjfX/VQCgZMcAYqLtdiov7S/KKDZsiw8A1OxaPqX+DO
QZhBhDFNksSWDkPmcV2VZfD6ZOZDQrG057hWM5rb92BFFUVhWlpeV/yQOQqTdFdiREyqeT2AQGT5
KQkWh0dpadB3PEVUiNU9Pj+XkBXHeKOFQZuoaaR0FpTwK1jmbKdkUh+EZWVodEXn524LZzKIOJu0
wUxrjDKC/cBl9LKSwiUhuhUjncnx2cBFuMKfrnBo7L1gNU7PRYP33E2SPgNPlmGaB+yzblF70LvD
2kdv+iHZGzsb4LzPqW0jxmY5C14fvbZvLKDZzIRYCcScsJB4T23ItMUBtps3mTn/7WTNVj+zttA0
se4wPwYUD6qQIlRXMHnQDk5ZlNGHG74+Ttdf1r9l32gqXbM1oj3sYoBxmZzHmWPfSIJu4ZWk2vSf
nyjpRJpxTiE41Ijmm7Ooh3fnXZhF6YQ88pH1qbMqCLesXvCXmgYrPKWPuMxqA4W17m7EJoyqR1cH
+/5fhbTcharf0HLNKi2O+/xCtWGJN/wKKTLlx3PrJxYxFcUinbAE1o3tYQAnsTwASQu7fzgDJiTN
AsZWzwgknc4N0m1+6pmcFrLR3Yadc57QZO9vEQ2TrJJalS5T8ICEgrgTE7tZTbY81sT5LelpckKJ
WwKILu4GhKdLuPrsZKExCgYMGD1QCFz0uC0+oY6ts8YafFbvrjCR0OYmwNMnGiTAdUnaf1hWJffs
V3xl/c7GDD35uipQpO8YFxEkjJuTU0cd/7sW1hgLDkdNXL2mvl/RZnyGG7D6YwcyxzJJe11V3w9a
DiKlfDOzlHE++Fh57KO/WSRCr0ZvYEJzH4idjVwpVcGEy7bmpUsQLjxRjPpSo7d5EZmKaqv2zDcz
BoWwLAS6ukG3xregEoHFWhzRjw4frK25gUt3/5Xp2ohE3p+g96TEDsoNVoS0Q9LH/FFS6QQNtvfk
7eKGHpLIzAc26KekumL8tdQp4JUmvyB1VZcL8MkRsCVaGG1/egcLlF5sG5MGLcgcNOs97GJSxqge
Dnq7DrDo4q+sdB6iUV8umBMZ5iJ3S63tXJwKup8o5eY3+uHeFjHF1OB7s65nTQIiCw84XoqFFo8y
cfGPHTQMzsOpmr4J6Csr5u6ygHUTHhNEqqNh16tB9+GsJ5tzwwemVcon7PNIji2J7JkkC7ihiBTm
MhsnNm9q/Ijr/PfNpEt9weQ4L9MiFomLvhmg1IdpRz2PjGf/00md8yMVPLKxY7CVqebSxux9DkME
jLWgpm8sNQXESHYpF5ZUQ75TmuDFkvau99Tb2JgZ4CxfyBAtkvpjxGHsABSiK4TiSHYOyjueqxp/
zk4IsBS1sz9dC53UMtNn5d546T4Tj0pZuRYh+HQ6rHGr6SesDmhg55Qp06R5rX0dmdnAI7vZjNfu
CTWuWy32ZiAJNFajYuOTD8M66VfnWiP3eo0gGpKPXVNZkoZOZ8lvFV9ArsAmFsbpOUqKMRewGDH+
1pquPxWbDqTYswZ3biSYXW88i72+OMti/aFQaii6ONMDnXM6VFgJTNDgQYWbCTF1GVTcnadq7L6+
dJHz1QuVnv2x0EMYatfc9JzWJddTv+TmkU9kTZm1wb7paeSoTIrGhhk8pxMvqmxhQiT4WNSxn307
JSKnyxe6LqeEwLBUKTdaefFZpgYiRhm0LCUM/UOkN+eJXItTcHswfAMlbMECjG+bq5B9xcALgbKx
K5O7zcVAd8i0U2KTikMsciiKAHz4moN1F05clNdaNLYgZJrN4yD2GP8EICndY9e5pOiihlFn0LFc
S4bLiQIbY60A4l1h//GQnY2xLVsttECitjYGNibveMPzYbu8H5e+O3fXug7rp51SxlWocEPvo4mW
AGJC1kQrpCVyKKqI1zNY0+s5hoXFAW3xbdbKAipjTbbVlCAK+qAvvA9pqkdOT7vnaboK4Vji+xaz
8BsLqSo9IMvTtcuKDkvLeZRdxjF8p7S62bXCtcvORYsyG04xjuF5J7uAOG1YQsUsDyDyn6G3eST8
ZJy+r5sySC/FCDBI0ai6hLlhgu99lIWFbhT3QRW1s6CL/1kSO0Pz+dvSA0Fc5Hj+fPOlGkw5Z2eK
T2DeLE5UkYnuxKJlF95SDLhgZKwQU71cK/C/8YtUYLyWwl+dneKFuDtAp4bieh+j4SJBGzF8l3KC
e1cGhBuqeWNsz1D6jJoRzVJ/CgPPplwAfqACaJkNKg0EERhzKNxKCR1rXqqjPH/xjIcUWUnh1gb7
M4cKrLM9Z5KFozJ8EkRJ9I1BdgBcm2Il1P7xpYCs5HE3gMYJtbzDnaNOVtsPPLcf+PvgIeKrEvrZ
aPORrQmmV1K3nsJYFsEZOYKVb4XNFgUdsPyWQv1nYb5qg4LN+uxzumx3+4g0qb0Vy+87MMcHqaOL
Gjd+FBs2XHNVx7uDB9ODf4FVE+yWnUEjsVzZz+SQ3QWI+kYgXLeCX3SYmNiiVQ5SZh9UhECx4YkY
ltGlP9r8xjGcVquxYpsZ1QMN3GZ8DCFeKPTuvZSUMQ5r6anEtrKzT14bAj5Jz3LbAHiI5dSqlvdy
5BSQuFSKL3LdWQMZmYaLX125Un9gdPc+03Br/qZtLjejcyb6DywHqjUqkVONgwZt1fSYYT+eTAzH
BGp1oy93YAAXdzv1XhItlnWfb3KELgtmj70pfD5CKCUTI8+OeFYcANV1ANUghQixcv/raypAX+tm
cpZSpbOcgwgnD+Elri/LMFCStwv/LoNq8PpCRvyhRvOnwk6Id0CHFYTV2X9f5RUOf1Y9QoHwaQZe
9qOT3py39qKgGNGoHg/PoymIgEKIDVryE0Fxm25DooGRYcYb6gcZy8Wgkyzqy+U57mZIVnfEnZSD
Y9VeCujcXCAaXh7jrqDpdC4LFZ4D+NnwvlF+GEmAHwtcbmrlxB8K+JsZyNiHoxQQU/e1KavNHqdX
4zudhABOsPTLad5832hlZSRz98m/hXmjromqNppna5fyp2vr1o6xLJmuBK5Pnej7gx2amvcFp23a
HH1SktD5oYVHbDjYwpFGGnEdPmmLkigOdKmbWP7ajJxl+2EbkV1U1a6JuIo+zp/US25Nk1pKvvjQ
Q0iqc9nViY7ZoiTbSsohx6pUo5jXL5RuackkFSb4GGE3JJ1uxqPgty00fvyDrX3vUVD3ReVdcX8c
+Xv8atAwQFXkHt60sJPVAVlYZS6ylb6MGV74FlVgqFlv9+qcP4d4PK3K6fqhXyPruB/6CCHzt2tR
7HkmzhuL3vslvxxKbmCfvkzQelDS8CyCbkgZ5cqkzJ/FxKJJh2zTT7CVbjEcmgcHqlu2t38ReYMR
jHho4b+DFGOKijANQQ7MufFnN2Bt0btIHIqrtTlkHRwn1ySpyL0bXbjRYYtzTXbPC2ladUisINvW
v5etptMpt4hslRmiNyUXeS36LrrgP2CJ9STeitel6K9FHJKHToXsYNFD60NQJYWYxB8PXbr3rHqJ
p6JvNBGt72AfMPXhcIhSQQtEYdBaffCKHVvNZ2sqwF3QKGx0OXVjO6iKsacOj51j7rSIHzJw4X/G
fB9EXaaWya17I4GIm/aELZuk4e3tbVRjKb5c4DIcE/nWLPhq/vgEnRvoEb/H1BF57KBbdJOmEgJe
c4GkUbiwEN0TUp273JNvXfTvShzqgDt1q1RJQBqM8LvFBVbxQk4QInAACBvCdHGmWkJrNgVlq1DG
tak7gKIS8G1LWAOULXddqSfeXjqQLyq/44bn4yyxV1lNkqqO2cVWNqdGacDyScx0i+QvPrwsmw8v
HxO7Djzk50Sh74WDqVXI58kDTGgAS+CwbOJu0PJRYQamHxaEc93+q2PAGWeftpR+VdK89GsnpoLT
2kJBplZkdl0kSZV8awu8rDeAeJ8Xrxw5q36Vc61PZAkD+cA/mj0dGlPyNRn3RFfysUdjeSUeZ7yk
lhuIzhrDOWcXvuQMAsYIR+oDdg6bDxttbo/UnfKKFwV89tToWzgvQTjKxQIt98mu3kw7xC3Cm+jO
ICQx0EbbgDeT2oPu52KyddGtJd6AvhDzECq9E2v6xaeGLOEGm0ur3+WYn/t0wTB8AJ5DtMdbLGED
WQ3a7l6w+JuRqZc5ofIDycaCGqjunmXo3QBjU7w/DKDdw4pDg3Uc0PYil2OczOsNtOz62QMleIMm
IwQeIaLgdsTN1mPV7lTEOYylquKrlZvns187fJyit0J4HR5I2aDK++3nYhB5sdNTJiutImJmYikV
+VDU5ne3aWyzLjz56dCG1hvlG6z0XxLcJc570V3Gt6VLEiJoYOJtkD7222IveIrdnFSZWd4jlw9x
DGxgqT+DfjEFTJzhQj+PW4TF1qkubrCgtNSFW4fgxI+4qb5+HSfrUIm+toGnTtGL9XUe3CNf2/z5
GolbvRKOQW/ZVHGdHZOsQ31ISQf1frvjMzT5MhECSFqVOpBMLAVmqHfrUwt6HINM0hpEf8Ku+Ue3
1QHBypeTiHYxdOrbbk63W27YPra8oe23n9lJLvQQgbB3bWLCxESYHLgYRhDf6S5IF1QW2yJZnb/t
flrHO7rQHiSVI10MGLZXgdqIrxVgJxfEeQe0T1KFs5yzQtfdgRbfBGoIs3mj2vbV6cfklQ0mst0J
WqHYW93OtfqsZ4hCFtjnW7itrcOlhATh9znHJUCegu8Jlk8FKVNSpLP4UgMgIO5p1xsiNQxRTXc6
bLs2J8UoRx7c17MZIdhV8lBGC1o6Vm8V5S+0VuVFrow1mfaXLJnYEl9WNTuj5gDF1ouSNyIfkWzO
F2InoCraj34UG6iimIHbRwKwz4O4W/SUZ97RRSXDMn9j3MLBtLNvo3ljNwj6/l0QYAbILoAYQGk+
CJoDJrPEGf/lwYkTkg0o1+eQRGyKXaqtY2IqYQAsFs5mwkm8PPgSnnyyK5LY/y1v7Cl3PIS813W4
5GPuODtAHOGUFo0ZAblptRAebfk98poOJXk+1dqd31PNth2GWmhv89VkH9NU94wUwL5Nxkm6AFUw
xjlQS2lPhRIhksCM+JIc+lfAxZ+O2dth7QPDgGDpV7o44ZIqz00yMMnTeVMD7wHy0KktiLJMJCcJ
5RxUNsHPP1qyuw/LmVulAGfraa7oGW/mlAzjT78Us2F4d9I6/AVf1wIcRlmzmgRAQL/xSN4b90M5
9L839VjjZpAIkVCReY+A4ctIqvMBUUZJIBP5e+0rP+PxhsCyWaR1Q1/3DCzKTXxZIdFbT95u1nhu
m9dndDVuLA94uUkvDD0pdQp7r+EkAMKDI9ApC6CN7S/nGOmBBTNEqsGMXfWUiKTfUlSryxHFdy43
xjxmpTzpBuV2slnh59ZqcPr6KGb06zk7bFc54KPVrUv8ULy9N4WMRPhNfRs1O6aomXIvCf0n1DGV
1qvY775MpvcvOJqI2qqX5dKJHoab/cKlUb/rbzVaOSvtBy2YBgkytLlUOUoqFFWtLqE5zMFBcOL2
cLtoiMbhhEfg/rE6ckxdcNS/GlYAuAQT63NiHCx65i9NtCaYwnb3gqadsHR1DtbFiTWSIZDCX820
cMzJ3Zndp4eE6yxDiBHbOByM6NCU+mNIKdH34C8pArIcIkLBbeTY+XSgjfqt7V9t16Hh5dQdaOcl
FQoiDO11z0iz3nRrKC0mkYLj8N+dzrLLK2vJUCjNQB1d/roN3pcV7C2FA12eZZR3QCnybw3l9jYT
nBBF8VZFPAZ3wAIbl6PIsLdrD2rTg5a+OLmW+9VPegnSOLiafiQCO5SjnCUtwPwcBL9cq064h0zS
02I6KG02XSZpqLvMoAZKIcZ0lzPClz9C8zRLDjjxhZuLdiy/FAakdVXUzhPmRAl3P6xjNVkCi83f
RhvLQCFNLlPCKFAYYUK0mKRuNvU+1vWEZoOk1X3tmRKfsZdW2FbK8zEwM0Z5qKBnpX0A1FLHVb+c
vA1s5qRI6CV5JUw4VaaNRhz7nQflgawuNiDU3CmCUn+OpbXs2hZK+KK4sEj8AHPgBe1tyXkQZ0ch
/WLjEGNgV7B6mRuV2ur3G0lxdnhpt7C56bkOD7trZGGaFXCAoxKpTTBqasC9iudwKaMIt0AS6eEK
gjyk3bSLRy2u+SKrZjQ329h3syWYR/4HOIk6W1P/7hG2pv+/BxEggD353CDI/1IAoX6HwKBXQmzE
p3Tag1vfKWDymtT0OAsPqqeEguhXkk+84rUWaElyOZKgb5wh7AHD/SB0LBDxm/3zZ2/stLZ/E+6Y
trcs+5eDd844kgIc5upJD1EqP5SYMMGyUGrbzJyK6QfbwNKNfFUwjiwszS1yyeI4JpbzBpwzudlg
FMTCCcd7mJVioI/Wzf7O5qdJJASPXza2r3EZJZ2ejSao3Lpq9ae/6b1Y4UFv70vrfUx7puVKnzSV
ZBTqkRiDdBANhf8zq3tD92FeWP3w6y4XG8nkc8ZivNSZoC4c3++0ulZhPp7niButhn6NQhboU+a/
FGIxpcRYUpIGyabRi1FRUZ8eChodJ67FwwzqPfRqGdIvIgoBcur3A88+W1cR/ZtYMoug6qHI6Liv
xBWWrDtWhR4qGQFLarEe6GazfLYCIk303KbABPkW4X/HQ03mAKiJDORCu2fa4H16/R99JlECn0Zs
+/j/jIaGOi9VNnHvo4bp/DTn6UGFCs++pYCW1MmbUE06CnhKMtA1ESRrN+osWljb8b+8/ZgZ1O4v
AB39fDSmuxpfbM8XBmREAdqI9UaK6Azs1Ndm3sNJbvRPod50aC0z1q/+OqexQyWDCZUVhvcoI4Q5
Lyf3JLugiWJUz+I+Aza0ILpxvJT+Jbr0pp0RurjXAIai36dO/NCdnXO9EhXUTa28DiNZO9PIEdvx
48Uv3m0UyVcyN7tJ1Tpls+5XAvs0J/H+oDtKnW163j+N+iQB7GKoQ7aMGAcAclUB8j7cm8VSEXV9
Szo7nat3qCJYmqKu/6rNye4VZyy9mimBSfUkePoP0RKsmSZmRoTV2dm5cIk1mtLAQEVd488G968E
gph8mQGnmDiZapghJZgnmGJjZa6Tp9Oz77MjacMMqZznIQLt6RPDs+PTqHlZgEXYeakQaQ5fGuW/
rpPqbNmsiCE0CZwcEu3aAtR0pI2t1dEpRdVJ4de+I/kWwRDhjMMSE1104JiGpg/+4Fg89dJY2AZd
FgydOZ3P84llGiur/op70I5eZOzj9V0t5zXgVJK7gWSTsC1pzIxInGxtcCUOEGnWQjGxBXm/O8wX
B3Q9/nHkQfQEMewY11aIxa8rdAVVv0OEgKzEuxGgXBEVq6wcecqRyobaXtpbSxxkrBf4bJIT6S98
RZ4WWaY8pZ9bBEGGiJZ+3OCgzg1xbP5qWGo5qfUYzsCx0GzOQL9p+kjAUooUUeoL8j64g4GfEQB0
MLyRipelgPc3AXBMAP7v8OWnWByKh3wQb9Mxu7UpR8D93mkE57lo0oy7s2hMS7tgXJvNU9eldKAr
mYMVufwJV15cfQhdMZi+glPg05vQEtJWEIZTncJjRvJ+wgsO3cfolT5vqi2H3GU2vsENyFzuSM+N
vPEL1dMxARPAUODJ3lWtTcD9CYLMLBQHlmHDg/IZChgMPgYAswjiAkv3ZWJUR0Xm0RZQU2r7MefY
MV4sH67NTbzr3XJbZ3NDTQPU91PbFZytxexjoRD4y+eZknrQWSjU7noHu8eAhQO54F2NXGVlvxOR
AkQgxLEUH4pNQtGEdWOICskjfHjm7+F7u29dddhyaml6KjsZRLTbCy4/xAMWrUSWvKPM7g98Lltt
DDuqWB4+p1B9D9Fw7Jwhup+ESH8jOTbhH9vz7bDKCLC3YiA33VBYT4z6UoV7PKdJT0fRMLzzbA15
5owGP+4KmVvE0MOHspxJn/c3Zl0lr8yH3MrN4VUHSh6Ycj6ndpJEA4MnN0he4h79DGZ4MnXRDbHW
JevZ4Dz/pePRF7xo6OFmwD64EqNAvREsQyEvOcdIhWyFL8StRpwGSZWoVeinyT38U1z/2wNzlYej
96wLnOlMA3hR5pdx0XILI8PhBmykOlEreUsy5mffXRa4e5PM/8HvWeJfeQijPlP+vpN2Z6FILvvd
wx+k0xgwmD5tCI2mbkwlHvGfhSWMvJeWerXwwN0X/sS0K8QKcLk1BslJFkGJmWnjjB4XFhoOHaZU
C5escLEZ2wSgQf4jnHTNpV2IO9DFT0ELR4H6TvIEjXk79mWHxqma3afyacttyHeCWD2XlMeJiYhk
OQ+tGcqqqo9SwbyVp5eYhOiq8HEsOpAkM36XGujGpCIsYPCM0ZiDP82qNjJlRQy98PBIBnV6L8gC
5SORIrvci1P/5v0KaA7jP54I+27PFey/Xycyy2Ya31M3ReBj6OZLqtHIhhjCqAyoQmpe/1cPtX+9
xiq3++beQSfdd/H/wdXI4RGDInGBRaCiDeUkg/en+h6nCBF3G8LnTMrF1L92AgHnjtwanumXov68
fAK/xa7mFJDQTonQwOpQmiNp1p9T3VSRzSeIYKybbvyFxyvUIqk93Y5d4o93fNm1v935pc1SECTz
1sMqYCP1BbUTe8Sc8Epfy3o0z4luvnEVvNH0BxKz9mV/BI1DzOCx8oUMgkdjO6LPYi0YtUCDM3MB
AYNQ0j0nns59wA6MhoVtu6QcP2T/rdSsiM85uCbXifUpv58wFaA9WlQYs0MQr4PXux8gcAzZUd/8
4w87t90e9FFzRoWnH4vvrZj3YuHQZcdBSVykqtFgVY6XFeFdnYH20YyduWHzOMHNHyqfv/oBpNy9
QxDUDcVecSctJSQRR4LDG6KXPGesjIcSvIsJlAB8RHCPo9lywceqqZOj2Y1QehDIgpD9I68DPUbf
yJF1yhXj5jbxZDWD+38c+o64WiQiK8pLG6Rywa30ay84JcxUDV7rddJ9Wzt0tWO24Drt0zdPIXNP
7F2svwblGgmJAPxvT2bZZobTd3oxlydm2AHykQCgIz7HzB2VKgg8mQUsMEsYRSpUkRBkfVRQASBn
KCjk6NbFnqDUyfdzL9QG1xxBxLL68rFa8GHNb2INZfN9rKs7mXtUxujlAQlr3HISglqkJw0B1kiD
f+/czC+QYqIS2NpyTL3axFoRrI8alb0bDAWm/+o4WrjIrUixT/ktqHrZSjtA+/H+6nYsu4OmgFE3
3GPqEZdh2zTiGhhmcrdz36G14BiBf9THEqxGlGGYzn/VyRDhya3nAfTsbUSvz9gH2jgCalj1sNhh
F3CXMeUZrzQLT0S/AS7jVIWI/EgGwGYR78wMc6XEc68iSRANkMLRHF6YQup4fHEpCqAKpWzoSDlR
cG2u8sWfDryrQGsFKKZZaqzVJmWfJMrwpa0Y3JoPjKqJEkp9GOo2R9KWOLSA9OtUrXN84W2nHF+0
uvwZlo0Ez7Zi+ZQQ4FkcAyH19M1j69cZJEyb0yTEXnxyH+AKA8cmLwqGikOr3P7g2KxkKDoBiecP
K3vy7swoj1ElWn/qhbAk3+ON3Ugjaqoh2gNvLOEAyGeKyHK8EsnkHYBTHF0xlgJvTnsVKAty37Eh
BAZcWL50gwYuKgG4YKI6567Kx9NIfMdPSg6CWUnwbzYsY2tI3yRTDo/juPvqehmBQOD02lRClN2K
tixAMsy76aqXitj9mjpARBMGO4t1QmO//nC7L7dZFcq0PxE6JIG7kBg3QM2y7FsaIR0s343c1jDq
WlmlDQWy9Bo/Ct87i0RGVpy8QJ2DSby0NrJ8Qktep0tD3alZtNDWRGGh3K1QIFy1+73DVJjfdbPv
HpqJUQflGv32ePYquFfiCmMjSilU8wfZFJ9IJmG+V7dOFDpy/QfB3yeruS/KwcPGvepMt9+GLWkX
0ydBnbybLCBBpIBMAKAu4CYsgqFPnLhtB9+7CxGte+dkUmtQvfJ9HAw8JHMIKh2zhgY4PfGSJfWI
8hOYIwz+UxWuxUCS31v6hCoad9X2MJrReQC1tzmakSGHqs7yLXJyBi7YPvWTBKvEcwAlHoPjxq9v
+HCnu3VIbcveMQhp3CoICn0tWHxosUuj0AmoqCoKMXiWUVZacewn9UqRb0Auds/uheSlsOiANpXK
hYzVZWSk9fq5lonDOkKtHDeBtj97JXHkRSjqaBE3BCgo6k6z2mGKCFbEFFfnxdJvnw+kCRaJltV9
U2oZ3EnWcH0OiTyYdsfE6IV9aS9PYPmv7u3AoMhbjrdOqUaYIpCNiazclxqFGGKT0FkmRRds7teS
VjKbl3sawjs3ozPDb99wrPCMBjAA1IPpqTaEbp9on6p9n2ABbkInZKvvztQt05lk4gUkgURgkBD+
cWWSWMZeF2CfyY0NduvoNUtbz9Xc2w5X5eRIjryrnw8bBWcVlnjgftAjNZoZyeJGh63gVOk5RVR3
u/UPSPgJmY+BmFO9WQcomOiI8GwCpfaTaiAb6WOlrmI1/cUAUNfxFHMEte8tIJ2xEWvNOpECKRYz
4jW91G0ge+H4ZIQwxxnwZ3nf9/Xv7qt3WdMAW2x5c+zG69vTWsOmUmTSj5IoPwe+BJZ36+440/eI
bTx4jCEKwlf6gEG2pbf0+nDmSp2yOUjBH2LSNeLGwRYtObcmyURT+qz2tg6xAIrfpNtSAkRJ93IG
u+Faw0e1Gq3IQxHNF5YfiLWnvVmPOalZvUgrMpVhNcAHWGyeLWg+u9fWZ83Jm/COiuDSgIgm63TF
ypVvlaMU2rEoqUqbr7NrGe/aO52XSg6zEXY548gPIU2oU0xBanlmnhoY8urpRGvGv19FTGQgGTOL
y/05g20j5bf7IUTXWVxUBIkSWBo3clD5HCah4Q0LEqunqo4OCnIMyM4txo+TOMlbX9ohaZsyYENN
yL201uQXBulJ3pMjU/C8Q9PB7W1R0M24Ybr6P57HgIluhBPLoJevRd8+oLpiNGhc//3nNKyfREod
b64yDOPQW+pbqcV+2i7X5u2o+d/c6mHsGvl+shg9yhvgqizIQsK3fdiXEq7/7yJv1a0KSs/7QhDu
gW8AdH/k0ZAl3l2NCuEu6Yo5Ww+5n2J3C9dG+M8EQbWEL5O2wvYttavreLLQrcvmeOGHpFEbOWjL
8NVvIFUDkasL2LPLa0EkCVceOvAqmHK4heBPZbgS5p9UG2nl46uKpQMtf6fGOR101uUiPiZR/C0N
8CNp4GJIYFm04ZXgmDrr3B9xrtr/nrOORooKrc3MSTZpfB6fQnoXp5NfgSUyibXL/8PDCvX1knPk
OgDT5CxfNo0tRoFUwowxWwnTVtAAW/Vci6mym1t2pj3GHcmFzYPVioCOXtwi05BRVtxz2gLYu5Fh
BJAwXo4uQPnD3pG6nN5YmBe3dHXISab5FvXxCGkW9A/CaKWLX7yh8x1vVsvbFgkOAFjKU0hMRS/9
75ExyoeeytPqdwjYO2NIxV2KegQzTQzplK1KIpwqQ3+UOcnnxSZJTT5QI5VhV2AKH4Rx6Ogo/K2e
ZMfCBVG5FSbDhWk3opL2i3MM2DZz0Hq1o2z0LU3CPGMPYykkAz+q5DwBFTXTDk9nQUtKMoTlLEQA
FAEQGQTUSjpeJNJqXNVzPCXk26RoSFimmCg9WI9Qy301a1r5FLTvJ9qlUAl/Er3DecOfWUK8c9zl
GHpEOFIkCX7IbQN2c0byZ5V7NMS8s0n+pyLBI+PA5SO/SP8HSB7AozD7b4rZefjPF/aiGJVdmeYy
rpNn4Mh9AH9nNut95QIHx+rOgITg8Wd5PP8VGuWOUwJH7fjvLamozpe8Sn6qwJWjwcSFZ3TK00zK
dQabkjHlyzXYS8CosJfafZyMhs54PJnfnp04tjr4UdGwObzeXCdy7cZDmMb1rmQQA1CSETRxPlyT
QOLCWIHlmmmhTwuC7/j2DQZDpZRsJeKc+eIqOMyuwzlwnCmblC2aRjmb2nd/pk3nTsfNDbz+1bfk
b3TVekGhTAYqbUmmXtNEuepy7fm2RWAusD1q56jMX7AxLr8bwBrpg4v5WejoP9H//DztJOq7e26Q
MYqeIwTdDbA5v5aAIEJ562bhUhjGO5/R/fLHRAoZjbT5xL8kd3R0LXvRTSwEuEL1NcN4DVIAjaoy
QLoPfV9g9TUEFmVej4N8xFeyxP5bxWiIi3DQGnWDEifE9LYE6fmHfcBKcHJFVDqbJ/sgw4rIRNmE
wHPtjvUyOOnOASq6HhOlHMxnQcQF+7ZyCuP8XONsepHmyHq+uQQd9Nu1VYdMd+ndunJXVpN7rV9s
G5xWW9Qz6wWxe9uWEWN8z3h5x8Vu2eqDU79wQ4YPoUBDXfGqFxnQA4Y+C52HZYj6k98nYdCeK8Y+
WxCx8AEwSh6EVNOn5BECKQYGvJS8scEg19BxzbHOa4bC05GGs/NRlhv1Ot5ZPoKC1HK4ngsfDKh/
B9rMkJnW/jsgtfHosV7BpMuoci7Gdf8TQfbcXKOwIAUTMSs6vAE9f5ckuYvovWvudKcTf+/M7Yws
ayg0LegCWAxp5AoSWrcXRMih6Gx+AZ4yfKrKZtMPJ9ROePvyL1ighVIw0ztBBrA8mX0Oxys0FAuL
ssNdkkUjJFUP4htVs+ItIcwCdXD3E1mFvnwqyyJqb4zx2va+nT/aEILK06W1mtNgQeuBaEVZrPSi
HubldfipgkFn6TftS/UFhJ+QBwmgfuOCUqnl8kGf2UAy5tdWE1nXhaNZ+6edzuHxE4Al7QOkIqL9
DnfCA3vIHybDcD6pdux0JNUzrHDcMnmy6lOQ0tuutK2cCfUt2tL1R2izwyL5Ig2c6Nh7+zRYsN15
uraNSMoSDP93n+zSEt+057Koycb4aOOYVSIqsPOhR9WDw+C1E46Km2jk49A2GelddHsxeBmZ3zjr
Z6Ig0p2bveyM/bxhg1rkS/EZGYyeCIWent7lpdtzwSdTDvWKpHYrmf37MWM5z0D02Xi0JtD94965
gD9B1uZFhvh2gu1hykSMYmuYxYXsKdyaEqUiaaKBBSkjVEd6qFoeVFw5HRRrcJns03adptyfRNa9
LgJ72fJgaFkVvOikpqzS71D32pdSrnx9QV0CAPy2KI+tKKAc9HTh8e7XYVqr5NJR7Ugf9DwB1hJ1
BVqOarwDYMeXiFA1eslgUsKxecNZbVEt7G1ZAdqOmzTdim98ofWSWoGNp0p7Cll4AmQi43WMrAmH
2hNfIkG+4dfDVR6xnMOE5Wwhz3V31azsHCB8ZOjDgJib0QSS3w3GBdzklWYajgQjtCsh+xy0ZKgf
h55Gafy26b7gqcNpRvzLiy0BuXNg8wVOCRAX5n8XEWfMuMho134DmSpHSt0Edy7pVgOlQi8jVjyE
G/xK6MOEENFwQ9WZqwbTUtYZy4an1sYbKxSLHaE6TQlKnFgildglLOZ27Kt4PD2EzATcyafZ6CoS
SdUA+7hAIeJ43Biznw1FIueBrO0IlGGHA8CPsP5xAdCVX/bxNZG1+9+7OT9/9QIrKfmhhPGQ1W3Y
ri7JRrMpPQoV6Qs0rwGOc5LHvj54Jnv5kFYY298DGKgDsksNTYkwX9TJir4bmr+RL/rrbaHbwMw7
TXh7eGjLk+PltSQPhojef+5/V63CoHtSXXgFIBsangyL2bqJSFsubt8zprfASsIEJWryK+t9/Cwx
VfMUUXlYWsofb4gTGw91KioXUbNUUP8f0Khv8rDtO8od++ap9whDrExgV1AhG0DkpbZKmrfV/rb2
bPUVyhtN4NHYDmxPyX0aNztElYMgWM9IrZxMND5BHdyqrzCRfuTzhBimFhibDjkrT0pVnV5zf8n5
8lozAAvz+wv4KSBID+mAlGlOAzg2fQ+aN+5QXotiXCG/87A5Ef9S+iqzzcfp4TpeKgMNE357L3bn
0RPmtNAXNHdkiKcePupQSCUiI26ubeoAnZToYlYPMjVYDv872CMiNkxJ0Ubu/kodivqGRV1Vjlwt
FDhSKwS3gQi9Trz90Vc3bsb4ZXyAWmsBL7QM89OerWZNvFkNiBDdbfO8mYCaSVOFpvi057OlU4xJ
qoRXN1MzTkuJsuwH+3iSraK9Z7yMWMWSYyyzmEyUCwRsoOBUhRp4a+tdCKH2zCD5VYzaBNSy2It9
Jl3N57782VkLkaDuoU2E+tq/Du8RRmA3xwzfwY62cJUNfvDFidmt5sZUDnoF1Gy1bUwY3Fd7ZZ6G
l9ZspdpwnV3eYlSahcEgrUaCedsaHyk2bbDspQ+AMk35gq411CY388OWO6pgB+lWGgTjYWM2kxZn
+jX5iO9tEbjeyfy30WNiLkiuOsre/e1eK6cvSa9o5PHuFXK2JJ1V9zTfxijUWueldbXAVsVN2SmV
5D0VqzcHNmby5H8de10STiNff+G9K+YpNI7YSwl5mgCiFMZAGyqvsWBmDWlIMdbULLlPONOtfnQe
oOZdxReHGBwoBAR+IPnPfFnHI40/aW2TMNiElTx1Vi9NwguOjMrmA28wnQLZZEGEI8iIyRKcOlAv
KSbLJrgY3S8/B/wnmg+QJ3y2W5uoS/BDiwzba4jHXLXpqGNOvIDjpfSy3cGn3nLNAnFlcXn2NPE3
K+cL38QclZ/ubuzSddQp5502KRWmCl2wsoLzv2DwofSImYA9U6dO7wTLYEw1Ou6bB5XAICGCRLGL
HTDAaSlDDs1b9AJ7A87eFzRr5j3OKWL0uR9z5cNtywN4F50jgEVnKC/kej/S4Y6pdgdxiLGKm3Sk
LcrCwY9/0DP4sz2EqsBOBEsrsvbSMtRvzr3k5HJId1mZp0kuLMZSTw05pdPbiTmxFFc/3+wesfsV
IZaqzxkIwbsfzkqYiHAzUpxeungrmACwINX2NgoX9xZuoeDOEFR0hjj8wNO621xRZV9BGiaZymRZ
wk++FBBoefihSbu3+lh5UR3yd/2S4VRqTTGFjSia2LflA1U4LJ9r51l5fECiAOY0bNLumwE18YkT
8vc6as5jhQH1YJKvaqkJOJr8lllyH0KFCZoCfeQpz0osF0+smzKUQHAcms3b7Q3qS0+V0DSAns2o
UiDlAHcJJC7CWbTFM5a/SP0gOx5PySaIJLzDxXClZ1rMy9LbbN3kQS539sZEZCUliYeZN4GJv3MT
bEx6xYfYAqAMuf8/HOXJTfKHNu+W3tFCyr0aDPQU981Ra0nX40OzbRhq0jAGzjP86+nCEQPxoT6Q
A0hGoT8HoVWRCzi4u/AHUeOBBRvexdqfWCnBBj4d23so9IF6gOqGlFC7n/UYUa3HEEW1vkoEb4u8
jJOcPZtpnhpLpfVI+grFsiQlni8HytePYp6fk9IJ6FzQHrU/uWTduMBuI7M3Z3rUsfrffCzQYA4I
xXTTW927JQ42XqjT2rowYj7gpiyFI4tIT5l3fUDECliIwT/lGSMG8DTCDGaUxPP2CujD490vLDT6
NQp6t7j8pK6EIGol139wF5hmzI/zJv1Nq/qJCpFBt0Tm8a7VA7/NqqmbSHaUt2gXELQ4go/37IHQ
htnRtb0qLREXx3FmI7lSq5HJZ0X2l6A2GjSKmaqTh+52jed2u+lUgYGew03a+kd5d5W0oq+XsvUm
/EKarprrOd6ged8rx+8TEQ4SBSRF5WMPpL42VdvGhQoUzYIs0p4+w2CDA0QnFrOAXusydfn6ycms
Poz3VBH4G1Q68r7R+WrmNccF3bpe53d2BUAa/gmk04C4KMd5RRWTFW5hZCJ1OvAvoLa4U9UWK7J1
UBvJjlMfagX44QmpHGXC60n95/eCf7gYLL3vlIYSaIkL4GKVtRYGoec5wzm4Moxzb3Zesqky1Xps
WICw/Pc1DTor+9RqR/3xcZp3XVwclsBzcPZ/dXWdwpJbwHzNWq9MBInWy4ynCyctktV4IraFrnM7
ydrOCqsC1OgVoPT+W6VVSqnbb7GAzc7kWLrQpy2CEJXkOhgtIBGuKSD84GX1xOe1m2iMM1uONRo0
FFJi/AJ0UTtxxxcnlfxZM6OcntBe6+UWWJAt9bkh1sX4/rfwtMMz9WpRGKbI5jSmaENSAuAYW7I3
GymJsbp2Qb37+qdNeIAq9hD6oi7GERbDIVBjafPH/Gv7Ltt1ZZ28xLcPAm53V14GD0v18hBbGoBC
B+7JwOS5oL1778yFrkmXYKmqK/f0GmmggD1v7GwfeuKOOoHYilbuIB3BgcNzqbeSqFbPSMHnGn8w
Hc62rGlPROKANopHA8cuSq8vkA6EQGBYX/cWw7yC0aCY4sYx6CvQkR+8PTEO3MfofvPhfgLfxnk+
lcOEKPFiFXoqf4WierWaMBonuFAsl21+AWQoIycUVYEuk1bWNiKW433oBu/bKjQ01kvVRkpeToyM
tYDkBz38nixtzDqbCXmtvi5PRG2Y3F1xTcdPYLz9IaddXPCNcr8q5Xew/rqkvFbz2aVc6IaX1f2g
44oPCBu9qyMIan50WM2LzpTyeVd3LM7Ns5GCp4STlJ7CAgPpQgYWe/CR+5aNZdeomC/KcE0+I+ur
hGD7eq17aJa+UxL2GpvaEEbcxGLZrp6bR8StescIKrtvHSBqa2k04iZxPyOasD4fj9pI09n8QBAO
vP+A/q7mGZD72tYXAio57VgsPDrcn5TTYaz2Zjtbcj++/WWue13z/m4zRUVJZL+Mo1973mvjkwB8
16jUGP/bW4huhdJ84VfCLObbKNgLeLPE5RoCXkqT11L9zJlZAIzmtZ4ZN0r8MDGyeuKN7EuqDN1o
tae04dqAKZpyTk7T1Nl9D65KQl2MXEzzUGrr2ynQpsPkjyIzFmi/FhaKjqZcjOKNPqgK2USwY3zr
8XCQ8m9WLkn1Lmew9ci8JLW4hrA8J0QHKD5bmmqpEVVSkAalizgeM9PkZlKmQU4q9ELkbSGMvCDm
HNJuxOMhoGF0EKFxXzrnaerk9hVJDkoScmY3B+AYqEIxu+UbZ6B6MBJ3+eeY34SZJYyCcDyND8x4
LrzTdphzokTgYoWlTcBhc0xmiMnCXkNko7Y4GmH/Exkduy78dzB/My2gx9yxkJvCmWYE2+RWv/nJ
x019qI5nPC8Koqf5KtYmzU0NvGBYGoSTC3F/sOgy2+03gZrDQAl8FjIE8ycLuqMWe2na8MQF8HPP
3pmlkFvtSHIJ4slcg2sJ5aQMaaqH436QUk0ypqX4vy3Sv3CSh1i/4I+yQGFo5qf/oW/MWMgvNxKU
JojXYnW8t7YH+nkmARJZGlubeVs1MQgoPnuvQXUgYktWfdv1RJjVnPLoinWC0K5QTqWt0Y6IaijO
tF6iuwD7cJ+wca46W8B8L0DEQz9XWUDdye0bSq/slpOiaBI6V4ixy8JGnhLbFbLYZlSBTS8FFZ5Z
wcW0FV3L+T/2Q6xpXVCYY/JTrkEQ4Nv+7Dz6DdK000MudkTsg6YF/HaeRSA4RNIdJb7LRS3+0wiY
GeVJttNhqBEidKKrLz9AxnLwmYii00728/jVNPpQOrO8bk6o3PWdf4OyeAciVypAVEc2DwTxC/Ie
XiYviqUOHvTKB7GMRaJ1CpYkyNx39d8QB+mJaPErqys6Dv1GR4cW5aL6j8oD6hxV1d0SNDJRb4Iv
PpMaQzlAHNyIuKrVaIgwmytG5DyAUP7TUYL7miR3R3In4hjNo2m9NGsUxXeUC6CdqgTJ2tm21UKS
ojHXXiZF0irXDths5AkQ7lb55JwD+VDpEdW1ZiOE/j4NiJ5x09t7Xf/Kj5QpNVS2CMqCszX2WezO
uZPJnH+Bj2FGMrCNWAFmIa/aZbR07H2vOWPM0L+9gRgcobvSUXtspPgFJdiZ0Cp738T9g/+CYj0G
ZHoo/WVb7EI4dfVOD5sY7vokEbCHc9E7/Ak6I/RbbzN1w1J4nxfHzhhjeMEYiIUM/RntTMwmJBsl
+d8N0UIGnLxs3gkJU7uJtUAdv+Mr+uLKoR23Dbj/mKJa1TIBNm/VVQctupa+7Ml0ydsS9MbZ6jCk
mdf0eVki/6TAtGuEq6S2UGjgkWzuqSomB1TNPvgI3hHkthxS6AV0Il8q5mLyze6HMJZDcL+BHU2Z
pWq/sGggzm1d/Rrzzs8gE9qYapccp1dXa+CrXl43XpIkguCWF8WdiQdhjke9sdBj1ZFQuKBTx+IP
AXboMMfI1QGRGmyKzgarmGwaZQfDW9kXOxpKHDR6C8J/impnalACjqS2SgrtKyXEb4zut9Pp15BS
vlVb0L86ZxVvOfB0yGxvB6i9tDZrqE2/e9VBexHhtfQkPKsE7RYTBJhrlWxNFkdkZswmCT5cn++o
TlHb61K70vQBTfjyJ34L6sAS1eBTM+W734hZZcMv8RElK9QFU9yxvarugnugP6dPXlCs4Le69kLy
EKqzN5H5azkFmNsktE1dXj7aM5+kOGAge3kgyN0iGu+zTO8y8RjBLxYNsl8TfhOOplwSJ4HZBgKj
E7ZTI2CkQ8E6Gf9kpYeUgf0/PK8HyhE6KjplB3jW+4Q3vf5cfR5kQ2Okyp4o25FinSS1Ww4q016G
8F++YgcL7/8MFFdnOg3M+WzMG2pkpOn57P+SpzYYi6YJ8/z7kRESKn/NZIBvsGeJANwngdNEBQMS
qZOMMDdpqGJeNkHPnDsHhv7tUMNjOZLQI7WYyq9+rVODxJnP4/Mcypov+AUY5Vyr8SdHxBk3LjS9
b4gaPVGOWDsg+QrI38e4OFbxXcS3DxkkErC9mQB7j72b/5FFYxZzxgoLLJZZ0EGfGyWo4b1IZ1k4
huZ3nXqEmYu2CLjab3/IeZuzocjH6UV87VAaGmCQhlITKNk7pICuUym5wjZs353ygE5C3yum9J3P
DJNn7I4BvNsjm+U8LTAlyfVhtKh1n4NqZg1xiu0CzxgRPqBKvQUUBx2YwUdV93kgMxdLYwSV6vCW
B5qAyy/D/utMW7G+HHzfKDCR1N0V3SdinexOuaBix3QiKSyyVowvCHFbhzWGxTHH/Nxyb24zs1uP
i8DYNpXAO+6v+oQNV48qanikoy9YTqyA2i3FSMEmBy554JFt759YLdNC/srnYI/aLlpQW3XlJ9gg
bSBvjELJDs4Uzchqd39LAd/wq0UtKY3i4+6Kg67im2vcrR7/sfXdj5NskfM4HRL3uHi/qJW0bn2P
l+3derCYorUYMnEaYMnlAAxLyn8xFD8B2Qh93mQjo+lztvf55KXaHsRtcqveMDeKeFiEg3PZECYb
8z58uro0qDSB5fRsEViD7yMMAb+g5ypVlEEe1XLGMP3HgNUPh/TSpxeGHFkYvVL+ABvyo7T0CgV9
WP0kbUoEyRj6HB+DJB47NxelRdQosRUY9QqLrkhXLDsgmCvfbzy5icaMJDq+r0pNOFCFRYga2Njq
+yomTgEYPPlEyp2rRIyLvwLGb2hVGVFuvxcn1npPH4qF57esc0WjENOLFHllOSk12oZrJU+t78mv
hmkddnRD9xsIkqcS0IKJUBFrQYswAuBYteVgZ7eZJ2SJa4Dv3E7icR9vgc7O1KykGcxZHtt9iwN1
2++dRnqsH0baf5AJ3n6qAhAu3pYoTgF3xY1x4bcBhk0gA/z/4P/BfbKLQDDKGMPznZJ9bZEKYWsT
fgx1cvad79v/8KP7fzPV+lDKpKhQzplsFawZh56Yu5vLY0RG9odS4eKa7UzGMg1BtOGAcxEXoWFA
HWdr5iSxiADff1Qq0wWoXC7eZN5WJFdUfdTEHfg/KBRLelMc4WbL2+GRBNm5v6ARcSVxcSIf9EGX
yJv/qwflsNrBYB1ND/fhcT8SQHbMNt4KaMi185WDKC9L9kcBbeIleXjdWvStmtQ79WuU/PtoJmML
ovpd2m1XxnEPk5w5PjY6K49Yo8KOvNA9Mtf7G3Phh/wEhbOu8w/XLrypy0JM9vDHz8H1R5R3yhRE
er8Yz+nuJMumcMyhKZGa19NDusEZZQAR2Nw97fIOYGlwueqIj0Saittr0NxyfqmZasVLUKxIdIX6
xLpH03qDM+6UMHLgustT/RHSNYJuIa5rZfcYU3Lea1OlFzx/PxNocxdNUoZ1rd3PLgQmq2ZmEoJU
Kn2KScLSvNjClZ/kvFVoLsO/BP+4PQmh71Q8jS7/moVpiwUjNSNkrxScQgO8O1vdI5C1Kb69L3dY
dNzCFym/VMs0xcN0ahAqiaxgd4Su7PB+sVf1eaarwxSpDwlA1L250zWbQNC7PKt7eDNm16DpPeq7
Azva3AHFj6GwyZ6Kdq4m1cajvrpEl76A1UcAiMC5tvY8DzxFDPu2fRc7Y//gwqbSZNGFVliTGD1x
n32G/is0C/5IYObqvagVZC3T8ioQYFBwQxKqJ6yszychIvP9BMZznc1spAw6v47BdB4nkQlwshVe
heSpSNy5iLDCElbmEGdCs0Y5Z94RhPCfVtvhhGWv9ivZkRAkx2m6/fuTtGs/zZZWxG2vOC337iIL
z8EkrQgHKsI5pVO8wb/y0965ofkG5UPmTjphmuNp85hiAAyMjDoqHv1MlKHvjklchtTafU1uI5i1
4Leh517czKZ1f3NCr/OaXnNYfaEAtnjqJkTb9DoaqI4VOFn6WQLr7Pti9yhKdE69pOdwZVMqhl2d
h1OoO+O3WmmIB5w8aY/7bKFSyzT0ZlL448K1Ym/PdumsX1pIP3DyuN3GfRnu4OhzYZ2dj6EGh8o7
MGilYh7kTvhcuKldTzniC1nRErlC1ecHJ/P0t48RY6Ld4mzHHLokA0kpBQqvXUbKEIQqA1hh7xYX
da0mScX4bPsmu4C3auiWTZMN/ju7wDjn2kVkMcaZnkBSmFmEf63dE+AKWa8OmIl9j3O2XQzAEA5k
STRdoOaRlSo8gOveIPp4ini0FX6xsl2Zfk8lvJmHSWBcmNEJIUrVbcFIaWN3xFwKQw3VTs041cz1
YoExUw/uiyZ8X2YqEMl3cGfAMjKauma7HIKs/LKLAmskN+AIRcw+KqTS/ZpSw5nDt/vQ8tnoqte6
wgoGClA/APKfdB289v37rS09alVg8vMSYRi46HfEv1K1eG1Wzz/EeeYKSqO0RLbVS3TwEJX/0goX
zzgZXE48WH9cbW09GbHU1JorcYsUWPfuhJFs11cqbMtkJyi8qNRv15Z6aWCWsQKQBkch4pmBeTwY
zkkWDG5zNTjIMHLgWA1xuvwBbJrY/M9dgPlUEFAfO7DEJKxNRwUzubNJGzXjWGLc3ItjTuOHE8fZ
0gbvpsWcHrmzpkt3GMsJ/ZBlgPCKreqo7mWJ+0uJL0woumqjyH+Hkrhg6puv1aOuSjH2mEscNlMu
C6edQ23f8sfWZM1sU9+058W6iO7wpLlKd9lhYon0tKQqNtXorbMHYvPKw8jq5zeEploatwje7pRp
QdGm1GukWgKtchf1Wz12C5m14X8P2Y2utLvFxgG/97dZo6ofTZ9VVODDHlowtegHxDlvAKYaqh/e
Xs4cBp1MpA6EenTh0FSGtdqpfp1j/McS8ls7dJdPlWqAjLGrZxbdoHcKojHVb/dj1UzAkAt3LQqM
P/NzybO9Q7ZyOFvTLx6dEPOT2jQh9GMu34tiywuzN8b91ulyFWCU+FNV2q5DPDv488Sf1RQOKRSC
HeRyoiDCae4bibx5r1g1ttlunMYIV6pnggyaQy3rLWpGsiRzYGs89jKdDtsMd23d/m/+jhBpLSP7
k/QpHGeQ611bgl1InM9fhPc/rYlBkPvaN37T0F9PD1/9hmmGfoPRkPIXxHCL5bTvgnuM7WoDa4qF
6iMJkQquaf76b2j4qAAu4bb11Zhylyn8CPthQct3Ba/dYDEyqC0KZj027zubAcTybrYmtCtN+zJG
1KXPLbQV2MYZVxIK8XaJ/Td4K3Y3+1EPWrakMRUrxaIQysaERK65f4Js/rj+pj1fSBmoRUkT9Ku7
Bf6tPtzP/s9v2or+1AXWwa1oGasbYcKTjrfJt/YSb/QWs/Q8Z5h4HjJ+Dt97U4BFeOwYSX3yX30U
0Ysvo67FGIqlAxp6Gvodjz2ZYRJsxgM8JSi5QFLxdSda4LaP4EqpJPk8Nv1TjCED9fcXdi6pqEUT
IerQTyTgP9U0mLa/6rOHYOqmP8LZ4yI98k3NsXd1k+17eYdaBnubm3FHOeY3mXJxgjYKn/V8X0tG
Ah3ottLGKL8BqkC68FaS5zfVc9Hwrh+Lrd6OZBhnPAAzfx14pWWKOzykPDUFvXHajSdeUliYYX7i
Ip3llbUAnS+YOlOtQ7QC/eoCZqblNey2iC+XQC2+y/jzRjsbG1j1a8o+ytEyXS2kKz513B8v4hrY
wfYh1ZKohmK7X5OG+qHM8YBEcDyTWWVnJ0jzz4VQQrrWQ5vnC7ZOmoenxih0XkHyf7o9cvzVdKy9
R7NgwENI2oyrjd+eufWy7teO1Sh7/+tTTEiViBLDkt1e2m9zXaOf6+LY5z7sKZ+Enx/TEQcWkFV/
+0+J56OLevnS7f3njlMZRPRDFZyZqwY7vrKooVNJ+gsvC48IoyENqGZnIEvdgPYwF8qqDlQD7OYL
Lumg1OGNIgzkBUUnVgRlIsZqfcKVo+FoXd3sYFds9MO/R3Aw3ychUIn96Eh2zmuupRaZW0NDOKG2
umvk9aml8XuSRuFKJkV0ITN+oA5EFXtitoZ2UMNL9GuU4St7UckEVLj9k8Hj3TyMltwlVSMrqGhj
63lWOwN1n7RZ/0RVXFpQeU+owBNvBQwg6TzCwP9CcAFzrsgnHz4LrEt1R0kwk5cCuFzHnKLup+yI
YWVDDHOgUuQQwYhdLeTDefZ+3K4Lhsaq45YaeZA7Er4HoOMgnq/t+FoTyPBF3g/1CcbjKOgLFOhO
rmkK71r2iVTpdOv6orC3JD14zqBM4UY5L7LjiZBnPkiHhKKK/OaEv61/GfiUtWqmGglS4EeXUKMu
Yhn8W7+pez1YF/2xWxJrIz9dx1fIQOEEQkeedDApBt+SOPoE3RdZshLgzCjzsZAoxs/HtUOTxx2P
OsJEmnOUuOtAufCWD7YRTU+Tdp4fZAAz95uF7hKjIIATiJ5/MUWSzd1KVW0oeDLWNsy2IIiDk2TI
HtbLcviB3fwbnxMh0EqOuEsyfzUDw1Cm5/CmDQnKGvEUYcKe9Gp7Sg35IZMbWwrU6YKgSioGjRrj
vg0S1nvhY5GUOTCj6ilQTwlXk8KRx8UG4fqBtvgicaiHXoWGxMp8wKa2l9pQVkO+0tI90qX6iDB5
bRDmZjDWC+EHfnH4c8udOmSmDejcgBDb1IUYpEqe9cggOepY0HYX88MzCxeTO6lmEdZ3Li54yP8H
MXx6dhisTkH+cPZI2dV0cXIzpsLQHbUhOC9CR4Q2mkQglZz6XUVuoLx84jAhxX+NB65ILvNztKfw
NVZkg6JICCU5iM4prbsbrKFnBYWbZwPGxchz2BovfzPEcY7URrmyaqazzncwi3DTcEO0Fk0nEB4P
DiPHbDksli4j3mdGYWTL5xBMqXcyLhtVlsMJfHztJ9CuecJ8X8Ewdmk1net/YIc3EvMItnwna/HN
yjGfpyNqYIwdvLFP5ushczQrybPTFZvM5ULfGLPRJq76ltLRedR8uqcJuOXv7OCfOhTcZKgqNVDO
X7XGicUbLBdLCSPo2jloGCU+XcUMTYuu5wk+rK7/uZHqKFh8KO9Ab/Vvmh+kMEulLB5YNrYKY2KC
Dnz+p6w8pX/l2A29qsf9q8AnlYtCNDd/SUK7NzV+dQlTcUG8gBVkl8bspA2Ma+jDlK2EwoUaAIuf
qoKD+zB2TEeyDJvc0uCh646PJ7pqR2rZ7FgHsDT3YQ+fxshMpqRvcFvvxnnGkLHNLWF5nufAzcht
QOGdREBdtXTonmZ2lSNBEmmgTZjbWcZp4FAlknyA1JIiVf4IU2QfQ70tL4XA25f8Nm+vZCQcYn87
7XtypidrElbGC7+5Dowqu7t3HS//MAl4eefzkyq4CetGmmYRwYY18K+L7vrp4SyLQe3ZSXIR89XC
W8u9swiG1zNVRQzm8oE+nRlYlP/FVjE61Nz/3QOdOy4hphgJ2SPfmlG0fT0l/+qxXzYAgC1JqOSI
Tiyytsy2ONbSzolOoi4Tdjqnpm70xFBEtXYo0O0kgR/cjA1/Y+Al5KOlnRwgygYeEBdUN/Qd67OM
9bseHGh6MEPT9cRR72+YMfOicAcg3aqQ+apnJfRJhSVhZOr1mZJle0NNALHgWAggBlrVdfOgzbev
UukhlcjNIP7RNcAa3bx0Wl4a6q6eQ/drsJrWSybPanQIyy6DXhYEGtr6m+mtmsQ0KzBbqVY4uv4E
VaFPLnfiXVHsX80vJsWzEj6Ckldq5hDvHA2pNSB9jFxEvz4XOd6RSnDAQAuUkerE7pP28nyhVmoT
uze8qkqxQBmkRPvlONs4wOExXp2FKX8UvC3RJDE1thTG8TzaByDAm2mRVlQmL/Dx7RxODCgc57NZ
7Zy4SwBq/opHCziEqG2HItEQEfMPxuiO9cw2l1HPPMNDj2uIDiYtF3TB570/5bBQlZ8WcQY/9Q3S
iihZ9M7+YvkKAoMMJ2N0XiUjs7x9XO2ibeh03HPWT1cskL929PtojrTpNHV39C324JHo5y9Rvf+O
fJsos0H5QUzVitJjNNpmizqCYus5Odw7W1yLTfrpVPHJ8rxUNIa78XDMVrV4X4pG4zLiNt5TMPAY
u8erYrzl8wMsP5I29PTO+SI3ZWkR2Sz6I1DXP3RZYxkov0B1Yu9j7pAyiPlm7taK71yBwhZf6qid
xviyClh7QbrQXNIgkQvu6y0B3y8p0BMgbIcqFyKgge7NxiaWnYb6Ltlh45PFqoaYH7z5uVtD4h+d
58ODVg1HvRKEtVykirSgzRqqbYjIyEqNgk8NQcsiak79nYCrLpEdaQA2e5xE/dJYcgNi8sR2Utlq
XlnCCC3vwSuxXeFCc9kmJmhEZrJqF713q0jacM8T/5oFgftBAH+ncVEHLwH6JyI06Ii+agCGlhAi
+29LUtqR+1ZnzIkIaM+4/dzQZmNOIP1izkKS0daHx43KbWnY/xIltJ31bS8EvOi2MNwQOrnc2mXj
vbao+kVqZRDVPm1DSiFkX6qyYrYXTGOs8k4Qrh3Nit7GQRfornhOfdrZ/9mcqNrrZrmv46XyS1p+
m+3qCU4l8gCrgF2wRpOIPLv/31UzpYI9iIqQgJk8Ft31qySZ9+5vH9lMl2Y4VZ8vgJzwfWkFSC2G
Rkhj+a0+eIN2/18qUm2Nu12OkMPc1qgj0kCf00jFkz1L9p42ZBdb+BiSBzpC19RSwXAefp7KlnQo
Ok/66iu+NFbMIIw9BkH/b7eSmSmKnW/HWDmOl5v2GKiduPd7pFaOgK79GL+6re5CFHvZ4ifsaoUA
TGVnh0UUM1PIleaVOTJFAWgq6vZMpbIwwv7SNY/IdKFeZtfF4a2hRhg7irI1Sf4Tf+p0qlEzDmmA
L4aKj2vP89Jd9MBOGp7eN2MKWTIEZiJt7DVaFtsOzmLJn20lGk7Th/O75nJHlVoQfPuEHYzjtza+
rDebtnWf0LLETWzqlxwVxJ1miVixP4V5omRVuyGCWYbPdN743MUs9BAgukLcaj/5yFjCSWaxEQWj
tHMqU6UhTy7IanEMPo8IiiQje2YrWRgR/YwNRmY2DhhJZmeYZpxUj35cMeU7jdFcV0/Qw2a0DQ0f
zZyjNntfB/kuDjtf/zD+kipYN5cEF0n3TVgaTeaAZHWFHg2YXOcFAcC24np6CElfNaoSd3QQOHes
MioHDLQFCmjDX8jYnqP9qpfz3pmr+qWgPkGO+yM2aBhlrW5bKz9wM23nMyoquDBMZWPyLyGrvS+0
8/kNCRx9iCpiDo4/jBpngltygxIW8x0zJOo7L0EoAAMsACUswMLgF9/I2u/TN43PrZfe5XUCbPnj
wLqWSJCLuU/hnqHTtH8m6SkK179ruM2jdbxw26NezVvlxmop3Z5h0CscCOtt5KcOqCBAb+rg2QXh
nxmohV0Joxk0z+dT83qEgVwBCz4tzGMNWWIGoLAC8rMAgplTS7C3BUPLXnxfUjJjFZsr5qyzINeC
YkAk2oF1GTpBsjBJJq16/PKJxtJ7RHzsTYTgkWxJVjnfUXa1sz4jC7XMFK+N1QsasCiV514suiwY
lmqMlBUXw51+VAJGmtYwXktnT/kNnusc7bChVXl8aABIdUtIwWmia7CZXId51eSR1zNDDC3ZoZX6
nPEWMc6nJHAdOS1KOCAs2y+bgvilFLFRpUtug7quUAXHSB9B/xqq9CQvBlQI58apYw4JkA2fR3F4
1pkcLxzvynxdnuMF1V9ihb/dmfQZUlHKNbT9toWmr6f2ff4Ka9pf7nlUt91KbS97KUNRBpWM633+
uXm3b6b7pqXWm1JgP5hfeHUjMB2gyVIhVme9loqx1DXYgpE2ZQLRzAA7b2B2JxRy7quWv2OJdK7l
fBDbF69heEubTHnRYqZFU9gmKiT3U3fwtlmYtq6jYxNWMU5XZSbkmzM3xe7LR4KCvbzn4S7fqOba
sEn04seo6gyzDWhACM8uIr1bb4kDqBJXtbImuknodE0Wa8J/ta1YDt5CSa2Dv/DawC9TYYyq9J8k
cEOahJhw4MXu+mfhZ3cHoBW900WHhK9z5O52q46gU91jsh2xh7c8Q2reAIZfiPWKA+oUsbjFjWZt
+cIOWjqUUHThgVPtNn1jUj4/yIv6DmwF+sdiBrOQh+QmxUpnp2CipZDi77dg4Ggt3NAR46eLUhGL
MwGCXd+PaHV/0HCGW5cA/3/j2xiCGW4tWauFaARprHqqate9HuOMYY8NkGHJqwPf1s/wCd4NWFdH
UfDNxVJfPJJMaBiyL5sqQOOrbRSdtm/soq8KXgxh5t+DompXuwbtCsAsPOdJcmVpBeOhQPO246wy
RNH4jnbkCSfSiPIN9N1Jhsx02R9jPlrN7VUru4ZIV4gKHvAerhuquVFaFouNMLmF5okPQDneFbWY
30sFoKMttH4fWNXUO5v0mK6pfGf2SPCb+RNk7l6jbGUyjWWV/6Em/bSFhyyW9BGQjNe1npL7oPsw
2qWkx7LHfDiGPn6AKBulxEIkDWdVlu4lVWbn2w8aKsBtvZ5qZZRJJ7Ak9ff2u0+zbq86TgoqAOHI
Tc4EqJpT11pKuhU+1wXhXfw9uwBtX3PHlidA99yplvS4ZecNZA+24Mb4SOxUmOcOIH4eYd5bUViL
u1t96bDUHW7AEkxOGftRI0B9RDd3putkpwnlz9yl/mV472BHzwIZAefXLgg/9cIvsEYtc56LZEiA
F3NXO7H+iIkGlhVQzpwHx+MEuR3ddAxWLQsvEjV7JRnyYPwfZQEijFTTKujTmOJtZaSBxUVdhveG
bLN3yttZdKTAs504EC4FJM4zg6rEC30yHBksBDBI6PGccV2MQ5zJG+v9jJy3jCrSRfiJqzwBfKVw
ka9trYPJUDsXbwJ4Gs2T2/7tDLYorNobBzhNjYXhICa315lrGvd4R2qwcb1JjcNi05uDRtgOMU68
yFgRMbUHvbw+Qi+KWyFY4AMcHA1MvcBI5Kcorlcy3iipDh5SSHI63Ln0D6u3ROuiE4FJ7F4jqWA0
p1ZhEl7wm4sbOGtGSB1M2vvTuHJ4MLgMFPzZSydIIS+3NfijTPaoF8H5ZhE6Eh2Ef6AkVa9Mzasr
QczFJKW+sIArsIvd2zc6BntA4j8RaQsOW4f2/mJg26dejLggUM2XuuwkVA2OVRwYkMGGOwXrAnSi
mbMvxRadjznSsRI2TJ1wHxdmzH3634+Q4PUSctpVu50805BJyK+wiiX/p5dVkK2JF0QPgPfLFHLD
i+swGcu9O9v2STjuhaN55cSE/4Sket1E6ihxjXSfqeSrILPSXXZV3xiIxPV4YP5lGkNqpne3W2Oh
wJGAg56x+G2cT8kJEoE5y+Rd2Ws8jTYHiSu64BgI52ZgLlJzA2SMsOEm+JHKjsgxB3wLuxc1zA2M
cPTJx4iW7wqcplNkLKisYfLT963hllJQfGeC/cfIHoAOlin+dnT3xAM/+14EbCnz6tsXsC+tbtOy
cp+bKBFWs+LZVfnLDbKh+lxvzsYVmzh+Kge/SsrnpqkLFP0o/PwZELtK8Us4Tgxaqn355+A4izYD
M33XUqULMU5lF08gROAK7pZvXxMnaF25z002o8S+tDu3ml54rfbSjITyhQRLAS5CKjQhOOvogcO5
DuASGMz3+oYViI5ozekPqckku+UccOxmEV8X6P/MUEQ18KSVX8Dsized8YuXyQkinU/VM77y63UC
TzkOvBFD9B9ZENssKm5bfZ7BqYgiiD/Cz5ypSCrZ1X9TnxJA3QSrDB2bdgwjaZCTJXuDWIIjhaRi
zir0rbKVLCearC+mA/IYrFIUjTN6ARZHP1oZWBBeTMMzBdNNSEdSXTy5U5Y+82hYBbBuxWo2sR4w
qOqgZA3QMEHBUG6ybc32JfM+20GGQLOTkCAKftja3ZepPtN7X+zhsGvgKitDbOoxF79kcM5oIz0X
UFfT0MZJ8ad+sTHcnpdrZlc9K4+5E1hmPij2mVD7CEmvgijJGFjxJuyTyQyuLF0f2RPDS5Ki1FPm
VwyOzs8cKW74BpPttjmPs+tPNlyk+ftCIRiINpuXMRWOJRy35J/CXWSK4FEjoFxBultIElVOWqpm
fZ6oR+PTb9ZK4xn8vGmD92QpAufxijeuTK/NUcOTWnjKsUOrhfVSnd6LIdnTmny+fnkpGTdQm+rF
WL0D3f35vljZcMIpA4735K/iVkGt+DGhXHzhQT72WZ/263gtS47YfVqZzeoIYSc3O8WV38vIVEJD
XLyx8UBG0lZVwp8iwaDBXvR5FV/piuAcOxyk3cyVFR6qrI/dLrPaqSxQEEXJ9H9eyDSsFmpmXpZ5
WBsmK8iw5H+pqoSU8xECyFugftJPuzjJIuZoq/JwDKgjK2lYc5GGbECnz1a+N+Z0/WsgVgxtWi/V
a24cObZqFomNFxGR5osRQ3+VQjkJ7JgTmmHpUPM8wUauU65wsxcV+1B+KNhapzRbfOqzqU4lIlZu
PAjyklIs7qsypYGi+c/rhfuSDjLFqEfS12cqF2pZhIJEn3QFJCa8z1TzSk4IBUtoezZ9zkRxgfWz
15YC2UH+5h6Cyzou42ETq5dw/sP0DDU9hIqREAZuQav07O9op7bIXtiyWoOigHufYYGy5kIHxJoF
/6ok/sq3qw70SpKVJVubTnsVHnCZMgzVuR56e6TCLHriR/FOlUSxNdB84Hh6Yha6UdkWWS0JKhIz
Yuqm+0uSbzMmkvlTsJWNKBssJYnhNvHzfhUtrO169YI/2/fgcThWce8f7ekamw2gqvijSf/eB4AQ
J5wsuG3NdRRO309kur12QVSEVyUmgC42O2Hs8MPrNd7jab2aKWlU5IrEHe6qHhBxKY+HA+Juey15
wT4kcDZxaFh0+Ul+XNC0wpsDoITBsEvOG6err5voisU0i0hQhE8x0aH3/0VwnKCGHV2paL8lMhGk
Yca0t6EUv+tim9ZjRXyLnLWFLtRE8yAdRHwZM8kycmqGz5ca+vnAJ3pA39CrAtHy6TixxxYc1yzW
4Bm4H+2rm0h9s1XlMTPDy31URPgTJkUIsmmmRUKPwnBm7dxA2YMH6R8YyPu39ohSxZLIcfCiquQS
yVGzx0z9WsQd/DmW4TaNtTJMxONXg5XdbqvkWqIxqeQLmaBFU+qpad6Kds+lZRJfCucAr4Gua1J3
papYctnirKQm91G9vb4AmygGr5AedSxD2v74zG/8QvcnDe0VzdkUdWE08wdLKm0OgFFNMbpkJ+gs
PK90DuE1TchyK78HM62lkfaCBA7MJNhxH8pgX5JqHMMLHORBmolFBIOvLxgraO4voZjDgcVhE4pS
uQKggCRulReU1MRmEw7AUpwn9NK2OHXlxh40ZS3KUmxvzg8cI/cjNaVhhQHhqyYDWwm2a3hja+mM
8Q7XmQ8H/Po74sK5/zE6KGNpP19Kkoy1b6hrvSXxUsVjBKjCxO6leVELhc8k6LA+TUN35H52smju
QI6M5y0+tAiuWXV6OsM7nHMxAdcT8FcKEu6j4m1k41N55+tadIQQ1FahbkiUxBoAmiD6zt254lWv
V1qhOXKmg+t+I+r6rPxXelSornuBHWiDfi2lme0ju7ARu6IjWg3Nh2PjmTRoCOlVz5zFxVovXvFM
B1a3C6s54HIaqPaVPpj3k0ffsQmzNxj5y5Qqsmb4B61Qp71nSfeyDJlUh63p2Cd8uPIJ/HHMqUaE
HtZqG2e7dcS0yefDG+zroPo0R8HLGaLgwaKIQNGJsx8J716byxCYP17bkzWdBSVsAnlouDKNTr9d
5SpBA0Ixew+srmPpC5e6qUxmyYCPwQIMuWWbn1gZmmupttPiTZgkIiBGRjh+UfOgizlZ5oQcZT7y
1f0/YZLVl+JMJSsgLFvWjQNbExRnNduUzj6X6ltyhZHaTgcL+97MuBl0WK983CFP4E9s/91v8g/d
Tskb+nB8mvg9IstKUl7IlyLQGOwh2Fyz98gfhXAqPm60xCw45ca6JEhVIREkQcabZP9f8XRn7Uhl
9V69/5Tqq8LswX3kkZxnnYLtYSjWGUCg6w5NROYkG8/G/j8iybyc23OfevXge3dVZS2rfowT4zxF
FivLdiyNJ1BinD8repeonsaiSSZ+IWkQd5DK+kojgJ7u4IMUIK1XpXriCB1GLOKwsqsjYEBKCmVw
JVB/KT7RKfpJp/BPeXTKMyvPZKlThoxdFv7FJDpzQNz//JxH8S81yXyZKKe+V3wey7jbHpK8S1Fb
jt7CPExvDTd5O660o1GB6ZC4wcVuhrRBAfQPL7geMeWalaJ3SEhbU6dY/JW+ViD0hF9zU5hwA6YE
Pcob8adNj6wyHEnW9XD9Uh6v9y4koykBVKl8wxZjUlUpfUmqOLJ9ytMcwMLgDNjDjFJHfrz8UCFc
EoMVvEeLCIBE0BECo07HjeonlNkp8D7xH/G9SI/l6bZ7Pm7fXs5fsJ9DGnqYPiSQCfqY+hEMfkgz
U+fQ+VnzqCzDhetwLGa6zu+/cSV4lb8O1sdFT7Yv18OmEcUfuAiTbfOzjowK2Q3ITdABRREqKsFJ
9/DLd62/bBMxu/NCZ6wpSRS+Xen01ZQA8lZoqvNtDDHHcGyu77Ptt8bXpy99+26DzZ6cgas12tkk
jPyp3W+z1YlJ4/0wrqu/9mVohCGFwsnbDdY2bg02e2jw2BHlQWaV3PYUIE9Oy067vF/Y+1oBB5Ux
jK0vFCJ+H9ctMxFesV9+FjW29N+vTojfVpnMq1G8e4MdLHtCEvdPR3uqVFquPXyGEEjDM7Gc9VMV
9EMx4WRBIRui75CmwwQotuBYApLBQ9W0MqNQkkZ+oSL+NhD685yPQS3D5t2xoECKJYOZanOIbOn6
8bNU04+GPIWEvcf4ArlGBdXJ7wNRNrRmkladkitl6USHeepNI2cnQWOwHSA5rq6UELq7J34Xupfg
+5Ky/A8ysrWGOQHt6TdkTMocqxaGZpHt06lePErjvyznwfqOatmIQ2DxZCqgIy86NY7rJYG0Uc0o
rFUMsG1t9LRlp3ysyP022QAVSuvFPm+hF16k1R6yk7OJJpb37k/eTdPrXj1RfJQ8DnxSD++2yi2g
gR7r9kKbsLWFEFOF1MBI79IYpEmQdJjdJQaJLIL8nBiAUZaAnGAlX157BOSOjuuoI5tYdrVccoC/
gDTOn4RLCSFWmOaoRZBwLb4kyuVv1KtbA9FLd55w5LDGB6ZyFc7ApGD3zxNg/L9deytrA6D4PgGO
e81wUTwXXIUvWG2uoaMFCUFuo1wtwq74s2PTOC9cSmE7nngD1sQV/b4qJgp//ILJ//SZLEhwKzol
qXHf32DQDpStYZK8XfibCUhNi9r0H5AWz1Su4J/ITmJ5KBssENX3Tq4Ggarnzp9HyAmmBZgLxNsK
HVLNQGQjs0M2CqUF+i9oQoVT4CnblgOSpM+gEB5hs19j1Bs4cWFL/f6s4ndxEVxPzqvkG4cNAWmJ
yeDZ5pYRjMUR6hqqd/HuhzvaWsZS7JU7t8DriJffw/berdFLKb6UakoiTUIPg5mVgAZvtYUZ1vsK
BhBLOGynzs4N4BCUoGLdqiOkdl9fVviSUC/a0nWOZB8oM/xVDmFxLCxZyDRGEW4DaFe4M1Ddr+E5
BU0v/Ql+Jp4unnmm4d4Ww+CVFccxEtcIrD1AqniP1cdrNV+1tBEDNaAfST+fGbBh9AdiGtGq2Uqz
w8wa00FLpsy14AmcBmpBVY8SBesueI/HtevfjXmFN5WzsOrPpaGawIKEGFNASttfW0YFv474PYc7
PWafPYyNqQkkzLlM3JaE85lasGJLDHZsTMgZEeMBcS232KU0Fo0uvZbLq+G1272eYPx0imJvENop
hEq63g0peGPKTnIgcf0N2Pz8LgOi2zNufIu6FS6efOpNsjl4tE25Ik7RcSMhLVzVEdi1yhe9oyHu
a9qycGUhSPZ/UO0pBaA4n2KCPeSVITJAGDv6nh97xDZ+GdffU9m1Wa/E2tibpXDePM4Mfck9+wDQ
7KhvDOnOLqyfh473G6QrfTa7+PIMMUHTDx/IMCX83BQGEBFMpzTE6vcwX+Oi8iaF6dlzufQJXC2b
1e0VHmgiwiG2eKmUMtB+JZabv3I53HbeQJmvlau1srSR3fwOasO6RKvSsnVURIdd2863AWcWcSVQ
fuE3i/R3yVqLRxR+BXegOuQqwhlhSPSb6xjuVEFyYuQXUrhYGblc/1WX873gblVzis6bhsAYv7gX
d/vadRrxknOGkI0HpqcUp6DfdXBcvnTBDFwv+LJLBG7ZVMNSGbrUwmohL0Hr7hYqWjyxHpkE7VN9
Z32BXADRDc0q9mee8Ir2zwBgVgvVMqV/UYA9+J8HfbG5o7B5YARWILGaDgBfoGJYY1dWy5VKePK9
RUjJIHF1CdKyT32ezcsRBZWbTENYF8sxrh5iCf3ZKWUgIFZMAL2iJPiDcY3G9Y6KOpbVRcGe6kGn
i4NjUS/XniXO33XrajNJAmUNTbxDbTwX9mYP1GEjihyozcJ58ahPdbXCdWbhI9i4Qot1dk92ezqR
cfwQASJFKfDHOlmq4ivolB1o6MGxXBnonDRoaa+POhAhcF3h1TDKTdsUksnCskKRGxOyTM7zNTtP
//gRxJpBV3N6ytr/6mPsHziwRgQXTYQirAsZSLRkOVom22LVZsOQQTkxWPw6fJ6n0l8KGgBP27xt
kGFngRAFn5sTTqCHoxkFTd1ijxAJGuk99MbSbDM7Ad/sTX+znxu33+wo0My4AoPkDTBWaILnlCw2
FL1po2ldK6xAwx3fOSh75NYy2mFBv0aeZR2aCZOrHDT74DQLolj0xUOl8kT9w7jbQZTk1XAsonV0
frq+RcHNIXmAM00clhFR8dvBQMqAY9o2kbLaV/LCSmfOU2m+uFql9fONCQMQIeOP7YTd/5NBnsAO
w8gCI7fqSDeMiNA8Rb4jTqD5KQp5XkLf6ygV4WheKCSkymZBldkRJ3WlnLx0+ivH/DYyZD3j1KFq
gUxBn7vci2iS7AsboMYl1wfv/cA06X9e/WCtzL4Gt3ZA2Qnv/RsKzk793AN0Wo5rz9EkvUFLbhxG
ZLFvOcYjJeTKU+hJh7G8Bqr5ipvSHT2O2e7Make7ydqcQWDt9cJp0oiYxTpUXF5vPIadFrke8n3Z
AiUlkgge7jL3DwShZE9EEIVm+dAvq6mYfp85nopmiJ6UCa8uGko++6n1hr6zhZNA7syv5Y+0f/j1
DjUsNAaMIBy+0kXDZSUfjnQ749QIo9Dqn2wIpk99PtkXGu+ugPgSkQuO7xlRi6ebUqAh8oAawGhX
tEhTrDH+oOSpy02EGqKNj0ZUtHfSADxOIRPs5X8+LRzq3LkKkR33/zLd2sFdki43t+WOno92D4UI
gE4Mx9NBOwI8W2e7Bsdd4cqahMIvuatqOMpH2BDMiuHRuV0GslpwlSs8w4WL8Nr3+pTsTab2R1zp
p83D36PpYyEVX6CdhTZNC+h8vBJnVVzuJbVqNVlyMfowgZUzcB7E2RsohTas23GGw7tvRqmZdpoP
ug8HtgtPAd1eVjw6Xa1azDbPqCkBC9BeK4FKWUQvxOio8HrH0E4ldeh5oGp2HWOonF/WF4vc8rwi
hd7jVnyawrGJB+veUmvh/VL4T/dhwC9UeakoGeTrVgGgYRMVXaMtor9UU3TKmR64GDqUWtsmTmJv
dCukMd3PyTNMwJ9c+/pwwjmBFmvlQzQ3AwrSt1tjFgU6kgRsh11np+dl9WVLHmPHxtnd+JzMmY1L
vbmVWhUWJ7yaBD1KRcbSCCPRuGjVuNHy+RTEDVz7N26/z84rSVcwk9ebaQv3Dc5CwxOMX+3TyO0U
b7gns+uYMMxNUHE2HOF/h/7wqYyMV7uog3fDGcJbZ85URKLMdQViIBMEA/qAUwOIcUcsY/JU01q2
YVBNuBDLFuwMDe7Uxbzxitu5Jhnv1Ot7wcnCdFb4eMAry6k3PW2uYHHKpfe4q04Gk3K3VtOVEhXx
rdpT+BANPFXUJLzwVyfpsDazDTca4CnJOcwONgPKAEYAL4KcVElGQThEadehwv8pmJbKA0QLnaya
LrkBk+6EcWp9GDB/Lfu5FOTzQ/yNBbVk3Ao4nyw4/ZG/jgTi6KAk/pagnZtnWQM7dfX3MwgAV07Z
lgMTKifzlftXxMCJIiMBnQsZSisiqqm1vQUIyOLYqUQwPsrB+Nf4kEorQUh7fBp6gX3tm0giJIhC
bkrdrAERW3Oy01nlB2T9azMndcW69DomGZfYtPA3VqequtdW7CPxBgbsgRReOlBU5KyOo7ex0ZQz
x3uvZ85Av5esyLQODcUXuXOBXMCwZUlI7Df5BsifiQfDRNH8Pt7NkmHlQ3p2Pd7+R+IsWdYl9Q2r
NPE/5MbEnl6mcAx8KjC7cQylf6qQ8oTi0VLtNH10EtZRmZ/ncGNxPjlUcDSyV8aG8ZRNr0Fyxy8j
+yzH4sfLW7CDfxxM6Elqtm2rzIjD5guU7W7fWsNjmiKMPLlmjMDCHVNsRRTAVkLAeMHbehiU2Fdx
xCkc9couRI7cyXbVUkDowvxu8RzZtdllwPj1jLs8WJzwc48XIDJoMvvTE5IeHloz1lUHr+oRivOg
ynEOHXXdFOQq5otARRvqvvGc+ntTL9+INTz148rZU7PRbegx5GjgzZXBxeeIMxmFR9M3+cbfKqGk
wluDQE7YlXu1KTIUvKbLwpsyT7bCzEpi8sSkM+K3Wjvx2HFmNOfH9vKW99jolP8K9LKpO+6htJvm
+5SCYNYf2SggQMuPBIgUPAIGHefuCrSV55VRNNHAsy/PXhCrH8n82zmLyBI9SUvadbvh3VEWZYGq
/ESUiCuSCplTE12HcUV/mssS5g/vByHZ7XLyYNOLGtlKbGOaE3rUaHIdokpFKkLivFWT9Ml89Xlu
IvrpKwty1bydPunn4L8aOT0J4E9FacT0e/4jOFCI7soEj4ZS1KTnufK+JlLwizsPDDoR0yDtZI0S
uNGqc2HjMkAKnCn9yWJxbWa6S4TkhlkLXFlyse0IgDCoki1CJZSFuMtW/CITzaxrTUk3CKsaojkv
R3PyBx8MSubcJ87WRWzpE1Vseq0Sxi4wZ3dKkMACC7tdc+EpE0UyMDCjSzuE5XKXjK7Qid6AYgVv
dB25ov+9l/F/Y5yQqq90wnlddDv/G04x8kIDsTNf9sQ+pG1aX2WMmm66UjpI9HZLxmEc0LBwbi9K
x+kr7ZyQu758iyWwotmuG1QdvC5ai/etRwZyVRJLxrQpSYQ8jubN3s6wy+N9mLuJ61huoRl1JVaH
ijrabfHvE4ftGqofLyy9l7Tw0L7R/9N3JIkkot/HgmM7c4UTQZau9A+AKM6qGZ1qBZRUALHw4E99
KP+xzRWLY1RwCmoK5ynnTXaLDVjyKhs+8HJepczVzjOqsTzkU5b1WcrbP8Nkfr5J9YLN6damQci0
5Q3F+hTazpZ1n+Ohav3jmxpAZlUT+5Q/DKYYRudDVLbqyQ5jKW6JWipbtBcMAO+eci7DlmPZmLpi
qLIOm997BEWFAJuRPSZpmJ+2j5tfbpmxgl2MArRxVddFwi5yXt4LeYbzk9WfqpbhcWansGAFjvd/
VzLrd5idH9AjIvVqT9vZUUcx7h3CNMoVIr6MATYtICvJFiGxDx6wG1V6iwqAdl+zPCkSvDDMZDUD
osSPT3q5DehDvhtZgMU5T/lv8ruer+g6CP0sL8Rp+DGPtcNuQLcohtvDpgrZfQHES1Ull/edm3yD
jgXwK4pi/vBhB022EuWkqYa+LTRt6u6iERJFKMzS3nYfjad/9KDeDbxD4FQiycrY7/V2tY08G0PT
fHLv4yExiebm4eg7Lo1HnRmh98DupZ4pPFbP+hOfIlDt8VDBvb1RIAkB6ZgB4jUEFSg493fCLNP2
zdmTXfcaeIipwTbKqQcxSmIH8iU4OtuB1pbCX/QRNl1ybB85OS654Mkz0pjeD5cnzMz98MhMIxAj
3GGZrXSZvyNkLBfzz03RdNA+zNVoSRwGJFUq3+RWZFutPp6I08UwJFquTUbSKVHkEuQGBDhSqCSy
0XybyL5JtR5fNhtmA4AUuhB3NZY5TcIQ1hklz+e0KBq1mTuxIsta4VZn24+klNAXb2HEUn3qGNRt
w2a8ufXjhdjwMZvD1wZ0SEWHae79uarcCmnR57pn1WUnClCXDUhSEMIgfhjr6vUFinckjBupPwT2
xdIXHO65xDxsO1K5Kou4xhZV7RHQHdxZoAQ1pUa2LNlYcM08XpRNVmY0GeojPv41y7srTnhBATRf
hcXjH3x/El4IaLKZy2oPG5a7JSk8oij46BqgCOi2zEqb7M6BuNh/wiN7W4zBGFNHWr7EWypXmCje
Ji3qykXLIGHKCx6wv6xioqHGIochaxfnbIPNqfX3jitx8x9Rv07b85dAxIlBs87GYD9e8SVzOzX+
0zj+pbW0skcG94VUjzxUXCnI0XULHSk2dmsGHbF0hxYcFZwKKeQ4zr9MAN3L4psREkzRbJPJnLjc
o3gY8hqp5e7Dv6Rsa7X+6mfkFscgvHNFTw8e3P+giU9s4MQnlpQzsqz6Deo/CgG9ib36kmXwLIpD
A+TongWRDqSTi4njK/fI2uuDKxcphqFj4BHf8shfL3J1+eW9c2XLofoocSIt0Dcvk7Vo1pOqU4/c
HrVfafzYbXPbC2vKf1GkEMo++7T0hFaCrWSgA1yQJLqOxCtGy44xSfQ83SOkX0ekTBJ+dRjkHrP6
6z2pqDqZFrfghMWOsSVTLK/1ogNwD5D7WSZx+mmByPYwOXfhMUMOPkGY1VR6a7FWfbM5VzufB+8A
3OwdWA+1sP8nxjkHBHfEY1QiAzQl5MXWZzT80Clb5T3SMjXHQLomPrIQFnpECQxuCi6+CxbZD9k9
dVqZ3MkJJpN+JlU3TxuKsKoV1TQUzApt+WSfOax7YThzL75NVn4SXmpKEq/A6l/6+gzjtFvkJGeD
TbA82QJmXpYAoC/soQsA8MI6T9Yok/2gNCbu5ucFNNA37Tk0aBqHnzjyGIX1v8EwUHTfmLUJyQEr
htv7wxuF/ZP7YEe8P/q322PYoy6IHXq1oypx6peKzJ+F/pK9bNXlUIQI+PirgaQBYJ7nXRhpHvHV
o7eTuNr/pEocnjjKPhdC8Lkuqk1/B5h9EzPhEzL3Vpu6JMyBzkI3LLDMoi8Po8UVQqDd/IvyGutB
p0ZLPS2JUX24uVIVqoEx1bBw8yYYuWDeC0u+r0rc1e0GKsKxVAfbCeoTUdwD0ZoHKsF29xPR+Dtz
G+DjBJKS1+Dr7DNFXuHuHyCFuSgEql5yI73o7L01ivpn+owDXc3fl+p+vOZbAvTqU7ezDDctQVtc
sLFg316QfBGzzkUYS9vGOfnHJx7W/7+DO36NKjMrWhAIRDqHxkxPNCXcRn26+l1KQXsKLxwO1edl
wEUeogcOfyP47WcpHajJ/RBzGKNbsdRJWP3CkEy5g+8ZVLw55UYrmhNDcMwxPnXj6t8IvprY647T
Nxv0j6pHmLR3tuvQIx8Gvzj1gjooYqR/nyE9k/w51VA6xiqfjv589+IRkd5W076GnBODS+OIWAah
iWgEYTLpvw+u568iKB+3/lgd5Z2+RqXf820O2TzS+SmKxC10z2sQe2lBzsGucwniUUgvJByfMc41
aiEhTcyOgak7/FRRNQH1Qi1m0Q878uPTI3DV6bYc3XgkTivQznMl7D+sWJrBrNyQWTvq6N8FwXu+
GXUMxSnKlqMGOQF8a8EW59gphCxEFJMoTc5onKQZ0Pk5LnJ4161jJOyBe8aWIkf5f0CU4/bsQ77r
txMFBbpNKhHh9M7gtp3lB0K1fLIwa57OFNoYsv7PMGV7icqkeDY60LosslvlwCrvba9q2IpghIhI
XIU3zniR1kf272bFpeDNnbjsibovvN2Mpa5SzQwUmBbH+om99LM+8mO9IgUemKTSt5gIdnOW9UfZ
zX6pVrAgRkldfAPGwVX6o01V3YWJFrLLwEwYyb66OR0rX5gfc70WWNugtz3ZVYJ8WmcbCOzS97vv
T/t1Yb7eZkuTIjUfD0AMmNTtwcDN5q/5qR/oQgTN61ng9Ck5qh0vXod5+tH8v7EWY39TQLC1gAK/
prPGFwFY0LTjL8vLiFitk+N7WmYO2YpwtRs4c0pCHtvo8UZm2mu8M6M/AyLUneyRgPYbRda4f+W4
eLjL2nd6g+g5bEMoNz5aLg45xJD0O0c8NxdAIXMRrZO4olj5vUfwnNMlx12neE8A975IhNKYDTXS
Mnd08nhL92SqWLhZE+03qThku8wSqrOKNz9Y2q3qlu5VdZseXH0dzrH2El75gsORTc7aYf8cr3dc
77p9/DAEkuWrufQbXTmP7x+obDAFIf5kz/lndlklIqTzFxz0PWDRL4fu+8eYKutWwzjRRF6pUEn/
IQQX9BqYkEa+bYnW6Ui4LZhujAWkxbNAbrDtxXRzjQaAmOof2whJUmS5xQ7PnVNAz3ZWOG8oxLEb
S1XnZ8xHEllXN13tLgDS4OnmyQars3KuMO/Zqi8atB51kWemc/4YvSSwHWGSEMt/2kBOxN/AY6Qa
BaRhrdXYc+VGig+O8hn39idtF1AOM/St6JzwLIFv2H6cbsOFQXh0+QwqXIznyvUZJa+jEnoLF+SL
T5FzBaCGJY2IGFIwp+C74I8Br+6WBas9tk+x1RGmP4xfsxkBGg0kLMCYOz6QGsOcfzcUzfNVuii4
Bappajx5O8Ge4/AaSyuelLMzmTrMApfhznrcN+EL9dVWfRPG7Wigv4HzrJC62qA1vpUSlI7E14ou
AXaatfNOOIKFoSs2rJgTnbBQiwhq0B13/y6GwPTA3zQD7BvO1UZFUFcvrZuPkfS09W1f2kf5tzJz
eZ13h4GWZxXgVRs/1rYyQUI1XHHHLggwAcONqzlvIobcgv3zWRDAcFs4aeaqlScg4CySrxPMn6W4
rYySg/OTDbBRCJj/q/8DNGd/o8EsXTmakH5v5yFdXA2ngUYVikpRYHYbLgnynSX290c2v5nnA8NL
tYPOJJWmN0/62v/azR2kdmXy1nmq6ff0wV5aMUnmBT24gUXMjOyg8mr1DtdGbIvQn1l62BP5OzXK
xn2WCBAut/aBsu7HOFz2XZ7T/ZQqAnT77jK7yT1/U+hwDGRhecY8QrhisXiLRLwV1o9OWUOyOp23
DRY6O+Mjo6v+UMD6AVnnTaf0YWQOItLo1uEuf+7Hm4CfwyM2u7d6KCFlSv3+tCK3szr3FfPpfOOx
pTn3dbxMjTmWanxldFyur4kO8kYVHkUeG+KQ9GJ0qNgv+PhBlXmdaoLX0mXmOhSgVMr2HtZmEhOd
26Bag0C1BuGCAKwnbl3wnvyQrm2ovVn242sqVbUpPZXaqxUZ533qO8fgvaiiYTisfNQnT5PD40Db
L1Q/kE31TZmnbGJwp8sHTOIGhZaXOVgPKPiVPZv3KrIMP1oDwu43EEB07b3jUijqSBjNEPKcSnW1
AJYaSHSp/RSg5vxLBag6k0FczUkrNPPI6+anLpEyONIPZw1UyYdRCix0ZlUZPp6nvoJJjIjsWnYD
k24L/m5Z0EPtFHi4VzKLeXmK4duaEQCAG6rBhhsia2ANl3xlIRZNsACwh1jTunrblrxEtpGfVeor
n6CCy5SxnGY4mMVlv9+L1jlBP5dKG8VmFGKm53f2ZcQ9Q3Mvl7ZvXQrdjr9LobB1vMctBYzG+EJM
DAxWnoo7t6jqzL6jgMPJTKW3VdD3q+E88eWgfa8rGpO9RC3e8WUbmvC1zKL7oSS5nhGNwq5m4bt5
INjak+tB5eWmPvbRS957dlqHTRurGotey0uaaBEBRU8fv0dpm9ajyLJwkjmXjs+iXDCO7Fq2vpbe
DGXdRi4n7Tq0KR7FnRwikgR49JmjT5JTtAvjd0gav3iGEMVaQsdXaMxv1wgYYqbnRnB+triyPVkW
Mzb/9IxakrcTdvUojE/o3rJx+fBP4ovxZRPjTcbph3jziyOzgpz7AEkgw+YuYYdZ7ZtPmWaf2pZ+
snb6DvxOLPm2DNoFa+sbhtTEwxiBRxIHvQf+Xxbz2YQdnVVJNxv7X4uF/Wk3d6Wt2f1TcFsw5BZY
gT3Z9y37yEbklNGbsdRJTakQgVicfkkV6vQ52ZpQWdbyj3HgYQNhXrnotXlX0RJU1C8nzn1n34qx
kHQXHdHu0dl3AizGyZ5iPDC5ShQbOYXWWIzpK66f5l8JES8FkQCUlpjo8B2HRWDUDFhgQeIkKgnp
tLIDjKCEatVxQjH8rb45MRw+R/zB64/Gsuu3aJzyaYAOIfXIUwrR1/Oo8K3lPYrnTnHTsFhHpHNB
kEFhfRO/C7cxbCoawmpJQ3sUIdI0vx8XzgDQO+Z68UzeyVTJsMjRRYzJgKDk3EBQvIk6kj9owIHo
XTCkBIJHg7GHAnLH/Y5VP6YwTuHijlIYcGK21YUVNjkmyKj0qKMH+vh1dHStzBJA6JfvGPzRHTYh
DjoEAeDdTapnlCPLYqXL0TqEi30WfWIAWhr7lRHyuNPRczOTl8Ih664V6eCrGGSv5hUPf5aLSlrf
qkLhWl6O2MMjsD0gaBl8gKGBhg4e7XUtqP/F7UQpm/xwgxGIeKenA350fll7ZTHthXcTfmvxlhQU
eq6GdcwEpW6VRUBCegavUyv4qQNsk160lXVfA6pt+VmIZJRTWmbCJHYLR0ialzKpTrlXm/UE/Znu
Rvg7VERgHRIjBwzQqQOsyhD5k4LnOi8n7QD3b3z+HY1WGJtljbblWfr1WYYIQYn7XeEh9m0hU9fW
dxlT6Hh6V5LOBf3U3tUHF7frYMo+mrRwrQoACtByuU6Om1kn0BLKjvu6hfoHpqio8MhiWfFwEsHC
GF9kpxwvjeVAFoohAxbb1YBjdEvFxIssgFGCu6pvv5XIr3JhGDOMfTE3EIvJlaPs6cJYjd2wcV41
XjQ+09azXiXQV45lLpyM5BtrENTDq4mhGU70raIRfPE+fcZagHqgK+9jFxFOB5Xw6b0LKmFa1jAu
AykJUyVRZvg0cwAHpul4iXQuWMJK5N4jB5aYZfck+BUIAsYhfl+Sr/MbmZOJGC84iLnX5RgXC59J
vKql1HvOHFHORuYyCRAtKYEV3l/QoI63LkdCAVo1X7lonzo935ptTLzLhgqtTllZbZ4W/kN+Hsic
/PWk/dfmtXypPWAZ+hX0NanSYzEyeijK/cK1PF8dW0+1L/0P+UjZWMN4w3E28lejcNi4c5Revlmv
ZBrFkocZWS/csiWHI1IXL8F1Y0HI9AAsYoCg4y8TmKJL3GLmbEzhulGjwY8kDyrFKHEr6t0Prv45
fpCrvYaBY2QL5I98ScCckm7wX+IIhdxauPXhCHz6ARdDa4HTL6s+P+kGGH3HAsF+1BfpWYve3JF3
0JZ7nVo5lcV+PsgbOXKbgczjMULaY9M9TeNSAH/f89iIZbOMtHilMGAC/kmgHu+ZXuINW4D6Kahi
KMrp/QNHtpNDXconLDPqS70MhCSDQxIxqJJrqA5A638unbpm+aCG84H/6E1apOV3lGL3qT4PIjbD
qsRuOKKZELx16Hq/Tw7iSA7JVgNygXaNVMmEFeWjavRkKeriKxviETCbEntc3AqpEf0SGxUaExX2
KGcrTMN0cd4oUu/7sI6c3qAyvW1NGbj1JEG4+0tuyqqO99Xps38MPClnMEthhzd+Oi6qmvyxXgxj
uKvKuCQVz3W+mV5M1A1QF/h8+FLu78qWqXFUetRiVylmmozxvZZs+2Nz/NBBye8vZZK3kHAyN8cT
+7o7XeZnSXFa92Gwn7HCtKyojyX6wkjiu5/NlLJEqdO/qcJZyz0UdF8ChGN3GDqK8Ee9h39ht747
BEj9PdHIIl4Lt4i5yEcKVQnsHDr2pm/B+keliIHXw//Y7VltwNe8sXGT5Lg19CWbuQMUMarCswUv
I6Gj8KpywvV2BMLJRhn/Pr7Xp7YCiqJ/fi7M7GETbhRcvk5lc5HlWCpQqZs3s15AAqSZgaJYp6zA
EfKh7ZS+Gof+91SFS5FYWR4F7V2u9WASs08mwzpF8/2eu9htvgef4jdiWTl4m9HabGezEfTB4XJW
VM3QEmj/S94SLJO1b/1t+Wr56jXaDzy8MjfTC2eV8yNowq469FMDjAQidGa7o6E7P55K3ixbCnp7
DcP8UaGEBgKDdbSXQehl1zrkBfAntUlW/KfOrhNeXgycUe/kagRApAlHbQD+jLa79r5ljVRmobIl
Oy8/lwfUedSqx6/jjdpQjaIC9agtdycLypESMCH7xEHI1qI2DYKOUiqmAN1C6h4jTBSY9vg2PlGr
3mqnoQNptMcRSHGMsRUELgoqZZJKU6Ce7I7DxTh93Kd/7R1K4sI8pFEmHKXP0y6kCWWbu9lGI1o1
M2s3NQotS3xLHQq7aL3GJhstrysaoEKgRDSrSPBBlUBKuy5RL0GruXxoc6IvyJL3J7awEBEZkHIg
sL2iDIY5WWjaApQAg68Uots5uu4Yxe4gWcSpw1houoFYsq2NntAhzpszrpQyswCfH6pZAyvoac6A
XcITVNJ+9WncXlOasSHmy6+YvVxxI03Z6A6lbwmrk/bA8oC4QbTzj2B0W2caMVMMGk0SZhu+UfFL
mvgNXwVkwts57kcwVrbqVmLvI/6HF308I6SplyJFSi+TA4TBU8zk0m6QlCTreHbCEJcZm0nud3p9
JcL8lQh7CNupHwmOm6/Y+a6bIXWhTPTF4s54YSTMM3DAQB4bk8Pjhkg64Y50orCyfa1xBKDIm/xL
KYyjwxpnbU9Iu7ANPhhKN/OurTY3T0C+9pwlSZDR/X5Dt8sUsFyZ8O/rnDgIXagG9PFMar/oqkbQ
4asS1ZcnVTnkCp5iTnlNiL3ablkCs5Uqi21xs0rvNI8Om1R02CwPERWYWOlptIlUsvaSx+KDR8yE
2JTrro4TcLAaSrecnJXeYDJDmXHZ9mbyp57iaJjVFpWqD16+HgSHQIUmviKg+n/EWsHHeMaYdXfu
pr0a5e8JQVHbnoICLVc4Zx0NKgzM33a8+xULpBaprReksWowrcREh9VWpXUlkuLHilhMNrcm3H8R
XQwgx8jjZ+Ix969kxKQAzItVJw3thiN4b+yOj6LdakbPSK1u/TChRvjrjFIYjICiEIV51x9Z7Y9N
xEHrP7pq1CXDvbKwnOYpSxGgny06eGX1MwWO13oXKe6vik5bRCpkrQT/sIycjyNLVD79zLZGPada
bIHP7ki/Uy7BNDMUK9sPg6PAsbnU8I6Q4RHGVnLzn54tRMTosGv9XhU/lbyqBBk78oWGmQDJWz1O
kg/qCiu8FJoYETAp2jiIl6pU4J+urAbO4ibTuD8T2jXxlgeKQ+6EZScwvd6H6G5l5+oO6h7Rl1dl
q+n8Lk5fF7wYE6Z40dRhCLyGHjdQ79AFdxVCPw2MNCTW2yJCwYJxkzniaqdOshZC1d3b6YqkD7yH
WSly8t8hlxzyZi4Gt7k1gWbMZeUqagSwDAG6TxmzKlS/kDPh1Qq/2vhTw7bfdBLPzzlRNtfHVGGL
D+T5qQnVyHhu9HTTltbCIYZ6ohuTGxrQQPSCvLylAwSlSztPeT60X88x6HDC04N/hEEl8Bge8eXt
DD09SoEFme5jFLfzIPd9Eqrk8kaY/dVloD1/Qe+bimNQBVdLaWIgKMTY5IY6D9yUJjmklrMqMjEE
YkFrHmPg5+zKE0CQyCvx53JVOK0xIlvM6i5nEPGCnvGESx9FdhznO6sWP/XLO5hmrueWVVMXOK2B
PITbcN7e5AQB/SmRan1Ipls4QoSENlZB01V2UM4LY27WIKOjZZ0ANvBm3znS+Q1B81U8hcXuM7hR
ZaieFf+VF5BaO5iD0m3huT5EvfsDbVJ5Ta5IA6g9P/HqO5WRqXa1m+46TEL9CK12Pw0DRhr/0QVi
FdP/WxZZ/AIuqyq3NNSw12lPt3Jnk5BSz+awbX+G9KO7UMjsV+EZc5/OHKNCzR+/fJT4WHw3x0Ua
pNAWRANpSwsSD6RH6BIzRePwhuTrn3QuEXbS3yQ3oRLAZkTYWr+YoJ4e1lphJ7fKlBowRxXYT7YG
CdoLvm/CwMe9QRf3ONUuhOfU00ZtOxQdYa/NczxQpzaW2UOHQO79IaPDOBJJrOKdWA9sMxzD9kvK
WNv5xlNBZeAHZbTXoSTxdbXRyqMsyjBb5qD1K4iozacyucD4MvR8t2tde6GHbszWxXlYpBZCOlPN
GAETfxE1gyI4D++Rv0DAdAwjLnwq0enDmazjhLJjUGA3QdKkWQElJ6hdv3q3QB3Fps53oJ4gYgB5
PG0l31zndJM7Zlpcm69BQ6m6g+KPrvfRXWDN0FzWWqdF71/gYnvj7E31AKg5d5bUT9bpcCGxU5ZW
Mw7g2S9Kxwc/xnSov3Bv12JpMdz1hW8Sp0Qtr8HvbejhKubZEj+29eryVhGrzre7/ByX63i1oMVC
wTeocpPrphQane0H8/iegeoour2HXl/am2pBx/88EdAMyAiSfVLKRe7vj0vwWRt3ykYRnZTRYO41
Urb7cKAXki8X9GnIHVw+HHKviGYP59Cnk1g20BYF9swGc+gZFvLuBnezoUAkzlhE/uQ3diyMQMnV
dGW+cwvTpRnCoVhuqTt/O8ImuDBPHNCdrfl7DLicB2+zpZekR0dpB4fe4LXd/XGG6UZ6lX1cNVYA
+g2P+AbzobMUDRyjVOp9oruct0fMsca+Qaw5mOY2viiQzRRQtWpJmaE/evJK1d0YKirBWKhAX85S
+Hp+YqMdnaGVbM2bDRJ2Px4XwQ+DPQy0drMy+dT1ajLQeurP9ar4d1K0mHSe9O29FwJ7syA8I8zM
KYPwUCkk2VQ1wxqg+sn2TTpaiGdc74K+8/3mWlH8Td1tZ0h2zcqcKa/PNWYb8jgba+MLwiU+l1xI
dhmXy+Ykw6wOJvyyJ+lpAQS+HcQE5XIgLzDpTXUovA9i1HYLs4eTKjOJBD/nc9F6QWjfHfm6j0q8
dJwTs8ug9ifG7VS5el0g6FnIE6P5uRl0Ra0G7m9pN3HiFVGwCo1Mm7HjtTuInuMNaEEzB68njulN
6gehsDiG9cOs8pJvQCvWG9jEn9Kh1TWG8Zv9SHl+v75a7Fn2XEQDzChidKgF/TjL4UEMeK1Oi2Ge
7FfU+ixnwVYCZEN/Y2yTQzRbkY4z6V1zle5gcqYsYNt7OFeULiB92cte7dxaJhAXOKbR2x2F1XKQ
koQZ7cdh/hzUfEu66vNZ73wz9QEq+JXn6oKDwkwmEQiLuC79SSolesP/Nzvj3wcrV3aKcyDzJKg5
ReFBbtEhuaAjy0h//UUZ2w8CiAhRDlQcDpbDErfUdn6cg1QKygYKMIb5zgVKHtjkEPa6CC6Mt+Qn
Ec6prbRFUj+Y1fVVqzyM36lxcD1AKvaLgZ9koAJT4iqtHiueinlhzJnNBnM5XFsmXKQEYZG6V61L
4B3uszDgPhZA4YPlPVbQIo3SEntb0K5QbPIBr6alUefXOvtqMNOX0sjk5XMp0BK9umNeZSgS086n
wORtlTSNco2R8Kl9R72HItTLY1npC6zAxyazLltnz/g9ywg8f7cg90Ku9kS95thkfUcVQkIGyBYD
ECpvALrylBUltdesthg1ciE7mskQDNSfdReacZbXaROaKHNa2veTvFb9+pPdR0YrZMWlsnTgvbbi
irBi/nwZIYspNl6WeTde83YJQHTsDRxp57AMhTM9uYzo+8/xxnDY6R3RRFSyzk8j+kR0U/EhRUW6
tOV2j5ErkdZhmTpzNzZ13pWhj8S9apJf9oOmkPPjSgzXKjpJifHDXd+rY+dp0E1lQxo6hOhMFSmN
uFwrnGmpfFyWOWqPdGRySQijWXRHpCrQwNPLIdDWnsYF1GZ0RjXRRWX7FLYJP0MLsv4ZDt7e2ACq
pW7Eqw+jis+w/zK3f7wUy/waMd9zOHoiJNxU4JYOZy8+mZATjwbI3JL/tYTlNRVTDqcyUNUWpopo
o1J7WIPmel2dDHvDbq5rS2e2iPGiPV4IDCoMR819iYt3X59TNTSOglzlfs3Hjs49/dcHcZK4zz/m
IjMj3JYWzVhRYoSgPB9kShXfh/+yIZd41QYuSmyH5Nq3w2U5jCVIh77n/hYtS4BuIbZhhKv6O2Rf
F6++6K1vQ6BoSIYnDhNwkCBDA92fFC5KiOBcGEyNd0kRhzzYdzirKjv9ZKfeYDfQmYdQqLMX/u3v
5tc/xOOy9+FMIuGT6PdIM9xn+rQzLLziXN32T7oGWzkeVt1lrZd/MhfgZwPe3Q7trCwu8FkAZ2RH
Z4zy/uhYUg6w6dfp3ew1hjDqqwayonPfqpEHkBhqoJ4vog0KRwIAYO2d1AgYTRx6pslNGA5b6wvX
E4Jc/SkMRasOHWbFWLbLX/DyE2a+PtM/UuoFCUVHr0j70cRokw3ubxOAh9gpUqs3a0BY1F8FLhbr
Brn7jgsLtmnUl/nBcr9vwk2Jtc3Vh5bH1I3Xmlt4y0s/BnBYZI+sZYV7Nfqu/aT6HeY34agWByd3
rkC6Q3WS2kb4OULsuwH2dsqfFIg8KEpv0V2bMo4lN2WaCr3KAkz5dh2LruIxrsrmQ8jEl+ed5ta9
dTBr4KQwpy3upHzqq4pGxXJEJ/RxQoUjb++zsU/u0z8cmwtmGcxaJq6g0AXIU1Jro3I6XZt2wOJj
OYUiYDocrX/Gh5Zy61ofUnK2hlygxJH4udnWiKdpntGEjxWJ5RK4FJ12JmCAVE6i7T6wVMfsFi7G
wBKTzMScdHpi1/LZAqtFO4qzn9EPVNx6iSXZQ93fjBPwcz2C6Fm0FDe6GnMXXaV08dhjv3kXwg+a
otHSBpLTKByJVSmnCdR5lwT5Z4qr2PNP2LyjDx48zqsSNvgzbNkCV6/P0mTmjDiJtKNNYaDd083N
poulnwpVAxiI8ye47EM/u56+qI2RJdLmCea7URJaYmiRFYAly/PI9nM1vAVzkruKewAcUa75WejD
dt6pix7jv32AozNzJE852SkTOMQhjQ9OXjxU434H+tJJMcGrv+ml2XOQCZvWBspetGWLbOJBydZG
vGQ2cEAIFtaETjLH7UA5KpBevW/5uYH03mZoI/vJzbQN0An1cvmf/unlr7moBwvhJZDDm8rQ44pR
8u8WILOLE6P8usaywXCl/od2PQhP4g90RhoBVU/0ba47uUT4dhkqQN0W8wHlGospAaA3Y3+8ESLH
16sMtdeTMR0qgFkUd0kCvhnNd+IJ+Ew7WSvAEC7mg1H7LgGHey5cLwVjGLc1govPdFprLTi1G3fr
Z4cC3cMKovmwBjC+2dQIW4xnnvFNvhbCLN3dY00xuq62HTkyfKwGZ/ybOIr+geQRCFQBssfVx5KO
v8BykqBI6hzgbx/3Cs3CuuKmVt9bUzJ+v0oN1t8tbH78otZ700D533pAuufZwzpD0Nr0ymbs0rA5
srCJnqLwOi8Dwo1NcmCV9XnY/6+xkb/6xetr0AAsEG8qzyXwppQW1L4NJsBeywHYtWDRxcxoGtS8
wN0o6QTrARAVHBPlO+DUtL2mIzdaAMUJNleLiAR44MGY9iHttjmUPkC8HvYNbe5RXGuOK/lZnca1
AgpmFaaTG5KGcV9xkrYt0X9h2vXIvNDdzg/YE5NKI8deFQzWirOrTQAD4Byxc7YmO0sUo14ZHtUE
siVj6MEcntLVB8g4h5PnBN8YEBtPrpfzIatmlwlSdyCcMWxhPtqCzqZc9ZRRcgrs3uTFA/v0zZli
rTd8CB2UUeyRdiP8n1EBI8bs+TU7OKz5aUTb30wnoFpNMyzDp4s7eXmD/tPmsZIdXVmdMFnODDQo
sj5Cpihb+ju/Yye4PZ2Mmnr9Q0HU7wBMjJXLzFkDyio4JmWgXbOG+dU2tWLUwh1KbkQ4kZI7DR3v
76FfLBdpm1uQIpSkOoVBoCqEHDWFxMjUGxSt2T24wyJGOZxDYuwi4CeVAK3N7TTv+nIiPtPW3NVR
B1YsPvSJesEW4KtzCYdALuJe9EVv2G0C5/yB0OChob8ibJao4+xiZFyrx8ZbSBVD5kMVxWG21aXl
FqFKyPAqIx3BIPzVXik22E3WCiUAMdTf5wlejLirmzRBgcWMwn8xGxKH1zMAkGmSNt0/QP7h6Pbb
aXT4TrkuBbc8uetArNVpux7Ri6uTAKyZL3C3nJEGWnPKf/sdjJ4CY9Z5SZNCNLDli93OxKgj6Jtg
/6WJWaoUoRn54NBCVnHaFGhaOrU1kNrvplIzY5CQJYlWaig9nRh8619PilsrI9VecU7wfG2f+DVC
ispNqCLakaYqLEBhE1NWNm/INIhxBOme8hpiFAgkK5CNCHOHg3FOALLYYvCPb2eFhtJvDXFN+GmE
IXSJh1qO/Jlu9dA7DI1llRU2yXLmmGUxtG81WtdlbeXLtrfxdDR9a5rMUdp/U9U+5ODbEGYiBSPt
0pNOu8lagoL42JLv0cCQ3wRMbNTVLgno4f7ADU+xPyfCEXMWxKSwc5bxgbo/YLoj119H3M6poBTJ
TrHnqCyjWJZiP+pgHnfd/Vs3WmW1ZLisQ8ron4oJdnob0vr8Swp0DMuCyTVAPX3FOeOmmablzpRh
E8ddCem+GZjDUwcTjs4PbQ+Hmg5/YuTfUdWT4npVFJIX9f0czI5ZCFh0hZ1AtZlqbOEj2HjkRvpx
uLfW6i1/SeAv6e/3GyOuP2VJkw+OQ1O0ud/mNRjq6ySABwTdvmNF/ARUiYZ1rhDREOisbGz32NDh
iI5mNtygMBrX6nDXf0Xhzu9fnKAF7JyBDAsnAI6Q3sgfrz05tffEB1unTumG9uYOs5bvMRKbzTkL
Mj5rhL7fIhRorXCZrfaFiCkzgxN64tTdr035WLaBn6RJ1P4mzPwiD+4oPSOxZsytgz3jsOj18GeK
eZvAfrsVfGkzeqQF3WTZPbHLjEOSomKb/MwN1AFMhUkGybJOhKlaj5xw3S9sTYn6N3+XHfg0EW7r
Zn4B4RxXct+Lfk0/ya4EFJ+EIjSk/MKp0HW1QFk0WLYBcIjpRMEHGL3cAjhqfH2tTTir/cMH4W4N
y/eopLEDZJUOpVxNmOf/rEA+YWPXqwCScrB9aJ2EvhSJkPH4Iw7W830g0ZdiBlvOmJMP3W4/AON+
vPXZevXkcwAzXGN9yJMWWW04MECasWTE1AiAPovnk+23DLhBnZb2TNX8/4QVB6GhO74Nq3Gwr7Xl
mqggTajVxiFzC+h/Pse/frwFjmDW+AfDIgD/8FN0k9wXFsRcVBExXKy/zMvz3RbmPF8raK3nQ7Lu
UtC7uh0cKnlEMC0460CEkf4m8oV5RMi8hYWv6REes41C8XFsrJWQGC7wY2C2SXl6nXka114sZRvQ
VXyV+QCdmSyTm1XvFwQ21rC7PzL8AgAMAHfDkxfiNj1kZ2ChoFy6qw70CMZserS/CHdPuiuLJ0cB
cqGV8lvf5TjfFsesu+t5CqAarEzuWYi+yCrDA+i551qQVmEpkw4WcP6xlYKEGEzYt+fK9mOborGR
6/5PH50iVP7LwB2ugEVsQ2u+1Id9KDQ9XLoRtgDS/kZ5bvG8L7WrFrTBc6vcLpZ4WUGeU/5N0nf0
cci0XM6SMBhf+5UK7HLBxiQmRYxZH5KzXi3BEWwMIyCKDofgJpBpjN+ewOq1vIUrMQHlUjg0UU/j
f0fBoT63AJiBDrgQOFHq9vYUZfL9Zai9juhwGAsNiUSsrARWVMc/aMeEQuHQU4QwsYU1WEhXPjqG
n4dNnTg3LhnIKvCJaBKQ4b2p1IgyOom8efAaImQpE0+PxkyHYlJ0CrdJ2IuFCxyTNvwJe+tCUobz
jpACc1/29MqsJ3U/DXxZ27TQ6KPe+edjiMTw6ockc9bxzJevYgOUzp1Nto59W57aczApI+xAgHcl
WcBb7F5LRxtG8kJ3m+oztvzQVBr9Nd/mV+fWQDFaX5LZLhR5YgLYq1fEpmhYFTZ03zaDOn5B4h8I
DVEiC4g10Jq4uo6dscZQotI/5ocx01XIIs0or6vszRsNngMl3pCHM68fHCrtrEFHAQD67JWa2E/+
O+1JiMOi8aOr/FJ+fhY7STbi7EhOuOmNnaSlt8RKJmBOaGdtMiuf4xObqiw0u8zFg0q1SizLA57k
qwkd4zVbaygu5/UkOvrt9JDtW1Xn/cf2c6nk5qM7lxbfRHtW9QbZyisQnB0bTfBGqjvPMPyQMuIg
6KEVB1cDRN/E1ASj8ZO9RJ1sC0J462SQT0b0z6XZ29X8Bk68fWxdP55Fk4DJJS21zDh4bEdDQvnX
xPo7DtmTWIo9SjEYzgu3AOTmh+VgTbAyyfotyTT7usatkr4xxDfy/KXQHc3yo2rq0mMoM0KdVqlZ
ErLxZzo96vscnMLTHyHJlSoeVZJbcg2H7l2Z9frW4276Au292IuAXZCNzMAQDVasrld1EeHkgFi6
ae0JILeOwcEVmDhEe7geyu7ogVNC9zWAMtO82p36k1Q3ZbZiapjM+l7x4+s78HuHEbogTJP/eiyB
SCdUUWTw46qfcCbjP6XqU/D3YqDwIAwungYVjKfydv46RerpUTePXpH5gsZ+n36DgW5LgQtHnWn8
9FqINu3tRMFR29W2cIuDbxUO5p5rellazob8Kp8uMliN2fp1tlOCtwp6OV6aE3k88yz4ilHacs+r
ch2lJ6UOboFwvAU2nKlNSi1AiOIFmerNtbthJyWRSqHofDWT1Jsno6/WP3v0p1e6zLEZibeiO1Wq
TOWUzG1VawC/EE2YjO8vOmQ9EnacwSfiqUVYsU0/ujBfEZjoenPo9gJCR2rC51GHOnqXFOjfO/AR
vllHoEXytd6HtoSDEizpqfEX8GETD3EOsCggKoJYapygxwJSjDm4EOPSzepbL2zFLmo+Kedf01Tz
Av/AsnEwD+/7lbAHTT/aLjSh0sXn5mLwnM53tEFSp+TIt+h2eU1i3cVVWH5ZWCziqbjucDLVuke0
ThK6H3aaLbJoS7631XJxOai/okzGf2MwiFKYpqyM0aB3kj2DSLamESqYxVf0a/1pNS033N7VvIOB
+nzbpnjXWe5VeWt+2h2GFGLcRWPT8/VSXxJroEBI6/bS7OvtpJLoYtNYH1eVaRtZVy2dB6WDkns4
enFA/iAtmI80sr5ejBl/qP387QSOaX9leBIF6IlveHDNKej0Ud2Et24pVy0ZQAUjWYTlDLqBJZZZ
ra+bmiQYg/LPanWezDoIU7/ya/iR8IS8GMQHWI4O65AJSwFhXeZZNimVcLKlam6r73U327On4oLa
gPN+XP4jBvdRk2KBU5A3rh4NFU/Hlmgf3ztdaDWxIt4paNFdCREbWDgeHO29yZUjqOR3INvH2FQJ
DqXc7Is7CCEetBx9QZCjsf9yhjv/cSnMgmPTJd3i3BSvMcntTex7V57LyGRttoJEwwGkq3rMYJ6J
YBg5avlvj9H7oxQGk3Z4vqMKsbukIleGUilmZZyxhcQX7G1qJWs5t2SJ7KXLJ7E+em68e78Fdt6r
q3ssoe1DFj3tJ0te0dHTR3gaKyBmc6iGcTBh4nTAiDmJckT0v+QZ9+hRUWEULhgiSS3LFabMQsja
B+TZHxvsTz8nM8jlNwA8Egp+3V7P6hXwI0G91gMYLBOMSqH86HOzJozFX4nB0Xi1Vy2xnoif4rod
xW1V8d8c1likpXfJWPP8PjhQXrqCp9b/9LMmLK7aWfeoUD2t8eNDB7lax17BwMH4cjjpviuK006A
EARQCZzJ6UO70wT+Ak60h+uw99n4pWzE8mQhK4BSd8eG0VGiKV+aoYcThebacHlLAQ6p1nt99grY
D/kMK9B+fzxioqkZ0uysKSQkAN3TsrmGXtUGwBoSA3T9MRhL/OauYCkBe7+o4GPaL4KT/LnLfxw1
a2GnxuCvPVxiG7prb4zHOCaOdikH9yg6QGZel4hoPDJCqraWiCzlpnuqKQLCJb5uet5I/j4EJSaq
SDzAuOhSvKgwhKEDB0NeunH3QBy7SO699dMci7b8RTmfJQOsEY47QQT35MAg3FLyJcxE9Ssj/twG
VtWJMo84Q+kf1ErFy8gH3noZm4CV/b65MmmUQXJhNiL/Z3W10+RLLPfQQx6+L7eomx1wiMaF1FHX
GDrfOIs9ymxdK4eM+sAid7gP1fD0kRLsUKZkyQhpWwkYlhcBL8aGzoe2vWzlR/KS+r534uvIWEOw
qbUihGeFNr0flDEtTSIwatXYLZIkpfTodyTgINy+Qs+6wY/MQWZ5lxLejJbnFYu0IR+oJogH5IPr
/42tbSvQ3Kws0lAhnQ5YYdjnb1aHl8W5qspeJKbQtCBt9hfEUdUoPzHjPjVduXdzs3zxWpQeSYfw
uMunJz+vN520smilo7+CFbQVbQEhb2NoDpK/XNY24+QnWC/PhTXgxuJmNv8lwVcW4QmifBjjR23q
Z/ALjuO8PSpY9liDR1D0qv4rB2W1dNzrfKuuRopZKO6J3hNSVW6N9Eyhq63YL7KmyvSCTLxVHynN
Hx061LJTAPGXWoT2SCOw5HQlyBRF7vo3mGqeqAT32EnlGZGCoxZOZolSRFzaLqtti1/kR2WLbjKh
iYIs509Q8y83nPrLDuwzXhQieuL+zy3HzXbdkfhVA6RVtogNGeAIjFLxc9WkToDTkTWBa0xX2w/e
hAXEp7pkQjur2WXsbwK042BoFoM9qSoHyjE9FksOZ+V3EHGZ2uKGKFGdre6H+ip2yYKL3sAo6rRn
BE+SXZD/EYuvFxQcoS+OazlGCzHzgdji5vhIomZlvD0z7XFywuREcLa5d/Iz1+AaPgW+wx/wrkGv
bAXvvCLkmlGIYQtkM9oWoOhKXRv24nU3AqARwlaNFrMwf9QhA1WaaLLDHLgHNnpnmxT1PK0pHt3o
Pgv/T2KyACI0ArWkfv2X/3Xg+95KikpZTp/9OTuFBDzB0xioq7wQ8JV9xLYOWrFcZcmMTLIqPU7I
HubjKUdZKbodju53BhA6aQSwTJ9tvKkibul8MU0LQeXciE3RBPHB7NMnKG3zQLrq5DACIDCVDBBd
u6p+bcIyPTwGbGpnX8zHXOQpDEo7OT28flbamKl0f9z+I7cd9ilBdwo6n957WFXBdqe8L3dH9usq
EVW8SAWuioYnJFHdHp0uE9i4dUtqltHdp69fV6wbv2TOi744OgWyKT3jMkOqvgYsrk0fZtUZujEs
zYrlHGZp9dVH6Ik4MGjyqxQZO2b8MBRwIGCWSWixCCOGyWHDa83jYLU6McIRzlrv9kIWGYUSV6HR
//r0TQ23ACToFuqDYXcj8gofRQmlf5pzHk7Yhd8NBr/Fpxfj59eQfXSjs1w5GrweGlEbKLlQu1cL
TK0X+KW1klFt0ZQ7p//Ci+cKlwA+dQ0/XlJC5KxWVNvz2kzjqA5+BhnsFopVk8cRXi4vLsiHc5Go
bR6K1rU7hBGbBrzg7oDkm/82rJn4p/xTDqwDzc8V0y8jtyKxPmUTAFeQRmg8R2aOSrODMGdTAvOl
ESORceW1g9xPHbwdPbWrR8kTSoI2E4rmSTF385YndWPyArhlc2A8QWezMyEh9W1EnUbI9QOKS3tZ
3I20hrO5KOFxxaNqZBoy1C7RTrdPUGo7y6RiAu8YUvVwKNTPaTifhAen2HRf2Kb8xMEa90gYqLx4
wC39SRoEHXfLPrrCgC5c7yArZ1W2PkswNZyXbsUOsBje3+ajRe5OVtYJtPJw55r6waW4Xnrh5S2V
VWOleP/2bP3pa0d31MxKaakIXdYFjfTJD6JLXY/n3DKVo/K45xIHIbZaw0eLkMziN/TalCEGOOjE
brk0tVHBN1lZLG9Rc0+LQyVsJyNZsSKoLZAFuAVMI+lw7+EaXwwAIZMrzqs0w78b62EMripknEiu
aiZXtiHmjRxXmJRM9c8LqVTOWpfSOJg9OP3b9qAMo7tQDvzfwLzRw73ZmOSl0a40ij+9wVTAJF2g
E8NG2BOsGlcny+KH42MUCHA7Ke5ZUE+LLWSN6JJcSAxx8OmPv06H6GT6qzqVfuoeoBsSxOEzxSyC
ijUNikKnK4LAl4DKOdNs5m3e0UIfQzqgDB+8VjX7IQm5OfnIhHAiVawZgiewMOzGeBLeQLmJMp8R
O8CTMDd2rBoe5a+RJUZJ57t5vGa7gN/SeHnHVpoBQJ7SjviZ55sxbQUAsKQkqvY5j06bSaQMoQy7
Fuc+06Qqpg5YmftqqhYfsd/tOSo2Jazp46FviWeVAWBaLF67Bje4eKq23GDtgSruxITECEf5mEpD
pQgEAs3g7nVSJlffH7oT51YzdtUnt9bLoNpy3OPsTLAm/OG4fZGOdtQhOWGdb1UuA3h4J83l5cu+
x2mcTnG//0vTadilvHEPIrNXhd9TivimXzG1iehdOpkKXaOroGeNunuwZlDWEFKCfI9BuTZzRRWo
xL+nZyuSYerG1QsOuvsHQRZXsKSlI1YB89Nlf22Zqbw3kll14Wz64iBNh9QeuBTOK8rl9CUm4Gfj
TLobQz2ECAJ+9YO1hQ45Q/W7cxkI86QwAbFDRx/tRqqx4p4uyIjCP6nlHsK95RkmiWaJ23ec4a6Q
DnXhq87PCiX8gjTr1XsYbBaOh2Ctt8TC2oPi9RO+fiaNsrAlkIiRj7CfCYgpmIOw0CVv+BMTHw0+
7Ie56rMbAJK1v2NXy4qcpAScOTc7KaujFqlg6V9FflNM/roMaSrOPV0IrjwxCpJmFhm8ixX7EB0D
ztHu5HURwiAfN094imns4fjjFJO8IiwwfNXy0iGtHSD6BFElpxZ1jY0hUHdD2bw+bjV3fNTj7hx2
/HUPBorpLkUG/unHK46ruII6j7xky5R1g/ZhkntfseJ57VqyAkF0+HOcBA7RzOW+WjhPMEfcz+hH
DNdIBhUPNNgqZJhomjBf5uTqOkgiiIus35lUYkQoi/AlT3LaDEbVq3dPeT1aGVtGChKcxC9nbxXV
94ALOJM6MTSUeTywvn6vn3FC7FZaNG5dqwhfvLRVCRfLOD7iVV9vB7chnDoAXRzxj42DgedI7/J6
VO5Sn7jkKgWyKwEF/rIjg6Pz4IrTpmBE9EtSX1AvT39cY0S2EH9NeoihOo8IrI3tX3DFKozgLn37
KOTzoutL+VvTy6PFQDGsCcPeMDxYAK8uqe4wfqc1iGmHLaS3DlhJDVogLHLA0a7EEAlV+ecLDhb5
RLrns6QuUPmQZZbAlOITnc080dft1erwa4XiQCottmADyUmPS50tcue6vHYdfIvyHGN6Qg/vndO/
BajN7AhYO8aFXszCDmD0hyLVcgnn6z9/TZatdFzF6K7plrIdbSwqRMDQtREebzsfRYCROZ2yI3XH
ibVpBPMU5Gm4KKkD9oqpmY11bcdi0JcxX0LRT1FTbXLCDo1vndF4jzeuNh0l3Rn+mhgmBbBusNM0
xPYQz62HQTxXc0zcgztg3OnxI2JnGYUX1SuVuSN2gqr7bFVHzZ1nkgObe7xq8KM/WHlGo4fo+irg
A4ap1/HOCIKn8eXOgwd063W5cciy/krbE7c6IVBV4u/haSFNYZuVbFgiLOalMiUNXLha7FftR8Ur
To8BVMgxnipbz+T1atUzoh/lgDuXbjEsaWI/5BuG4poMDJ1xGUkmQCcL6GVLMuZ5M0Vut7AEVd8j
weZs9wzOWY1IUKaIAUXt9L0fNehz3zoyQPMw45U9dukBaw8hvhP7eew4e/ndkUQ2uxMaRRDHPxwa
OPXb70JUNyfLuqLgyV98MqD1wN/gFQNjzP/0Oc2aRJxoP3aiGdWWVIfuMP3F+8vF4BX68muntj0d
c9GGT6Ov7j7DkkxkI66GGCWe+Ig5yrDan9EqQggXTW+hn17SzsLxswZJ1s8H7TfYv1HwfCz4D+G+
tZmHu8CXFuo5f9SGlxgdAQ5DXCECcd+2C3rx4FfyTeoajp53hBcB3FGuAetOcw45JVQns5gpAJaA
mK4396sqKGbLNbSOW8NpGdf+6E5EDVGS4QcLHqoc5vpFrSK2hMNNWBeOokIPCI0RBU/ZeF9LBxQN
Cy3Wkcpj4TCXgIyrg5jtYCug15lDHges+qNKAPN61ac01EoB1ULOpWK39rBtakQaFeRw/mPduWuF
h5dLOFv0vtinsw5H988wWdsLKaSC0N1WPD2t+kWZ8xx5sX0tLJ6qxx2VqsYduFUDfWKCXHmcuohX
hYT1JWwXCYESXUBLes27qcE3wIZRYnKPsBuh1ShRE5ET050bH+WtiNVOFmU1231Rt5b+ZYHGBjbW
EzMNiM/hjep4vWixeEA5PavNsnejJdhsAn7VYrjr/dROQ4V+/ocr9BgJOUdYq14mQjNt9FZw9HRC
MXDu32UlwCzCOs1weHqBFqTh+gMpAkphFqh9c9+DQqm1quNBQSp/KjzudZ/DMW5wsuiclIi/aCt5
1V7u8TI1KYe87rpX+T81nuB2+FmHpIxRLvL21kqNjHy0Crx5CDZkDe8ORICWCqEMYg4954WlmOlW
BkErCBuTghHzhrtPAtkL3MHYwsxbTq17b7BguPt1x+22IMHzhYQPuRGyDCyiW+sQH22XguZ/3cck
cUhSoNQTaPN/kGEc2JAATsaCjJ6eNnIbnDGd8z+dhjjT37cRT+lsN4921SQ6HTR9DeTG0gQ2+dm9
l5XYfUPNsvTubgz6YIYXGc4oGBVObLcDJm9kaNC/BWAAuEPYRWcGQRxdCq8WX9rrGhlLcleH8MOV
usLDBNaAloZovpAEA1HVW8WLfniB3YyEk+c6fpXI0HKcgb2m+9lqfsdFoodz4mZOrEQYqOXgL33F
v6OC43b7Y8MEDCBRlToHTq0jv2k0lG6Iu3gp2s4Gyg4HbT8DEk8YL4prdSziYHwipgFpwNMUKuGJ
3/MvIjGBx0HGkEGRkJPUMoAAbziZ2tDd/+nqewPyUKgDXEf/G76YMx9X5u+B8R7lU63NaFNKppy7
L9MveLaIU3EH2EWKqWeYwnYQn/YUPaPEYjNw91wYPhPSvjWJEPfdgIFlxaq7wgkoJT70xVjVjLnZ
slKOheSFyVKdIMHMpEvagp18exEjAHN6Lq6ygxIp8Cy+MKgqukty5qczms0MebyYb/YgEH0LEJvl
wdfSokeVMKzO2k+pg9J7TtfEFxlirTtp1oRO3SI04A5ZOG2wnNYsRI6gsv0dfAhZ/gezIArsJ560
Z5I+DaEub/0nQln6JYliTAN9bd79a0g788QbkZQUQ/NK3Sd44y89XKabEooHssjQGEvDHG46/UMY
9083Jv7jKNMK7OkvNA3Y+6VtvqLiXcdH25bfS8hHFwQJLzXlUCD+eEjVv2wcFKfHq87N8LPZsPdC
K8qdFUDg+N2RW+L3wg3wZB+iOoxKzoz7r3WY2VVbf/MUvLraP/df11+veB9w0Y/rjqIXMUe0L6hC
nfG8Fgc61nL4m6bqhNc7DkkjzWeAva2VssMAqbm2JqYA93Dcm2qigq7v4M1TDr9JPEcKoZhhVGgt
ZI7RFlhpriLLJIPc9DHvJDCHBV0DmRSwACVeug3BvwN+Bna8LhViajOg+CJX9f06glsV20T3TQuM
FmX8HE3/Mwv7UUlUmGfkZJ9eMIkp1+C3k1zm8MvoZ3UcCVQTHfqcHFMBRF5VtS8GrbiexoPULixx
m5hCTKML8GNlAlN2TWo5lofofLWbziKJB1sBu1XHDMlUpU1si11ZXKv3UCxljNdba6H5ofyF1YZR
aQtHV/DSMO3KeoooBkPs8Z6n/fnL9kgmFoAoPrc91zaPrj/IyLyAIjRVJ/iJ2Hgs8Aj69SHYvY7f
nrvjHnST0orMJ/DCO8jF66jgcd5aoL793DTtcxntRGH7jP55NbsIY6SZJYYRPUaagFu/Qpk+O0pn
TXS0YsDNq9HsAcs+Xzx44Q77hbVN6YY/aOIWnyiYsDNffUxtDGgVhrnr8hNFq3cm8xvE5JKO1tqt
srDyIQmAYQKlEooIKXlQthGW2sxe+dFysKqY0/rhOM1KWObROCXvjq3ZBkV5/SncwEK3kkZbuOl+
EMYUMZNEZen1sJ8Q1pcwWr3dy4g3U+1x6NB9QMYYfqt9WuO0f4GBYzVRJRK9kMhK5CI8DaLHW2SK
oF2s9RNxSNikS5w06bgl6Wzd94DyW0MpENM1T8tgOPex/79z1oLctqGVWGdshu4ykOsA8LNH3LmK
uOQ8KW8AbcUOiX3mv4mROvUlAoV5PlRwr3XswuyE8rb+v6mVgFyCr8Xh5uTo1L1xSobY5rQWDLY1
/pXwSFEXflB1yA2FfqzrzWNmHbAyWCfBvPtnMtUcSnUI+imwennxVcMd5WmkQCdaNrnrOr5sXBco
HEFdCBzOIC6GYhQm3AvyfGK9XirpJZCgayYe34bLVJCqEuqTc0sbLZK3Tqf95nacDFVuzLgFJd/r
xwuisvJO9d0jwVAes7UYJMv/RZiX31N448YTIPtkgdN6uNv0XSgoC8U+7xqP1DkcZ/gWICOuHU/9
6bteI8Y7jpRDgACf9GdghNRnuRtS/he/fJT0nHJdPCd1Yvslv6gGbvchyhKWubrQtiyLC0DER12i
wYgAflPzWewMtt9UYBUY9bxJPISdD0vBWTyWjaEnhfYEt7MBhoAoxPUWQOGAwGqm20f5/gQKQ644
HeDnQ33t0tbUd+TpDwbsH/1j61/jHY6sDAeggV18Cg0xnilMmSiLOiZtYqp/PAvwPufxMRjH9vKm
burRGlx8GVD3mms9RPVGm9xuEAi4ZXR/ny2RJOtB4RhIR1y0+v9loPCwQqDV/ce1CWd+NASIHojc
W34DK0dU5YRGVvMeSc8xYVWoejsLUbqyZJbVPD69dZxmoxhGYW6jGvxvWlIxFWSsUf7Ly79WSX3G
KKcZcH8HF0LU67uG+QLimy5VV/IxX56mYblLGEAc2Tgf16xexyfr2+nNZMsOuemcII51fldUkV3g
NqtE3GDRjB0zzHvogV0hkVKhUAoNqu5kJ7ZHY3FJN85o7kGJPQT53KNWkWfB+LhQ6c1l9L2XCPg6
3smjVuw2BhG+nRjuhL+5ZK7dH4dlPF48eQYpmXxGw87YcKhqpMUO9iXPr5T9x45hZOEpCZif5+47
nCMQxkIHsqlH1I83uPAi9foEhwQU1x8yp6RVafldjoBdtU8PeUIIYWtY79YNFEVDyNlkvn3+LcXY
JmJfDR+UVUZKMMuhp20MXQiRvref6q6XtTVRZmEdMuJa0ncibA/pT9fIfLNUy33Uo/jncGp6qd1W
QYMXEUh/sWvIR+S85mdgo/WMXItIcYuGlRPW/VbN2fOsJuNxbZeqOoueVwDv2FbOGG8XC0o8ncP5
VVcuI7JDloJl+O2Mm6FGVMxwt49NXhkIlZ71YfsRyEzS1evaIg3pPSvUJZOxxBIpzROHhTSnt6qJ
47YAPg/401CHErkR51nKkwQL+uqWJP6DKLWfZ+6H7Yhls0F9SOEVbvKGNqfiPcPhU9ByjNQUaplr
ZQX89dQz0X0lWUMZ5/iV4pyTnZCVuROxu30hZL59mQcfT0cCrOsQoB/xGSz0vFBSYycaBBkHJpF5
Ecps5MVDeVm8S7WVdyVByY7qH5olGZ9J2Pc5EHjlnKqCpm9DVkCOgq4ioOhKZKFOQCqcQE3Wgmws
R9pSzaA+En7xLNhx/7i1kPgwTXU0mM39NlydEqQVRjV1lqamnmr4ilOIiyQyuHQe8rBDyNTWKq56
jFhBD3c/jL+f/X8gjvqorYTZ2i9S5SxD8S4mIYR6DppzadGR9yPXKYAYN7E/9KFY3k+VyDTsfEdx
Lu12QtW/ufOTsryKYHP937cETonDIQqZNn8acYIgWIRXFeiLRKQV5W3Sctfo9fngeiqHj12ByHU+
kLHuo1b+oOXmmHUUAlA82Eer+4JdJv9FJatQMMwgAp+7uYrI7H8jc848gYXGIEngxFOQ3p95nzx3
fJGJBnh8G7hJFb9gWP8ggD3XHqxatqne8ZPAfctJgCt4QlJZfMXy74hDD8j/rOitKtlA1Pfcwa/b
mTYhz0SF3hHQBYAWV4dDdQI0c9OA9GzsuWUOWv+1LsC5isL9NirQSEAP789SxzCuaUpU8yLag/To
2p8jg0/OPgU7OriLjW58JmqEHOWAOblVrNVctL3w7uXhUJ4EU+fgTSEnAI/qejB5dsLYX/kNa+HV
f+EUn68QfTeUnoCdOvHJ1yJ0EDu+n2Hm2vSlegnbA/DL5VXjkUP0REZ9Hbx4PSVoFG1I/HOOTIPi
IOC0BLGun+VE5y6arib3q1vm43NsRqxvmBCer5EcEp/HLMXMFqnFZ5envJZFqtUw/gzEv9SLrUGu
3JPVdG+PkZ6l1T46tfHiQqDDEyskNSs4yQnAmgcSke2TiTisIsXeFLG6VoSrU7qghwEV9iwY5R8A
RqXCiw7TVWAxtpHHIIoDh9yV4K+M1+vyft9X+x8QTk/4GKfGDB/sljDkCGiN9hRO+Gqd+ts9/9iU
9Ykqni+GhXoA0AxOqnD2wFYMHk56xHdgcGDjdzTE4E5Sy8iR9prAhc0A2MN5CbJ1RHhnkIJZIEa3
VX6gnbNAmbHZqCHvjUwHf1PNbAfM2pIu9S3R44aZ5KIAB9nrwsTXfAai27ixavUw6wSYhByxuPeR
GjVZVe9P008pWpyh+FEHcfLkNNKAb1mf18tOgtuqOFc7XwAf6HQyn0zYz7nWJlwLkFwHZ+Xb6nmq
SR4mmJcKVYyj4BdhwyRMjs4LuXqvkl5jOKnz3+55LDfq8JXh+lVeiKyuLnhQwy/1Oz9cnBShNuq+
klXDPMKTRMV0eV8/p4QuIbQ6llMI4mvyNvjwUpwFRNE7mZ/DQWF95FOiOGRQ1vEMQ8pxlfPaCNVj
8uiic8GOWCWIquFIhHsPBL0q3x/vMvCKVB6YKt+E249cnbJtNgEMSnq52/cXesulGpC4aemUlfr0
+MBelb8XJ9wZYaNsHhO0KcF+vSgCs0cFDd+zsBxC6q7Qk3UOgKJALr5/hKvAmN1kgLaccVss9yLp
aZIxrrbcqrTtAOFrQPFzlHKrRg4lOmiirfaFb0Kb5EeGfZq0oAHE/z9l5NYk3k6ODKFpXYXoRokC
AxqEMxpYUrJr98hohV688SRB2JdsDxEESq459TmTDdMc2tpgvxL/WIfgl/NPHBbVvScSMdBdFrU8
s1hXQKNBzu1ToZ34FBo6fy7zwcpF057DW82ZA8JPKngigzC07ZXm5M36bduYcdZgjjIKITKaww6Z
OVKT1ubEoAE5gsPy5pLv7Lt5T1VSZrs33yh4I3AEpubyYz55Xc0JqtgXx3uQFxyyqmC1Gi6aF3BT
vKOLO8dMCqffxvsRmVUgIyNfGnX+9grUWUua5v5clZqe16nQZzybw24MXrvUjH2XBTPSrZQAokkJ
9V7EW48/OGtffCrDsbRmB0dSS0M3KRBjn6tkewdWrbzY+ePsnaARWKclXsW2Ee4F9dBr98G3KsbE
HZQv+04YBdzxf69Mcl7h2cYz37CkXs9CWHWv3+t3XiZJbRE6/sIm7Ts6weQUi/l5YeNdEPg9nWWI
uhnZxzdBkL4G9/FJ/vB1uCwOvpQZfd/G0wrfH8FC/SzviP6Ddw6bRxq8pUMdHw3hBgyIjLIhy/Zi
Be9Hrv/PdLAc8MwqL7PYPTYV4Ti9H1TAyoi3DLV0b217x6UqSW0Skhp9TFVaDbgJNZ3CEpa8xhCN
YwEJ5MeIjrClhNEzBjsNAWsiDC3y0YrRcssChgcgIRU9xrvhplr7cN2RJFjv9KvUfDaH4fplj0LI
L5Zm+EzTtKzOTRWPI2ITQQFUukPqJUQ5amA/8N1jpY803coV3n0gqS8tQrUqTPNO/kqnaIqIPC/L
O/oS5TceLFYu8riJdsTlfpJOAJgIICvWdjoO+AjkfhTQhTAvKDl7OdQyEL/xSZhjNDjq8YPUyCTp
/iIZELOle1g9Cje/X9Wf7TJ7QTcyN3bRsTwhb2TDe/jb9Q3CQg5RRg/vumT1GE4qwCsF/1ojGRMz
YqP2ea+pVXSUI4OsSxVEfO58OvVBm/WtGk4u0cFPC/XZ9L6qoG1DFhh881f2seu2E3fzBhRXPq0u
VETCdDGrF+6EVG9+UH8VMedsoiQ9PNU9FT7tFqc6qoIqTKE3Mrwv2YCshCapW4LhDRdcb0Qd5mGe
kECt2vCwt2d+QE+IFOtCjHMO2JTrbbI+TI/lz4RuwFBGyS0gt6ZDAk0dQR2asR9rzpz/MVN1S1HN
/ePwkSayWbhrcm+WL4+7Szq6kEErxv6S5iC5feNOrZL2buMSQmEWvLHYcnBiPtz+NcwBzN7CIiyN
bAOVmnr5E16CnfqSjChIBuxKBdLgSn9BEh+8gcWvE4aVDjKgnks6GcznuRGHQxRz/MaoSzuUuAus
o2P/B47u7Q+8RZuxOuyGs9cahtQ8Ca/7mNTfd99GBgDJsIvQGnXxlqxj7+SK36N2FbmTW7O/O72d
qgte4NCZd2bYv8QyxHW6gq6i2Sq6eZ4WZ4oxTw5UKcAUEzKWMZ6aGhEF/MW7X6JfWycDis/k8JAX
KNitEKr+mFBXusWfQyq2NcAcCrTnvW9UtkcJGyyC8gIbs9B6ZoFqBXOgx0g6mqQ1VQxWVyYMkZyF
dmQmf+Q76oi/812/p9fwV8v2qXI7VKNVQCY93J7FThA84x/NsOdif4Gd5Ekmevt/n2PERtM1YbYY
gNOfe6JHyZ+RzqH4vLhH+tKd1xXUTZI+IpXftKz9o0r4DzRRCzlvMiYWcaRU+nqqxVIcLmkTtHEg
oas2CTJuQMmwvMxyIRsbpXYAXFlWBhWa3q5rHyndr4X/6Ndwaa2emeAAb+PyFs28t5upUCA/OtpV
TwgWcuV2xyNC3WGSBgdocE5YBVunseiPG8+H7gAuxWNKQmk16GbJ2fN9+S7Qdw80qfrNUTM5oFmq
Fz6MRyyhX6CVqX5ejZzAbdx2wUszA3GNZuuXEJrTEn39fqDHsq7L0G9JlU6JtfWcHsryX/HJPS2b
pKClCXYEIa+f2fvL85gpjzyL72oVeERKEhdvDpuNAylk7K1LNsA7jg0eExFC15M22FKopGqnk2uk
hUtJEumPFNI1WyYmJpY12aJ/7WMUWgs8Hz8jM0QBvFZ30UM+0LlFDrJhxY2hm6ma273qO5u0r3ic
a1K2nIF9fK//orQKKEk4UZToP7xVn8+xs++stWAgtsfloDYoYKaQO2c7Q7S4avXxidDkB27JSIUi
VNr/oxj8i0xcmpwl5ild43jmKCQxUV/+d+ZkbDQA84yO2FySyBcUGH+zArIzU+6ztWfhjg6bFsbB
3SANaxrEHLag+J7xkIX0woGlwTEDRlo/JK2WPCZ33Y1ZBk5o/iu6OQnf/66mUN/oaBBr7JfA/dY3
ARCtj2k2xZeg4TcKM49g68MVVCQiPxqLNu12XilIRCCzrX36r0WAJI3HHKHZh8uQb5kGFSJAQv/z
wUOnW7qrVEqYC/tpHM+P39mXbhFHvCyFH7fTzxYmDga+4JEW8kQJNZQWSPya9vCO5JEkcszTPO15
n3+xTAFqDSMT/BNCwTWbBA3Ce2UL0kxJWWw6baqvXPCpgA8BzJrrmabclAzDAJIN6DE0HTg0IJKq
XMec838SZRR1sOiSa7WA32CJ/c8p/b7sbX8/yHNc/kCpCPE5PerPi/ShgRuhXACu3GMBSFmbgXTu
TpQjJqynZNth+J7TgKVXGw+ppLUEzjfFxR7NdouRY7sNGbTxumROTHi+WSAWfzXbyDfMlJk21rET
oLjPISgt9hrGNk3xDh+46sdERwV6HJ0EGPijN3iSBdMjpm0NOH635sOkG87qp+RCZ1A3kN+VwWVS
vYVi7unouNAlNqxCcJpgppJlO9hu89UkhewuFjfyXfay0633cvFNcW2kSxsdxqlinnLzV6Xz7QgX
W2MCgTMQwufuJ/Lh8VA2qarLyj5ed4XfC7ZqFto64xPggDRqR5gp5GALsULx+6evMI2Hml5zdoy1
PiWb/jdU52YeVkGCBrKc1dzLcYYCiNNVpkM+LwOlMQTXwQ8gkdG59LLHG4LXmv3mgXo7vhc52WfZ
moB1jvxKVG6OjO5fUAKVbMyE7uTXykYwLoKKb0XPYyZ2eT0KaXi+XOQGpJPRZDAMQ9OF7M/mnuUt
n6Ag0jS0KrblJn7NDeO7444FzBsyZFDBxISc52iarVfPyw0CjeEdwwqthX46DrIOJzuclWTKZ3Pq
gjJwXciw81zVOa6aXLCrGlMl2noriaQthDfovV/7n4TY1+7Lio3ogsOlcJQwrUvZvRtOGsHAzpzb
DaoiSGgoNYZZpAEl6kDEfb3fCSGVaQKZO3BlzraYukaUzL0/vnIzjTN0zCEY0EjQq+BDlVoD/et3
2nU7PKZiZBJP4dU5ml7Xsx92/i7oDVymvdsljNnA0yiAdfWOTldzu9pAFlG1vtI6LPGA7j7/9K+D
G6E48rM33LNpikL/2lWmtx9ZIknbxHX8Y2ByZXNMddVKmmzYahNk7Uz+qUFe7Ml/TO6dDBDtUWXg
OZIHG2N6Dx184bAqgtwpx3q8AuHJshHhmJHh+pHcUXJVRfR4gr/3xehefnkvcL2m3mgs5YQdJu9P
FJR709N7N4thr0Kdez4ODlBK85e9b1wm6bUQowlgsnFO3RRKqJ8WXL53Pm75FfezpHwUSZiuuJKU
dG0YsAZHTKBAUWQxvFKes2sRu/AcgKTGNQafv5q7TY3RjsCVcpQVhCBfIDcIldDExahV/Lfn+Zvv
6MpiwNomkMdEjJKGbUgQ0VeiRNTAdoKdMbPRkh3qeM3k7ZQxalgLKD+jzlbW2FF5rj1ldq8OxOy3
defW00Q1zSPr0nU73YMD7JcHXN9aAuL8boILJvRDIvbETypK7SQOmnbe2S69BtQBhemRQQk6eN1L
6TmG59Cn49FZU6nLlbwhq3bcuFuvm1YjEs/f7G9AQgC/SQ3mNqVqjIME/d4ecgW2B9qi0MYe1llM
Gnbh/1NoK4JAm96NlAZNmjMaA9mLJxnyEKoF+JGyEzkpRgxj8GEpVcdf71zbdZ1gPGHfKn93eBkn
nvgodYjLBPsiDpGn9hUlyNwgGc6BYSdFGOaFlu4CLPvbJYrGJbTWjD1xqqztaiJH98ru7pwuP05L
bTpoO0vvvYY2bw/ypkD7eMX4qkqSN2dNU6QllNgFHBZZplW0t/1AIOqf2pFw2jsnX63XqcOI41XK
Wts/ndW42ErAJbDCOQ5tq9ZY/TpAo0giD+TZSg/ZJd2xYsZJcmAqOk7iRDYHH6BTYn0/RFmCZZSc
2FLeULeLsy4AGM6g3Vozc6otSJNkalZU6xdYdIpqkWcMe96WvqfQLtv0BEPeI9DK+S+EHQ3e7/zh
626IORuCXv4IlyTdxR+q2VLLxFllca4tdds7gnTIVhmKjxE0qP0hu3h0potePsamIA+eGlUO+7Rf
st96yMPJvipUYv+delQLlki/PoFt3HbpA5KBw3/6RZOEDJOOVn5JJ/7qeBd2Z19vdl3cSXBQY7rr
D0JA1pXyvEwZoXJ1rghk7uz8eTgq+lj5oQx+IawyqeNw42QXPM6cpOjqDtaHp16pzgVL4id+Y4/p
Ur0oVMAis1DZSUDKwStdeYj50uXA0AdWAwD8C9VRbnm53RC5QOrd1um0qWRVpvHd0/1dIeZPVQc8
Q51eYyRF2+u78BmrN07+xV4OxJJeJKSwp6AUTWz7+p7lkPlDwXnj3yJjNhGjr1WVv6zVUURO1yBL
5u8+3rGL7n4gVknnSKyas9GC/v8awFlH7LaBI3udZC0xiR11oWbOnTWuZaKyOZKT+B7xBlRjRv0P
Tovk41nQkMEXQ8pwg0hEgdW4+8MMlaXmLFONrLLVrjO4wOBM2aNMaAc3i3ObOMOmtYuETlWEZwgr
fH7CaG7R4CGRzJP9QyNPoGhn7Sm6a3r9WjQezrPyePZJR974kclOWHnPRwNxObl7mJpyhKrIcb1L
EZ2nEt3bQldSUFp96dPr/vNgdF1DvKu73bQnq9zzgZpnAKkt8gEx96KZORYhRwQSD0Q3OFzGQArQ
r93VRJZyCNgCrpdxmOTPhwPuTTJkJ7YTbwuuhy+SPCLpu82ngCEcfienE2EU9yR6prHQ2FiI/u2u
ktuuIL5uMA0nMRACHoOIwiQE8L50/m6JAuHrd414ztZBE1k5RBF9hMVbUdLzBhr7XQVoEQQS2kTG
vFaJ5dTXWzjz042ivwnWdlRWwZnVHQh8BXFO+GgJoPQt6DgAsXsIUnpoZOpSG/L57+8dewHBLSaQ
uoSuXh/BXbqIzg9gBIJS6/LOB3/UTt4e+3Sb++zFpfE4HaR46n5nuBdKt7B25DHD5HYKl6AgstLf
GWaotNuBgGY5J9qSYbJPlomgOIWXNW4e8fGnYZBAjj4C5JxG9mVdoyUjZ9MFYGRAOZ3HXMxNqqXi
v4xvgkA6jOrkIXaum66jgeujDIhyK0GEhciJDlRDFNnwfAxqoXww5FJU6EfyVWVw0kK/jXQJJoIp
PZ/eSEttTuzDxwvmXnsNBVIqnDheWEmTtZnQvWoZb61jd5AnYVF7dQk/o16Pzhtc13opZevBmQzZ
byqOn70R7Q8A2xdtAH/5hwPb9+626nns12THGFIugUtmmBIH7v1wCoAOaXz9s6EHHfuUVU0hQFh3
Jx/YTZ/yiPc3qpm2bmG2aMLEaOhKIOtVeuuhQ7aswan2JSifcaoxbd/f1SKrmJAL3RAHWQlESkMn
SAZyZiZCt09z4Ykg2Yfa6YIRixOpzcRAjEE9z3bBfJP8p1GKvopZPWdgzJ5g1J5af9wUr/UH9aed
mZeZu/cVTXssdUZq0LW0OTxzrrMSta9KyB8sDbzfe71U99ktOlK5tSSCt2jbS0ityypP/XIQ0Czs
7GIyWrFf1yRzpQlxzuDS6VAvFfFNaASE5MZCCmncLJOT/G/KAGP62zAAli87vNwYCoYX0FlO0OtO
8eUwLPP1bonlFgXj4n1IJcFHIE8TdT0w9YJmUQemiNtSLxBxpGaRlpQ8z/7if8zwDe73L5sIy15S
NboBBf1I9Gnnm1Ig3EpiyUBu6PXFB4ddot78Mumllrc22z7phcMUz8CdB8elEVRHWA6qTZ6juAM3
hK7TTiS69V2IY+aHZh7MZWs3MuAuQtjSkRs77vEF6FmacpZgMlrBNraweJdt7nAAYvUb5g66i8ED
V2dSzfvMAroZv4hSp04ch9XPjwFu9rmkKr/WZ6nL9lrMQ2b8VHQtgERc+Tko0h9JnjoCOhFVLnJ4
0wprrgsZfYdS8dob+KMLCS22Io3kHhC4gqPUrms77IHTheuS23qf3ytw8fy+rK1CeePUKluYSCeH
OLdSHFyNDt7qhGvISabNmJKhpIAg7KSRNen+hSZTiw3GF38b+SaamYw6uTOx17X/wIJAgk9GvF5P
jT6c8jgCYxei1GHYXiqZWPZErnZbPqrw6nyYSKHIMr5W+2zALEcQKIr8vYQd0ZWK5RR6A+BvBdPM
Q9nUhviS8Rr/9RM86MIrw4/0b8RjH6HCXtetV/6IGpCAJbEvcagN0ieRSXM+YiF8UrCAiEwWhLpn
8m/Wf4VZ86JDEsjYGHHhOw6tFIl9xLdQgW8ll0prxU5YykGxTQNkuffIox027s8390YqEuQhTgoh
iMGWjJ3tBcmlrQs1igA6evAbA4VSd4371ZPCVBuTsoSzj6lOXCfYcRaqEJyqygSN2YWLjoO0/V/5
HLcmmfoUQjD293SLCa0HEaBHv262r/y67mtwSzGhmDGXPWdZR/OqJUi3T+y/HPCDsxZNPFZI9UMX
YqhN/eekg3mzYKKhHLIC+871efHeEM/KIYtkOvDS4jcZ3Q9GYNZX81CpWhlkTiWXx7H2KpdTBPzq
78vzL4F/yIWgvzkDaVyIWELuEcQhoTi9u1VhX95jCKSvp8x3TbJN5IL/3yX2VmOHNMugHy7WOjdt
ROoLzDASpHaT0d8fpjGVpQICVxXxybR+b1plqP09QJiROwS5mIyUThyBktYmcyO5fciIVBQPYRjh
jIoRHf+zbyfoAqRrkfzMlwSvwqk/Wu+3dmCUw3VN7aW3hFPqjDI0jNpEBEy9bnNHRKvHaThz+eWB
KUZc84IcEjtNFbbUak8WxsYOL+XyBgXxtglRvu3he9NINYauWps516nPjg5pz8xYOyQZdNMvNqw+
IpeZgGr0ed2XMF5P6f3EMyPGEWkvgVA/r0ee+gVKmCu3IF8Gz2PAh3sbf1XeYWAVCUzDe/i1OFM5
CFQ7THUgvCUYOk7HKcGdLp/LPnnDRaggvecg67AznMLtDvElip3t/zSjeXpbstOK/Gi2qnyaZQXZ
sfnIwhVGMV9SL2RjS+f2veRA4hS1k40dlzx2AyS4GdJKByHUfhZQPKmUV0RArkCCFD8vmN+Lai/Z
QJRtKs8VMCqNjSOrEDW3TFfgYKXK+ewtYlzswDMC19rnv8d/3XpSzWC+XvM/u7nkTzzdQ5rL/Ovh
3BAe+0mlEAqhjYRUaB3hCRGziO95v5TJGEgyswXdOrP/yCBR1c/FQD6tUWq12iffFQ3QvC81pBwv
+vnsVUY9nho6ovPYDo2H70uDyy5W/f8kVSeJLMtJBzul66XoGr8QquuWglC7mLMD4hALBrB8Tpau
xoVCimLl2QeycnoGyT3ITIhlQ0nRqZpYbdyePsqmESySqFG5xGJGFxOhb+F6g6kMnNXl84Dj03gj
SsihBPQ0HgcKVnCo0sV6pIonZ1INpEdLUlNhpzJzM+gqxH4sT6N5ZDA/LfX42OH9giv0zt5mSWQB
ehfaEQurue8I5pfAqrKaWN9nYT9PkQhnVioxOScbAObncd5hPDIaA+VzvqCLLOookL20Z/w2p0dT
CNz0z5qqQTF5DB29a4Arssin55zSZEjAfnGjyQ6LWfJUhP8h7FMEYFnzqTjmBB0geIH47/W1UafV
jtI04TCvCvhFFEtGag61myZrP5xfcdQzEzrKkDXGz34ZMno2Q6bcGFyLm8wfT4RmVvziq0ljnFOz
4MIebgMYpmuP3BNGI1cOQIWtmVjxa9K0AwJJaMZhyx8/9POOEVFcZiHpEilqVDFVvixKCLCv/6vF
DhJ/HMisj4pyIGiXBa/dDBJXuyjllW6GXqjnnDeHgfyRpMHkoP9nhwEnc225pEYcAN244hX+1gzU
XEmt3GE6spp+bMkjfBtyr35iNP6rQQfzFa0ZHI5Ab6YJzlKIdXYmaQYqo84B6P4O33k/2d3gzN3g
0UagqnkmgsNwfURkg5XOgVdI/KuWekAQrEP4l02fln5Uf+W8Vl8fgRy/ycSaflXLW2pRCuZE9RUo
dueRWmjq8s0Ij6biSa4AGKxa33cxunM0OM0ZVwG2QDcms8irWpISlnVek/pX31N8cGTeLNcXQb0c
n9dBeawbelGrkA8dnX/eRoFhccJ9fA6RKxEe82rgekQRiGJu8149JTed4B4XiYFfttJe8OgvFHxb
ns+dJG1clVE50TzCsgL0Ekde3FNaTqvl5dfse2LAQhbzUYMyjud3uH/9bz2FMloYRNXe89u8/Hts
4PucQbEdUagUiIjYtKyLGAzIqwvDpYzTiDg61gkNgOR1AXgr7zAvvHGfnvVRXNXoUbmqHJWz0ZNh
QLseXSD+6WksNPtNwsl++kPI3xeCld47vta76vj2Y3q6ADkciXjFNdgUb+peeBU8FcF/vRU02JaJ
lgyDmNMZYwvi6URJLgUQOKRwDbgQqT8CzBTvatYJS+w8XfhlROBKMMKg5x0z1Eat5zTs6JmnUeCQ
MO1cItyorigRRupl59shkmxzw655MRHfAJSf1nwu0VmaAEq3H7nRGQJo340CI3hlvZXH0+F0N5Mw
O5Oej7UbX0nm4j65SsDQaDJ/cVt7CNlqoSlfiYE8gczDWMbMDp5JTfpUCE3xKujwyrXRIuAlXpZw
Oo8OY/cqH6BQUykzAyNxXrlNDUVq/TgRBqz5NYjxbYdm9KMfFt4UJMYgVNVg0q30heLVQUCuPby1
1O/xwRddmANclXBBbuKXyy6zrzr10VqtztL3LKE9tdPYn1ZszFhxxP8Kp2hva8fisqMzn219dWdy
/kr0Ozkf+0QFkPSK7+kyimJ46nmJ9uIal+AsxB/qpNH8lImOGR06bxN66RsDL30Jc2BCiw7AHkqk
oESg8gwTuqWXHhQiybVkW2mVsZNLMoseXE6pFf27RzmmmwVlwl0XX3dhLRI/pbCO3SAdNWWuG7K2
eRaG+czy60SxwZDbgwzJXQ0GUTZjx2LTN9ssxbEd13gf1GK0j3xrN4R4PRW6xWyP7sRRe3RzPKD3
Q03nhg5zn8b12PHMIJfxmP1W0QCyqzQMYKqOeAzHP8SNTRH9GNC3GIi2MkBw4foxRaXhpsdlYk0f
27KKYLJDnHsRg05zxhbsBlfJ3ekCln0Hul1JVIBgXoDOt47C72xSz/08JL87iJ+G2S5qlzpdSFb3
ExA1ZYa5zBu+LOor6nYgTJqo1w0RCE6DN5f0znmE7+sMVbEOV5+NGAV1QEcgr1NUYFrsnTI9CkKE
9ju1H/rYqb97IHB+ecXbx4P7K6YmjMo63RznTmvBbufK+pWMaQM/LPf60iPnfIcOYj77q67Hnr54
/4+QPH5/sHpKEdl7KwXqurfc77djWyGFISgCodf31pm10bxEuHltbK1jE9948P0j2m0zf6aT7Oh3
lfaXaS4PvoK5JveMHVhY6JihLyGqsMyq+9UwDOE4dSqXG9oWBJSKk4355bso8T+BtgdV21UpVu97
FVYrghB6MQv20yimMJAODaP8nlxilwsXk1dNihxF4LDTPLHJsDjKf357OTJYBl75gZybzjN1VLHx
/vJtT0k+NwAqLcSGALE2tSoHDLPfE+dB+z+lgkisI3esfCLOQ6Un1A35xZqm/zbKKTu+5tPIPQen
qnNBb9ZE78OtsqM+PLg8ollIJ3C51Fw4QPnlyLT/l1wZ1K6m0tJoHGzijwbOC+nnpKEmJn9WdLnk
lbr+bfMv3S8sSXHHKaFmbg+0FN7gh7TlVdb3eCFYbiu46/ZUqss0AZ23YQ3EsH3VwsRdntwCEit0
oDGxX1Gv1KuwUOjy7K9J9YP6dZsNUyqpqSn84hTdO0myGqRHzBTBj9wrldkOppCjJOZzANThtBJY
Cxq2Bd5LC2lJ0I96X+vKILRrHECZHUP2O44leQ+d7jxi4BGX7wWqhf7Y/WrJZjW+19v0RmZ8uDH+
41to43Na03AUfiwjMKO2bDfD16Fv0elivt8skfnnjbOJD7K7h5Z0lkhFMXugF51S698pHPlv/OWw
BQ+ZYsJHop5HHv73dJZ3s/De7EJ6X0dX7uOBDLkg6DmgtKL+Hh3wTlRcjhjE6XemBLDHe6xrq6eQ
nRaQfb1vNQYMYJ0N3uZT7OHXT6rRJsqMzSsWtZDc6gnDMWUgGgY8hFNYQp7FCPj862eRJhh0nra1
5qxq3xK1uBdKxcCXVrxgAAQtMUbZXWZvHIsH/lQU1JHaaPwgtQk3DkyBYPUQrsVFS8gMT0CIFeLP
fUCq7Cizd/VEIEDPH+6yywroI6BiyuxQJaXVRySooyJeS0O+9gJ6OZ0uw4ZcZyPIPOTblSH27Hzi
gyGfiNCzdzO7PacU7ik+EjzQOhg4V29wXvNJCfCGsqxu8WbbvdfVD/7KTlEMyjHiTkamWZtxVHPp
de8CLYzoG4B2cQOSe2xaWL7F8RYdSydsW1cQMlDZjYW/zCn7Z2Cj1knNWbgvxAYTkeMnSFE3MQAb
0Z1YuoWHrdMcn4nhZPjKGL29pEcpM2De81Kq2WXI5eLsNpfhAoMfk03MMh9LwmgZ0fBpN8Pnu2lQ
X+5QamAO+iW6+swlWdnRa87anKzGVZCLI61O+jer206YRVy1w0nF9R2hAHSHyyqxVoIk8jcmRgIl
eySFaMDE++WY3XkFsEjDNBkNbCNV+oe30pKaSePrHazX6E39SUrwhbTU9OOt87j9vviQGZJzzZiQ
6vZM8bNwSQHUn3+Fxd7oDuHpCOrToCHXcLwtl07gtEMOac+6d6jm6D+cVnDz4/pch+gVg8QoS45o
znyX0bAyFKPF2YrbOF4jKOBJKemQByJ/6st+sHkmAvZ7GTBePmk2f+WyWUTbh8QETJp4ctNuoZHk
59lZTVP1fl8gNN5SmAG1BTwybxecGA9TqjNFknmVwC297MH5tY4FDYbvNCHKg6GiQ1DofazRBp1s
VcCxgYBFRwNAvwZRQoiWmjH38nlxtQLgod5dPs+0IeHNO5Wfb/PZKzCTx3AvFmHpKFZ+hMFebcGA
fMGZRHDNRAk8NQxvyV3t7GBlgWlYkvWuEsiYPxpAHa7ytWILm5BfUJtpw+UDVDwUJeV6s6n7VFbL
DVrkoGCSOiaYno9SD97gR0iLlUz/eczPMxxnCpsaxZXAL2h2pQlx4Itf+hGPDBehNGAZbs75a8hx
D6xfNAnqMk8/a/lZj86DjwPvNlYzgJKPCL3fRfEt86NYWLy3Ea2FLBre9UmXoXF5iw4n66oXrtsO
Z/3KeILv2qfZ1aj3o400wdloW1Wt1xHSW1TxtDRRJRDtNrtEuFXiMYfzw+qalDkiSF0SzUujCyTq
dEqw7rK9Z/yK5X3/fFBgWztTLQ5bx08D9yDzUEy7tzFOKZZ2gvpswmUjvQHWtz4PLvnW7ZW8EoXO
YUctmeSTam6quqEz1v7COqmeu3ziwVbIdOX5RW+AuRRmIkJk1fu6Y+b9z/nBD2nltGyfgdK/dJxq
tOB1FmEvk5LlYKXxNStE/YCA7g9g/8Bo00mmnIaAJg6yoxpmTgcS1n55TyY2jeHddSTV5UgpH/tl
fPUdNNn3Lrd60mvRdDdFEdhgBsPRMu9q5xRCMJKSNR9Dt0tnuVKaE004NrmOc2b3D52MkGZMc3No
nob6Me7qM4QX+kM+x5f54OBNDfiFQeoGecSHvb4B0q34DnLIWwfSUG/Ni2e93UD5QkTipUC0N9wh
OkIznJyPD3ly5eRSdf1GRFXN7QTpqwKw0+FYL9GyepGC2k94ekNaBLfu5rffJl6Zzb/3pB+l+Eih
Nm+9Nl1/O9FwS1isJ1OWIUO3B3gDjlligsJ6HL5A3oYweRhte5jt7Zu7hyUh1AcT/gioORJgnMJd
PQb3tymNerRFoJvwiODaYRm5HKCPnsGbLLu9QK1N/Iz4c4WiJdc2E32mtNl6AsQ11YrtLoI3y1cl
GljU33duAZ3ec9VHjTMrll4ndzMgelZWGOKxEuXaUBxZF8yMexOpKenjKGcQkLp7uqm7Q7PS0H4Y
BeI8czva91qvQd1XRZ/+L3WE3YmJxgpL+TZnCA2143+jUzkVYpF/qg10KsA7FjxGAHua8hOpPEuk
Wk6IGhFzBmkDoU8yGT6zWZq9q5Avb1APrw+rA92dn7IH3WcNX5wMMrzmYWN4FiO63vlB4mgbe7/b
lAMlAXB5A4dHFidsDY70DqYLq0GsfX/fWBrG3Hz2cMNaJvS75Phxs9byAZTmtqqaPq7zMWK7qp1D
43CCuCIi/eJd5hZB2ID1DRRLnCIIMhOUX4qiAH6HAypKi1tKP4z7AkGWEuY1ZLqzENZsSLDD7f+c
knIJwGA0mXGsJAQ9Ddo6ORceDJfgSqfMfkogZI0roXRW+wGCF1z5MGU6jODczi2sxu5HISkZjbcT
K8NMlSRjNf2crwvOnGwQgiyhHiVH8BOgzOZjuO+qgcREYhjWihErLX220kpCrB+/WnETWllEjhVW
CQqDz1liaCBvafNp1ZFnOaZKbI8lWHo4kWJ85ry+LIviWZ9d+E0oBd6eIYS1/Ec3s46xalaBmNTt
CLlgge4PPACkV6XGQQAR5dKHvFQDTZ5brzof4WJZ+9HSbbyeNfvhMxJtVSD0N4F9eCaItovs6mYh
b09Moij1gzaFBHs+2r4NeG4WlXUdZmMNBdjSCJqzmHwpXIiBNGvRVl0tcVAq+D4t3o/7O2PkKnn6
gRymJCxYKyORcGMEXt+8T/mwMHI/Caxa7qQquEFV1tFORYu4xSA043uxP4747oBDWRv39YNzEvm8
RBSm8++7B91kuUbTHhNOthlct1+iqUuZTScV/JaFYcvGnHj2REqWQopJmxMmqgYtIZbnB+769McE
XIR4S4f7bAC0uuGX75m6R4SfSBzVbsZwQI/qMNOmVfJR3+0DVXTR81DOp3HDBF6T3cZWbcd+WYcT
GLgu51VaWiuj3KcnNTDntASb8CweZXV1RJhrlrDwx0Q77cL4VhgbuZuDaI3Mr9ZSZohatLG3nI4M
gFPWcIt3Al1QHGvX5wUI6tY9m/P13XEoDwOk0IHP5TPYYqA953EWNiOYlQhmLJtK4fp638X+jn3J
GY9N11aFoUY2sfZ83ReuqZtdNwKTwJWgzDytF+K2vU7MDvEDSA6MRGpYH0ceJvfG95uOMTZsZjfb
h+aDeXgA5W1vNaENtYiEugX1TWIrHpUtwYiG9VxNQQ6uKJGZC9AHmrEEcDeT1iVQXUqGU565nMxN
RIBhHET12NO+Sp5ir1UpFhdxOepygD8vxR2tk3Y8ASacKZs1inQz6J7ftwpl4zIvdsRn5r0rKxJA
UAlJXrj2BLzKR5Gt+VUHFbKhwSBDLEMkCQuduiDvjF88/pZFfTdM/dCoidG9vfdo47b2ov0+L/Dw
mMsKbBq4F2ucnGZwctIbK6Vt+aOwcYOjdBt5Vaqu93PmAlyNGq5nzZ+E3GvtyXAUeGKNVrdeEeXl
gvDaMwhLUwyZpbAniQvq9szlfoew+K3yJ/wQFQeO1ytOMDqcrXCrEsSykwDcuONC6Mu2uBWNQjTG
RGqmGAW9nmhO+wsxTgaprFTeyg1IwaIB1pCbSnVun/ysTlzWwgASYCvqy3aE9rIIJyratuKxmpMv
hvVbUl71abScSg4MHgxCsAuPqdwZOOyFJXjO8j6vVm2BHybwcI9SWAJgqDV8nDyIN9WLt3znVSHz
zO42i6rTPyTA6oJSYRMgffuSfrPO8kUItKmvpNGfsu/aYvzJ5kyzaZVZ7j7THoSRjQxJ+mBN4V6p
8/T5nbkyuiWLkFj8/Xx1ibnHrw1Sb+oIELSJfrqVkfI6RQLOUwGyL20mpX6eLMNXDJDn30U67D5X
MhDbpx8U7NMokcS0+Juwqwm/tJvUk+2SDqRvkgLWAgWF7IZ0rAEBOxJ8WP7h+Ks/aXRoXYgFh7VQ
WwP6F4mdPwo2d8bj+IssGqT/MgAIeglxsPQENekkx1vjN6p8JqsCqsoDHw6d3+ZlGLJrjSUEiGTH
BtnVQQCsgVVW89IU1Q27Xru2dh9zikc73LiW/HtFIGReoGhNP9p//N+ADUo7tiLblCIRhZgRTFv9
lG/3oFViaM5UEzpCNtRIVGoxuqEI3IFWZ2k94UQsjKopBbEgqZ1akQVXc/yu8adXCf9RyNlVTMD3
6aq1xq4g/dqCUW/kxetK3l1BmbUEYnFuzikvVr8/5ocER2b5jw0UJECjthssXAE6MHhHBGsiD31S
hhGcoZnqGfdprcPjqYPBZaLMavR+4EUvGRt/8eLkNS9jdtUAl3I/oNaa28tMWmho2GxpOOT2hkmD
4t7MqLrqS6bNFSOoonngB1zZuBy5/MzXSDmQz1dVJFXMhKQRY8l8ikomP2fr5OiwZW4VCM/ThVLw
yR48H1unzSpZAmhKuH7NhKX1DiKlJcvCRv8f80ez1HQaKzZO6jN/41xm2TLxZXLT9LHRiRGEcIHr
r2M/5UxWF03vdFrcMlStVhX2ZmLrG4NVVU/YvGGAth0yJwgiNE/7YofCWKIdmjDWCZugLZwa2bEa
flEE/VhtRw8O0TLDDCEG+ikLDcz4kjb57xLOIozjVqkx9QK1Xpk9amLHUxsI6+F5uLPOgEMO9dPt
Ex/cHZMHLz03MGFiiMEcZpBkM8HKrXQ+431z/FtVL+aqYPzBxWw32nuIG9wJj8d73bAURLOUQT56
c0ldsQsvZB5FcQ8rK1DenTucDQ7cQcejIELVTDuPxWTOkv6tRU3foRq0cko8UfjTVntnBjPC/e5l
Vbx9QaRfwqdZgtNRLNtIBccuaA+wobYuOs9z3WkSpI17aURdetnF6rCtxjldKcBGw/tGwmDQMYqM
b0t3UO9HFfisWGiWpGo96ueKGBZ4/34/KOplkAWph3OYR/WPS0A50OzgHnuZmwLnjncBm4S5ZGNY
5yzYQ/L9nzkJMBss1RiEc7P2pmt5kIzGuyUGmN6iIuaRvgYVvaCOSVIEhhfcPWGVHYtr/2YB0LXu
uewOALycbJYaZw1CvtpLNdvDSJm6yF0OJtuiXwxcihM89fIp03dtzjzcLru7KCgqdupc3OQ4SYqH
WtY+Tnir7Vf2n2VxulVarJvGcyMVvRNscGj41TjofHuCi4E68UqljoRnfQaxO6HWFSl6xJ5wDBru
k4P0ZZeu0r8FgzlHvD44nvcP8wN100zs6UxTwYheipjJu94xlyt7Y3WleZW3FNckVVhJfdEWknr0
3mRBNXzyZ6M7+kVNZiTf9gY8SY1tPH6mznRr0EVNRcpRl4kdtq+jq32nVSX3E8a434kRG23y7Qf3
3VjvZy1scVTCHkJAeq5HmNThrORJtWdu/G6xH/8LkKpBTJNRCmlU6UQin0Ks7VYvU/4A1FgKkBJk
YKGCgcskHBRKynqhYrB+kiewAWDlYWYAqF0As6VaLIK/9seqJMM2w/x2Ma/mwYflaEtYhcdohX3v
jZXPCZifhN/CmUYay8SoedKd3q2tintylHNDQ3Pw8hjkA9JKGeJ7klNObbL7jVVyks7Z/5ZMgEOo
WgGMuyS+54a3i2ZQ0ELnFMGdcCjnX9fXsSJ4E2cIjzAj6jTjGWVw/DTVuULloStgw/k4Ksmgizsk
9RckuXMKbsS+a+8aXqmdbZD/Yal7NgcavFYyboX52bS0DNtSrh+FuIVoedAU16coBQXmi9WM5bn1
CiUj8UPCXKjdAU8ScIcR3qKai3piAlS4TdBB8WFerlxb5JVrFFnKKSz3SM7K8trRYQYEaE+yW+mG
vD9je9Rvt4U2jmoXdaNT9lOW6Zcj1CcFuUPbJ7u8dNeFMjBn5eiX3deBmp/Ox+SXifhYHlSPFbfY
6lGgIaaO7LsQcWt+ysSSMtikL6wFGXDqNFpBYUAPQH2LC5i4ez93nq2o+Uh0K4lJDvvunkNNdhYw
7KLvHn8SmygA7vRTitiBsT9o1hPH5WsnMRXv71x8MWBuasKbQ7mWKwkow02ufKb7dhwRVU16lp9m
AUTUOHBzGimtaT76HPQTEixm8PCkGMP0vUHOh2ud7X3DzJEiHbJe/Vh+QChuQj8/txUawzApiwez
2fWjPQ7pI5eiDfTx6xIMi9S8HqKeOPbmCiLHXsfL4rU87vngg9M4zFagCR+muP++cMRwZIvhRVqO
v04yg60z6/FzlNTfnF7zM7KLebOhTvmOvcM8LIy7K467LF4H8UAHHVXCL+uS+7H3DmE3OBQAeIAS
89Da8u2/ELObX39T3k/HjcKQQ+SAGTaNBU3WuNSb5Um4pPg2t5KK/x0mii22KfrqdUmM99+prZXj
1j45jhAeetbzEJaIUFq4uWWQ8WfvT/if5d5+8RfaRHS3FmPra0fdrhdZapfbInTUq20kvEv2w8xp
EeaN4BNed2R7efVtx48q7A+uc2OD/Gf+fnbSzi0RAfogBM9qTeY2WoN/KuXH/1vTYQOnCvhotjh1
dJe8s2Mwcb1B0pv0jko6jsLI8p/B0jL3R+TeJxpoZdaAT4WqWJEj4NlIM33pooYpRTYw9iQ37GXv
9G5NPtoHs/BUNuzjEPeN1DRnajW4g56A0HCwgdlvdNxbxQImK5/2ZdQucPQzwWTOh5kMfKgqEkdn
Z87uHkQYwn0/d9/F9JmTWYzXoiu17q0EYGvT74bezfg+YGHkAEq3h1DMvaJ66V0lNOFA7D4yIF7w
pjacOkOkd8f6Dp4Y2eMyMDcu0kF9egDoxoRguDWuEAx0tm6evXmK/QaVVzpt3MUIit6iDGnaboF2
pWBzl1oG4EzXp8iLwOGtOPIPwTkceXEHzM7qppNn5mvY4Mc7CrkGh8bvbLFmSLjFSS1NLjgZ2ti6
lrJrxvWd2Raus0DHRaonzJYKuuC1yclrL7bjNrQB5ISN9QqodrOSVPcCnOCNGkuX7potwAy+fXF4
Cot8M2mIHkEzij3nsobYL75snPLjtJ9n/vzgr0HGoeGU54utUWkdBBK/Dtl7bS559/89qsFKPrvK
vd4DPK/zNkfWvnjZzixeIh17DrvTrg5dNrLpta43ed2+BTcZbSq3af6vnKoF3gsCuIrKcYfzRZ2c
u+0CVUn1pFUwmHOp2C4dgH8wakGNzHNZ0MXnvlaFJ1SUJm5GXJVvuH3d6WbgtrXrJt2xHzroMSmr
37uMmgVGt1aklt8KssQ0jpoUJ87qAu2ROBpwsqGq21pRInWvNmj4VDMw4RNWbvl3rE6I77bFdtWg
PEmLPBUxs93TbVmUwhCzfeIX0ByWMvxHldNJuLw8/I66tHBff1obYpD4KsVLUaRiMHVmwSHW+Kts
9z7ZzZNRGW8oL4vNrXaf0x4oteKKwuSBBxawyTO8sG7A7dzTPu/g4MK55u5J1KLA5FzQ/Q1RNbkg
WIIpfl5SDkJZOTrGmjqEGRT2/EJaR/95B6Nq7ALl+aM6LTMGJk3oTJhUOvnce/Og78DIpAia2kCL
QQ6REiChGAoYmCK49A5RMqcSeQQbKW9CoswHMDJ0OY4u3eFfIQKbyifTrs5++7ev3yjc2kTasyAv
Z2ECLoXPkXSborWwTz1Ehns/Fc+hOFW5OOBVu0MWweVic+78iCBJaQl0yGgQszFxEdkcE3EO5K30
SKRebNC1a5hxDkDAfbeY2pdsHjS8laRXwGxjyccLZh1AMjX7V/FVqbFnKUL0oofWj9JEW3+76Vcc
nlixcfQ4Q2vAee7Hz/F6Z0MemOya/ZxmKqGVzrlPjm5KqBmzxTS9lhfqefCb9MC94vSCGEueIYzK
U+LgBT3/ihvQottcvqe6NB7luEd1TCLrwzrZHRrDWOCXV8wn+8ytbp66hN47N14qN+9wlhol9GCv
sT7sAu7J/zfIuQssIJlOUbY1ZzfI4tSnsmUNDa6TfC4RTMZjwRrarpMgBvGu2ompgkqrXERfZPUL
PIuNCPoCax5BYG0rx7xpkzZY5xGILIsvHKOOe8Sgoe3kcijqcW4KtiQgIBdcp9ECX0sPRxmmmo8J
bJvOakGcaTpWWJtbQK0U65RmnLS5U7lZ22DY+PBB+WrrIkSOxODssjIHiJuIXVoju1+RZEH9uo0M
PS8kEcskd7gM+wpFRuKSkqd98aniwdhH0N4kacs+1Saf0LwivH4LLO36Al/45v9Ay6mgvvVtq9x9
UGetzm/jYR0sqRycObIJDeVzUmdgR7No7flQUFSfrLyMa1UWDFCfIGUaQpxB3hfwPAo0twL2/TKe
c+MDpLlykKrz/2fo9Eztk4pQ58JyfNk8iP5oXn1DsLX1EqXVzw6IeNeGABQttCwPwVrLGnHXB9n4
METBp7NtxiiWL328WPvHvHsNvcLMQ1lHcXpL8+5FoX+69/7cfGrmOpOPnM/RaOH6J9QpNceIixbV
DD4ExQwf3mwosdf8RFl2kFsX7eagKzVHiy7OxJTSmYYxbyD1AscKa8cQxJfRa88MNMhXRLBjFFKE
MVYcIGz0Pi4joI/qRARGwbCic9cykuU2ZHvnwSioTdAIQU1r6xMqCp0rG70crsyl0xs9KWZR+ngR
9BpLJ+9yfPDEOTGrtwLtsVto+b+IhgJ+t9YHPZ4XYx+SlPWG30nUNairBbGeqj/aH9L1q0Dr5KRh
3IrxYewkSTH+vda+brRVnVfDy3QOrWkQxVksvW+KeTmj6OTULK1j7V8kzJuS5RRTTSvxt5UJFviD
1kfiBXtBUr6HCYXp+JYs8qRhAPTiELE2ETOv4dbwbeaKgE3w6ftKyjXKFsWoevNGeFRGwpxWHlyw
ZkKAfwJtpJoN1rUKi0yRIxZ3C9WXQrYEZcVll2PvjLDQnvYHmg9tmjhtBQkPtyNROsYD/5OJsruG
Ar0PjYlb5nK/Eu3uDzDdnM0eUKVCcNsbCXKmwhbh2BAHeZHLw2+cL4lyQoPniaphMlFVTLThnrVJ
V3bOtkpCfGaRq6ceg0o/cPp+3vySrtOOHWR3IDsGKtVcNopqFwSTfJHczwm9A9kv5dOIVvNU0x2j
SlvWJ+Yh+bNSjGEinbiqAKChNjCJVUezhiOEvohES3p3UWG7AuSJ0BkxzRnliumro2gQJ2qJuUjF
vVA3T/CCobBIGan/waad/EuuYdumb+rlEaMt12pUEzNGFrJvfLK5XxEhefFxZV8encUVzkWFAFW4
Herpkij/Yfx2YRpnnqMsCE5ssoMzAZWEkHFx88Fco9PtG0cpwIgulqnChbxK26Fnk5xzpuR+pgRJ
nxVx8OL7kAdPg128J+ohw45Ev1vU6k/K74KxUwxYVHeT7zMoqMsgXYlg81PLP0/LLC33mkKJmlZr
sVfmHNvHQO/2H5jw8qgFNzHwnH0dne2B3PkOFU2FFYeWNgzSTNmTl+Y2qdyvCBg3bB8DEJCug/CX
MK2hNy4wV0nmMYsH+GbfPUC6rPVea0khqdlOHNXuVMo+kMR7nUz49zT2Khg9GWw+O87cNV0DnQzj
uChPPk+SpaRod39fP+TTWKTrHNfo4I7HKnDGfNePia5XfhxmWs+0l/Yz7hBpzcIMOXX+tBo4+sbH
nQBb4aPqWPwBUbYyOuAHJ+0Av8Zu3AtbgCQgPaWPMVHCa1fRubemy/T3s6drSPeYQMvbJRnn4Uuv
Are2ktElxx0A+wTbNnaC41uekhAxJp/iiQtiVVnYXuuKFtzCP43V/GODtLZvX5T83opXMI0yNZHR
9K7SwljfaBAbLyJOOLE2Kew6b3u5ZcwwvoWi+4cA+X6LgrB5eU9R62AvdQUUvKeCWAeRyqd7P3bj
l1vH1Vf6UPWuT9BlEZduf4JnECTGgoNiJ3Rn6IDSF1MRTeGYjKDaHig9FVF7qR9Q1riRgSxlgzLe
V9vC19EM2dCSgqlXdt1N2n48O9g9MKRMv4L01pNfkhGI6/H2GtSCeBBhTEb9RCCfF3QmHaADeyDE
7mCqf0AEv2ONqOG5hFX1IRV894UZKlwyvw2ClH6Us5abbQcUzi/6BfwlNEY+nbN262aM64hBC+zm
bOj+ZMgQZaTzIVa9qOHRJS4f00nEH6xaIzsy20TUlSE+tAPsyXSxxzLnHcE+iw8Q//mguuSwXKH2
dTcDzjLJwwTobzMRSTWH0DlBNPHapvtz91TDVkSDb5edt7vfojQprgbM8nzUbR/24D3SoRdngaV0
5vMjtZbjsczPyWBIqbkvizB+PCEoqzSlqb3TTTkUvJgqi0lP2y2BZBUFi/Z41nzkJoGxNwXl96xS
swuLf3VbqspWlGunpp7dL5qRM8+eOMoH9dcQCGP4p9LGBoQ6qzFaUi/yPuaDUD1hWJF5Genk6waM
63M9afCpwmg8fMnCYvmvITdEsIDtJ0WaDfh7gvOwqLcddFkeOEsS61Io0l7RaCE6s21xgCps5rsg
EgjdzTUYWPPiTgiNi5WPwBGUn3xq1GLrjf3zHSRMAgpFMQ7UZG9FrZkFtHx0wqfvU/DsbAuYVQhp
tSVuLiTA+F5uTf6HW1M5DWS2LABUPjrx63seKzXtM7tKZH/gNJUxBDX+NGnM/n6wR64fIEm5BPSA
EmcZJtqirCI/Mxdhfrienki9vDmu0aA2UGhv84EvwtxrK1XKzYMRIU5HpT+1+x/WP+0Bo9fPjGyp
QQay+U7sEg1rQoS6km9AHIecVMbbF/H4DQSlp/PVRuajmxnVrCvpiXUozf2Tkx2OsLDRhsNoqIGE
Ovs5ZgAmtP+w67HCKUD7RCGF0+9S4iKnDhdQZIODLZRLqTpC+R2IakxutgQquKPThKU5IRRyPk0h
PDsW2tKy3rCM9+oCYIS+1WhlPKSTX/QEAe7U2tWpT3Xf0png3fqc1kFd/IHOLvUXqUijAMpfyFWL
YNTwIPc3PADt6Pyuzs7C5rzTkmB88YeE2dD8XVUKmp7msWwvJ1eIX1yEuEP58Zvh2XE0aszJqJvO
IxEQwIHwjfUc0aAIbdzO5gJS1htbXlzM717vQUV3a7w4J5F4NWCeM8Mu2nzb7ytxKdd/HDOqK6+c
BgbSgzPZOfOl3Srxui/LNZLzY38e+B7OSwVGLS2ydX01vQX3zkdhb+iodCfgxYCsz70T/UjjO1A5
ws9XLosUo8LgJtyZASZgtoNpXKqdoWqXMYhvAaDHFAMcjvx79EW3DObyBugqb48fQCf3GO1ro2fp
u4SW3YWTR9vSahSWcu/hFe47BQiAZYOxYtXdfBu/71dh+mmw1YowmwNSNWaJqdThBb1UOuPlrojR
taX2GD9+5YH0xjv1jLZxJbULmn/et2YVVg/59WbsjvZG3TJi75I3un4VoCPlpa5g18kp5WT1LO43
d8ljeIM1IXMNDYImVaNTiH5Udx/l++523SbxD9w7uYoG19+3pieE0WHLE+pEWY6bOxqxjGjW5UaR
AC4Vv7dbdQjsI6d+ysk6WzRk1yHM4VT0fGV+q5T+yF/q/7UUCJI0pzqABkDCNem+3yut/GbTZ0e4
yTWdHwZcZ5RLFhTNcfDUNdNK+2DIIaqnjlVvLNHPZPVQiUOVRzlNqa1bLnNy+sYSPk5himnPcNTC
ZXiS4Uj4yVNQXG79ulWgdW3xUl74XUh7ZRKMKhi9+i/20bMzBpsimdJbMeLB2ffWTZn8LAhwqiD0
5s4b0ZMVRQoO5IW+RNWtcY22FQPmvEwkw/JMoOHdOtsK37uE9cMidFq1rHhbsQ5v9tTnX0kgckFx
xpmMogH7EovyHgzUbVfy7ehu//bZgKLyMUjgj6sInlacDubRp7kusxA47IDPrqh4HcDJhtqjNLtg
TIjxatEv7UWJmiptZPZC2mkgSu1LAI6150AO+93oEPC6/1tGqKX2zoIyFS+WJ+2IW2KHiQVETDB5
TQNbRe32OcUb3nkuSrGhUpoKjgBJNqQRCIqI4+cAPggBtil7j0sEU5DZeNaLXC5PiMf1HYRWA25A
eHpSxydPEyHgODejU4zdGyHRlhp7YzLSn3000TCGys9IZBuK5Tw5ed+eLvCetLf4fjmHnLizuEDi
fc+xxYLjyxZNDAq6/Pqx+a4ubo2Mpeze2cKOqxgiHaeqRaOi01yV1nB61iVHyjHJxgFuazVN7cyM
3+/YNkqoenUhjasXqUWuqqr3QnYO7bTVC6rH/ploWpHy7NftNOIlsV+zM+GKDRIojs/iN2o7/8HT
DUXIaxR6BVlMtutHwHePC7K2FxtpnbscnA2OA3dnS12SQkkY1rI1Adi+ZcUrt+8SYg/h9nw4dg0K
AXt/TpWkDwtOVwjqIgm4d7pLAz2oXLOpJxWhOQN32mVIPZq7FnV1bPX1GRWJNIw1EhEIyfKER1iC
sJ4pz5ilFTqffQoOzRRA7DWlZbyNWMwZQ0oPXe48fnR1BZIEaXLYQMGebHdmXea13sefGnLMzkD/
X6DAHS/m2wRatkwA/SPQaaklT45OnhIWYdGHpIjW6W5tlr3r6Ir8c7bgFEtdL32FDL34cFOr3Fn6
6mP8lxQzprDshNXuwZxNnIgu3mu3hh0eIZhRjd/genUxL2gv/QONFhqDbaM/U3J018xeD/iYw43I
7iJc2UYowh/3H63lsO6IPmjquGVdNQiRmBoPbPOXV1ycJJ0zz2YBsetNwBUrAb5IGhrJzo2JwHd2
Gir5N0nT2PGmZTPNS9IaySI+npX4BlLq5JzEE0XMPWKj/kF+M/CBD5cwlxUygZA6nrFoemjrTYfH
fVGayUnVuc0bo08NVtPFaBv7HrM1ZrLAHD2WOQMthQvIiiUA4Ut5lE4Wwjus7AOTcSqSsC8zr/jk
FKahNGCaayAdK2ppAgpaHfEN7iynkZ5tvzuwq+bwHql5mucr/E+prrEHfijwKwCNkz5hQWsTzpH0
SywMNeo/G3RbCAhGyCI9U3U9X+xgi6nUN7RR+r289Z9d9zK1tJTnjUhYBTEf7rrRaAgkRgttjZ8o
7zUuzEa2f4vV6DMjwwwHJjNA7FXb9lJ9Xtat+xNk0IadgjOrsJz98LSN3JUxgRkWpYv1FlOQXv1Z
ZF9sHImSpDFl6Fdj7BRILCHce8dYsVLAUEJJ9qt3SaE93MjotHjAKXQBOoctaapUorbfxI+oCRTH
hK8ZmixUojxsglANO3gzzWjQPM4j3yM4VrQQwBRroRLy2EL31LG93Hg04LRJ+dm52AnyEmtQv45s
C3cPqciSYifwrlsPVyOHmvNTZMUgoMvKPXSUWKkNZht1H5iqGiGO5vw2wSDGL5QowNj62gx6Pq5u
c5riJdKUze1FWIIF0D6aT3ocqlJzLEz5yZ39k+xBmFz427d4obHdKpZ0GVPVTLpeDgpa27NrltpW
oAeAzV6Qv8F0k0ihv0Q8WpTxtWztIJ39qZCjdRBX98K1EfMHSJx1/UxTqOz1DJFaTlouWO4RRmZk
/F1PcpXrFESdnY/XU/p9WSg8uHA+Chr1HD80T+yu3I+Qb2Cy0hGfoUq5j4sLP0Pv5mOYLHiVag8m
kbPez4ias6g4G/t/vegdZXSv51CpZo8nSmRQ6m1vfgmDknZvPc+N+QLBgiURe+Il5gYLC35S4Xc2
HBtTDOvARjQdPWl1/Z11g7t2CBP2phPe9fNnGXw9x7t4hjm1LGXnv/rRqNU4FOuzFSbNpMe/KPZR
fPgSpj1VcifkncA3LhDmSYw6p9xAi/VWFUoUEpaXnDWsiF7At1NG3FjAG8yQgtHK5fudMaTmiSTR
E6Lm+88R80m47vKmUJIWDiWSwtTs0UvYiPg2xHolOmEiSOxN8PZHzdCuca902iSZeQiGDuchSIiy
RdyvtTxfdJXg/5daDXBNknnNTepNANqowqNPOZlYRLBmSMKg4Q3UakLaJEuy/BIedqymMU94Vfkl
72oa1A0D/k5loCiDS0AorhY0WeIyZBP1tnQk9jL43umG7Ar00x8MmU0GIOc3g/1KbkYF8nFe2vhZ
jK/x84qeMnRsjqqAy8+37oO5Cv48zsJAOanW1zSHUJlvnM74PwhQzyDf2UTtuLbaF8jw8J6w3bsy
GRS1KWvBd8KDFLpBbgf1tCJ0HUnuQySw4mZUYn8r+lhZ3wx0qeQIICycx/fbR9Mk//eJvB7ro4J2
9R82vjNwti02xmrxt4Usm60Rr7f5XiE1O77fQ6Ck1u3IYLJ7rVkjEUtxayZKjQGMSI26JYwg9t7Z
oEB7Dumxjwpx64/H+aX+P5dTfaqq864K3wZdOct6sgOa4nyHy1/Ou3tbM7ogfQwF7qrYF/X5whpf
Zh3oSzPwOVWVsiWXoE1wWY7IAc1QhduZpIrVgQNwP/gOLvRTyFZ/VSwGZTMaz1ALhyI/iOIC83MP
q0xC8IGV7PDTepbKp0eF2ine1rv8ETHjT540A3PrEEMzLjoMrXyd/5QoZ9nVSLIPnbcwUnwSZI3H
dp91xGNzxEL3SYYm/mhfpPo+V89F0iv2ZfHpNJRnt8/mvSXG6DD/pQRSmo/SjUyeMD4fuyRf9Hlp
LPTtumYpABtL2rwQR1XyigvVndyR694dwL24OMhzO+uBO9Z69czJ6mmHQjAG3VbRcRuao8y5rVtG
XbadCEW1UDiIBzu54dkFjgnYr0/kMtQvXPQ1upImNa9tNWtt3rwahuj5LahoRxSxWvmEr1+/DgzZ
LbilGs0j2+L6+8aWy4uJxo7sNQg3BXEgFhISOBs6Y/wNkflCBr9c/zX20s7fLc+i5JkNZ1uk0ueB
rvlGtOz0jFmwQmhk12A+VPvmDU7wij9LpWQAfYtHrCnJ1oGz+8pmViXhfWaNGbbEBypsPU76FI5D
ten0KjGEaOPVCRAaCfQO+uJVbFVIYYTMNw0/OB0v6rMSZaGFBUvpC5L4puHDqJNgwgEee0/n4xRT
VTPFwqS+39xxZHmgJ91i62yU2kxsyIHgQ9U/jRLJgRW+gy7x6NJa9JjB8er8WWXS6QY5UG/Gt+g4
R3w7eKB8U6S0ewORdB4Pbu1pRiQomzB3ZdO/rV2uC9mWdHp+vPkazsw6y6BIqq1ZeeZe87LdHYuE
w0EHE9rfyMJx1DOrtxVLhy+d4+Rs4VduSjd+xdgz4+8GkzlibpQjl2ISSTc1oN1T22rr6rr1Riyb
Kn4MbzQaVU3TU4hgcBr8Lxpk9UKxLvgoA2B6BPG6RxxDsCU/3hOcK3T43U+9TgV9cEF7MGu684og
nPf2kzdUEL8ijTRpfwfd9wRJ27DdbDfbkBcWzM1RX6Aa4hR1Zl6h3+EB6ERzLKHuukU0H6HjCQdz
TjZio5qJ40QKRhGsEFERZ1CFs3TLhRsboSEi7eFjVDsau3Wka1VsXjC+H+HcxL6omixNxPLduWHA
S23j205+aWiZUqJZN1n+wrR+sJlaefpJ9NIZMaf3loBDq+Bi0WCWGsWz5i6cykkoRegKVhAmFUCr
hz6tqKfLhDFMx2Q+SrtIXFpJw/KVzmZdLELB7R8S4r2RsC0ADS15r0A8FfHZiFTeNo4eWkFmUWMK
72b2yem/bYGQQRnv9Ue0dh1w3nU1yDFDZF0RNKVNAWJ/bHgB02Yu86jbpbZBnTzZbxmj0JJIck8O
3EcOw5wmAwuL63Vx5NaQ2DgyZvHX0hjFCBxXHK26EuYPBNsTXbwN/ylOHmiT7Jmmiq+fO+fT9N7o
evjroYWzufVekY9PpHeFNwvxLhipLS1GkfDFeY61R0hzOu6NeWg6yKZACdhvJAFUH98U145MiEO8
0dJvRn7CXjYWfXld4fP9Z4Thiwdoz7Y4TL/ItFsPZANjfgHqbF8zBIyuzqre7xChJi+/2rsUc6z8
zrR6UuPuU3IOtXc3p+DIgBF4FePgIIQe3+qobSSerXfyqBg6aFAmxLWn+4GxnO6AGag9vy5mEEnm
3tjZ0/wX7HEo94kFh9uqEkBClju6Qs06l8/YavMcbNFH+32znUR6a8/CSdua6LCOBptCDvVgRKBf
LTX01PPaXorB8LFQQ5tN3gb2sJncjZ1AEfD8U1XjMy3tF3vD71V12s3S4ByZlzR+764MsweiTOEK
I1PccImzk59dpZvliJ4Hq1fyp1+f+MuaG82TSwhxgzzGQ38Kp7qs6aFiasgO7N/VVuzL7jJpw3sH
28wWMUvuNjqqjUTXwK/Q0tShDO3K73Z3xSfSmISAUguOkdYn7c4EMFtr/UZEX7q+DAbA+Rq2T0Oa
AX1SlNoKEEvPZq/WUbUa6U7o2ME/XXdzcgW9B2EFahDGEVSYttd7lraOjypQwdYNz9mwo18Hq+w7
Ks0/M85A0lMrXhzg5pnIl64VeEs5BZHgt5zFnG2YtaKwbrk8b7eA5kykjtmu/Jg8qFft3Z5YjHvM
zH7PS+jc0BbjY6guzbcRJBmfKby2l8qiRutbrSH+QyqBGlUDuvD+pDv3xJOymBExkDbXJmBmLb1R
AUKl64e62p6hBjJsr3f6ttQIK9OD95j+zZT72CHLGFqnT6bs62NTfBlG6lUfeA+szqGjLh4lYZoP
r04ceq8M92XwCAgwrCgGjA+2aZWje9MfCdw+HOIOBQFwW5zwpt8p/wXKXgiGGurTQaVvTrzfmcZK
TpotC9ngUb53j+gwsemV4QUoJBJBUOkiu7bJH5tMmHUfUJIUqoKEaTQ6f07KWxlMyGlkx/Gu5oeg
kn60n2RC6MDtZ6JmUvK5mXFICsWWcpBvbC7HQmYPqBiclSE2yxiXSNfOjw3Wuo0d6Koqnvc/hRMW
60jo+3frnKn1ZrAJnelvf9jn2O51HdnfqJRxM9oqUAixWhRUn0h6pBz6nQqdNIzvErZpRbPyiyuh
oQRH5HtXuXz0JmLOK8p75b/pf+PD9z8YzayakC7OcPoqNldiuBgvikesrdB47szUvhrGIU9ZFucy
ndZX5vXAQW6gzdL5IEs5ZwJ2z9fb/8vPHt4ifYxKW2eUAspeker/m1vpOIl8PoM6K/452HnGOzAX
luKE7Bvqs2daEPprQVEt4cKZdyucM5rqMEo4qfxFMwHRvjbm487FFy6d9hxgFQZiOvQUCGda4ZfY
oDXbinaC/MxuTQ3zLuOrvSaRANvY3yq2yNJyhhLxt36Ok6cm/nl7ax8FvqY5eKwFR/N+o2EFJ0Fw
mGQg/V1xdum3JSJaiPceqzM2hHOKoSMAvDbxPeZLlZsUcuXuFkM93D5yk2kaVGmQGWhvJFQ50QWI
4urv07lEUM8PGRbnGZ+ZWON9w2jWi/bnChSpI27AuX+R55OOveTfmg0Kj8fXmamQtGMRIGyuR2+t
TSMwaxml1WP4L860A3TmiRvggQRGcKBfza20EiWAdCy6231MYgNHjl/OUp4SMGDr+bdFPJTAcR7a
IT0mv4j3hreKURL6W6aksEW8Sozeko4dFZli5v5xsFW0e0Veoq3sMJSFY1vAzuluKVM9r1DckFZQ
FwcP8ez31OjIeiknrghTiK5QisF1N/9zEhQsGgjlqw3wXliCblTiJSI6wvnqTcFcx2WpNYuQLXRI
6p51KaYDNqZ2PP+1+Kp65hLN0IaUauXUEJuQhZ5mNXCvGTaVX7V5hW7etVp7OqWSwREYPqVo0Nf2
G3MG+bwyOjwKpt5MeD8ecfb4OmAqKY6LLDI6nx+pP8V0x4Lkl/vUQCKEQIDSu9G1aAmi+FIpaU6k
VMB1i93mF9L5Rknc46S83+oUpusxaOk08JC+/+47A1yqSAVF/G6IYau0iCzpwovtVZddDqW0MjgE
wkE2++ILp9C9YfGOIlvqwy8KyPaW52i0yKfQBthnBXjL9b5OH3wt0GBs+dyDQywl+qQ6c9m8205B
HWhpyyGmaVG9zIuj8jFwhIwWXWhiBw+NHB44AqYT3awXz+WSxikRuqfVqvgfF5NqMEkp48mm6B3y
QGWKvLIpOpo+a+6hjv50xxDpmLNZZvqUZD+HYjhdMYoRysoYnLXEFA31Yup+ZHK7hIMhBPaRiDRH
T8+1IH7xhq98wln1bWx46fZX6cfOEvHaf5VX7nNUagx0iHNtt2EvrFGifGNVlbqujQaBok8S9pa/
TyGHCajHzgbnE4KvLU1tHdjHtpnT9zvV6W6g4bbmKn9OoSTUYQubjULcojc9N3Gm9mTEzbKGqAbA
WSQuwUR/d0QRzjv/ZcMuHkWF1PLdf9AVe0ENvgPP5NnVONFJ+rOGqueT92E6u1BztwRfzsXvneTu
K/Y8qy48ZYk2PugiVK+D2u2sax8Z5GiB53+HCUZHwlZ8O6pt4+nbwBo9kBdRA7vc2EegrIFprptQ
xXumpS9UWNrGdyX7sgT6eGXj9IU9STlBlraZtvRkO0d8g/fl6fzb01Ggc+QWYcHajIV0FdHG2ut0
6rC2KcZp8KyJmHkNpfMbIO4aQz0WUu4tIjT1oFYs3zWl7qHTFr7tph80ah26aArq9XKZ8AHpS8Zp
ZIdMxcIGhfa+Hf3DqRaoR65eTCdaPFSPItkMcG0ZWZ0a2c5NvkO3tkdJ4pJ+VBFIWbDFu2+Xx7qC
8j3az4SpDVQUxunyqWJOCsO8KU1JEWRHOO2X8t5yQlIUHXCsOBUp5DYavjpCrngXnroXHZ5A1135
hUTihdndyIIko8e5rA97+6aJFPgzEaysJ/MiOEiuNVlLo2qBakVw7XLGFTcNsTTELkpLgNVSDzwh
7hapv+9mNomIiJfkUeYfG4Va0/s9Pwf/r/yEZaQIw0c8j0m8784wOsZSL1o5aumV6ArQudl1bK3a
wf4W8kzDhGp0Z3Df0IkSclvuMf5l04oOt6JW5q/1bk7pFEvoAHr2vXaPUx6bN9ddnn5Z9rVISejH
k0yMf150NYmj2CDX5r624AjPI1sEe0Agp2h6/SieSv+ZLMoILcIoeuaDIjjXpt07r0anpqPA/AqI
65qV+Nqzedefcs5y9IU7ypDzSvQ+ZzkSHiY2BavE7bStXKFParE3c+0/OyckY4VI2u1rjbsaiHX+
uhZ37jKJm3EdGbCT49hf0mr4HoTE2sT4xfp8Ub6SRnx8n7RUbiBq0knlfovSqAGH59YROVisw/FB
SdtmTq+p2Q+RClqRlKxChJtysJ7clXBoWZb2Gt+8r49swUEwoi1J2AmXaA2e1Un7L3oQzZMBxq2r
Ctby2r9vudnKIyHwoADBR8sOvg4i6yxppCLPEw7VWaxoKwhNeWkIt1jn2NjM91vX2SFPpMCyje5t
sXEhLkLLkIUjfeCz6vAdJmEVHOMVRxdKSa/dCgAdR0FWq0o7DtN4uWsCoIXNJPCqISGAi009SkV/
LeJyBWGHzr1GzOblCW46Jl7jG4S+hooq3FQiEOxIjq+u9ifKXRFMst8sT0WS9XlE7KUWKwSn4/Pd
uDLH8FzaNSkCvD5o3RWqDArCOP/MGpmq8PZ2TCM78qPfy6qWQLltJor5aVrK2XCMDq6ESo+lBBz2
M3Xmxx+eUQGcnUa90sAsmF99X7r9Mv/DhrfFVcxSqcz6OuFmuV9GNUaQeozYMaLTBrJIbWZIgK61
HNpOjkv+Zv6Ai3Hwy6vUyq75ReunPHejx96EHjMuXCchn7+J3eUEN+3V1rHMKcx+h/4gB22IoMuL
+Ce8gbrZjT7mCBaBaPAkQEdNqoypLt83m7kaZiC2LlxsDb/iatlCaauhQv4hVWC54A/B2PiPntpI
ykC/pk0EFRX6TZ1XU2pwcwgy+5dK3i4HbQ1dnm8gWoTuU1w8ApWZVUY9wnbFuE6BbJ29v40B8ffo
HpBj6u9MdvEDFgU83hbc/QKrnKiHYpFZfTvaR5GZtbM8Drnjh+ylgJZu/8Pk+kE18gJ5ULqtzO5p
BticPCiwjaSoYHP9IoReP6KTf1UzlTdvbKSJWRz/ck4BtmGH3trxrDyIei6zDnY7lhbo/Jd8RC93
0mWcBpk5HGtK7UGAfFPJxwdruLw8vTX3FTEzngJRwtjm+fI90zH41tEkaq6hVhM3tnMVUzoHXnxE
QQOi2PP4ssCGub2St3pBh37aShhYqETji/XiI9rM9MZTlFXzNqa3v7+3Sho5Jt/0CFeM0lKAB0oZ
yQLtJ2KOQqTSmUS7ZvWacCWl8/2paXYtZWs/ZEBPNC2iO/W/4nWRMzsv2RJ5/hDqm2K+eo2XBBV4
8oA+RYj0c7jblerVT+SFwfqmxm/UwAYZd5I+p3PgjbUnkBz/JtML1ywxO4T6jJ1UzZWDztwWHpy7
eWNaKK1g6TTWbTG5YE2zKOXlTjVBKYQJov6Xs6W1xIlMOEVa4lUYNQ1sxB6MXHUZyXpE3kDd8YSD
EZLt4bE0g3Cyz2E8ICi5chhl8P2J3+XHAIt/78BoaI5JOC+scScfy+9JuQBvqVUTUJtVHlc1cyOo
Jr5cE2Ek65Th2bvr3K1ie2JgRoHdV+wTAdsaB1XmqsRsfvhqxRGdQyr3pRNx6OfDv1WfG+dJGwZP
Hvr/JUQdFUh2hyu0uqyj7dULg7wtVzfQS/4RrDYtHHHb28n2XBSzkWk8mgq22cqCNAszEMrfc26X
+Zn6mYsNr02i8XqyRy1O3K/RJ9tuSOajrXgNvPifXP/ctG2AYTW83u/r+vU2s5tylQ4H2ZVh2EpK
eNchMskU3q4j5+qaa1ThJHWj9veSIJTL9Jv3iQXRsDlv6XTaDQHGj6OGdbsQIVF6+saAMwhRWrx5
jOatk2GtCoBP7L5rWUQDeu/4c2WZk1WDH+J+JsaazIA5XPTHCDcsUfP8tZmb741L/C/kzSGEFh8G
LYKyu1ywVYdfPXYBhAkTjzv3vgOpj+WmeNzaf8Cbv6fX4S4jEtkPkwI9sMsm3Wy+DxMAgChcKkeK
j5wqVDOv1jl3suq6KDCNuds0JQH8OJpB/TP8EuTGTbBffIKM8Zd04It32SyV3/yJG1gAzV43geLd
xDTnLDezUrA4LIiEEMtlSl/mj0raubRpboEslJNkKDEqlhY8rCU91IyMgBMRhYk5LsfIj9PHmkHB
SdkKYpGaOWZextKz2kIVQJMbUg5tP5Jc0hdrU4dxZgVPaKzge8Kt3E6LMf64s4ny0FGv6MM4Ue60
8oaGXObGwQpMB73q4yuxh6o2WaI3d5R7QB7a2Ju8UcFIACTNCH/1a0IQvSBOSUgDNvLULjZ3qSVa
Q+WDhdNCqF0Woa79I1AxsGxQXegCGUnmZIk6FRwYSNcxplzRA/8CpfFbbfQzehnUEZWPFrC4RZxk
8q8h2gEThRczsInwoeaEcNq6OORp/yRykku0GOeGYTDP6PUel9+IypdUkMf0ijXOyM+axgF5HNZC
50ONOvcc8Evi8KUbivhdk4zh8QeZ7w2BNxhjB1TwslUJpec8hQ6/zh1w7dfzJhY3gtT1wRlRj1PK
YLRpE+vxNLXXfaqJvj0xQZYV+cTkK44uOPhq952rxyNdtyFe1R0VANtnq3oSYn6NFjQDJSPguyql
8WGjFnaWqy1+vA3M04qqi+7jyAQNEldzbkIqlASnBrc5gBtFnJIMbZ4H0IV0g33srNUv9I5PJTh6
+AmWeVo1dw4GauM4vLyVz4nEveK3PfROxrQcdG8GukQFnoYRahKStPg/A5tr5Mo0NVJ1UW7U1rkg
jq0T3dC6cH10QH6m8VRwSuc/461i60RofzadK+loA6mHe5FWSm1Y/PADbQhGBbiSgDFZBMZ1SdW9
Pr7E4sWdyjfjtLqE4G8R/YaeOA1fOBDzvGQDQV9Yt5d5YIoQ+SL0Y+zs3FHXLXJ/CD6ax6BTr+zC
oqMLT6IoKZUcihm0KZ9cAFis70Xq4SZJpZNNkwtGRZmjr2djFs2C2xWk2vBYvDOo6dULNFMZftGP
/PRmermG7cAkQmOvhOUDLqyD7qtXNsMZFxlC0dRqjap1kPcNlnwBTCvhVBhKNAPABRPR73uusw11
V8hZoL1Tog8blwMbWYz8+A70bDj6nazAGTwRZcvKrxKliWiLPjvTmkdUVYD9UcwNowZa+LHIHzUB
eDvzihVAMuatx/J6E3yRH/fN2xvckMYJMEjCVaH80YkmckKdLdhJ+cSGlFVs9MyepM1MTjPeDkn6
NgDhbSuWnG9vzgwbcwsI2+pEz48Bk+OROZ9IgoyGwDoeR8f/ckVGAtVc1Q5ATpXUp2AMsLsqWSad
CO2D5F/8wexRbs8qnytJ2t6OlGwHsv8UlVyvwZMKfqzbm4xQ/o2V2BQSKlwvFaAFhRRIv8ERrkDy
OzfGGmZnfhUa2AMOWu2RL3JU90xBcHZM2pZfqZ5HN8v4sGphiXWySKjALdviPoGw6fahPUA/dZ8a
1yO4jHPGVhVbrXkUC+U3eiqmuxPOe60Ee3+YBto37GqZQpKeGAfzpeqgBaoeTiFj7FE4dkd2qrne
VklbD8WGsOyh7xchvoZvXW+v6lq73VZ2KOzimvIIZXm4GO2RJGTaY7adxSxJU2orQUW50EqnpKUS
Svun1sS/E/y3e2+iZdRpK/YZViKyqKcgNt0hBR0BmA0EJYKRDNYyikNZXt2zhs2mthrHECeWdg16
/xja97vHgm9bomfV/lx4PI8XH0MW6kQc20YNa6H/2HP4+hJrwp3mCyVER0slC9n3x6P+BcdMnjj5
HnAlRnYA3a64XmWtO/IZaXHrSzOOBg7J3gvDKFXOejeCuSN1hxlq4PBJmvwfa3t+GCp1Ay0cCHll
nX0fHKgv9H0JylLrYmWanlOCG31pzwyy4IO7F1q4aTP4rqjYiGn0UDrnkoHWN0fl5byzCRDlFwXL
fMwZ3QJKXoB0+SogeDYsGNdK/SrmwF6YguTkp4JBWdJVzZ9kz3x1JVRd3rINzep5tToxReqGRjVV
9Kq7pf8+JZl6Q9XRzWjbYusfCvqC2VBz1CPu0hq1mYyRhf2HmpfS9HAAvnYBReWCXF85pU9ZwJi5
nZc7uBwwc7NXCg0O0Dw5+1Yz5Y7xsEXcevzXiI0fwyOlL6DzXK+cibStHgKo+mDUAHsvhaEAXEwr
wmTPwC/nn3fhOPfEjDalUHTUx5UZJngKzgSlx2mjCvwqfkvX1tVCEpToR/sFcdAsUaR7+5oARthR
z+VfaWE0ndQGD+TOIQuMd/8prY0+6Z8y8h5XVHAhqC11x6lX7rFhKHwhm+0AuE2CGTeEcl7wdFMQ
oZ6iGCFxpPWplQfP84w8/vF5/47F/wRrLX025Wc3g5tY4GotA+zuqYEo2RPJJ1lX2chWMVbd4KeV
fSmY6C01kraNMNDsSNs6ljV9CDZla6Nuo4mVUN6wHFbxwzVNr10+t5gbAfdQbv0yDWgPcXmacdOc
H52nfSpSFw30Dh+dL6wbysysOCZ7/wGBTB+ocy7sS16RSoC44JBnj+3SRqJFv84V25FE9Kue7gLV
0bP23m9l+rKdXZkUEgng3SOghbTpetD70CMWPm3wOBTc65vnzyUea4brV9KpoAAenx7yJYLw2bUY
sLBNrmb4uMMc7AmaRsWRHM12N2a7dFOQlmcqDntgD12TskbAqBs2efYfatPofMue8FYLyEQcZm5u
j+9Pcnz7NZNfoVJpdEQ7Ym8RvjFalR9rI4WJlsf/ngBFp1M3m4wJxBtmPrJd1m3FTZXvKAzaPXhz
o3G81dCPh4lPXNTI11OBcJnADDFXJ9Ixi5qkPRvRpK2fUh3M9YIpanYXYYGsgefEPWBlYZZgP5pR
UfDUPOQ1fmPQU0mDOZW2+RwWqW4AE5fRF/O4d0AtBGRWLvgugyan8uKcv33EBeiGy5n98SXKjq/q
1uiG9fyJW7QIaTdmCy8fghvvXskV9GAx6y83ROu9Peln4m23JEicK/AP4KY1DlRVJNsov6E1BXaV
ci4oODLzlAG+arGqqe52Mf0UkW8yBfH1Xa9N7xbzHULuqobRQZlp+NQ85CzDycMWWnhFtPluQrI8
e5PuuVWfPDm6aZgaN/6yKn4VSuESYFBylCeB9vop+ifXE2yA05XrvN00Bh/A+FH3Us105qsd7PTC
K/sJpLYTDntVf373YDbK1vd7j4J/pk1E4O1Ci/HldPocDkWwKkjtOxVoFIHmhVakYYvN9Aze2Ljb
NSrofXFfTl38lKQ19BWiyI99VCghOHy2l1PRfzANqOvNNaALDauAfoqrMVB0JWxAgoHYAYd53OJM
WmFyEwty1HRhfTaGO+KSpxQ13GJizMpP69j3iOP7GN+0wiFu6HyKi3ijtVlojreLaERSBIQDTHTW
1EOYxEM4iTs9eFZL0suv+VNci0uUOvLwPDbjlkONaO2jOgwJ1Mn8Ga3wsDcxeKpuZso2CxuwsMVX
IvPUUYQKu6q0SCLefa1LeCumX+669GTfcUI6N+ytFjAtOS8+iNfs+uLgPjhJS3CTNlFnTgtVqDoe
9HRQKCKs+MpOK8qnKPXHMo+6lQCMwZyov9nC40iflYrrLHSjSkrYCkFX6tjjPETl/6r/NSQI2q6d
PhJg5Ur1KRrtVL99FSbbR1VL7a4d3FHu/Hngq7/H3+rRgc5sehN2UrXDtIwUAUOQVRkvm3L63AM9
SEqJu2waKhNXWIdJ4+REqZpre0drZm6yiT2wt6GTL2buBRrg2RyHC2F9HHCmHU5x4y73RmxP6rpv
+oMGw662Byb7DgZlmu4Ll0bxClVmAdUYGDIiRlyolzOwyUhHJQrBUvj0Iw1wsD+hEggnVuXTMvDH
ItgoDS1/xlXbnIKEdQ5BSRiJt5vum0d1i68v8Lx7cO9+xmgJ2VHPP7Bu65EWXQY6Td5bVEP60ysQ
xQTzYKo63YH/NfuTqm7jfR53sV6StZ20Uc40l+2nVJmxsrpti4uV2HE1xeDSvuZP4l/LxjhmDT7O
OkLilWfujFN4KZ8eWAqHyYbeFNDIsTXGtOnQDS7Cy/qk/3rRg5TlfPK0jTzi6gpMMKY0PnSNYenH
WPQgh3QBK1pRAuIuyJRagGl7MhM/P589Uwrg3G9ZlDJLwuPL6tROPcMC+uW+60ZwcGoK0a0F2S30
Ihag8BfY+EtbcYiLzVWPQqBeA8F2m/rBkQhSeLb2aG5WMBpzLTi4Ia/cTgqbtIwM5ULicgJVJu7x
dNtNRjoCa7QeaO1whhfRVID82y9MEbp8kz12GVDtEL5quOQySa2KxufBGyaiAowZjHxOP2i6kkyO
yGsPhVPzh5YvirxSUNQfX2vebCSaNYN0btkg9NjNR5OKgs1Y67fSZedlBA9NvsmQCMi9xpcWNxYK
Cc0/qoDRF43d3LrOvTmVVEnjGCWtCOVbPMcXiTSIdE3wafno+rtnBLloZwWHkXHssgQ2Ojl6BK+q
N+HyHi5V1DycfjvPgFTkHswB2hLs9I3oRIIH07iWLLyR3/ULqqFHxd2+LFYiyufuCtGWsrcphgep
yoK+FQm7AGOFW9znSa9XzxoonC4QeJW6RFB14FyUwCm5n85r4rXXgbmIsY9lknivPbLwCAsAQpgn
sQZUyrWBvXKH/2DL4McD1lTtzUYH+3tGX+qn3fLnu21V6ZzfRGzYqjKiHTPfHMmGKZCpWEVeP6QJ
ykg1IEzhU50VH0dzBs3OTAka9OHCDojIaIsReH80LKxDo3AJBhWRJdwB64UwAajPJ4w1sre6ZRns
c4do7OxZuxR1/D5//3Lu5MBQ27vycIo+8YHDFvdvtrZFYxrJFYv2NuwsgDChQTvb/mmXv4LzgGXh
yorb4b8Ax472f4LLAPEq/5KmxuUzQ5bHBNKo4vy9gMnzq/ZnXrdZpe8INjz0uniYu2iIpaKLPiQK
mp9rV8rywgMoOErgKr/fmW1dRlgHPC6NEiDho4t5i90zxCAX7cFUS8jC1Gg8XSK2Iq8oa9FUAcgD
68q/HMjNQv8KusRFbWWi5KSWd4f7gLAI1ywsBsPhWzb+GHp9t6xkRZ5j8IKVaZhXqP96Y63nM5el
XNrWp/VFcrq7IsXDgOUNkTmC3ZULOQZLlEGjaOCYcGKuvKsZ7cSpQzDDOBcnHlwNcU/utjQVbgqj
SZdGFoM/Y+AZUKpY8PsA11sPrE717ukEnhel6zwP1ScKoBPN7NPMaWiP4JZIyB+PtUTd/pfnUYIZ
OEseSE/rJlcNeYgwAGK9/aI0bztVFy4jl3sTRUT6eBq0UKoHbA6cbk5TbS04uqfq4ndUPah3pRPA
uiWaq02OgCQUlkTeGJ1FDB2QRkxPPAFFl8qLlYhkzpBBxfTTgSrQ1Q97yogPP1BUu523Eko7Qn2D
XvNvGqdFGYBJH6jimTAV4cQKI8WlTArAJHDMP9nkjcHNXoaY/riWor55Zy8b9HOG33KHjI1ZXffT
MIBxlJXutH3a1G4lt7gC9ZV+esKanTL6RhG7+WlzwY0IV0mxlJoy8g2qS603CxKi7DMpq8IwrEcl
qIQxdhfUT3YkkCQEMTLMzf/Wpsf71HjVW7lKcGuS8E7Hy5IWeknQ//Yv0Vydh5+mMCeCyAyxQvTC
NcRjDknsgmCJCH2z8NE31VLDG8nGFWQmzQlfwmvzj477tDCSwXb2VF+R0eRmFD+VbwU/upAnEtW0
6l+TI5PvWCMeAL3b+JzMbeUV+AeZSakhvQdZoY23RRO8/v72Ek01WCYDP48QVlR/dPdrIeBMRPe2
yRFl8OWmKVRrI/U6pYvrNn4JcKhA2BbfzE6cPe5l23L4bTYMCPZbhmlm5dE7dOncZNAekrxKoveE
9brE18coEeTvXTvzUwXhNzL2Qidf+TQu8PJY+sLmui99N0XIWBegFQOHEd4v2rNuuya50urDrAuq
aWl2+ThaHXlrClFkdFPZOvUC6/CJ1OEZodPx+k0h+UZeP3gmJjcGEjQw5BBHrNn+xQ7Nmkuelrfw
07FaB4gSHw7NEJB0q5Pkm0hRl3UC/LZwwPFLolXUxZfkdMfe3LOKHfJLyLo+SbshZjmefHC3ekNx
fKLl2v3vaOaZvIq1YTAz1broQkXWG+P0N1XUHJZEGNiETLm/1EONPMxudtQnPy1sYV6ChdTGV8NQ
rrZdKGxxx6+V5ZhIwMXDxvLUOzjQcFhOul0/0rE6EXm6CV+IS7boSqHAePUGiFAtWAPQoeQ8Pj68
BDGPFIA4X4lBLgFgxpH4FGDLDFcFIKPp127U/38RkKcjxZuYyu24POT6NzqWUyHYwn4C18JpHXzh
Ow3kyWxya4/G2nPwHeku+kICK7jhbTu3mZjPC0ysEUM+1EMwJo8O6ZC61qI53/zVSealbJsznIQ7
H9tC3pKFQam5XX9laYWTPuDr1sgxwQd7U7f4YkMmI4u9XaqesCOhTmU6DGA2iPp1Jh4MsI44KAk3
bZH3jK/5NfdM3I6Ol1mzSxc6V520lBYaOh/kq4ot7Wzt6pMRxBQ/t7IQ3L9dnPiX9EAdZ3Vx4ie7
NbPkAz7S8ZbDlhtvfE5c3wkV+bPYxODCj/KluSbH09suOKS+FYRFV/OgSoBR5M7hJKhduxajTYn/
2GT8tF++CRMqIJm1Kdm0LjE1pevVcbnAP8/zf93DTXjabSC3LnAGiG9SUlfgN4kPypPmsfZiDqP+
u6TN5jpbXyrU+sD4yNfApkTWhzNfkjXXVDA6hIuEOjtT0AMGf5TihXMBxFfaj/isDNsYFo+Gbes2
PTCxPuflgPz85cWfNICDfKFIQp0tAOjTNdP6Zr/Z6UKIX39K0xPXPvbJnYai5E7r0449ZBISPEAo
MWSuFOsa2Lwrsl+seUUwBk6urHcUGyE5y6OxR5uqUPa+rsKKiqD23W/HKFhQoAWcFod+N45B+9OL
gB230vGKjvcMEbHMfGb8D/LUzfIyxppPdYHvREP01iqN5WavUJY5Ng9bjgae9CX8s3DXLt3VXM9l
uRfs7uhFdjdyKABDX1oMFlYTIwmzTN/WzRWGGy1TJtTCkue8pCrBRixayb+DqAP1kJIdCG+0v/Hc
KIrG1ZUVxtk7YIl6dwKYe8iMWuaW3lcc4ULYN9OiDD5N2iDOMWOeXG6nQCTNNTnEiodaaxdydvEC
dcJP7DDmlbeTgGfgM2Dgb2L/U1lqreozHPvZ3drr8zgZ97cZcvOBu5TtsQMxmWQkC1F8IZNEwh91
diL5EqDg0w0KFyos/4YEzcpy8oN5gfZ8FVmYADLHe8n1irN+U4NEBR1i0BKUrQj7tvbBD1qPMrc9
0q4YBrdGGWihy9g7B2dC4FJUva1K+6YNKmXW3uWYahjmWbbYPuBCp21kWs/jMusMOkDnj/4MP1eA
V4lb7qNZaj2dV7ZECFVLd1hQ7Hsc9LTOX1s6GsG3jlvmL7PPNZEAYqUXsZ3XiFpu/uKMc4+c9Ogb
hZDVebGXebbAdksLJZu62aynaoRZ60AgBDssjDOPm1ixsjKHSjPhgSIo52SHzDs6uYKomdpRhr30
si+dnnaMTZ/jtN1cZe8TZ82n9mAHs/1LT+7GAnjZHMTpjBlux/81bbjybeM2cfmlADtln324lLJ7
+YZ1jzz7JbBQe7bB4UCG/GAuCIUN3MwRcLw0+ApboHTl1j7ze+CeGwSDAxjJyjHFNAtnR2/30Mka
r10ulp+XkHfzgj3UFeeNB2+Ca5meJDH6cTAaga0jQ9kzpgd5NTmawUbsXVGaY3PtTBDqcgDZEIZc
U3O3G9m+0oW6Bd+bQTJ4fncqHKdmJRldPEN9F7FshkHqFta02e8PrtyzNxN1qN854duTmEXEmJZS
ru0V3wFRnyJRVaV9sCXXyZdwoL8aMC/v4eAU/Ta2c6mhJjiMHgHfG5XaKxvlhsV5JSxOCFC/zf5x
5NR0wuxvqLuAnWV4h3Ep/YUlawmvbzBqQJlkViZ9CnMZtAO52LnjtT3Sp9tkEyFixDes6TaZif/J
VSJPyNsKcaxxuAPQ1YVoG8YIf1v3ry04Ek8jUNtxZVw51KMqr7Wjs2AhtkvRkzL0PkYK99jrgj7d
/mZNFTovNmWFG4zhq34958mAYyqrUBjP/Fm/oujIPbZvSKO1pZJs03cvMZ7HM0cA/Prd/E8/QDtl
LwX5MnF/orUG0Z/9X/WyYUKZ3oUKZZibgaJzaRAlx2gm07bBsbHPPHx6KLqgPckn1NQZEsxs5Lrw
0MszEXve8so7/pyuXvnZ13C1fWlsfyfG4JL6GzwHJgqifro5HwmgrxLdcDm0nTzM9TLK1ony+SG0
ej8+2o0850ly+hRRXc9kDLHlUK5A5eyZSKj4UInLmwrtzYRunAz/MylGRIaHHIPN6mu8YDX5KsIY
wEXdTUvA6zwvTb/jLYKGEaMmvTPVUQsmVa1NHhR/aZWS4OuCfZM8F1q/OnJ/4eDLx/QWEIfAy7A/
7/gfQNGO/BFGqlzJ1T25FU+rWUp8cCjuFjukWToubZruYiMof7wEzErm+8VzfGNleso7pN6PLg8Y
6HSo+hQazLh+y8dhLJsIzM6VAE7vZ+RXdcQpLa7dOWDXIzeWqfgdLAia6Da4PfSo3LOy3AIoes9K
wEL6rob1DpYFUUCPQzyLRM3TfSr82EaHOmpBnvrg+upmRp7ccqW117Tyr3ofBC5krvulvvbwM3eQ
MRrdRcq2EkKR/X/h2eNbAk2tMKktpmGSYCmKSMh0A8LjU+miZPlmbCg88SbKLN3q9ywWcgKbK/fr
IlIe8/QGWCOZZtpTiGfyXUd7YPAmUeaS+3bxt1UQmtblmR2lsbcu/shR5VYevwMCz7GK46u0cvWB
8TndyxtXwtBVu2tO33MbBfORUwbOpNhWqsyAvxYpOrijzCm1hjeW0gXKcT45PrtcT7DwaNL5qQzr
6jwO6mrtfxb2wIgrRwKW0W/sdpJe8CDQLFeAIO/3JPRNj4fl6luxwkZ7ZZJimr9c/DOsdEpKAM8o
N2n0fWObswIscYqQB1AZgJkP3AAUK3k5rWK63RqGDm/WiJFIqg7tnrY1PHyfSnH0pCSmcEJZwxTR
LU8+eyDF9vZIZYVMhIDjIlVxwxOH+5p9AVSqN6+s/O5+Zpnc+GcHHB5TjGSc9H96FjEy4SyR1Ue/
BvQLrlYaaA4er90HS7J63BbZicRiHiRS9lu873OcvqErDD3Sj8AFRo4gsEOCVK02WkQTLpqHyhZx
O7j8oSECB8GJIESI7pXT/RFAlOf+qcBWlGgQW7+sou7kLWGvVQphjzRj6vqTCe7V4xd9P5H4fP5C
4MkF15KT/5Rh6ziestYJk77u1CncXDftj5tqYDoz88RGLiYNkLKGHK0Ta8jyeQ7IytzR2t4yBhz7
G4cPXqhaCmJoySvN7RhmQ07SEw3PjoMeKfYrlZosnklYegxqKxFKtAfA63Yu/XxUYf7mVexTPwCC
wxLfjzwcAgWeuouRKx53eKeiaA7i0fx3B4ABOn4APUAtwVB1tcBE9FjAYWI/7EDNfL7k9fR9IMym
WveBIOFbiYW4ZVPby/3yB/+4CbCidhi5DuuR/1lhSlAQXKd0y7C5uYsjdF9F9W+iATwEAjSUB4Zf
ADNOiVK2prQ3tIABLm+6uxe+P3Dr2cSFft2IY3efY55/fOXsGD/HOt7dLAcgzmy/g87O16t4ZuN+
cfhtGySr1GKd1JW884TBFB+aMfnmVp4vTjMFzstEqSvjdbWhotqAqWRcj9GFXyvP8q3GS5rVQrFL
QAmb45Dpwd8ENEORZHa6UssoqwdmuJrDP0B+9pH23DJZ89lcj0rw0fbn5hMaRZ6/qyK1/BJZI2m5
IxopwEvPCIOeiyRLdkUYbtdoLx/ah2gV+reyQXc9F0rDCDx2lN0J/99FbAsEPSq5ZLojRLqlWpGd
H8vJtBnNGRUTSqduQrQGSwrQJSPN6rS/D1vTXg18lie9doZpW/3e6gDPa0tNT5bWJARy5FI3+9oO
OetYrrgr78tBt5sRnBBhw8HSKSMOxJzoELixrB/+qpxj+OUFqWDdrHeAzL7DHM8MRuAEHCYLgnn6
h3Jk/rxxMnYHMerlJv++rQV7kDpkNv7u9Y4R25IDVxM0tti/KxDLzjFzi5OHDXZ0hW6p+E9Foqgy
qgnxbgi59sRrWg8VEKhmaizlnPGTWQNHP5q2imTC49yRb8FDNZjYPkXIK9jmGwSMOZwjfQonhvJy
vVHa/z48uPo786xpG6VF7neReYdNXC0cdfxedjIjt7hcxfLYZcDbQ+5rrnf3x7cR+wEn4h+yxKJq
uDIIRGe5TfhL0MjoZJ7ZkYfahwsgEiNzjsqPZcsAFmnFEq0j55fUdcBTVx/tiSFpL+XA7fZUh3Q3
LpGGfsrUu1Uw/bTL3ACPLaHNwIwf9h5mv1nBvuA7GTiopGJfGDYH6I/V9pmk3x9VRD5RR/9SrHZY
HjpxWaAO/VuBjPdVzAJSogNCEWQ1ngF3bKP72GGM+ReZdQEdMtxBhcpKYCJ1MmxI83ZFKx11yfMQ
VHMTW6oBJdEARwgGAn3NnWKjQY8iJrkHCWDy8iVAvjSXCJg+xNniaxfI9T/fFNSllG3FQMHOP9qR
lA4bCch98vMW3bgR1rHpnof5hBCQFSPB0/4T2wNkBfHqlzQnp/TfteqiKyyyxDx912M2xRJRYZgh
27iNErPv8+iX6BiBFZNXaVswKBlLCHsOZHyvv67l24c9IQp6Pim4xpUwpHGkIvUNPLjUpsjSrE26
MXmUgxNhcTz6adQ9+5mcdLghBFus+pyfPz5SPHTOgf+Y5bHzX8eo/zlHljVKe1bAFpLuSH8wT78o
MCax3JdVcdfLwK3X/2r3t2NcXYyxAHaOpxoszFWKZGquinRN7H09W7rxqz6BMCiIhpwD/YdudRhh
rfspRnJzJ8Gmjd5/gOkYjEug5ZM7NtcfawoiBkjZgLxTYsq1ApvDGpue6CX5a4UTG3DGp7XmK0Kj
SSiaWL+IAw0LVImBhPWmPOy81KkK5mtEm/JCjroUDEbR/4t3qOdku+xMoImZt9Rq/kradpHzoCBS
u3usF75UIHSb4IyzwwZmg2Igg60u5q5yccujX1CfqmbeUWwZq8QBjx57WG+6gOsd/gjMU6VRbsef
b+kH3UqhUbnOpcM+baxywzF4XAKnAGPMgAannz9hOCyQ9rN2U2qhkm8bn8j3tkJyRFGWynXy9t1g
2fIOoK+BywsXzU8Vau/G+VbDvDQGMVfRPqp4e/55DkgKESmGRyHQv9QYTsRdhM9i75+Zkcz/CiiA
n0Q8VE4nYajrCXxB9M7agbLcrm2gC/acS6GG7tWpxrosZWXHgq73b06fgnDMk2dSgL5Csd3hbJyB
YGSUEdguh1Ktqtam5QfxCtT/BdvMK0PVrwG+qZVjPSK+Mm0v6iy07yJGq6hcN16qU3tmIuMklrQG
5dC9Ik9piVGv6uqi0DMIPYPFexujwj6lwSJZ1GSfpJSUimR9pUy0Gi3lfi4mST15viLVipUaHvBS
T9Q0Dv4KOAsObLIUeZ5tvHtxFEj3RRMxlU/ajpX04Bdcnv1QGHtYX2YcYwnGfY0OMUwX+wGZ1zXT
Xuta349hqPV/kQktIGo/Bv8/RHUlJjGwQnwGQbve+0NV+cQqUQuqc0U4hhwbMBjYLoOVffXMVvR+
KAtYK6GhTeFtbnxytt2/Wm15m8rQJczJW4FL1b2l/B0hCUAX7HOz5YHWW31l+TSRzdUnFHIHEKun
NkslxsAS680UaOM0CLTXD/h/qgecWM85c/lS948UHDCvnDz+woUHXXw3KW3WToG49SQ4o0/AwDRW
6i3oD2oO1pXcqf+viO0iJxhUCmfe4O1L9fP91Brgl9w7g/ytP8xXBra++6/u1COcDaCRsopbqkeG
cnRHloA9pYmh901Tl+ms5nUp+D3jdVLTJQKG+zZUaneUxUp9Om7vU7MNELF5TTrjBqQC4cXIK28S
QjU6QdTJOK0A7gCdLMeIRnwp1dL/DWnyNJ5mtbSrGQxpekzIXeEdzFuYWxLQwG7sZZen34uvOtjo
pOSE9jvfZMV5JfoTOSi51N6bWHXCIZXtis6AiOTph8eUMuBzIIwGjjVxPqoXUg69S/qtrG9Pc/hk
nVforI0roGGhm+qw3+iHesvLmBZle4M8jmgVjJ25cgrbgHI1gxQyX13DKUbZ5ZGhsWN1Ci/7d82R
8y3WdrzpRHEZelBO/dy3AptVkYuFL8zrZWX3e5LljLdK2imgBcaisiKQyoBSPwWWNq7E3vOx9edA
/Twr6ueNxgh6yfI+aES60OF+oeeS/g6wcYR3YZy2JjxWGCN9d08FzivsTb5VJ3exzwL1ObcXnYp9
QUangFUPkQIzbRwYTqxmAgCuqlDwOF3xboYIzUOdh4AYDBXeEhR4JbsJVDHWvS1m0Lrlmvv7FWTc
Hai4vF3MyU669jIA7IMJwGV55boeGWdbb69tP4TM4Dldi/W4gQzK+hutIDCm4Qj0blVFDCNMtuMM
RhbpuQFKvCae310iZYNwXsqqXxg1gB2EaiFrr3jird9I6sLT51s+WeFWMVi3t1xD2KJ9/aKOTtnx
DTkWNtXvAJVh6Wy9ObcwPByKf0uD+Wnh9hSRCLE5xCENW0iapHTMfJrsgothxzzr5bS590KuLi2z
TcV0agEZ5RWclly+ML4zeQ8GDQyelSLKmtFu9s1q2Qx9gdwa+WbJGccZ8RtOC7QarqGci6dZ5mGp
BMC82XqVsf6RyNtbIj2MnMqV/DVS0ZckyGAJFF/Oy05epKb8InPs+h1ppt4+EwUgCKc6huLgM7A3
eYeJOhz+9tP6A10Pzg0ckiB9PSQSiKTQ7JjOfg/wzC6dcXL2pSHP+UqtcKs1Mc0TYOMOid35mRjj
At4Ty9jP9hxDnoMnQSkD9/gtLFev/WEz2JYVqaAhigJDX4rqcFu2G5Ru7DrfwhDoNN7kc0EgRWIi
cBgArNpBfvcRiZbFe+EXRioK9FoEN8ndfO6cx+5OyqM/ylHv9NGYgVI8idZOYANxJ6YbyOK3SDwB
85YJwZR9XqB4bQai1LnU6RuC9IuN6d87e8IugfREeCAEkPW3xzZSwjOfGkp2/26brxhAATkuiMFN
lQJa0x0J4U/zbZfNYq+o8dAb2bGBSTrVUCflnpbMJF5Pri3ZKPoM35oUDsjxU/K+Pf4xemuvIbek
Jc7gUhvxtUmUA2IJyKwcIR1yDtcavdQXptbnj1C6vKrV6SNtEW0rqiFsgpgkQee5bU40dfT43jbw
ypGfxxh4n0Sb/BrpK7Y7N930Mb1wPIpMQqzcswccadp5Tb1JANCByfny+mzT2YbYomOqoCuo6Tr4
/ECivgfjg+5ZaWAZKTtQwWdqnVKmg7wcIgg3V0nnYeM8pxcqgHRym2SMU/g70pPkSgv4ehQupkKY
x24OXcjSpVqNJDDaNL0JtstlX6x8FlCohN+NgIGRxdVjmmNKkjYIRswgNHB7Fsl2XnPLisf6sIA8
pRJ3NQLiqO8cQ2jY6PYeIdPYcXPhzl6xPl47pZ8P9fOYyupV/Z67SapdX7hzmApt60p8Xo7kOd/u
KQ8tl4pIg0TR5y0BzqrlotieBCukKMJ+zaUzxq0miLLnxSq+4RXfqy5i7R+0bHKYPPGm9CCvf+Jw
n4lUoJV5Ld7930PHoWDxNzSdq9zthOVhUuI52P7KrWtQLo9venJ1CjHPSLwnLGUyIuZ/cBIHX7um
TuOvF3tkTIFHVq13vtEpi1lMcO0K3CAfi84WK6ZuYnjab3gxrJwrTUexBU9W52cP9vwtXsBJYaZQ
HqiBiVmSC1BXfpkVjLdQcJnup/Z9MafbSOGGdyUgptTbtjkXPoXD3+++J1Vgh+nSqs/SD+qFmQwb
Oku13OyAXKei8x2Kmo+Wenc/qNYWjJBHH+/X2paAx5mM8cK/v0MqH5PPHymTIujtjcIzbCiyY2/f
O+lDUPyLKHobRN62SllA7zp0w+gX+Lg8Q4+Pm+4FXztWqoQwkEd0+vSKNZe5k2M8jAHVkXmPeLhp
NdFEPycz2IsQG1HKtq7Ht2Rm3ZCWZ+wcD6L6+BAod9uaVLphNqNF80VJtdkyMjrXnv5UK3tMlJEm
/QXQSxXCGlgxCvSaWlXVLenKTlJdO+fo8kkriE2zzWOmHr8i1uFftqK0eMJFYm5m2tdQPuSwNB1T
pcLTf5Jx/XdUjgeC3ZTPEGOga4u8etE8zF5zp18IgIRUhFh6WVKfBIG6Wd9JzSCQly4wYUK2JsMU
oH988Ub8Ef+QbE/j8VaOd6kI6EmAAovq/ecmU1aDIhyCZP0m9x4cv0asz3rONMiJHo5diPUJWgAn
rsNixtdYx7ctt/BttCYchWdnVpKl7825kPJe04ChdVeGk4EBvCfu+90jB5C1I4/gebFX6Rluy6lh
K6aPqRuzxfH9wTP9a3i8OpYdw6l7WVNz3UBCu+EfyxqQFiec7Mm7rdSio21s10rcUnXpHp92M/Zu
vgFDBNceT7rohMo7/CKIXQCgG9MG8uskcUY1StDzNsKrjv55gSFCkPbG0/kvOggV2J+R4xQlJK/y
XonysOfHPuZwtjt1/iYuM/p27cCRVceoYJv+wAAHPi0r+qXFEr/jK/9YKqRT+lkKtrvrcIfjxhXa
8zfNRWzgR2ilEkGt8qt4wZLWwZU7SRnsUROXG8lf9Bhwyq2S1/xZPGIcn3IND6s3zzRuDBkkbVhT
m2zErL2vCSvVZoow+5UaWfpgQK3PeTvxNxKM13zZGKcq0DiChqRPT+nGvg7H1t+F405WHp0KbM+w
BMEuFZIhW7FlyAehGB122DUUmFKolL9qmGeoI5rW1zEr6NlAxgtqXHAFnom4zcLP9Pl5Eup8jS+8
DfFHuHHwLAvwaYDuL8pRZkq8FXGSU1DG6gp92KBZJn7z1dW2Wkyv4qT7gAModA/FhcgWRYpKf0Cu
WNCZX4CN7LZzDZjTVVY4Dlpci/pphxuzExrQMs2ooOEeFQ7xs+D8YjZu7PerBPMh90VNymVTQt2Z
Q1FKSDTnenue5bbRTcNs+VdrPuroCvdbx84OD7ip0PM7eMXTFlRU/5doA2Xs2FA5203X9aCXCD1e
2+9ocwH2e+4H8Cjs0TJicxMQg2QUgI8ZBm50EbRo/8m6WGrmsv50UOWDQ4HuAUAsI/diB7WKl8/6
lGs4hZ9v622KmSJmmhU4zCRiukdnWH7qMxDeJv4E5BUuRdp34/k3i+G1sGVGbNMhlYJBdH6ZHAq7
wMibk3Bu+ybsku5mGKgUta9WJWHrRS7vjTPVqcEWOLvzSkjJ8SzGuQp6+OX1JqVmrvnGcwwZC/KY
RjkXa27OGnK/Q9IyJL6brr5u7TVHBxk7Wfwo4rFxrsB10pIHah/V2AdMcqt96xyUAhcr+M8ZwF/b
OfstIsA8eR8m8lIx06RVjnwVXTA91+DgTQdgkBkEMj6PHYFCYI3kDw371Q0m8Dkfdgpvh8jTURkD
gfJPlt2hHZIbKPFx72qAH4HSJTh2Ln+VBE/+Lbs8q0JLh6JC3OGdJ1+CPvRtpKyq2i4xrVCkgiQa
3wZdcXvQBPnXLgWbLJO3AgiKJr3ULUD+MYSVvFqIRGwbaxwarIsPIQTVBF5Nvwmh/HCyPNuUvE3H
7Ut1OQnomMQ6gh5FT1oA81tGBun0SxKEeqpXh2qv6LIllmdRgxGatHkyZheiI415Q+6Z3mDwwSoD
gccILW9Mm5lbABBroHOqnV8hZswBI9nbqVyHZJ0M74Ao7GHgiT5F7JY3esWsJ/b2JgDlj/7NqXA5
gKDA6Z2Yg0Dsrt70DvH+OLPbQY2XqcpbX4RjvBNYGyVfCtxlnYI1uxV4oOdiD0DBWMS5UfIxZfEg
3VAP1ujW7m6jORNSxVBfdVVOcrafO380FC9Wv2xmD8J3t09kNTeiWUvHscCHVHc3wqQgDn8y+m8I
TLz5jOIvQ9Ux1TAVF3UtkO5FWB02wFtv/C9MRyLVD0jT1/+aFZOAvNyWja/O0ulASpfSU3UzZSBx
i3SHPFhkzJY9kSnQtqMN6qvk2kF9uZrGnAEYP1O/zdDUvoTpIG7tqyUfT95NptMomAhlAOBq3u69
DKEIwq5htCvcVMFyIhUT/UDHSauMMJZSEQauDF9xAaikUu1QQWC3RYSSVbw3kyd51CjDeXHs7DyO
DUcU7qFrwaLs1jHG0mmD4lAgorQsL71oT7uJ+//+EuTSwx9CY4aCY1uxEPl+yuVtOjz0rcgmPb2/
ak24Y+heF8kxYJEw1ZX0WUIQPI9gU3Z5+gfLDYWXNCaOdU3Wie6reWioPkNLpJ/vIeofb6uaATx5
XHYGVRDZBAoHlV2M7zuBk0RictiYKlVnx0XoYEiz6onNE7ZUD9hUSGPS9WF2dhSXoB40JzhwwZ1s
hXQ5ehxnRsCFEsrgPdaFKMgvakfRJhysPur0F9JiXstxSOjkbiRSjwqnTxILppvN5wN9NTTXUxQ1
PZGUOzWhk50pV4hBnh1nUYfv3oOkHuMJ882jK0rwosfrwwGU/+q9+Wfb3bdSmHBmVGhBP8hXFQfY
M8DvtHL8B47k9x7e3z9piPPOc6KW3l2jE//VSxjV+ElcEoAqVWfouCxVCyOg8NO2V3lntMwvtN0P
KHsljMiYeWd1hFaQl48kac3x3CMgr4V39Wxbz0WfN6wnnWiAiv+Gp4ARlQsgQpTGMiqY7DfQd9cQ
vYExFkh+IxAIPfjK7kvhNPzb+t3G7nhAD4RDtNtIZKwgDRVFVyaTjAR5dCs4CQezfx0Z4X/1pg8L
fThKzI016iTrDdyi/ZRcHP0cDQvpuNB2+u4wB4/x6NSEK0fNfA096X9755TQQVUpz94ulGTQ034v
E/p5Vqo0aCygiFpVVEMB/HY0ZFcIVDafhqlHBqOpN51cSi7/gfMBTi/lAg0tddJdbLx4wvL3v85/
YRqfjro9B2zQ8ey8FTyi1RXP1Ea+iUe5fmHUbu1179zh0iUwUuUg4FgXtrCteJd7jwYD6RqkPUXn
kbl538nb2Y8Ee/7BWHF3ehz0/7IB00IuVKsFDj4EUVpCCEwZYQMBVkC2AsbXfaAHkh4yudUsmXsm
nt0eDR6caYPkf4jZ0Vy4Xpb9EXS6ue86uUyuidQokoU90GHQDuHBu9t84nJaU7hvKpFb+JAQGlRt
oU0bHTFNqEmoAPB4OgcdnqNx4KzW2SOrvj03d4HCTZKmCDFytyUbiuwaWO+dgTb/nd8dfzGyGhJx
Y7wXyGI1jemVfU6oR+7RVwJP8Mn5lmM/NSXZY0k6/GpNIglYVpQLVh/Na+49h8O0WHq2tZz636ib
Blw4oMspoyDCcaKdeEPG5gPeNwrTLn6RI/R+O8jAq71iIlb/78myjwkEW6V97mJptFYwgsCfsAeq
yoofEdbStzzPKGFvXdSxyGxoeLBct+PD7/bVa95CUlzwcMF3dY1vsl5u8Q4RpdWjfpn2DpOLx1fC
dsbRKnDglWLjjU+6+B6EUb8IvDs88pFlmRKfnGC3W4PY29ewmR13UyZT/+sWPAjCT3BnsP2QPZA8
kDicWsq3IrPsc3smiMKp4qcNarBw2vhXrHEViQD3rkptNkNPXR2CCk8fH6DuLfSoxevQrGUaLwFw
UXLkLZQJN8iHGUDgZXLlkdUo4wfjL0fTHIY7Wc6/bsqjPHgbCF7ou/3ALEPGaZS+JsHFOcOgMSIZ
FNKS76I5kQjJ+yHYfBy87j7IqckSspxnBlrpzPhlPoIYteJUdHkQ8Pbl71NNSNo5+Cx0kmOQOF30
ZyJQSJDozXIjC0C15DbyTRmNbUe+yy/7MN8jD9xatz+Bf/IA8G6DfhpAzAZ9fyTQ975UKqCeWMoj
ubqdZdNnshmgQOjvz9QYsoAcw/Ef6BERQ5rl+Xmnw2sfKZwEeVutI9qCT5xX1MCI6zXK0Dh4L716
bSfTuHJA7O7iuvBkCgQcVTcb9bT6nLtz8ktl5Wt5i1ue/P/jsHzYI4/9Q6A40w9PYXaZ8vu3E3gy
x8g7KeZ0PibKIMT27gIcZAZ6CgjC1uwmqO9VC5EWSFCKCdPqpyaqx9rhQ9H6zNOPC+iadkuf4k5z
YawLyL4eHOVMZsg1+vjMRty3AVa8P49XZxW4NqUv8D10EY4mP+rU4KHn/4CnzwsnP8k62rU763mX
qz9N69WAb5P6d2D3bjom/uPQyLnG7VTkgCYzBxyqGqOGjva7GrqyyNzyxukljnV+lpSiFbvuaNvf
jyQxl947M2UNkBwdPqzhldy6uAQFvEUKd9x5GdhUpxpKI1swd7TVflnu2/2bVyYEtFHOoNeAv2u2
PltvOad3YS0fdQekuLwhhD4zNF6+WyOCAesZcgauuzBn7/4FX3kBlA+NwIstfVUluFZ1dXPAN2uR
nQLhBYeBmdNofCXOYKR1lppvNmvjnU+uHDlh77jSgzqRsKD49BP1TVvYikAEj5Msk5OYy7qMfrau
akF2mSsEquIXEah+LHA/WruAqiZT+vzdDf0j09V1RwjzfIkUPcT+saLUWWDryVkdRsLykSYK7l1R
rXxojJPNwEQ5zREH7lzdrSTqRrceaROmhcZPK8xxx2AHyAmakQR6vi7HgbtmmsfdRUeWtjQxdWNk
JTYFECDaVJCyhurtLZ1PJX32clg9XwNThIgaoGZsZbg7fvqyhLPg7kh9VDPh93bF4RPrZGHTLDnW
aWXxlVHCxP942p/4eAMHfywZr+lDv2ouTn6/BVsf872yTC5qpDUtudeKs4n1R/ziP3Ozkz96QRDh
Ej+GxuRcVLj5Wnu5LkaU7QXDbp5yAk5mVOU9w4z9dvgVS5FZtUwneHTY8j37FMsxxZgUBXYrMff3
eMGxkIkOPJ2gmFguhFT3KADQlzKxmBl5Zcn2TcNePLZsaoZKSZrQPtKYFJjb9ngVZNNt7Dnd8nv7
YEfj70U7KucbhIeIDl3TPGt1YFyiXlOq8lSCID1Lp4+WzZbWFsiM7YTpaEhPLqSAEL9eOAiuG9UA
fFW56nghoNUyg8vO6wwJZ6YW7XCWhUpQM5NDXkPWEwArJ3TS7F3Y6KffHw2Zmd4NVov8HnIjzLWP
AGtDpqQPXQDQRcimb64WNTtrFTB7l0jGiJbXCxHqiuVjn0D1RJvdENb+dRotbUCxHyIPZ0jq9PEN
XDo99W9sDTak76o6/x57m5R+o002zle5C/j/wvhCf9B03hhiYSubW68TeRiTjsihd0VZC/TKZ/w2
cXXVt162e3tBy1LSAHi5+F3u8sW2tEvBB15NijbQsHRKMrYQIvNvA7JLHHU3OuCErMyrrXiWfJzS
SbVBaFeJJNl8mMQzGaUUY4x03+KNAB5cPnjA20tHWJqxGBkfQcPM4HFSRC/taCWAYGA8XLLV/GTI
b+E1fWsZztLZBTenPQlBKO9pyTuoEsKp/KQ2+8ptPDV3EOycir1yLLivpRQbAGNRVBPXsuU591lF
nc/eKrKFLufRVwzDZoSWjjphNvAlzQfPoZAeS3IjZLdRjQu5btBPsxqKTft9XTk3YqcdLQaRRD2I
jmKNj6qRJkqXm7yZnxE6c/WN8XrRuAErBiPxmv8nPMbf9VBkjP0ZUf1jk/80LRh5b0vL2CwTmvKJ
VAafSWRXkjEVhnWjmPoAbVrhR3GpfuQb410gDJT5+zefgRklJguDZHjC3BxfeZx9G3a9nQfKgb/Y
svDxZUzaljmFTxgn3HbBHFZ3EINRkINL6us6aMV1Ol+Ofp/jRWcM0VGvy9EtjyP7Kj7BmSRcVJId
o7hio4d4YI/h9QQfe2Q0MkO2BiQMNRyRmXZ+XCkcj1m34bJHTsPKTLwOSAkgo/j4KHlKoY33lh1N
YykeHN7BfRRWU9jQjXvfSO6W/zTtNLq9W6UPwQSmUMJp4M8d1DcxvXNmtc7W6CrawzuTjiSDELom
eC51rt2LEMDekLQXrd1q1y6qy79BTLT+sIYxpF6NiKX2WRZDjuEkdalcESQpzlSTXoeaRicdNE/L
qFxWxt4jTDCxCQdTW7LdEXmdroZR79828Y8yh4ajdafCdCiBzbRDCgRRQb5TU1AGFSaX3ezwfSJN
AzjPHAXsZ1JUVCkvh+Ep45tyzhdaRLsl8fyyVTX1CIebx2EiGgtYInDiEt0mRUx1TJruPOljGtOq
E6EvcR8IGBUnHj+boqqxhf8X2dKEw9TOseAWBK5ksQHIyMhZ8tW0h6rniUSez1UhCxS9OKL4FzQK
6soxGwpI510wjAWZR6emR1qYAfrfRrr33HAOkwjwnKV9xBAvphuxQEHZ3s1AOjf1rC5pfNpbslQG
f40wqgLqrDQwH7yFWxKZm8HMnHk+y1QpBXieMH5GHBL3GgiIRb//BF4AHr9Q0BeO6cnV0qLRfGBN
Qy1eti6EH+/xD5V0CcXp4ttcBg+NxRNIQebkP9LDAt8oREnGkMVDDJCtqDpiLxJAlyOlAkZ0BKAW
b7PgBuZBv6YlzKZcYb31Hg83oQOLpfdTF80GZIOgrdTTmmCfg/w99x7DyJZc9RLWRpRfljPHlu1U
gBtw11iYPB2FWL3Dkji31yeSTo6ik5sme3V4EQGUGISu9hXiMoL0xaJokHRj35jJ3jtBb9BgOrBU
Va7DE5v4yIg6P/o7cUkT3RkNm/jx90k6XstQkTvNaN5RFPPqvZ7UQ4G1m+OUxDKQEtMG2QrO32Wr
KEgiQwgsau+fvaavTh2FjdHR6z71B1n4re70VmVs8hMsSgrNZ/nOx9jl0Y/FDAPmGHes4dTXP730
glIRFGx4l6/oON4aTQl4ephxjJ7q3O2wlXAHGqWWACdvwNaPLzDcTG3rTBEkKnCo3rBXOcS8549i
Px6DTW8vL3uHKMVbTss5DGBp0/826s9U6vimID5mqlxRy4ask2ONr+vtQBCG7sEXXsjAj1Iig5f+
WH2sSf5e8y1OLxlBLQheFW6h//Aq6Cjc3tGNJGxZWYYIElUaL4yeRbpG4cHDU3IzAEozdSvZNgYm
7JBCnJbcwPuKFZHquxwMh/pXiwZURJnBIXB/XjDA23ttIcGeHGx6tS3WMvIfaIHuxvEbYLIRPhNR
UhhBLJWa/XltMSV3De4NVNa1KWItE2mcpnW0ZBYlA0bPXo4Axs6UNEcucNqoqEPl3zMKvYgUpORv
raSpPebSq82GrkcGLMMFpcRkV5mPN8MkHCgFr8k5WadZnsKvLfjCi3ffXemuKKTkR1QzGBAI4knk
KXaamNci6I5/F3iMSBsKM3p+NFQonbtCAEIf/JIFAS7+N5tRIQghwSSCg5YnSuWjsuA6ON/L1pBr
9ERhdeLuGj9U8Gs0W51C3wc3O7m4DL8RuXdy9U9hIfHH2oJB4AyjpARQtmeO/TiVUDiug8XhAdih
pLaXt20k/5GUUg1ii4lFPQT2TMP+bQ3LqdczKhpw79OUxO2FwXVoj/lBUp2LTZlPGT/WXTXG4uoM
zNt2atwcESAgYmvupEzkuTqQuBwBFl/plLAuUOx17WC5QMr6V/Kj5wamBj4r0E41E/AwV/7CSbEG
YZ3AWFagdIm5wsiG4uUBUhTW0sjebuaxfgo0swsAotNg38KP2qywXeQFhh4UAZS/PbVCnMZY3Kis
f81MLLnByIXGOSzoln3Pfzt2AoVfM7A9nCTwSDBmt94p/y4pvcCHF+77i2xujyOdMNGyAl6L/d1j
B9oFmUvqyVzW5rQIegBiasV8xyhCYo0C3XECUdBZN2cOXVJMwG+lHmvx7AxoIJxDzhI1R4zAh7YK
LouGqZMNKyPeUOL5/Pygi5D8bHD5tyHtZ4/vWGEdHfU6fpguDuDA+V2o4f8aLPAusl3zLwDeYeC3
gGSx4K7O0yba4V2PpDxv5Fbo/tYMrYbnPAG7AgMqnkt0HjoswrvK7551Y+frf5ADWyJVlP0ckIoy
4uXkDcZ8gO8Hbhdn3pe32BKysaWsr3TdVXDS1FeDjl3eiKxXouWpGW3Jw7+WzZ/bXRNAgI0aRc7d
4q7WPBXbgg5qDjDZuDxbrFOoMBohY3G6aL0q/19wJ8hKj7qeuyjAQ4KVz47Gqnan938/dOGhcFFG
Q/6rKD68LX14uuwO4j5F9TQIZMyj1RUlMYgM2+RIkcb4HHy+Swbs0YxDQTWE3PznDfBBfWfWRtSO
k/RO1Du4yu972ekoBPAWs3B/HWimoBQVCA6irY3icOwDfd2mVAqNbhCIKlsL8iFLJ2S3KH4F6pXx
0eWcm8+EwISDXMgf70/7bkexyyyZNtG+HQNXXAW4ujzSIKXJ10tZ+0dY7KLgSFHjudY9trxlgFOM
Wcb5OzgBAlgf/8khtewxDq+A5yra1ODHWlz44jCpWWdvSCWqfnEHpR1dz2QIafc3r9Miw43rSOAq
No9M9ccdn5NNH/36WDg5GtloV9C8twE60cL7ORw2UOtqcWymZq9w9cktzcdsqZsrWcl7HjgH+AWE
pxomEub89eMOo9UgPNJC9ryTNO6eMjWjv5nLl7IFzvzUjdO1g0YiZfHenhLheT2TH5M9oxGmcoQp
K2R8WA5gfVvndf4j81HPURM94maX5Fg0XIlkCbfIQFoZuQb0FwY7RCa2pMe5WW0y5Jwx0p1HgF1n
p/twYab8apRKsae9eFOGN9qqtp1tcwwct2ZOQ+JTEQsW/A0hiRlLz1M6/cjX2iWuTSBhcEuzokyt
bLjW9qOa3KPBwqPWk95xEmiuJvhEpHP7cuxz3qXkBy/ds7cAdACF+0277E/tmurVMi18519gkypz
rx+BepDEbbgWm0kfuJTP+GK5+tuIPkgtlX63U8ZjN+mFbh5aNy3SGtsfP5Q2kHLoJC+3tnrHjzEX
QSaxiaA2ZNZuEZnci09tKW7zSxC3GiAkLoFSoFhS7+I589q9fYlMg2beODt0SNlpIJtEqIY6GZPu
P5SLFpI6MUl7ND8x62TsCCaqHEQhX9T7Ocqj+7BLUhFfQD88tjjmqC/Mi0BMEnN752M+zO7QzBH5
pbDXdjZWGgnl35Qd5Dql8VaabZ3IQl6weUCmzxvbCeNFF9+vwWYQEn1hrE1kFOpeoMGC2DWXCaQi
NY/O2+V3a9Q8bY7rs4LLe8ExRb4lO6CaBnxGX938HXFKC1v8f1k3xdJhUEyM8oVmUi1FICTPCupd
Wgy6u7X9DWfG96LzwYzFq03fE6jbHCliKELVOanFzFnWNedMsY+8FKnG7Z+rWtuTsMy+xxSBktqN
E+WwAn16cdNzjeaNkKL6efSoSFnChS2JXDm7NeL6dMnnQOtWiedOvUcV+9o5KrzlSIkgOMCqFK/A
2dEKXwyhr2C6NTCJBf/J2bqlmeq30zb+X1RvX/c3oRaWGNGQkNBTEC/Lqd/mZEYLlCP6/ZHf+ZNx
aSZvHn/E4zgxEwgLrtTsFowdKEYcaZlRLkDA5BCoAcCydGhUcPvtY9SznT+kb05hVyDA0ODfFvR9
vcyUmbbyGzKSb97jPC+0rLJgw3NUQF4kq9NmF7D6j0s9UNWgOCKX4FTYmcRl96w33t8xNqx6uez4
j63dgEbOVKE82JLarArdFUyBci6ke5ZZ0y1BNmTo2ZQ2Tn89CXsN6Yx4vIUvVtmD8SiinzB2hWJ9
2C5hZwoSnc2pxUaC3AUzuz+PnKwrCaTWY6zGy5bwjUfyON1OujseCjVLuYuTHr7jTaz2be8syPSd
jwPLgHHEhGZzJogLhFAGv4YQ8Fnz+Ukxug1Pl7f/b6A8ZQrcpPiaZykrlhldLh6jKgq1t94OFY2C
eNHjRK0fT1SoUDzxqD4Phv0LhyeSU87WgNJDtOnx9VOncsfOU5EZngiZEkkfEgKqoCWqmsIdjAat
KnD/uqOGEuyId9YWmPo1/ndh46DhEpE7F9y8Aws9NfZJ7UtWfyOy61K54fw9G13iA0KvcklRvYkE
Fj+29sI+Y7+s1SlMfqvKxVij1L+oDBarcaf/xC/l1/LVga/RI2zeFS4rswUXR1/7YrJW73w3Vhqk
WttqJoxlk4hkHe2EeIHcdaiil+wckzsfHpY3NqaK0Gy5TT313orDqvUO5lyxJ0MaQOmk3X/QgxJT
fieG7O+IOGVT4LH/OKMVV+Cx1buIIvbcIHj07DoHDZ8cs40LwyQqfOJAbuN8RoVYYVabdeWqOkWn
KMCq2RJOJTVG90V8tN9+a8vnUjO//Q5olsRdgiv6roLfdSkxeDQhexiZboyk18kIUzvDyWlI0jqk
GhtAgxkGkEbo1/rgk5HYZ9QFbIuMSPGIphUPF+LcwItSHM36ffDYp72EoV7m5E5RXgTpwxS+DVot
L9Z8g+a9K7HAGC1ME4hxthL8QWO5fSzNja5tfU56cnxbfDPExa9emsMaxEKEm4KfeFQKmSHNHwlB
3yLOUPQM4aAvlbw+/yHpTTbGxbGK2AXSlPdB88QfojqteT5rLl7cvMTxYSUTI77eFDSxoHg9+hrL
xiu91z1GozT9go5cQxyBQoin2ycJych00gLp4d28qXBq8c2Yivl8wXXzfba3AvqMXyQ0razSXiPR
BmDBU6adJUSN0ZW7C7Gnq7TGD1vPFCWNr3INibIIIg1knOTG/mVpyEat4dIReXQ7d+4lYufvzFlk
IN6fTZq3D0bM0seDf+u0u9sbpKbi2ns7DBnnA3AQkoV3zytGkA5YbN/7KJwg+Aa3kj1LLdS5DD3N
852z4cJsxy0iZj9GADeLUT46qO8Wowr2cJvWtdOSUrdEbuYkuYrG/1TLlOYlOuq85c1bYVqGEIjW
hyTYhapCL1mMih+vPkN/0C8S95CpKgYettjadYgDCNLSw22Rn/8OvqfjtgMiPpPORxqZFdREpBWx
N8OxUoAyoNe9OJ23oVAdzhTbQ3LOeB5jWCnL7TWt2aWf2bZKPNwLe1NOQqvzBQ32vGKxE9i++HqQ
6VjXYHQUrZBZ3Qud5xcRKC5TVJa3584TbZgBpg0Rjo0KlHik4huwHY7V8pgnJ2O4aDGyMWz3912l
c8clNrpFEV3gWlcq3UpKCQS8aqGC7+kNS8cIedihR39SRmSF54eWKhuUmlIIE036rBBPuP41E/m6
nuIvsF/0orA9qO6sSjJIECIOVsYj1zJunIDi6LN+4mq2cBrfHFgCgv7VIc7gmrP2ZJhfjJnU8jtc
tn0yF3HfE21Lox5Qy2U0rzfd+Sb/S9mqtErn8eQwnWOJBPJWInBI5L137hL/1S5qnQmkmm0Zngfh
EzGrvGFnSSx/ufE1OoKToU1uBvj5nmq5cZT5y9lXG99oLxAtgCP/csmL3+8WP/wl9S3TNngnQL95
KwfRnAXagOMozcEINYzXfW3ISntGg3iecsLm0v0wmQu0ORw/6vjtbE8NLABa4tjDSKLyBcVoMFP/
5ik2ue82Z1NPMTlfSsj8j+iaPNNzpGVK1FR5IRDRaAnaMpLQBvmPJR+lZrqZ0EdsyhTouKa/rQPq
h9vQcHs7hMi/SBYsk/muqw2poXWdkQpWp3vjPgAWj2EPkpzSSakL7D7bkqv6WG+M8nFEkMTUi7n3
xRCc51QYy6DjHnTxCMa8cTep/CMw9MlWb9A9xS+qqN/GoREvKxSwpKJ3SJKv90eA8a2YFPnKS5gG
lX2SHgGUGJ92Ic3eXb8MLOqKeOu2yJFYL5Uh7s7qMxuv8XszbM6gcztGy5NHGWdg2A+NrrLuvq+7
mis1MDwkEXPJlXU3JB3ONGrS/t5zWIYuw87e6wZzYGm44GEPirHTgLjGKQI8r2rkmuFabouNRXet
bVs7LXu2+j77unMNON3oIjt/jzJxqkMNuiIx0TwQGpOtxyNmr0ItlrXJtS4pBYCuBm1/5md2VgQT
t5Mg2g8LNfXKTYIVTmHyX8I+Gm1vcjWl38L8qX02oTUpDjYT3Rps7fOWcU43eyCli+aP/M+8hAOL
ES8kTpDK7r9Rn2f/BxLBuQ08ddel7SITaL04hV1F3ZPBig4vvsnen1Wt7aLK5b3trXgzcrEuIF4A
PT1JCaHl+UqdMSFCd8+uUM9/TW5izaYVa7AxBEJWJG/+NtIG/M/+mY3tsgz8wXrfJFTOjVB31JZM
Bnkq7dkpI3yWevB1U69GEEoFF+uKe+Gie996m5UGqBCGMfsZvib3HWUqqpkDF6J+uwmNpjffydy9
4lRiFeitSUwerO1g+fpHtfK6e6bOgrz2x/n8bz/ik92DSzYpO7H/yaZ3mhZ+3zdDGGz3HU6y5YyF
Xg6QNTld/n1pDvs+aAuuAfjsCtdOprrJATIl0qXMqn2ru0rMVPLipLEhrgj4DPcbvA91lnVD0L5E
w4r/hnvWPTvtw0AYXPMW9FyJYLmSP7PeDfdqDgysIOvv9qnFJmYlFm/gtA1BsfgQrE1amMfAtv2d
vu4ZIX4naT34z3qBkiC7b7kb+WU5kEMFAoApLwjDkGgFhiTLTovQ+TOR3FKxuy6fO2kbzMFocEnM
ZAtldona358RkpB6Q0kEnv4yospYuL662ymQ1aFxen4b0rj1XmOej1joFIhGLGqr1o+S9iGoG59p
XO3yVAWkeR/Wkc40pgLR29EFsmc6RFxIHr4jqUhZpMMxHIL4VYA64KgC9jVljuJy1Rt8zFCPKk/4
oX0DSLnikuPXY0QFFnI0/BqE5lL3r11/EF4W9Q96ci8elixijA7U73Ad26A4i4kda1Q+ckBxWupx
vd9lwCKu6GseE1+z3Zjpyyf7pPaYH+GzEulO/VA6qV+mQm8o+8v4umWhVMUd6PQD76xW3g/gv6gK
nvnrTpFVFdKo6x6KrPrJzCuWusjiHGY//If1FmE6SU3g2R+MzdUrmD+1IICyC4d5wVk1KuIipUbk
wxAYSiYjuXV+hW7CcBD2qDf543VeHHCSN3/144lP7XoW5BbGgRnV3KR8ekVVb/m4CfBsJHemCKEa
qQKTiBF64NX1a+u6lDOIRAQi3LK2L8utVr8JQndS6dg78JDg9TSc1HKS8q/UMhycTcVavRW9Q11n
LFYRoy+P9wD8F8opKe6/LXd/r9ZqNkJ7EtT2mtU69sj3APlzf/C2W/sWf0vUvC4He3QgLGxHwpKd
0wxl7dEJ6D0yUx4uwgywXyiy30+HJdbqnD7zckQfvOkZiTBJir5BzwNGsXLY/2QKWC2oVjxeB+TH
Ej9zEDUrFbh43yWsHqWZjOCUb6AzRjCtCHJ/wYxhBm5K8WyeCB0xNTeCk160G62V5Ohb1nr6/BmA
jK+NKX3OpODjSd2dNgcUz8drVz6KwuKrHAx+uUQKL7VQl+cphtBnOKspFZkPTvbxaQ022KA/h/IX
4yZN7jkq2+AHFR6ydcVUWWRlAl0ASpTDPlDSb1f+TYp8is2w1V+iglQH20dqXKf9/cMPhTr9E6z5
5kt23AvdZqQGf5+ZcTlYX/EYWF7oj7ZDQkAP7TO95xBIx/yINz7dr182NSxam5aPIMjGprlmkzPV
izCHrwi8DqQssK3rZIXrHCA0AaQ/UBdMhOOIvMSrdAC25I+Z/Lk9Obbk2lAAHZ6JfDcscd8Fj5Oq
exSyfCBAMi5P8P1fyhZdoobtqyXY+ncwj5SQCnvMNMFz4XjRZ4tx+gtBpR8Jx97VzVM4548aLD/A
G2tuBxZByJjkEXik4aMIpJG57C+CW/xjLdr/KPJh20WfGEcG0l6+XWxQ0nx+z6ktka4uuI5eFmcj
/+9PRh2oOlMWbbsH0vTw1i4yqhqZxHZX4MotV4oQZE7Y+yAJDEKCCo0kHEZpvuTImGFCVzDtSiAf
jLvtHJv+5AG3gMX68NZurJVm+9jq5+jv7bwirDkAAjK8W30rlVRp99K/JZMeNbY+lqcoNDLK9179
hYkMI/QctIo9ufs7+A0UBde8Ja4mk18VwtdVPndJ1CUzM6RA3TsDP2U3pe2VIYXoEaa+lLvPBXos
1aUTYIEZ1Yub4DexrnuyoVxy1yeysV2771AW8sMF/OGpyPdVPmnMEoHi756OQcLnaVlmKSlfJSnS
NMU4EM2MBTqW8gC58nCcI5jrlq5VLETZhGnS3vgbmhJPz41rQLJQ8kLgeJKJ6vnysxXAevaVciH6
tKYS6KRzUpwy1ogVIdEOJxEw71x4zmk7/JWeYA+q4zsliDfiiOBIabSuw6cKoJGBA/Pfvt1UJvXK
NrJM/HKvZ69Ie12MDuDP5cssevyGBDQPea1TFjDXw0DhOGNH5OzHFKiKMxjURBnXBZGCIHsX/UnA
Sp4lmY9O7jdX56RUJYErUB0r6813KcEE5W5zQ7Num73y3aPQNh+CIhF8OhJLklr0DMJtx3bXAdFV
PGpnqP1zxCzXC0dCgQeH931YdqBLTLSoMpjD1eE234fBLMpD/sbb95VjNxnqGQhVQfghcATgIgZp
fKT0eYoni21Qz4AYmRQV+YO1osv85LVacDITtI8tmjN4VDFOEKW5hZvBSnu4gULUTMx9K/ZYJ21A
gCvS+6itLFcNDPdLBwKvG4AVxjf3zcBiIhx2K5y/QE5dIt3CiF+2QzmA4PBzQhNHvDVj/5PHX0B4
L1Hrr8nu3B92RdcRE8jrOUyW4goUm+aFngK+dLHaQA7H+M+1xKlz+jmg6GU0BcIjrV69xeLFQSnD
wDQrAKGrNK7hhxm7caoptyS7KlX3S3GdDTRoleNmdvcq/DEh+4pkwL2DT0a0NITXCtmhugqa6j7c
YhIpuWp5BqY9Borzl93xmEZMu0mOdC2oqvmF7m0afh5sLtGjc/pbeULdMsn+azI52gRpniPTLHOZ
9f8wNrCixrHlSfhqRE40E+HKQE3HAALyqkNX1xxTmow2lupZC5vzQqcAmGg4fQnD6EQByvUHVLSn
QiDpRiLxmtYPhzijoPYCkoYkZ0p6RFLEqZTlYh+iUjtxltoCniyek1kaBGZYBz6NO79dk9uqKqg6
wGnLH7LH2oYT1d9CQVuKz6sqxJWDZcjq69MSh0Z1OlAR7BqzezaHnXqiHgY9UAavKgcdfYFhB1Xv
4A76QyaAjbX/B0jZ1HxQsizBmG2SjQt2DuL62Wt95x/oIA7OVaoGDHUV8r+RGEnhYmueu6qwcsaM
uiCgPdptXzwvL1ovEsP06PWi5n11rNU0mBVMhidUOlm58TEjiyeJBSfiyV73NS8YS395oABRvHPd
kidjm4t4sH+rjHSp0V6yBl18aYMhwoHG7uzQ8glcVpQrhn3WwRxdgkU7pt7/a+blvnpEsqRm9UJK
2AtGDDIuCsr9kIu8AW8KaPfnU4ICHdJSO+hQ49oC0bpqIakwHIky8ZAUfn3PEqCC8mAvbuNQHc3K
T9BbJUiD+ECyeSfLcOPwcSzFdCftxc1q4ZI8zuZUlDUJYDodBC1746xhA75Dw5RhHkOjEpnAju90
xGIwAX0dlC40nGHvjA75eXGpI8pd3CgJ0WD6Vk4tjY3JDFehYGYVkcHnKrt2twQvvXjMjhk49kU7
gZzdZkA6rII84uzlaP+PmhiQ3vGdmNRevt2QAdZeWfn8R6Wxu9JK7iq0GClJG8vn+q5ARJH5t7k3
sQwo/aJuCV/2WSDEnNJpBjAJrPsaq1npxR1BUc0UOry4pYVQxNIOIcqzuMlbQ0ue9NvCHHLHy2Bb
5aTqni4OfgWkOksBBnSMNm6du3aaIYVeq7J962P9qEt0NuvCiURR9FgnhqiuGaz/L4cBgcQrlNnZ
p6fBoiwg2JTk7ebNQVds6gQW0GxEfsmXdsZaojxwSNW4Es36badm5m502RcdRrpXm1HTcwt3eItq
yFfOmbILITHKstlK5i29FaZXl1ob5EF4RyFAJT6LXTu5peeGeyumHvPVGWxIxarLHo0b+Ps0uWuw
xvJb8/FXm12wmgoHgRXWYtzgqRzXgAI0EyMG+M0Hq/fIWlgMQvibaefdIuNLa8j3oCL/3PUstYXy
EjrwQZpIeVTtdfQm1F1bOu0yS3CeDNH7N6U6dg31Sxe+s41XIcXCtbruRpwKLgwRH5mQfyCMjNUE
UnaVu7o4/6EC05rAWX6Ku4Ca2NaeaAtbDH3Uu2PmUcnbtCxtyIZa9cTK8mWk/V2NxgzorM/PC8Tv
tml2g/0Zr2Qx0mL259zSeaDuKz9NLG/6oULuytlMPinhLhen7PTHXPTTP1HoLNlS8HKHOjeEDPYr
kizEc0g9HzDyM6mNNhxA0/4Q/fPe3V0iKyRROQX8G6bGbsG6o/tXGLoNsvRNg/oxnVjyoQeJbsuJ
jcZSZb9jgp1UXGymRUjCzf2hm1NOv+Za0OC28Y/iBVqNA3nQiM+/+SgDh0audnHQAY3NcMInB00i
XTye3fUu+WHbjjUZdwYxu2yCsGTNmV4hto3C4N5fnPkNTavf5IhOx7tkjf5hnYb7i9hv4+mEQH+u
NqCsR76d9fgapRWDPqIou3hF0V1duW52q/siBSOOdOgg/pDuyotc1WVn6HmLQIKz2+IDoRqXCre2
4NhwhCAzofK/m/faehn9Mte6Vdqj4prpaGA9g0ag7ri+SgBmLzfGNM41TgC7roMd0m2f1PO0Vp7S
sRO5C7Q8vYSoqPb2OxRy30hDgsudslWKLWVkh5dX8faS6oyEt8dRv1G/nkp9LkWAO822Yi22o96w
oGeEc3blvYDQv9UXJsJP/MGiasXv1eTJlvcqesW8VArb2FVhKEwDU90DJMuu00MsO0j83FGIlybH
EOiTC9HURr8P+sal2Q/6pkpIDkT5EXqKLdgwtPPu9xlt5HDvkmJkqKEgukddunflQFuZ8eK2uY8G
1jOG31xOsukK6I/QLyyAj0OTWdbvyFhtf2/5No5jkaHMck21Jf/tfo71dxFjbSQXovt5Fa6MQVbi
nESc+rTIo5Ia86+2TLa8P7ycExWJlBqa2mut7CZrYIs5dT5quUEpAvbb+0GsB4HbNh+TjKgNS67p
kWFlfRtjd25fIUyPsfAp0X49Lqf0S0wYl4IQ/rXlzYmuiKPxC9IhnNLnDhhoihelQJvYvFkxgvMm
uzyulpU92IupY+5TQGA6gsd6mPGEEwUADFNwKSlLoT/2TVnjCw/2igUircjtFErQ0mYB1JAX2urD
utXObuVl7UFQBqzg4k3XYj85nbDX+QsmexH8zWT4+4LwtGTOCc+9MJjrDk3tsbe3ifKfyJSJ6xkI
+wJgnk/HDquHC7PO8z2+oXJP2DCmynCRhOuLYeqzZvR+I+wWQylQ4vNqZha6eBwPPR9KTHWpQFTN
ZCwRU3qe2tAk39PGHk4pA3WxYtzvx14h9jfwNNyuK2dCCv2pahA7TTMIp5ZV+f2vJ9Yr7RwyZBPr
abKqj5QDPBYxqVU7XSu3ZUdm2AXq/tofvvl1lyh0m4dv/vuBIxfsU2bApacOzvy8SXOOA3bzlQPz
MG6tr/dtA0hK0knO9bR7pp6SQQPRX3nm/yfBd3pWRq/CeafUcEM7uVkhqUwXJZBkdSuen+uR1298
kkL1g0rC8rN86CUH9ga+f+fghVCxg/+umDje7vPxkN+YecTislP/iwlnVskewdFeij3kTmLQrZ1K
1Xp0bytoO+rk4EZVTrwd6Uia4ZlJBfvu1bKR90Bt3fbxjGFDuq2jx345N6pvl8o5d2+1W2lMq8L0
Qunz2mcDiC4gONDUZRG1D7+3gurlyxx1mndc89Ge8iTqv8vifAc4gXiqJEJgL4sq0g7WcyJvnMqr
7prCed49RCkqKC4OaQ+vB+77O3bUzN/jE+KlLa4lctzf8eCfzMn2dgxQwRnexYYf9Tx0NSSKJUMY
A5XmloQ9bObRwzT6ON2zskdZcyWt/7K9awwjY2Ld5cgx5SLmXTapfNyr384cIwK6Im7tauNqDcX/
IG5pSOlmoMTTM7wboFXT3+kyPNLMLTfp6MtS9Cf1M4RPsk/rBRPs98IYqijQMtOL+5c/CIKfxPAL
JWvfogvbBmrlMomDFUysaDmCZDWA6YD77PuczjAQHRDR+rqx4DxPwX3/eo9JEAwdmN53/KV9DvlS
sHg3W0oZ3t2/lJRgXOv635r2X2UwRdNF+tBQmWduQu74qheRgUaBwPaHU2CZ1U4hB9aEnJG3gbsl
GT8QcW/7SPV5PmsjQ06FURfiw+cuYnhDd5B4Hj3/ui1thvON4onYleHNblnQv1STOuOKfluNiQsN
cQ7D6+HLl438/sr+jRYG8oDuqNuDZlTEthnVzRoV4EqJNFyJ9Cif+OjfERVtT2fYNgpxHK/h+oKg
z+hxPDds1HgJSxufwFrrshnZ9B9VYxc930522BDvKEkjyrzJBR8/RkK9i0QW1rsKYpgSJfpYY0l4
eNTtOsBEacL2lTIhodd5bMp1UIjryh4mOwJixv58CK1UUcQlqAL1+B+JICrCIxRFAf+YqEfkl4G5
i13HaoBzbjyLGpV7/9keD6G7jX9ZUbkU9AR9PUgzz+MCDnosoztGPyAu0VLn55TbWNiviS31IvMs
UGEt2pctOo8EHPD4Rfz5wznzozikmj770jQcmP6NPDiFmx1nN1gAd7OO0zdXoSJUzRzI92zepIeU
2cOd+Tf3JMOXYXLENR0MdkVvMWHo/S1c3MBqiHUwBaEvt5NoADBOsVfJtzkwsShmLJ9sFx10Inkt
qU2cG2kod6ZxE7DcioM33+qwZIm8vbxMImBAq5YzwTAKhDgjlkOOX4y4Y7jYXpSQi/HHiTNQ3ib+
BCIUgAcKw8bRcI6LKdaLUmgf0ub8kD9hVeDHKxY5+YKRsDRgb0VeaarrPUybNMsGVB1NlmriAQV9
tmQhO/sOCzIt/R3Jnwa2j+qg70obdDVOLo/2x6CgV9F+rNRyJ4NQE+3MtqONNrM+pAxlxxpQmRL9
tbqQuApReSCAaw7y9CCGN0mN3abAX5sQO2vkvVJiOaO0UyWie9nXDvWMQXvY8aiV2sT2M3wQyEDT
21BctL3dCgpC5gng+l33kPKPzaoVB8fIwiCnS+jA/ObYSD+aBT6aQOZxY1ApuhAzwGINgtIzeUBD
x99cbJhW4/Mgx0iAlHpfNeME9X5wWVqRjy8Qc5RrRnb9y3uBD+DICk0fdpAGirIGjYMX8kcsvOth
CZEq21g85aEyCNlzqeOFSBb2z9WG2l+kFyu2KBXDjaFG1shKcWJ+gFc90Nnk7ml4Vuzj8rGyMDHt
mNNtWsyHOaqRFi7pK1SwDMMb+ULxIEZTyucW4Vu6et5QWRwXf4nqIgtGVyqnKeLqd9oIRFZFCYH7
AtFMBWLizKc/XIPuaT3QGQ3M5OgMfEcdLROzRhAX1ylNajJwffVar8tC5ftnBTu5AfLXvo5XNThg
3LrADmvgHNEVBa/hEm/tDCWXl9WMaYFdESls8kHrwbg63PDr2JW8r8Avv775ko8M9iLn6jyb1DP9
UKOguCTc4yN0bhn4nxkrCLTU5trfWQN1uP+Xpz8kTUTIBv1FZ4TXgGjReicSPyZVGjHKpSypI17r
+6YqwSwRjU+K4EmoFdhVLFkT462j1B1WmXiPmnUddBUf0Gv3f+3owFUDVfHO6zxT/q6Neh3peT2m
5QO0mqnbQLZ6lLZ9PI0HjRZkktv/M3LpyXwSkSkBi4xaWJKS4VQUSkfxByvdKpLFNN30a66ONHOY
bExopdCWNSMZhh2H2Pib3qzeju8TwiWApAipNn5hwWkk84OhWzb5Q7uy1YXTNl06VqA+YMxR+CUJ
TJPUMmY9lBQAZotB9fUAcLD3Acrp8vN8EBWcJpdgXHdBObSWX3WWJ2Oqg96G3AUnj3bHqGJ1fnZs
+renj7zyGAvfeHUdvno3x4VW0MFFJw00JOsY55xN5ndhe5pz/BK/Q1i+28/4QV5Uo4VseQkeKaNj
JurtareZapk80TX2kOBVfR0NEOsby/1NoHt335w+fX2hXNzKFk4MAMLwBINw4JpICgf5HoyccoqP
l6So8JT+5bzeIXYmYGe6Wac59MJpFpMo4xm0x8yVdN1gLOENaZTF0GUeD5emsf9Wzn8zOsUZALwj
u9zkR9S+mgp6vizMcu1pZsOB7iUNpYUmHhFBqWBRCFJ7SwGh/1r0Rw0pbrkRr4ppfLxVEENJnwuR
clp0kgFm2fl62av5qQoPl8zpZsAmcGMXyMuttG2XFQsenFQCKZbwoH/86YRrhiqOobGeKz3LI5QA
QPYcJLFII9DbcMCyNQQv5Hoj6yeolsF6krIdo3gFcorrR6/9QQ8ucypJ78Xsq+JCZXQkYDaXfUPd
uDFEAu/h1XoYh6hX8wQmjI0pkYUR4a1czkreP1Xh3T24p7QMXlVcZ2iVltv19ynmf6oF2ee8pgz3
bprTs9c6yuBTyQGUIH6Ywe/qnVDZMPcl9n7A3wGAkCt2yygZp/lS1FvOu7y1+nf5Pcqz3jIXf/77
wM+CaY9tuLqgEnItRc/ronPG69jenfa0JcHL9jzxouO6iJs1qkubUWmtdmL8s7RiCSQxO95iHfuP
lYgy1zSB5TBojM9azihVNYvMdnbFVGIaiB49GT9UfZuiKM8hTLKk2EMM9bOp3xLL//4Y8ssGsRnt
P60wz1aneVqJQ0fEM4wzibGs4pQE44jmkjzI76VhiDO2uI/zChi9Lvh9VR5wY40ua/JV+xJVXzLJ
Xab09Z/9XE/JYzyCP2ccPYapl/KB6MRH1sPx2PlaNeN3Neu3ufGwnBKc4PCpAxb/u0GKtTfNqo64
3hHIE1/Jc92feg7CyJkRZTHBCOi+Ye7l4uwqkHn1PZn9ArGr1GSoD8ALfvUNtz84iOv6dzbm5VhP
RPdlK4V5bxBQHrDtvU8+uWJ13PZ6RcaTZI4ND5LpZncGds4+Ep/kAvdmcngL+QHvCH6SnMjcDDLx
u/NZPH4mI1UJavgzESMhFS3SpGHG7uozyPrcD+yoGPCJD9sQXWY/THpABQyvONQWKRZkeUwQYWky
O7JEEuOItyxxPKcabZuTrUE0oS6XVJve1caeQ0GvHntLkq3slwN0O4gY+OHz/3rvndNjaS13s4U4
F5NIvHXD5lwa11vKbEuqMEQ/tNaON9BNi8mAQrNuF0Hlj09Vmt+FHE0RGTvBQn0Hy0mutD+jjYGR
+F2wlN9GJauG1xfo+LoonUKun+T+p03DHIVYPhtBUYHPu3PJX0WrjPOy2xObcFUjt4jGzQpgpimo
X4TpMlQe9G4JA5eMasZYEEJSOrGjKj3yPLYZ6r00DjrTjqFHsuw7PomdpAvnNP9wudES+8kL6HXY
E36NbEnwmZSUHsuzxs8UMglA7ombCJyVw4gKxITKaObWc8VukLqN57v0Uf4/sWfolz5pN++yCaPM
Z6L2aI8YZbGLksvcmW0v6wXiquONYOwJ42iH1DaZR+o9IIIrHe2oCpR2ShSKpfJMUDFe/duF2xwe
pyoAuvohVd8QqbwYLrNsjQgXIg4nWwexqLNjLu6REfVKYiUtAADH0syaaRs21YP6FWxJMNhhAQkG
whRPSEDvseiGz5gOSEebc4X+Bjb7OZfqJJ7ydi2JMJ3Si2G0iGFqwCAGgrI0khLAC0LIONFVwRIU
xSzZ0a7VFyZU+xJNzscOjkiHORyFfQIARV+0q24LxJD7X7MVgCW0yfHrJKwEFn0lyFMtzS+IhUkz
oeKPXT0YXsZi0jwSW+eyGOPG8EHH9dKjlZ4WXI2Jatx64E4aI8WodCRhp0ityRtQAelJO3mOysuv
1kDk5Djg1aTy9F/5K/6kTCRo2vJzmxrakt/r0WhWPwsj0rNr7vXQD7Ugdr6vFNiplS55S7fSPBdg
zCVMcy1vNjy3toki4KonCGGzRAaHNX6psYWOP27VRc/QH0gsWKJLWzlF+ES39k0XjfX36GaWTP6O
8DTrPa1a2ge3jWDxDu4b8GAD1humLPygo3Zf8MqiAt3cQq7rmtU9mHZ5x6BrdFUrFTHgCrycF3Zs
mJ2cosj9o0LmceHDH3hlGwp103pcRf4U5xew0bsLsoh7nvoKtXwRjZLeAjB+HId0Do3Uyx1vkQXe
xdDwVs8T50wvzjnf8Q7fP96OOni4TMpZUTUekv2Tk8j9v8WwLPXJpz9KCoDz5G2h0w/Oa5ZUrLr9
Ig+VurTzb7aY/Um5uabUFoDhdpOuNF7HC3ZiZFmeZLmakS19DwdtTQ25xOu2/523+vsOAXT0YHbE
2fIuVMWvr0GxMbyuDfXkD+mB1gI5r+zp8kTd/1DC9jgonqOO0cq8nir7f4IAoGyE0RdqPW6aGPCm
QiHJjhfR7ZALsKSCSGgVphOJNX7p6A/Z6C7uXvTZ8pYhLkTqIAVbHia/plQLTaTFZebpNrIiWgyc
FccGJsbWemvRVsGY6l6oLOhnnTrJmZpiUSCn8Or+AONUD0saYenLuDpbMg4YxMiImGhgYX5kmAMq
EA+mP9keSAhKNzgVjPMpdGJ0ynVHoe31lGd8YVtY2gEjS3v7h74ts4MeqSd4QzfJZReIehbN2GT/
9PV4IrcR71buC1J4tQWbq5Ia0XOCtF1JG5cHij6up3Dm6wsr5LTm15Kami7zVqUQ2pO64owwteVR
VMV+dearunH2QswzewfxMzkEt3CNyww+gLsOEgdjhpaixRReVrYoAiRihPQR7Jga5cMDyY+/54hE
oKqT9huTGDYQyAr3Bylb1rcOidEjDGo+T9K2ygsroXrgGrDIxuUMngXOVUKqwXsPhYFYfVgTJagg
98KuQMUNq3nWnOhXXo/KwG/jYJO05WGt1ekCZUikFtwWmewMicCGe6+GUg/3PrcynbYkFwiaE02n
t2aPGHI0Qtmn1onGmxLCVsrlpG1dmxGiKE5hDNsiFgjGobihRpDA0zIR1AZecQ54xwkE2rx1bfrl
HNWYvkS3LdayJNHDN3ZS61VmJU8LKlejGgQ+pN0xVEv9hrp1/TxE9Stu3WslDpzlEuWSfIUBYJ/6
KTL6Howy5G5RaH01vVe7VkqxtXBcqyNyVTyFH+IXKLRHEcLOamw6IqH34YKPvLnUq57Z1QGvuoJX
Z2AJvOjd/kw0C+h2IuVpxj/Sl7NDuNMYEzUSCZ1ERxvxfyMLISADnHYn26z9ik5tkXlGKuXMaNrK
JWi2Te3dla2Hb3llnSceAZ2/+eZ+tm8TSElpi0TIsaje6YdcZfB5oiwA58Kl5Gn75j6fCKn98UYo
4t/a47MyejIZQc8VAAL9rJrgkaGJS0MIO+fWHg2ur0+CNMVaxsy7HxJKYa/+EMD0EQ26f+vtXW3O
j8Vxc4ugnQBSN8iul1k3JPv5BdwaEkRyKCM0z9sfOO/hILxWL6HQHPJZKife46AXAH05d8BSEc9Q
TnZZcAr+yIcoH8SqjsY5eTm18ydgXQthYQSQ9bbuHuqePQHXCncsuV4A9UdKRElVZdEypCxO/liX
9Zpz8TnbfG8PQJrXI69iwD2R6XnBZ+Lbn8BXIHEeAIpWnHLKuhy/9b2lLHjtQNju0uoQVwp0kiHB
JV4HqN9xcxBMsOOFaEJdfFCylU0Ql5m+Yo5BepEJuAUw18kkCE2mtNoQ/5sAhi5mIXrTsc5AxaAA
92TkBP/LaIA51AH5ip7qbX7l1aAP7H3igKPwYkZEagK8Mu/CbKdZrcbJGICCmDB+6Jt3khykXdOv
qASbqnu3f8APspRJX9rC4egs659KMCxV+zkecpYHSdwweHJfO/WMjOKHWkPMAiSXvs3VHROqFq+Y
AFLnO3GxuKJ9szBIwJzf0pRqDbSpZkrRyrGtsxuFmwBc0b0dSUGrCwiRNwU0jadEiosGScDatzeL
yG2H0rovORnlK4ioGqgUDfHQU+syYl+n419Ixl5NFOUAqt+LX2IBSfZc1HBWUSf5uMBihWWKNY0E
mO9ba2hxfDbeNky3n8GE2PZd3zgzGWgl0JshRl7qL5Dgi0D7/crSw5ZDVFmk1RxXbO5Ps9zOVOON
N5denfOcLxRcQFY96Pz9p6zfydpTQTSE44s3fAXITAcmLim+8AY8InG6uX7UAgXpt4BmXmsZOZnM
/78rcZtzzCFyLC4dpT9zbVhFs1uyDY9BrCvTVtxsjgZWTCNkhG8jZE6f16YRtzdSWW4WY6d+zFLJ
cuTMykxdAAsU2LAp7AimtRiuGTg5KoM8O2Vy1qndmiNBkr5r+NpKMjItUCG1wTQDOSmC0nIVXfvU
lPA/HZvfja4zOmSG4MAIiak3ev58QroNRl1S7R032lw/CSEPoSoEsfHpz3j7hNby6MzgvPn+zdOW
UdtDgKNbEsfQDqwrOPPggEKY89PNdafyhXF7uSZVtTkmx1V5nFbzqW0c90Yf/CcqbILIgdqado54
emkSD1A6kkY7nLoNWYSvEMq+2XZBLhUyPdGZRqUYw+x6vdkEMgwhYjMqcaVlrtgm1mJHzi4ddLC+
E30rgoaXKDgeMg6Iy2zZbbwFyxgLPd5TqcacEn6qtX1/6bM+x0EFZHZ0hBlVgTW9/BHB8o5MU53B
B5kI4E8S+tG4O0pV0Z6l4wUODm5rJ5SQYDJ27etJf2oMEd7Okx0ASOSpthnu/pm9ONP36VTFBXKA
+Ilscx2fFSh30s/YouX7iSObbNscnF41Z1sW0zEFHI0OLDd7h8+uKbGF6nArSdHT+kLctH3LP+lJ
ADbqxK58bAhgbQexi1qqd73oWI8EhOp9aJRikMM4sq+YvF6E/g/cofYDLXOARcDl+QzF3QDXfifp
2RdwCCsJMU7jciLWG2yKaTbNZS7tlLIErDWin69AZjiwfmcfIDQaS4fWFvG3npxwt8P+9YM/rGUh
JJvii/gmV9PbMNdYmjOxpWUw3KNiVq+5+NQooXdQzpSMMuSusQilIEIU9DooDWrtVLBi40Sbi9gt
/sHHRvCcQZGeSfB5TIzyZdLuoIsDEc7TtDaDixlHo8EMYwcZvjFmmctbw01K6f2vZJLC5z4S9n21
wg0+/SSR+xIpdDV7lELlERpaiMwUwGJKFQAxVmrHaCgceCDUWZzaptq1SlDQDMKhVJkqiQJ4JFKk
yiTx/srTzYjzBHCVxBBLYvLTaTN3z6OBapxIZ9TmkWA2jM62Ok9eDXo2V5e69Yoao7ZuqikNybnP
gF7qB6qaX3HNGxhFr/eGLDJZ7Tw9s+Gq5bvMGDeN0r2kj7OpSfk6BixrXE4y+OUX1Y1KDuz0aa9q
xI7gojtI8kjzw0hms2WWvRpTIXUTbmX3OezgjTGswkEQyEFtHxXAcErWJERrkebY/ZPBby4EdmOi
cKmV3i3i6LAU0xjXBVnPtYxShNrK+rYeRGx9B3vFP1AhMpwkDK0bhR0boZCD5xdaYfPugtnnjIf8
VyxlRuf3T6/We6Mj1d+WK52WgCdh+X5/EkUnJ8AFArGSIV/QZ+LQYS6lG553nRjXOaNUIppl6W83
Wgnu/zf3Cujwcb7+as8F9eEcVZZuiXV/gYLdgHKE+CksYqoIM/fgybxgQPyO5HDXUspcLAjzJllS
xHS/bL03gdRwcyyD3at/F1ZV+Tfxx7u5GZLLGinDa4vEqvtc05esLtzaaOUOUioWzxaffyY1Fv47
/F19O7XpbVutYAMgWlIH+Z4eFXwahd8bN5nC4AwAgU311EHBfTeXBjzfF7/Xzeh/sWY8GhFmmHWf
mbkFm2ScqgcxYog544RR59IDrt1jhjkzc2jp4+3+W7tJS7AMAhlbvG1cscDt3p1R6ORPdN4LkDUn
0HbUZ51ItfXP5dXDxYsfgw57Uv7mePKRjS4Tz9fkjJmED60wIUFXj4oR8Ls3qVkIJcnsPXoQ7Ayy
qp9eQ4lwND6IG8clL2eWb/klwMi5pJLQElWY+mV1ACRo53IAYe0n8wni0rpeWRiujhfwpIFdXIDZ
9YNr0rViFyI8ANNv3utE1/MjGUhe+qfIonfyDJzg7watHQtkqDVoACCYP2MxkK232kgc7x7IHJWn
C4ln8BNMogt1VxdSt/1Pe5vMysYCQnAFWPqCQrR2HdULBn8kxYbTPsrvRQqdRZJAJ51jbb1ml8EI
Zr7em0Q7C8bBlUCJuPSny5ghLjXfVsIZc/gIpe9i/p4gAJ8BCoHDVba03LU+6YzH6IxOUM3PA+xy
Z4vrlLjcszveGpnT9d4s7SZQmeuDyWcXkSevA8VNSnMAqRffYUl3K8Va3ECOwrk/iuhxoP9dQLl7
F1a+246xjFqPwZRpaXHhRF7HdG0HMSa6SOfYR5WAW2rtoHBO7lGaackt5yoGU9r/BH37BjcrPopG
5wHTku5/BhpLCqN51dpGinbcYam/dCh4MTmHZuJP3e/bSCISi+9iXlhqSDA+ZK4mNMP8OS2gIT8c
fGVgmvNu+ZZuK2e6Cryl9Db2dWvrVGuEaJ4FYBtJuSwuc1DRe8zliWK2S7J2/F84SBAvrwAGsI5b
LteK1dqund0nZmHAGkAM0vjBtxDz3HYBZheZvz+vbH9e5cgAyAsMFnr2q9VPwOFkOJZ4Bh5fiIy4
riIiNirFdFfsuS4+w6A+mEYvLDg2kM+E92l0cLAD3M7P84enqCK31SZdPn9Grb1UAnbRWs6L1HqD
i8FB/jzCSHHL42AKWjTiDcOMb3ImKS2+GISfEiVH7CrfaQysOPOc3IQgJ5gQbAfwrloswEKlVfXK
0T02znb0/BX6/RIZRnJMjmRaVpm1tOJkiHNL7iGwhUJWAbhd7ZV3CluvdKb6JDyoNtJOHhA4fxlA
+VD10g50OSKFkcW4eXiq/Gp0dkaWuUiIyTPEZMTCmbZb6/kHLQxrsdwQ/MOyRY4Ql08+n/d0ob0j
McG73MlLZvPNA0xZLyejGL2Baxs7LDciffL7iE9/RW2S9Gf9PkX0gToM2iia6GFf/L3hrmxam5/2
3KGf/ozfPchZz3cD5HEUfu2ld/0aNkkfXt3SLiA20v5fYIFdlL/E+GfB4k8ZPriqZhd8sUzgE/L+
k2+v3wNDFUSFI6lwmnWYSJqeY7VMvqWmUkil0Gx8DTIRAkoyXAwta/YpbcNSdoYpN2YPnWpjWmaF
jP4YS2aeLHgwyevEbxvGny7M0bvKX2P9J6sWABDZeXdgBoM87GtlQvoFaw8ZXZrWQJdYAyJIdGDt
UF/Bc+hdO2B4MViroxaLBE7Yx5zTT1AcTv4YOqPzZ+jifPNm8w+LYjPLRQ+Au918U7ksAo+CVOOz
ez5Ih8lr1QHIYqjOpQwZLtJQXTyO8fkOTg894SDD7eqsq1i48WkcEdNXZNEds3dwyWuS6+MU1x3f
nTALRRTT1cszFooBdsIhDG2n/f9PP/TPtku7hbcUzs53yATycYC94w1+9GNfIZ1W8fUja0mDHQzU
+rGTsqUxktR34/RBS00h6JE0ruez869EaUmonJNnFOcTemDDtzOQD6//jR0n69MvzmsNuqVZp347
QUYEw6RcHp92jPdiGGh4ATkaO2Crtw1mMU4EIvBSY7IvwKLLStuD0SaJ3VhDGhB7srqO/U/wXrtK
Ztl6fspvFLlxcfT64JqlLB9zPBp54BXbL2HoTtzXcP5dfrENUWOZvLxlA3Mt3TPo8dO0m6sBbwuk
JimdxT9tWpOLGsIe02JaTfTWrZ2T2JyR46IbG+K23JWoHrV1H7XDPPSr6AT4ZivQ7NFB5nqamHSf
lByCCBnA3H58NnJg8OdJuULq9M5E49kCMQfKogPC435qtzkUPzw77h88pTnG/eKEFMOnnn0JgWqO
BevazL5DJz9otBmlZf47uHWwQhbYEy/2Mb6CF71flMODSHDXfivsUTTB7sEFcpvQQBjQfNa/heAJ
RA9pbHIADAN3dSIdGTzguKHV4W1nYePz/gn20Gj37z2TQUiPM3Jow/8rCBiWKnkEuosO9u23FYTt
9ZTVrA9d99IE60GR7YbtPSg5dPeSAmQDxx73szD/uHZGWJw39vNcfEfLsG6xAGTCdUp9ES5Dg8NV
l6K9BCdB+mTABduZWWFZVfWNJlZtyqnq6PtH4rHVoPI0cP7c0c5jU6ewxxpKydydGiAx+WCFxT5v
YGGC6LMrBMhEnvzOlqM5uzxVvmfQGVbJBmDzvbsu/vdJwTG2OlnMxw2POnXYvj8Ol38ApVz/xKOg
1fBx45ZFVOIgvaTXfCz29grtPoZftYE5AvLw0tibPvjGBOjDouu4TcD2fBBd52OebuNRoq98j8wQ
+H5p6UD+L8roGvcLVBi1edIhDHjVh0J0gFQ4OMus+LXu3Ilw8dknpe3cgQMvvKv217NsQNh/MQmf
/6R/5uxvyyiB555ozYu5MBPShxiVyxGyHSLzc1/aq0Y7iiZkX0Q5hBbXrJZPUP767Ab5IU6ryyG8
4QE2RVHHId3nlw0DybBy0HPfFPR5URj2nUBzmfK9AVk1xfBMZuNpRrn3s3k0eoYHELxndNdSnXGe
uuQJmEG0gduDcAkoRhehIVXRGse5/UBwPr0IQYLJGI2NWy5tEGv70lmZp+upFQT8No35yQ0o4Ebb
480W6ZkR4/mTmpSp/dqWFqvcMFT4youw7+tz+vHiaw4iUPHz88+E81v7zTLFNACCh8koUz/s2KJe
tJ4TIhm3IkD6BbkCEoUWppkpysTsuo4jFJ/WDm/ptqrCle8xuFXC53Nxy1bz5yyF4cS6K4gRqI8x
GMWslaQ0qmW+bGcRa8VfBAybYTnqXy8/Rzh9GcBtpG63zvvsecx/8zakTylVSgUS5V4rEP204/yT
KaSXWKgGPBybQpJLreC561WpvTuzK26Qz9RD5YjU2qDsZoALpwmuOxxFoxNCftzWJkyxtWXh0tqZ
d5r4qEq6KKtPIOgvyzla1prNG9o4QtERbyAKWAQsi4tbfpxMipUuTqL3ZurjrRma9UC9mQ7qSzWn
dD+b9SBIUmxLLkHjQW3LjJdPK0kJRmx0q3iedeIAbsTEGHLpF1yuYjXur4Yx+dqNq7mTIL4nJMJI
pTTfVKPmCA1jLUYSZld9WQcTn8qgahQKOiOMOwecqkihGo7anY/6pxzaVRMRMmUM2/iuoQAnmzxs
8rUgDvGPMz9ZfGXnRuFjBRf5Fk1yNErGfIeLwRUR2Dn4ZKEcCBrnU67EK7tVQ6qsMffC8dCm6fWM
TUVO4jwym3/pg9lTVWjBrw1J3T76tesMnq+lktZyGkBXewMmZAWLDvKs6TFEvdIuda2mpyI9K71a
zOaTLTOYEiqDAGFjwfH1+KV1eS4kxNB4v4R6iU+Ccvi/Wb915X8wryMQr9YXeS4L27L0UNA0YkBo
i8Zp/dxlARmGoD3wiuodJQLxskVGANqv2LTeVqY1XHMHhQPP/K/PcPoWRCMK1Nq/+E0oNJRaPR2U
vIMhQJ0G+1bOMhlL0Eo/NBeM03gL03NQc34+X996zDRJLdTFE2G/KuXnOrBrZ7wjDxOx+MSV8fri
g4Z8VqXlwPPN9ZsK2Sxyff7oFnyDiJPUoL+DlLCdgVRDuqoP3FR1Cd5uh8fTso65cKwhDmiiKVvj
IuE/hYcgeJMimpfCuAj2NE5nRm7GJzB4KhB7C5OxlvVnQmCm3Y4H24Xe6s3cYR3mwU2/lkpDdHi+
znlfnAbSH/3cQHVrem0Goo/ehLBkLbgxdCz/BdGJcV6dLyNTC6YSWzC9e7JjmYWsWjOPlZ6Epurf
VYEcr0nAUIl7hsszHTmtYR8Dz9jQeD0H4UOVV9y5IFFBZ5GbUivA10re4NsYwshBpvqsvNOFR23s
f4v+TZXPmGjbeXROhFy//YBXAfqQnJ2pSqX8+HC1E5Fw7yY0MRaiQuBQZ7A8dAt2S8Qxr0kN4XHA
LD1RVLFMHug5sRtvPxbKc4Fl4RwEfWxEpDScZkWrgov7n8kR1mCVWR3QArQk6ptOU2gMMwv7HYMn
ZmyCEHM0ATnX6dASJ2rIxgNQU618jmTDul/qReZpFbA+cMjKt72loyzCaCVRzDUvLL4UHQhVPADY
RZWJzN5HSJXcetQ0VryXDvxHcgejfXZzA8M6P46fCAf2Ezhtz3wvJKyDdavswbO1gBdeRIMOTIDB
0SilIr7d1rgzPAOnNEOSP1D1u6RpqZllKwfeDiLPDDB5GN+0oCAi2ezmIoO1urAIP1p/1jaN4ko1
pvwjRgNU82HfpuGnqtzhaQEKo+u1IW/aOP00hiSYLdhaCAxfuXREm9SJNiTl+Tsu6Dygbi0y047r
PIQIl6UWataVRDx5oYdXO988R5QSn6coCXwcDUQ2ssye2ec3p/URSE/KXnBu91r/jFC9kwhOEK9T
XepnMKdJ2/x3J8tLBdwISZezZLBhkfabMVKdQPXusPIpSXe+/Key6v5cHtl6VLjM6Ulof023fjxr
2D3cWNPc7XGNOwxWMeW6rq4JMZJYkEuFDv2XXgmeM5Y/4ztvWxR1Rs/p1C1yrn1r8LPpC4Q6IimV
YXYU611viXGhV6KyN8FHtcTNtufrXiuAywucgAdnl6FmoUCohXjckPIt51BJ+/Ld0kKMToyCysle
R6nGXQMv+KmgHVhTmj0IypvP90kXIvKpnaa5ODqTieutHugJ7deZ0UdZNaaguQDQj8tI3vJFXp1J
OZVfDZe6mXSDIDHQkJ1M9DtMpwaDaiNCPnXkyQsME/PukHwRscpl68yOS3r6+EdlLuZ/zZ7cYEzE
Zc1EEHIYwPO7OXnKeuqUiOQPPOIzdVvE506bYYQ31FgirJPAldneHtI0ci3hdJBkzK6bJ8F7jf0d
qCD13u+BAgFFycAxfwvJzTc370DAzskCeEgMHBUQTxzm8sA19gQKupc9xa8cjSdw6jYqT2XKCGM3
AQpKjjJTEMY6M9OYUzlmiJS8idJh5vfYjY6RDCgDUgkskr239/tAbuQiqBGdxAELFbWPV2jQ4iLq
q4E4mG2Mpe6hrMQA2fesjjArQNSdc/3D1JRBwjYm7kewQwOU1qvEDsqfIUdkEdStoiY9ZKEsE9yh
0a+xttelDkCW2bvSHfdEDS7V/MVHrlFcfvzXuCByvQw4DBpml19TH1nVvNFMR+4JGkOJ90hNkYug
pW+beMLZ/FYpGXMWCAxOsV37p6/NM21osvzMYK2fV1WDGucZmSyrARKzvT839C9DR8pbwSILuWAB
oAN7u6weD6bLQTSqZ8STuLwcDTOPuJ2ma1iM3rI+R4bAJM7/oImK+cZctSApgwZfZQf1PpwBMdt7
t5HvgIERRJJYVAWzk1FEMmd+4hwHDWfqXal+umsNYE5SPu81DtifzfOiLwF2na4c6x2flmkOABh1
rh8HKAWUQkW3MELjXmbq/g1diDC8Uq+aEjxxOXelxl08MhNcdK4iEEHLkVfju1hWLWN2MxuK+qUB
LeEUdYPWbYZHJwQMN+2y3taQOcMZQ7niuOBuZGYAc0h1TGJ8BJcn/+bmrTjelpfQwxDu0AE3DTpN
j92KV+KVMAEQWN2686AkmI5fhmV2k85DzvlVH2VYJcWW5HGjawG/Wg16UEBY/ZW6807fZ4dHtL4i
U4LNCuJufG45sNaizD0JtSIl+Hnx3M0dWquxNPiN3qFuLa1kyrCsvXe97rqTdoPBxAK1T3RVKsVk
NxyPB54x2czl/n3sI34VVBSAKFqT7z7asfhqRUGIVM2dxCqmj1da0pWPc+gE55XQFESQZboxAagK
Yy0NIgZVIW5FfEbJvgr6gosqmPPYN7eZnolHPIgABXj3TqJxMtaa5zJNFW8LNv2K66Ev9pNUh+EX
1mAOit9u3NhvXoTtA+wdLPQRVhzCmCy97Dn9aqKOR1oXvDQQReOfrs8EprpkiZSfaSocJEVFthbC
9c6FkvyIeby8WHh/ivgUelC4Qz+6K99GNMgRw1D35cJXzeBtqYd7J3Cm9Lw1DYWsg6R63vrj8Lxr
9k043qR/G2bsebupe1zHMFsd5DGEHevZ7NTV255hVR3OUScNGcaRv9NpZsA3hcNJA+smvjenkX5y
3MtPGbDZChmmKMklAObk0hY7vjBek9pZRWCvGoaRQVUAJt75M+muGvaYUxFVjtQYDwbkuRzs3hfl
MTOx9R9DEKuqBWZjNmf5qj/ZRQhGnAoYALouXwKMQJfvn/4XUeHWEjZFNNPDzqd7YdSEMfjVhF+0
+hL63aq8Q45wp8eLaNgvGSaCXmKl9qkJMPEB12RS/1t3+MpKs3RU1f0ea+PGluQhlhWKjrAwYW9I
KfnOVsovf4qgkg9BUzYY0CCcf+VoQ4eSmfhLmHuqcNd3+H9Zrt1KZsFIhoNfWCKhmIcfBztgk7NY
TuPjrfkUcnPLnnZ4jZzgLuKHmsh38UY41XbFpHYU47sLtI5OW8oDeWB8iEKJEqUPulY+NsAYUK/v
C+rcWk7ZIW4SDjZrb6voD56RU0drqmHVeXfh/7yFp+X91YdMvDWk5huseR/24e+6lU1nc91wZl+y
taTl2SnBJSulXQ7k05AkGJFzTUkFpXQrNzt6qFb6O5tQMT/T38dUiZ3RQYXa6j9fgJCY9wYiRMMf
TZGz8hftIhTIBBCCqisR1aRX1+3niqIcmOHw1YPGyqOshkKfWK2Ql/4VZ4bV/5LJaPcu7Hx/CRde
uZW2xhHpC6KZ44UzAapir3kvTtFVGxC+4UO4JT7Fe2KYUMuvdTcjVW3e7Ah3BYdYzc/iddbzTrk2
BSTsguomD4XypeKbB7xFdoXlk2PgVowELJEIujKuq9VMLtLu3PLE2MyPeTyD5FCttkNZejwDO4D2
7SHEIJhig8oc3uBXF/37e37MVa4rvQJqBaG6eK5WN3jW09ECM3qz9lM3vG4Ly5Tf2u68/oGWnV44
XXHJhuBOS++ggk7IsJlE591mR4L3EwGC1+tpIMgoJMFWpZbWQMhfwprdIDIbVkbUgnpi1YHZkwQo
JW8ik0pxWi8ihVnkpW6PX35ubs49isWGrsjGN7Th3IRVkJme0V8+PoL4cpD5IOKg9awB2F3u1w1S
Z+1zIe4+GWZXA+il1BoU+/bHyXmU0Yg2t3iIGQLtJ8hXT25m63c3HFMuC5af9srmoWVVjj6nVqRE
3C3QRf4nY1jPsEFguxLlwrgmx6l1kE/vvMJFzm9hTO6Qt/RX9+YJlL9R2xLgSO7M79kDCkFUysU+
35vzOtnJzwC/w80WHgM7FyGj5XqOAJpEDcXmfDxFXS+VukahkVphRPi065cE987icfV70HMzPPKU
qMiq8dnixrrcdSoE7h8R0SdrRurrRl3VsvNisH9HRbAVcCZp0AJVCjVOES/9PCOl75XKu67djJGT
QP3rehm4BHxWaY/E6NqXcTaL6IFZy3q6MMRxmJMP5BygA16wVf3R8fTaESmUET2s6WPRW6sY6fNg
5/k9FSBtvOPwj8Jq0vYaZg4M1o9G8sadZgGEJCp18mfexWOfbRHyyomjPMShi8Z3DAduTSmPvy8V
i5SATfhhVgBgSJY0SepTyLsEqVyIdoooN1+IBmrCCtaYwesaLHCGHPg/jg4oPaAJq6srItzzWps/
YU/q7Bid7l+Q2DgW78JmNwmaQs4nF5ayaR0H2xuN48WaXoQ5KlEWp8VKHqDVnR5vziWNRC/SIBN2
bID5U7eW4uQqTf+Delu2psbxOKQy2wKvIKFlm2E522DhD36je0qLj0Z0fPOAusEMWNfEpQaGUL4o
fOsnFz74k99ZDX16ofCFmxWzOi5GWl8esDbreDPURl8ZitxnvvGvF0xdHbclKzpC/AjAonFc660h
UvAWZTAgC5ARaH7ZPOn7zlm0tGnoYT9hFz/eudg6QycoT51jy0noyzNObcUUGsb+TytXr7H1LzNu
DguzPggzKAbDAtu1/43QubZeenbpqdjCAt/Usk/rZaCBOROx4ucbqAZnnos/AWjl1n5gNo4R0d5t
gHJZ2uwnS5JcH0jAL9BtIFi06ss+icqDEQ/tV6qTW6Nq29ZSs3VDjZyWVplSFlqcLN34Y5myAUqp
s6LNJ/O/PioQT79Q8VxM/RTg3grKMg58yAf0rT+ZqzGhaevNeuWA24uF26l5RwKd4GaTQ1o+ZShm
vrnKgnZ2biOk6YVbzugrXM5HU5YaYUSnJFqVNevLF9JbC3BiC9r5J7QNvsRN5dD6se00geIMHdnN
E+64aC0YyudmTbjPUkXmyUdnhxZDyvOLh4itbgBV/zQ7M06Qp3na4Jqdmo3nQN1uWlkPELSfBtxR
1BQpf+xCckiBFtMGfODvYBsUull85UJ1fReF6UM3dr9xtgNMXDK29pGxcTiwVkX47qMKZaUMr2lZ
rOhoGSJZeDBC2jpLcvhjCWwE8vViGGxSV4jHnGh+e/FpMaNpEamSiyVybjCAdJg/V6pvjJXeN0XI
3r/OHMOiKHhp8CQUAkpiWbTWpR9mbS8klo6SnrN7fD3St3k8dohtEA8LdIHDPayFD3ndedsWYdqh
kOBJlOlOFrQK7K+D4LhcA4KH0YoVnWAvMp7fvAZHpZpw/8eCznLe9PqATTV65e301WqxjGaohTKt
+oSaTdsHc1Qc3KatA4nfdA+2IWegfHQ3fEBjcyk+vKl0TPsaWAO0RUUc+Q+PhEFQLThNLoTXVOkj
bsQXnsAVwvxUenJj+yVdqzKhkBP33bwywpAAiobqNK5hxcNqLwbvbZFfWL7EcSV4bRT18nk3JuVP
Te2BHD3x/hvoplITZPU1X6laVG0Lz3eL1X0pGAujOB12SUCAcOYQufohm4tpJ4hgue1Mwz6k8ZI+
hlDNU6B/Am4YKpbVJsjxl9i9nZVO1VV2+yHl3nBps+nXufh56kS3lKQzjWzGpy/v24kP3xfqACyt
CC84OyaYzkJUhAaK3UrT0mAHQV7wt1YVINXPKcXm9VJnvLxxTjtfoLuGyedZ7ts5NFNPbLJ+91yM
hRkByHWcp2AxQFg09cri5flW32MaaALb316yI/c79fpsHwwiN851jXMNQRe8bku2eCaLi4H4bxoO
bY4mA6T0cLOq/WaQ9y/ehFwsuFyXO97bIHLHZGp9XvsqptRcPssR2n6pIINekTnchk4TntRZ+0BO
y/nat21EXlRP0sRnSPy7OISZYxSNBJjWb+ko2J07QLRh1Xj/GBEVJXuo4CNCxbqQe8bTcE8fQiRl
qUUYqNEuY5SA1+cKMzW0ctS0hcPyHodaaypuM9tdjI3QvOs1pAzENa9QKFq6YmsPbtQXItoqW8jO
tZ1JNF/6LbqkLkSxRBnP+X92AOQ4C9TTIFg7NonEY+uZaLL7fYoXFXhj++2PwaYU9unANopHA8ct
MuepNurFGhKVFOYrLZYdwY0KLezPBNJf471yE6aMCpfGfdalAF9dWSqY2S4PkWE7Kq3Z7sSCpNol
AETYjFm7n/NbIrO6eFyhENkb6V1L3WFpBcOAIrVGzbVecniouBr6QYaBz7hVnn2Haf+1cRuawRdx
99G49jERRlSzrULaK3s3PojHkw+AlUMu3B5Pi8qMktid1qda6fuMOwh8rhZNRhMj/k99lKAKx4pj
OTgbxMRDFz58+A5+Bdca09qdHvYY6O/h74cvpVawF6C0yJ4EOZOXwL31fUMEbI090Y32RqE50Vwj
G1bueCU63LJFnA0S/J1HvkwLtUaXZnwfb5dZfshZF5MRv6rkIE0DbAVFj5aF8GprnLqQuD86eWjY
i1n6L+vY4DrD/07ntqTlpM0BQta3qfgNvcde1jwLqAcbutkezNRNMPYJVeki5o+NvgkqhKfg+eSu
kI/2jiUC9fNGcyhCQhG5MocivdqIM9oqgVEoHPcg0E4/SzucfU9FATa3N6Dpn/BXlwQS/Mlo4nrn
tA2i+VXokbLSsTlmzrUwwbeawbdBoIGd5V72s9rPNcov8aOHCpqr7r9A6/Xa/IoNW+e0Ca+Uo6pv
lpVPy2y0929qDDxEIxCloM9Wp3ld3lIlOqKgfZWr6ZqJyTUAHMAG888ihN+wKPJYdH/eldsd74rq
3j62oogbX/RrE+JWMCqfggYDl5WBL3Ccr/3LiKnVEm8lC1pREOrFa/GjaXrd+47HfkksCdP0vior
tdfOeZtFnbTGfYQeKj0vSMlNbHrYtDzHJ9hWgAVJY5VTmecRcPgy2uC2l5H6a5J/adcDG8Fw/X+H
WDowc/IVtUugQSV3JqA9zlqrFUNhhAoMstOiLTlCw25+YRu+MnoV8EuCvyQPZyiHCV/aaL6Nt5zp
yr/fyp5L75GYz6l3vLUuJgCC5fB9svBrOT2mIbLT3eBDnkdfLbx1TNQXoUjRwhnvhQF8uJcUGmD7
Hlooz9Er8Z+V4IUbZNJ+WmAigJxWwR2Kmyj4ut6fu3vqr6F5Ml19fc020+BDsO78OFpN9ggTaDVT
NYJhDcFhVBCH0TfxAIwxFqHXbvunIk93KZ5TyXdiUonUtH11k6QtC8bVLyrEbpbmnZfSeHNz70NK
aKolqayZRXcVDbiStEQUJWnH0Qu3LaB9yRwFNL5/a4m6WP9mBm3Sme7P+XvHt10jcy1bmTnsevpy
+44AHdGrgoG8u8eKohJsSlHHzhA7HExDGwxCbJ8Gfz/vu6cZRhWtKyFb/MjKhQkM+2dKRQsXulDc
Axz6Evv0h4NLly8UB85lXwuz66AajnK/NCrOBDrmcR2BCFhquiKqzdBbTqhCAG0y2P+JMSVPU8+S
JRi8ePtebUMbaE+nF547r8IDaja1mQERUKAacmEyuXzd7yHwPcd2N6fvijDqkSfwa1+PmYRh0SnQ
7VsR46odzSDIPfLz3IGm32CoJ5C+N7s7O/yJBCZhpIR1SNQ71W1aIPb2adOnLYXgpca+ZIYXtCoX
EGfWDz2bYGjBwRphE2JhW0Zpp90qomCCFMJVbaibwUf3JPmXAfkQGl8Z6dAjalg/LCuTpEQwzKBG
DJCcoavitI/iJkS7IIEcHmiwW/Zhlgp3YbIq5cOy88A6arM5LcDKjOfG9DY8S5CxOZjuUb2PDfh/
nUMsNdweZh5RzOk5UFdG0lzF43YvgKQW1hYwh3p9PyFl3sdkTZCpEa9DVqf9mhbqdp2DpjaUDJL1
f6gcXfdXrhJ+Ldp8e2lnQ7TiYhSllHeD12Iuu2FDPOUwaSqlZ7eE2X/+ODrBm9FOvxxFnpS8UEF+
X5SoZGzxQBbVJZPgpM2zDkRNMKb/T1j/BsURURSyUhBnTbwTb6/+FcpooIvFGUbAJTm+x4hje3Kq
Cp+huO/jW4Li2e7b7vsJKZ97GmVHfkPqNtVPlk0EfHvADaxdWFFStxeZuu5zkGjt5Gw7VM5kSaHZ
MI0/sdZ5sNRR0DNy4N1lTDztvEEgc0HXc0ut6YAnZRu6D5LaG3H8cvS7TgcgGRM81b9lQtuwZzZm
eE3jsXkf4yG/Rcm2x+bzhwAbN6qO/8FfiAOdn6OSawv9goqHIj/EjB1OrB17Iow5u06COmfFXlky
Y1P68Ta8NSg0domO1sEkp2LDVx+YVc8vj1whizC8TUmxx7woDTaOk2RyQLXeqeVKAEyWdScbJz6O
6dh1wXNIZaDc9NIUVszZG1o534+pj2ccr/rtDKiIk8l3meeLPgjPX+edNksXKtPrec29BzX0ISv5
eVT/C7NeO624Om4Onyr/22cVLjFZutzxEqmdX8gW5LNYpJnplz1h9Ey0lqMzZDzV8yLS4aI0sCOC
NTtNTSKgU9Cjmw7N8J9usK8LUDr+her+TVOfqD/Mb9jia30R4lPhgbUDJWCg2PlUikq16UFWjdyL
3u/q7gChNSdKnZEZSQPPsOY5daXjDthRNRSHJbeeYZwd9lE7Bf5DvX+pu8XSk+kRtke4VmFDM/pX
rnVwUVsmHMtqiQQxDRMXIl0HOC1WbaqDNOcx/9Oh8xqJmtgQtjjVw7D1J799kv/XSRBwYcoPInzu
YERDEYR3xtAUP8IXzSgSFqZasvSvae7gm91kPq+plM5YfXIVrBKNBRmRhI0RZoRNAP2p9qy6iJTF
tIL9Pce2pKQmo4NhxsWJRYughpSnb4/hPnv0isqtxUCg+FxOBs0oHF07sEC56wx0cQaFQ/G3rwH2
8rvINw3y6wndHBoFwro6Vuy+kZktwaybJWBGKpKUF53IC8fQuqbXXuWkUQqZkfBmhAxQBx+OxXhT
/cuAtIy+O4ovQkMuX4l7UtR9bgFF99kd0F4W1q1f3gfQivSrZy8B6r9H59/fuWLbvzKIxQcyEx0r
I8V4Ygz4WLhJDtHLcptZN0oTGAGlVcbJwybIK8NfDgJ9LbxX91TleP4Y5LffXMDyA5l6OTjNSkQA
PKrO+8mW7rs+dJxNZPhPX1/GKg3O7LQe70sQuhoVrxZ16pxqReTByngWz4oQtSbT/+sKXJcZm5m6
Y7gNkTYVa7LDPymcrNcSuwyytE3RjGMtAQ0Lu/cOcemzFJYFoLxZenx5LPRD0v4U5J9+NJ+ay3ue
Gh6QkRCF6/wLqgqxQwt+3RAQXh2M3Q5JWER3o2ErSPrIgRE9iJ1Sbt4ICoJh4iq+xMtmnmO5YPZI
ChKjoQ7hG36mJAI2/56MoOQoOJqOPciz5Hr4BqvukWKZiY0Ai1ekl1EjXuvC81c+sbl/BpNwlI7F
KZD4opjzQui3Xjo8tTp23OUs4xgzs9DtpFG+ytnu+O5U8xnRW6mHTpm2OLjzj8w2cH+NWfiDLjhK
DgcMfTuZvEq64WgNSN0wJ+NMfbWoNmIeqJq9hauSRs3FiBMFh/IJ5OraMgNiaQ38/58Gr3cDWuiI
cCSnJrfmh4EC2I/PZWkWxE3CG2Z6JPdSj1wcg54Sr7qhrk+/Ahr6X2OU1+l5s+cbCbgnpPjvmCA1
+BfMCrjHUaGgoss/BnKIrHy2vdcgNS2RBeJlCiAxg2fbC//8wd1XqrIF5AIbf0xP6YlPQdbXQ5hp
G7Hx5yOoNICc9WO8etWWfMKlsY1kxTm+becD/iuWhd9tIFOnPo8vy+DoRCrexuxDIwflAKwgESfm
1BqPgKR/eq/zjCuhenChN9THNhIaP/lbNN7KM4ubj1uoHAC6DzE7lQP3H1G78t5RqEgFE9TURG8x
tPnNw+Scl2sUjfc3kYF+IPIKEs0EUTe/wy/0FLxdQH/nZUmD0lkaa4gbQjZGFhnXQ31sSLDVIpX8
OqNgMNDIZDpIAYnK44YuZ30rPdY6U+eiyqdFvruH6usqzTJsxQ9qYMPwwvlRYE5wCtO04+MzBwGL
pz6arZF8fGNJa13fT0Vu5udh6tUHW7mBTTEjlyXG9NJ0NfkMUXJBVBy9r1w4J38lvxNRJZsjUoq7
Yw11MekO7Yrn2mt/zDBK/P/gdNxlmgVPv4nD+0c2A4oFaXPeMJge7uSl7alAcNvdJg900VhzAX+/
CyOgJzYLhIm729i/2BxKRLykrqL4RtLgO0l0hb3c0bY9lrAxEKeOvwzn9PyCt9LWsFwhNXIIsldH
+KP3Bb2ea0ldMD9DSdhI0ltoSPL036UFUsgcgDsCiTzXIz8A1UhxCeMGOv9RToKZFAMbfxGdibmy
3SF2Edf+oi21kC6Dq1xqTiOA3/VYZ0BxbvLnBi7EDXOdnWO45eyi70m8PK4HpOh2j08t7riNCrbe
ZcmcjeIaxJ++gRiw3k1au8Kwh9SRsFd5SOurGPVgA8rd5Fx+kF0/H7w1SHiityYT6brInNMmaKwy
Zh0r1OnWcGQCmRv8/fOOn+QqZnhDa+JvAMVp/AXnGhLQbAAUXthR4h5l0k2LgpDkb/kpGRNCGP96
qfgE4lDQidhT0v3SHP8ysrQXiMfEGu6dZIHKw0UVsjjMTWVgMXaWGwcqKrebQw0g7M0uSDV41bYk
60zbyLM5OA0PG3CuGjEWcYSyhNq1o3IrxX4MZKYbOHB6eObASLhYcUI1/wFR6OXDibdXHW3rSD3P
XpPo3ISeb/Je3pwbXxu1eAXCBzCgQHaovJpdQ3AQOt62ahr46s1lyK6TDvEYL8per7mkGxsCP94g
xANX4sGaDcCjYqLlzeQSXJubfosInr4aujZgprLXnSu8rMJyMg16ISK/+whmUjOo981a1qVzBOjK
UaAS4NCaB99EmSPyULQfDNfu5rrMAkcCSbGBOnETgRJhmjcjfjcNYse6O//y6uKLKJ8hncnOm07F
b+o+hgwuOO73Q3pBdKxrEeQWqUHI9Y6cVLTLAWRdyTymRMddY2031axWqCKYUug96a5mpRHdcO3U
57vuZogxtuSt/1ZG3EUSB9cl7pt0A2im4v5Io+tmcQiixtGWAOWdgVSoWjpRs+zjlYKNXH2trPz7
LcPLc8m93X28tVYl0IWJmfvP2cV+N6iRkzHGrDLKgrTxjXAn+1VhWVmbfBcD2V6Rq2FPIeJdKtz0
inU/PBmJeTKsKgxzENKa6c3qWmt7ROnMuqZWwKjzDgyzPCQeivdINi+pMDOndKHHCOUB6fEYInjD
E4Wf0egs9gbCU4/khO9iS3EmdLMKleTRhfOw7hv+DcMILvQVM30TktZAjxOaGzK0P71P/LjKyxtf
m2SQdKnY1LKz5RpcyHFoceuRsWiCPUkLe8MnHdpsKTLA1y+V6wbru311cKnYC4gdnf5MJXGJDaT4
cBOFUCSkf9ek/HTxOtUGP7hghDLL+NkS15Ave9OlusCktFE6D5dmecdn+RgF9JURWNvaGQWh7LV1
x46jSxbUUn175N/dQmeTQw2nI4/5LnvJENKDwy1R2or/1ReDoOza2+6pOwazhLBkcaKV6FqfMkIs
uristhuzUTYTjTYzmxYgiy+12SYjrWyBCXbTG64UHnD4cJ0vlT2WT0YX1I+rFVsUTGZiZrrodn6t
k31f9aD9Wn9OorIrqmZs/yfo2h06UD3Is0yRhSUvsqJYsXXxPk6ctHLlaDOmVMQ+/uoA6DpRQVUM
nt877/ispk6oC6TWEZpOuVQiUS6SOc1lVRIAW5U12E6by4Uaxjk5qX0XQTglV2GSVYJd0hotRzTb
Dxqiu0C8+RuLoRcT5ee4Mbwe3tlPV5f5xPucui0sm3NPmL3gBCwSBVTHARercRSI5k4O1jwKAfoi
bUN5XgtwolAEB1rsigG13CvWGSUV3QfpCPRIwul3muWWUDfjkuLZGzGvAnUHmkg04ucoPvwGIoP8
5VFNd4/dqOr6YThwDJChNLr4NunnMjbsOWaKpXDgPmUTGwrRhVPMsQ58dPpD7ySwgeVFcnC0l5Z3
EF1Kz8mlW++t6UxxbIPgJu6YkMaG/b/TLFB6qAnyaClJR1+YX5FI0qwpehL1IsL3L3OkO5SDuDE8
vZ4bEEODeqTB2wHToQDZENdq6KvVNjKREMx8MSOw5qSpLIF1l5ZPZCC1MF3sIV65a/pye5H2CA4E
SrZDRfIjFZ1zTP3IVtXy4B1OCVO2J9BZPpm/7O6AuBntLyl0/nAKyw+AgxaUPANe2Ru3NDOQNo4r
OKXntt7K9PX/t8hbcc5GOtHqOEs0hOAcTkQfvx5/xjzJ7qysOvR+vAjmVi2Ko0gjQvoyNgZE9MgB
nheo0NCR+PZT0DSUdBwRriqLyNUH4HWGyyYXpi3of0lkql7MVrjSWvJMcmG9uhyyQ94vEmR/nia7
raQKVuoV0JCtkrQzPKgAHN6nqoVri6z/fdygSZcZ8VLxMiUYxoox51bc5KWWOoVJWC9vqjoFdzN8
ivJ3pfChhG1NP62Z1QKJwUp5ySCDV7FI/dCZ7VPQH+DU//JMV0FhsvgxNS18OiAjC97LO8pJrgiW
uazgwTOvHGdpKiTLubbWJ9AslUhNE6sRNkBlE/wxE7v9F5X69q5jVkAW9Ecs1ICOwPkLC3JDKPHM
wMerYgRUUc0Atwtn0x2/I9K6h1SDpBnlJxO72kTQH7Xv+Upq+kLg94vTlBGSMAaTzZ4Zg7l7F5WQ
oxyhyu9PUFqbXZVCmLMQpAiZtZXGTJjKPjSv/d5DF4syCJfQukz4WWt4bwoYQemB8BNzJQG5E+lA
/O9YI3tqJtjr2LxodskMFq3xdWlN1XQWcloMOJv7FEfWWXLEJubh+WVCm/StJf34nbmb2+y+lHfV
e3lmPNukCvsQ4aXaD4/Bp7NCdhTX2WY+fqkquHWx9xDu/DT+0GuJ0Ys4FzlvDX/+FkXqDlZD26TK
9eQbklU0sZKhNCXOg0lDFUxdUvtDa9Fq//2gSoURgSiEknu4ixlS8Ovqa7ne/oaRIr7lFAHmNrod
la/VTSlKhieqC/72K1+72QHD9+T1DYEHwT5mOnKNMaFQGqKCgvaR5uyJdL7+894VMnNSs389LO4H
ZUZxGZHJO56ZIGrWjLtJgO2R1nz02OWW6FWWlphdOK9mS5HA4zCrRJ9lRGH3CJe8FPJ1XgBJzFLx
tHLUX9w1M4w8+hdnngC5nA1amtme0J4u0kdkNul3eOTNsrvjZWApE/QjpfvfJX+XhQtbsqIJnJHw
G3j+13z3fKQSlk3DMa/WMG8K5Ljfm68+VU8EY1Gp2dc/m0p5hd7mcTZJp5qW1J+OE8+P2dLXH5Ku
44HuUXHK9biRRLFp1/yaNbilRFgCVSqIw5X+nFNqsLbpysms7qjtzP6ZGWicmtCkyfSyhb24mzTe
AJQuYgC9t5Vu7YiBoz7gdhuzyd7HpDdxZ5tJOIlfbq6m7JvKZDKGmWtEvDJjE/3zv6cPVmZYaxc5
pQmFyxFQ1MGSpxyeLli1/Cx8y+wmIN6hkUc+dWjOP6oZRQg5DDsz8LZCB8u4/0UVmX9zZk5zOj0/
IPA1YL13EbOOrGgM6tNbjPNc/5d1ittQVWTH82lw/ETJXd+2/0JkdcqtaEAw7dTxy25zlwOGu/yQ
MNMkwAuMOPTZVTFtmmPqD2a1jeuplBVKl8/qoO9CuN3T3q9sQ8tu/qWxZCDNcodB0nls23/RUQ9V
yKtfTZe/twPVS7mFAPI+TsaLdRifIyqiFFnePkV0yr1wuc1YhckDVhCnbwTN8LSLofcCEgFZIw0z
EIacD0KGDq7iszkJVZ44ULtHKwZOPDjZ8P9ISS+4F6yn3RdrVrKOC4da0yWP5JoH9zegWhydMeP+
0OtXwPrgMRpCGUJvPPzwpwgKdUpMYHZ9IX6Zk9MguV8IOsqS3nRG27Uv5RNc1nyGpJ4ABDG8lN8t
QWqgzdOvRBTkV4k0cWFvg37hEqEb/KOokUHSH8ELk3ca37B9HW3OFzc3y9hw59ECgDRKUFuyisql
GZ0nD2N0Jh4beIbEVLuTYxKm5j4UDCLJseBX1V2hkaPWE9ynSsfGjMrbweB0etQ0eXXovkNVciuA
6Tac0721K37bUKnka50UTx7KVCfhFqJCdlr9nR3WjEZKlPQ/P0+Y1gap6FjOriEfYU26iAmWmzUF
bAC75kxUyzDWsWr5PJ5B/eBT5J2jiYzTPTp1f25M6UCpeAq2nkE87ZxDog93isA9F5g8E6EMsFqJ
rdUqC2r2fVu6e59BtzK9if7J4AF6qc/LWZjOpBbcxWXgSAs7HkDKAHCP1czj+1WgY5noX84obSOB
RA8uouv79HG+wVhRPspFuy01zQPcr0uYI7dayzJr5qXV8RdKiJwqJwGXcjU5a7AAZHp6pyxR0TJT
4c8/URXyC6fx/KJf7uBq0lkpAStUz8gSukdAepmCt8V4g850JsCctDpQG2DId/2qAC1dGBX/Tcyr
UML7RaO5FyZDgFiQqm/it4i9IoSJhgoWniakLd4ylXQura4kTxMYgUcfGGOnftrb7eQw03HTo0Dm
i62Rk29EnIleVVFlcD+4b21ucztNBBecDJnaReZDLwKbCWpeHnNTR2pOXEQjYS8/6GF4yzYqf+L1
4/9iNIiJOvH+xBCVDWsbFHk4eMSFl42qmVL9i70AsMJk7zVGfJ9qmg1XMK3xcqGtmS778bPRl8vp
WofnXTMpA41pKblS9LbwJ5KGRDvDPQSLMtFqw38NhJjwpzy/Sg9H/9Ys4ZBXxTx5G08va4RX/YSW
baDfUhSX3Dwyxqw4LIKr9uWr/z6GRqCGlqWtHVPC6pvTok3WCA49Ndx82nuyEqSZefEeTBaLPuJx
kGjPdQa/UN1FP+oZId3Txbz5i7viJvU0vAxoLw4C4G+XATEzXwR9/6dzK1Ff05RIgwXfpQhKsU3c
3J0k1kZHyAl+HuXiAjrHKepNhV/BQ8iFwCx8MiVYqCCZSIzCx/imr5Xt+rHdxH9qIPWxg6QwD96I
pHq7iA/VQ63np4lGQS+lAwtg9xZ/+lSY/cBfbWfDGbxKCTM6clSxkccbLPuvTjDibt3b73R4hMAp
+V8XiWqHED0hpPvzYFeWOXfPF0VDS73IWoVASDH4YMdKtgzsVTL5hRCSHz756NFwymOdsu8FU4PA
srd9W17cN5uMe34KnWqn9UotD2YRYvCpJtiu6cD7Ypk/PFCWT0YFxsvPtJ8IxR5rF0CdgxEUn5e/
+dYg2QfWv36QufW8i9g4E5jhTpNs102OVPaLen51f/8NKmMsGaYTG739lRL6aKck57INIiAqmLoz
dwht1xP7koMOJ4tiEuC9XcZ4ur6BiNIDMoYXtnaY3kzXxHjAu9R3AMc7aE1SO+q9RTebaCYkMrtF
DKpGyBqg3Irdu+IOK6tOObNNCv0k7qfzDnJ30GA8LeqnXKO/mJWC58deOolosCsS+OIY8eLjL6UK
647g87B/HRdDyOuy4boiDdU/JhI4a+SzPF7EjQ5LlKyCNUV0rbfRZm7/pMTQ8ka9braRR2bWCXQw
IGAAUK2w0pkbA5xw6LJ1rMo5eNFRphIlDfif8o0VWVfNJ9ouLHGYw1DxMxP761U/5xKtWMgZ8VEc
4qdmYrcCHUZCpQg+KQHoRPNVTymyNpe5Zlb9EbCl1Ef6LFtMg/Z68U2bZmol4kHEbyLvh79AGZw2
w3hvp/rr5zTJ/MwSQDJ0Oq5xgAgr7zXNzXkhUZe/UOBhcCge5T5zUKJGjxeaWCX36A4RmRLZwG4F
/hOagrtXnIFm6YihzYZzd2BNbkCixzfkzUR3lUXIRpAo2otKdGS+M6+aPLFZHcCXPZClMP+lLN6x
svEFOzz0liMOM93KEGFsTGxf3AIuOrv56rdLw7Ei2XOegdF8cm4UeS+iXirWyJOjZLh48Q+HBw7y
meAEF8JbPZOImtW1Drl8J0WRVuw4F2wNflNyWtNp6b50nHkF/X8zlHH9iOMDYGSghjLXoNHPZIar
Q6zj76waEvObl7Vxbc5QJvjpl09iz7iF1pf0M4IJD9dRonNdA4DctvxCCjuppvRkqD1ulXYxpOYX
0Fqxu8ArBNsuWsI9m/wPhvvjk4H+pIxRsDyyaPlHGo78SA5+Zd684lhxC/N97mztQO09rq25kddu
X3yKNGkenw9F+ggaAoLU0MC3UeqWq8qIClPeindBkVWAG5VAlwaKL0KJVq2quYFDP2ERxgOgSGMw
or9OGxT4jx/ZP3ZIBtpvr2weOoG/iNb9VfVPJVFkte5WfSu3x5et+1Qq3QujXANt/y5dl2XP6yza
hakWl13KuAl06JBfIXdLiOXfzS33d8TXUaQjJVQuCIfsKz++CcA3co2j6/ek2Mv0iIg49nxXe1Uh
0X3pUY7JtzHieyIcL3tAlNhiQfCyjHNv4WHF/V4/7rrr8xsxXVF6DItt1vxcIfGbPeu0tZQgidTn
dA80K27zOEWwjk23KVFnJgXhipL5f0p1I65XD96y84FZ78i4REBfIPK3cltb5cw/JRfScb4LgFzP
DqJFuhj3d6EwfWIvgT3OsnrG3fK/rSQ8cqYfw3MNCuQ78bcbOWbJlSdejxzaCb26n4dPYlustjL3
ZCZjEkBYDv6V0gVoVXrKl2rRPZoYKA5KV+S2K8wejEUDXQH1ftGxbGbpXMbG+ya56nLuAVqOwJis
PPo8mHbgIQ2yTCuujshJe3H6P4vbexh4XWucGFgXu7UoJRV9i/zRV05lZqZZMPqMLcFhMSwGdAbN
PtaqUh4JqQBCGUQL0HuHNNFkFoKZPfhYQHl/MbaresMG54gEfapV+CPPZptZDTED1+UvE2b9Av20
VBqB5XFwJIp9q6wwt3xJtgdNiLEH26z07C2NKKVm/N0qub6pmdknbbYptcI+BXeIz6XCTOkui9aU
C08hK9CjLxERjcYNgNkCZSmeEVBW9gjhkx2UJnq2w5JXC6UiRPIdhn8ETUaXzE9xHmrBEA5b4tCw
jelIH1dnjxOXoxBi7trYj6pOtpd27IPoKPzjBkmGMvU88Rk8QIHlIxSVL+Ujw6F5QG8og4jqGDAt
IuULJpJHa3BBZ5bVsJ4rm5HETwmlQ8tU9OctRNKihe+1LlnhJBv6/wKP3s6eVMoYZrBerYjlBgO0
ydE6qzMQ+0SOSFBrGU4P/7M2vaMIQNMxjS0j4cHTSUkfRIUy0ai5HPA+NWJwnAJrwyt92X/TLUBQ
2vhvRqbhSwtlEbDtAWVCLy8rDRGrjdTIEVSrgoVSbgfchl2VraFDcKdKBrwvkKyemG9AcJjJ3WV7
NW70BQOzw/hy9QFNpNMzRBAGcghh148Z05TyVx6GgzziMzwLHN4b6IFf/HXqPj3/oGNYUJuKcP9G
DZuf/uUp9vzDKZzspPF0czmj8EYLj+mUUXkRX8p1f/5VPFomKLKNBe4VtqmFfTi+vve7Vqj6tmA6
y8654jRb0MQ/Cf8/Af62SljWCSxLrplykWlmJdE1rj7qlvMbJg4OsKKzxefvQ33lOKh891JbyaeS
jtEtYfvFA62AUMCbgbupQiTBvBlW+AO/23GYvrNaZLhRAhwl5jEaf0Us7QIFW4V6S95EdbP/PPqa
6ZHPFUJ89ODZkOZBpirKrE1942BP4VaAK4C0Qe/Om0mDUvMxEsgsHlQj2KjCV1MCSXc2JziQnSc5
W+PpNuTbPOyTZQeIKEnxEkJWdzXK+kUFUJZvsjGRI9GOrAP5Vl4hB6uT0HSaBR/Kk/zL/z5Wn+vs
1y9rUr+Ci4RJDJE1cV5PpTSxQEbZhkMJoSJJwUlHnPndG9M11vR4R7ryWAI6wI41Up/JG1MTlUrJ
5p0FmrjwDCj5rahvAI1YlKVlnlrcd4yAnA/B8Y1M731zZpnsj7Ho6B3gPcCjQjsCL67yRUQbqVgu
xZk4d0zRw1+0teXcLDi87P+yOw1iim5mXYKnoCJp4y9ir0rCxGt/AYxhHvAj4ofe9nPDfmBrDEcy
EFstHvu6/cbVhC5K+5aJ/LHp3hy8XP7Nb5Xash1CeGb+33t6UU+EwFIGxVPUF00xQpj6KMVsRVR1
I7vUDIlzsOk3qjPl4L3kJr67PDquzXdXyFxAaU1xbD69LlHxbLTKgI05XA1n6CpioCUUL17dUGPy
pnAuBSUwMpEbAX0c3/HviIgkbb1DcLvET9CFL/5qMw4qSY9ctVO4YhvQfXHRiqDy1BC9T/vP6xcE
n6UbRhZg1NNQoyiYORslTu2hNDEMYTStkj40gd21OCJcXP7PR/pzdAhAFaQ2weP6BlVMVLO88k9n
NySubywCfpoP3+yAiR5wd1PpYjyCsE1VpAKqRBIPsoXPRDol1DTlOzJOwyvtmw9v0xmkaYKew7KC
SaSxXtYcyec6RgpF8cly124iWOLJcXPlVpxIPBxMosKljQJ0t7v5wNyh2evlMHPTI932kW29v0Dv
tKfFTZz1r8YyIP0Vd0ekxeCP1HKWolewdyUmICsZk5rCOcj1tO0Z88L4tfyrH13UzbqI7eWdc38p
8TN6oZqgZg7kbfoTPp+4GHobvORT7AKtpLygHM+psS4IHnp9f2G4p2lxFu/ahoFaFwi8y6Z46cLm
BmFRLNXAu/ySXCBUnzpRC6ePTlzDColpJV6KH5IvorSYaJx2p6Ph1hWXBUzIwMgD+YdIlWHOktn6
csIR39nACrq2bCu55vndDbxbsKzc56krqWuqkIB78Z+mQE918NfpZMP3F4hZxW55SMiWAIMAFOVq
EFcK5Ipx55FqqUPw56ENIRS35M74OIvBKngJZ2QmZqsCyNS9sNns75SY8hShxbEqV8HUPsOwAX8y
+DMRQCoZQCEOSCTBwbHtNpUgcRDaDux4ZW4b1AhEKO8LLlGTLu5PebI3HCBKPnk5mcTMLHayc9D9
aoh5Mew5ubhbJQzCC5XFXTNQW5q99hX6rwXoRtTW2EQ7LvX7xaVhJrHjHXmDkQOA535VY6bA+Kfd
K+maR0fjUDkFUfXIl8eqvFvo+zNF1lihVjsPwGx0MQJ3CMOZd3inaYIXYl5GM1QxeRMUAwVMfBBF
4mndOZnNR4C8JC/HzscEwoQHo/zGzz4EYUgsARstdPcz4yzTw8vJG/6W/LpcyzFYRamKwqUrRQNc
5IqPULCphFyN74qUZk7femLGUiSHWk6weac7dZWQsDA666PvkiWq8ujoJz2z/yw4veLEiSAmNZlh
BXKCvW1gPj+Z2M1rOCKb2Wz46HS64urR8/XhLVqS0M1eW9SZnzuN2CedeHAok7qbhkv4s1/CvYPF
XPeAoC/5nB6m6LV3iWZ2FZ8u3PY1yx8SXVM9sGhAULSKo7B9HqMlj372d2VcxRC7OfmvyTCu8us9
Zi9uEMgewMya4V3r3iQXaLojFXtzxQaXFBb/BFo7CZyVKamTANc/8F8pPJVCBt76K0YlXBpSFWtD
X7U2tpCbQsevGWm5qfdvHmq8k6O/jt7Zl/fZ7yISHC/PLIgPPuUzp6nAsxUHGYkZjghFuGRTatQ6
Mc/IJm7JAtGlAghYoSYjnbo6gIJLxBG8tj4WnCZzVAmDCXnlCQl6jYsEFh7pDWx6aVD3lzvCxvAJ
t8NmBG4UpTY8GBuVpegXbZhn2WIW8/KBv9NF8+yDEFEeCmHh0Aj/llaTFyRn6TpHaMhMvnFjS1d2
0A4bHyitQuADxiT01SjwFLUS22pKz0TRE4bfegKAvCBhIQ8sq7i62sRNIj29O1aYZYGS1KqkTNjO
I+IIFYW0kJNB6sjEPwmwD8hNWcQhr2EwRrKP0qLnB7b0ZObjxH9Ovomg4eLbJ33OozwJkLHSahlN
n9BkmMH7YpzqJiHHKyw9UknWeouCj8MgqGMB0YdOXv/JtfHIimZFFTaVIzcTfP5McNOV1NOmdV89
DfvMefaxvXSVs3NAFjVai3OavFken4cwDBJ6pyEshh4PGCUtIEXtLQtiO+HFKxImlpTWqiEUyXRt
Z2xbp8YzlyfoP6O3Nx3oe0OnDl5gWbxF8y1z/Ex1PkglF444arqdO+ExzLpFJ3I5iR1aLKyyTW78
lza7FZGcIj+3rw+Iku9upFC03F5K/qwYfSE7yFM8eAP0oc/mCzyBMkKBZ1gReU6cSnX1JT+qA+E1
k/XQ3hWVq0asc0Wrw/isBFknAscNqHwfRpkXXaPiKuH9LMKvJflggWlpzsa6uBNcEXgv+vyQ2quM
GvjWYdpQr3KFXojYwqBNNvketMFs5QmqBUelf1465yxD8IxkIrpiHN4b+HzmsEERFW5M77FBdhmB
nfB502moMaO7InZVn85qp6rj2qJ5rwzH3LxtmwQSyk92LHgqQuT/rtU75xHSrognGb60jrUIB9FQ
nr9DowGa56CxbwWKcvOPYZ40M3e3bdfcWJ76QqpcOj/we4CQ1LyMefwuASvq7/cv3mJHfSC5pku1
SH26yFRdOk0qMNh8UFC9fEkSryKw6GiwdHqa0P5NIsBi9Erolm66c7Lq3sqPHRKwU45ECRwC/3ZA
0TnT4DHwww9WG1wq2ebdwuuZYkO+FZdQp9q/bHoZE8JiNgpBW5muSC+R5eHn6uzV+ptS1/ZH8pwC
VSIo/d3y5d2Nt6DnCKh+Crrmt7ccAsOWU2bMqzHcfJQuN2rSoLgr9LqyYUQjYnDMAKHqsX9X910C
uJ/ec72aV2gyvW2GZ+o/+ePe1rnSZyXu6TjHnmoqPBR7UfRWfQsmE3sqWoP62xPHBff/Cf1sfhGQ
nBR2PUoEVZ96/rKxQDIbsI8CdRL/tyfL0/XgquA4wznK/iCsutXCFcIJSL4lZhaKdkn+7EkXlaOE
JcLx9Q/LPzG4f+s1IPDaGIbpWW5orGa5A8JGKpJ9KeXh32ZT3ZUl+Tj93PTdUgdC1mY+RhJEgncI
UlZqGMjjKeOYbt3VRaV53kg3PBCjblFAq2t+ikY94Ra6sJ1fvrlB01SJI9YgG2N81wCl9W83H5TB
xxS/b7yQbY57NQAoVFzQpAl+O0s6LI+2AsUKGwdWOp4LRQiqegu0bXGcFTNcG3IbVwJ6ym9/H5NL
0ipXQjrEnAYHIr9/bC8hKkIOAqg2DGuO2WG9ymGdW8Ud0eyMSlPQiNa/z7VmM7NnSAJjoww9nzMM
i/+YI2yeo64WEVWJ03s7gxkJ7l74pvprBgllxPkGhAh9a7SfUVduJFQivBxQy9FXUvQwS9yOQGMv
Gq2EndD5qibpAMhvMAb1wv/Hr3ZOQLh/L6l5mfgz1gLc3LisF+xJfTD8SEO1cW0j2mFCcVZ1Xzyp
4CHQ4v82E/6N1q5AzuG7kZiwhbJf1OVlQNKSNdBdzfG8/eP+Nkv6ldP961bF5gZ+4VCnfSqXAVPk
QD4mxKImU+cs/+5LX45cSNc9GADmIdOT0Vv8e1yylTefRLwUQwVYKmDSTfs7fSDCpIod8eIyMVXv
bS6CDKCWcND67vN4LYmB1VtQswTJA32Oey9KsuA/Vf+jrv7qIpWWbMbmRvj5jEFNO7dcluDfgO04
LEKnd16/mjbeDNDWEpMszc6pOF+vQLkCPFrrfNnM2brD/3NwMxH3/Y0wXW0Z0YMtE6OZlJR1QXSB
MIs+3xY/ekmtisrqUp4q6dDaUPZW4d0t+ktnYVPNEt10uv7rRLGOaFO+YTbuVcb1YZfxrff1/Pif
sGaJ6KlRiqTSYWDOmzvVfPRpG2NnCxM/ntfB5yacXkzGRe2M4DvKkZyBdIjhgCO90ltS0vkG4Ta2
Zuy4sJtnX56vcZeVRcy8XirUhQ/bRjWQLcCsG05rrGatUHv+/VKFgBMgxxVHkwOPXxkzYlvaUBhg
v3jGgi6EKKTx8oqq+EjOyn3vjS3y+ib/UsCDUl/+6CVeCcqJYXssRFhvcr6Ho1HDQzhcKc6euW6s
Wju0Lci+9w9OOYTCg6MIEIQNE5qpGTS28q9i3LMaTE7mKDdpRpQSRIJ3Y/W0I8IEeWFcDo8KPcD9
ehy+/L+QVgqP+rG44NO4z1/v0svIXyOJecBTCsqEPoPiQOW/QNnnPTU5F1jlbCMIA0LnAwxDpo6d
z+Y5twiBwFkrNeAko+n+dlkpXThfK/AeY2Htm/0GvEqrjPrjZTqxheSSpw3LlJozI7BWX8HZNgxD
T7EfRlmejlaQpwlOdv8gtJsy8uiIpRVq15APSDxbw0KOqejG/v9elmtaEH95zCT+ksocWfNdBve4
BYMeXQba+68aoclU6KZalC5S52P2ZgfbR9YCSYIAVXZtE+NJqlgs+1WmddLWaCXeyTSjxPvcW/uE
xRZ0ynJD75Pc971TLfV9Tq0lxlJXToZE7sQ2AU/Gu+17yMju5JTiRZCkHoBwW3iRaWl3yEemE5Z2
+7b14hiI1Wo8tTmFcsSCtG4f+EUVciHmUh6REP0NkklDXYMpAffmqKQsSkWOzhDobxQc1Go7VoWm
eBbQ+BVa1Xb9Cvxmuu766mgThIoYtgEIYVSMI9tyTbXO+HPH1w+Y9gjnQABVMAeyJy6gM7VkpmCe
del4TWJjFNicEqHZw8I+vuhyGqTbyhdctxVa3u/ysQSRobnERhaHRq5w+O4qwS0kaw8VxWNxVoKF
bKtRl9+u6fgnEby3+TzIbvwUa/ATyIRaFHi4lqaHMhQlbWYJErBJGt+gGUH6I9dbyyd2OzZSkDfY
KmuiHgRkPZukjA0MhFuiE5leScePK8Hozq6CLjOmLn29UQw9ECUk5PFqL7cWDsbONlqfJ33fE13Q
R6Peyxz6LBjpGcGSbwhYwTm4JGVk1ZveNA7Stm7AI/9tbP4wRvjWZn7LfUaHDqZuadfuOW/MI/04
X0N/foX24jhPwqcODRAoQD8lNUyVPqk+FjLwMQDdtWzT0brB7UQp2BRJxm786a/RnIObvDNCFPwl
7Rg1nGMowVAIniruziNC3RXSL++O32XGm1+rCh12Hy7JTlB+v2NynuxM0tfK4DCgPSC9qUksCaLM
LYgszqpk1X2h/BVcgvjZRdph6NCBm6OTSL96geeT/US8Sqk3yhl+xSWWS52MCOTNG9N9WIpJttMl
gmcQNWcv6ZucnLVPp5MAzBJuZgCDO8T4LZ3Y+BbcI0q7hYtSMjujQDgwbp8pGvwYfpvIvpHbM1Y8
I+351jqxem4WkDyUSyw62myTbFQQ7CU0wjJrMrglQSU6XHNDxVXi0MibUifB7T6I7dW4Yug9Yvkr
fbHynaVGRU+k6LDpuEx/dQMO+75cnCc0LiQz/ieOykKmM0BsEPvoqNDL4zQkMa8OmGq7GZgHNOs5
kSwM4x5IKZ6AVpGoIarbi1NL07iyRqtWV5H9RG9c7o4VHf+b+/s3BNIiE0Loo1gkr6+veZMSsFXW
gaaffOsYiq2sTWR4eg8mJmm7mPPxNZmJIUgEW73qyn2iETFDu1ZCkPvCPaMxd+2tsaYuLDTQ15uP
KsaAO+w1i6nt3aB/xsR7mL9P05/gMGUn20T3Cw2AKoTuU32aIqfWgkSSavq2yfu/dCK38GE/xB/D
4E8xmkTdqwXRHC1EMqTRjKGljXLuA2cl7XGmNIUjN8nQKer+XJEcu6Q3HtymtjaoVC8prqgCTQ1m
+h5kvmovdjzw+WGgcY44x94HXMjtGy6n2ZvIJkm7XxYQ0F4E2opkeqxJvecRIVQcJbcNDtsPxcG5
7SJxlNXSmADjtnaraC/vw7l4qSNYu3WcC+w0o7bV9URYhNhWk8rvkH9KR49Ha+4YCreob4fW4oDy
d2UVsZRpN5s+lGnDHtec/H86bdLMzQJfqUtq5awDtx7rr0B50EzAsQl9j58Fs/ZhZ58TMzk9sk/T
zZ11shKPMdreFL1UIo8WjfiaLFzQnxhbQf9oqGct+4A2GBw3gzGXUCSk4m2rxqGBfoCEO7HLto60
c7jKFZ6VqIVX2C6uVch62DK/y11Z17BCX+VIkKBAqKIcWPqudz/e+A8jcd8VR9QPa/xMUfSAqdDE
VD8C+XNMU/sb4MtCnU8sdn0ZX6F9ZF46nhtH+FU1pzkDzAWvR0Fu1MkdUi7gX3BwvxrjRDPwLlD/
HzeTxmovsJXnZkip2ndrdcbce8laDKqld8w5IiYR53nOWIPOw2jGaOyZFsbHgOst69fJmxbSthrD
dRNx5UqFD69Iv6cPQwHKrJGrz3sq9TYAMpfu4fMjB/BZEhhXoqAgl1RK8jzqFfkX65JzU3pU61m9
P2W6wSmCyi9naswFRroQchxdcqUdXsNX5cOK53IAVT+ZlDaQK3T2SlFf7mgCFz+p1C8xK7Hzi5A/
BJiQkEEkBflrCmrPDRvmaP11LAq8xKTty8c6P9qgxO494g9X76nAGRwuXGkR58CIxt1IxjgeMqq8
+UnRzYmLsbxglmJ88HtoypmNz18qs3i4hQSDmpLCF5P/Hb2IZc3gpOf3SV+Q4tdOJo6uIEftnhTi
qthrMjAhMRg2dBFgZCq2Dc46KRlh1D37DJyw4BRsI8tn8EVpUMnAuGXNqduPjsO41+ZROyJ8ACjW
LAtgUBeitRJjfgRMVWHSn60XbZYfp05GRbqPQJR+Aq3KqxCoEaaESzGPORsU5/aaQxgz67hWS1lI
asWz1bqlf2eXrxdtNf9DnIVcFHI+MJgeYqbZXRHPsZVxjLvid4aznaYN1VRWsUflcq2jTQ8FPrki
0lftDQowSKxSxgYzJp84X0P9dCbAXQFsjlA3vbI6aXk7rBebuYsaGVbDOt0AOlwM9wVXhwZo2goK
bLfNtO2S1T8IB2VlWujo0F0uAbZvLtkUDDwNpQIJSIlf0AIfRq4Kc34h+lFvOmUaE9rDeXZAPzWm
aapeNUaF+169AtW1/k+mrQQUGXI6uZT24f4/CP+vq5Kb18se+rHJOxuuwv++30yuDkJ+m06f9NTg
V/g2Dl2I2yKhY8Yxozn/rDyxDCU1uoewZlstpQzxT/HqUdf0DJPOe/QuxyPN8uE++45QRZegGmZB
LnisY5vkv18VqpBtxtv3QM6vhB5fLM34yO1pvqGk33KLOc8KG0KGgkOoqj8tkC5ViN1QPwDnuIY4
i3DZupm2SzlZQBUynIOftOHazUp7vOC5/BiKddDbauVvCJE2yMPvJjsf6JUJ9A6bu8sprv+zTArC
Ya1KvbRZBwJUgumvnkz34wD0tSTSX2V1k1hnedKn59ilOGfqCKrSVBOx/KcLGiQbymwPTs+mcdMi
XtMFgpDvW3yVc0r53VKQu4stppHUJs9IFjhrGvferO6ZSWkHuQ/Ab8dwRAL8QRYUyBKKSgOVtP7Q
1G2FQg9NDHaWOz8+NniIp3vot4ThFRJ3gGH1DubcXFgSauStQ9UKC58QwwRtTeZvJc/gIX17K+ZI
rgIE8VouTZCQQHDQtbRkjfVia5hTzK7yG2VaJQimFmj7xg5NtIc5niU5ea90b+v6+0JW0mbj3zES
Xh5EojKFgb2tXD99OnhDAxZinbnc7wMiG83GSRxUfa4AaKe9Pbn6hq6/zDsbiHYbIp4HvfP2Fvrd
kekMK2gO5swkUALmKVtOgzd+X5K0yMpHHmArHA5zw4iKF2qj+/LFCrhMP4TmNRtnQKGHugqWvATY
3bJ29yThm3+ydXKNR5AZgyVhBMMuwDrh5hCfbVX+iFy3FPOKELFmW7aGqqamRwFUcBy6AluVVUdD
cETkYAuFyPhD26hcc9hDBBh+mmaE3OOg9yw6V+iBssWW/tqjcPocQryKZ3WkKsQq7HSDKfXIFLr5
zi1tpwSdcrzH7uAwvG9k6hIwYDiI2bb4h1acAC28TwnCpLq1uSHh4wk3BgNVdGwQX5JSt2x6K4Pj
vmtr2BtT8d+g5hqo/EDvpD8FcAZTOtQrDI/eKwAQWJX++b5OBY/4E1euQ4YJgJmyXB5dHckdryOK
8hgCTN7dkSObr+uiQ+V/aj1A7jz+uOVyS6C6vlfqbHDWmZBIiSyjF7vYT0659K0eI4+EzHZJ+0eK
KGJWJeyQBmKf4K9gfz44MszDB2LSxRH/OfnDZLf0cWA4Bp2FC93Uxcfp+QitQgUtzH7RsqS4m6Jl
r9K/kTuonPB2LdKwqLmL2kDsa5CMj1XQOU9/75qae7Xx73Xd92BdprFrxWCxe5uRswudtUITeUFA
v9wolsPESmOZG0On/lwwq6o7eNN3zxy2nyk/vyQso6C774I1T57XBdXCvyMTsv7nzxXY0858qr7r
deCE6XXUbnwZ/a4G6B0DReIKgf0fTpxnWfKHjIOBO+hn8vf/tofGBIapvdYWG/KBPgnIG6Dl4NCP
JcbDItVkD1ibOBf8Gt6iibKAlDq94chrFP5V1lZM1QVtPiQ1KEV8YlnwgfBPFfAAYWjbFI8SK8c5
EZc9UeNp8BG/iCZ9JN1gEz1IGcRKSAZBNEYPo86u7DWLEUOm0dDwb31VB3K1RH0Maz/xwHxu8byv
A5qjq8QM1xGCR1YtNi23zhflWCivi7H01hqkHZYCY10OyI0YV5ZfUHrfo5biRAm1lPwP1WUMba1x
msoz5yWxo5JmaV2olASM0ixwRbSenpC0Gyu8K8RqIIGWH2JsfRkdrq4jvXuAZbmqO04XTWkQCjUT
NwGC0cC9sQGrOE/tSswWc81szZo7daD8JUuOT8BKG/6V0HsxS6LE7M20TMhe2P30OqUqVTHzDqfl
xL7S/XKYKRaGfwl46712qoC2tOIUYY62SV1TuHn2xwSso6Qv8vNZTZIa63PzqqFJ2jhwDN/5M+Bg
GB5W+RhG/7IIJ4bNnnzKVfF9XBV92CWXBBXBMIpqPgruJ/anJtrbXbjFUMyaldisM5F3Vnz+KIrf
848DiNJ8xK9kYCfMXCVzZvnsOH0fVItbV+tjA8vD/iUIHbPswAujdabLzoga8AV/BYHU7iK/lpel
WPDNdvxCzR2b46oOx7bKq5EE4zdBhxPPhWtHmV0SxHLrOWYYEqRNwMyXs6TQfYucrsalqrc0vd5B
4+gQHAsZO33TkOpNF0FvMCp8ZHkzzXsoCMatWMeYPD+XP7w1WRwDa4AR3DZ+rI5wy2feeZSQ7JuU
Q+Q5xyULfa+wJrYBTvkkHylOfoFCUiSLsglkuO47PFsLlt8DwqvpkFHnBE3eYIDHuvmiAe4988UN
l6JIq/B/YeqFpqxkEOTk5c87IsZUZIDTaMcm4tJ7oO16F63Ck1ZYOjRoyHYmdrNueXI3gnXlTe6p
Jvx2zj0MygGRVzc2SzLLb/59pTY9CVtkWpaz5E10CtDX8gYKsT8R5oaYmT18Vv0Oxjao2Sj+7lGO
UhTSdDmYODBK4SooG0QAN1UYEjtI0GumWZjG3sp1SCnKmYuiK10Q9bFWcZBqjbTUQtp5jueyk82q
wRoG35pdL1hhGfOnHdrhheUpg+4GWJWXNrDNh8UDI+FptrRCMDKD3GkrPvmLDQILvLmCOjBf7lP4
W7k2Hd3jlq3JH7SEpL72LF2M+7c7Z/I+b2kuFpCatof8BVQCY+jJJcpmNlkBd3UN0JV7awSCAUqj
P1PFI2iP55X81GtSANVqGFYVUgJuZO+6aGh8VdBPr50GHbH6fu7zjmsQiWq7t1xT0wSCWLudILUo
tv6X3zBgALXrNX/o5+sPd2e4kaeX/nst00Gq7p+wCwI1sqKND13+fY67Ip76vDH9F3gYNw81wJon
HGkVyvk+/IwDb+1Xdwojt0Tivn0J3LQZUi32eUxe5tCiodCwIHYPJsge1A6NlXiZ6LvWeviIbGGp
UOFXI4g+DsAVTlzUrq/nWkA9MUFguk7dloZLfiVayHpXFHBswjK+24C3HnLB43mSeyaGBXrt6CnD
9uHK+Td7RdT8g9RIrr6SoqkNLoyU/IF9L0MaUPNAeM7G453vg2mvPKn5+ScbDef1numPGRHS+Cim
M/PYc6YK7tKcoKm/pGGCIJVDQa/mhdKFY/b1kRRPlm0KcaK7iZYoNcL2m5syVuz78IzBEP/eU7Bw
Hkk18aKEZWocNiDTCUtx6iiQdinfO102Ud0pT83g0uHvACAVHY7vLxBkWkdO+FLJVTMIApkxABx8
PvbtvpxyfdaQiFDV3pkXzEo5gWWh//u5nY+ay/gzrWJJ+xZ1lMkAlJDoZM8j0svIK8zveB7YXl4R
yWglL93aBy5PS+QRjKRoSWQ5kqhS7Sr+ftbTw+JLqOUNx89P3tFeZm3DE0y8nOjE5yPkcqN1/rvW
F0Vylpsy2pZ++9eqqDo/hK32lO1i+oaLJuj7MEW0kYJsNZrugj3nw21DZxTINKeDHd3FEcYY1QQc
NMLDbZIIiAi/GrM5BDrVzPooUY2ape1MGBaBGvqbHZJLX/GRMR3I+iNIv1SN9GSTlZ2VZMpcRsMk
fDu9gqZf96dud2zAsN3bkbCDRKqj0J9KVGd1ziXEaQ7qJxcFQJYCngXMxnYEmKLcJsJdttvgpLeX
WR1023n3wmtnfWmibpF2wqwnfIevksaHQMz2Rm7ZcRHO9r3+8UIbs/FD+M+NmmZ51zq2kq2F5iru
nX2faPAyWISby9ubHdGmMvszeshV1Vav1M5ACW7tJ9kavJ48WCHBBgaZgMRPCsGkoyOP+Y/9tEZX
QBAKT8rH42EiLziXFQJDtaFxtpMpdLjOekjT4mnqkB22GAn8+2lujdDfOba6ZoHYCwNV8DiJyIBx
UgUov7FQnA5/TC+0ruOPG76a2tKlbFsj/J0K3mCGA+iKinjmkFNIEmhv64UGbLrJc6SgXLVS+/83
rTjGC+FSUV6ovn+RjMyUJ3qxDgSvRtVyzQmUhv415ZGUiAjNMaf6+IrwEj34HcfYE3S59W/SjMo+
TsYBlLyxhdLilFJufBfuQwimqAfU4tmc2LM8sUvrpZwKxlALCND9wzJfh4OtJmUuz6s97HR4hTD9
B3Il1fKXqIsRyyMypEOKD1MHBtH6rIZCSwx87D8QnQqs2DELMaoQc/x4dQtScy9E4v+bRu7M79tM
X97RezL/LE0zZg1w3qFy8sdpTNl7E5Ht4Jz9F1HF+HCKqw43/fSs9m8zjZBakcnxx9Lhrmbasi0f
aNXqv4PHNuGrRokGjn0AYi8OEzAMOwXB/wlDrIzXlJUlfPIHbNTpuOVbLpDX7i7OvFjaDuHqRf2e
7cGrsx+nzAZnmQPFIHWP6eEfid6YacOkAqTFTI07Mg4yTJF2GIUq95S4CvUM9Fss6v9d3vg18gUp
vnZtnDjRzUoez6MGUDvze9bw6rBO3xnNCA0p3cHMhR45pyQ53o4/mpO/Ckx8THOIpDmFwziwaQpq
em8/L0epI6DdM5OrTGf/33kP2tN1ysXenbnolecoudAi9IJ8g+TCg0M1rUYQ9K/LFY5UjCfr1V3J
U1JZKcziZv2mkFlLvS0idqa3AWw+Puz9xx3Qe9KAhhJtEkf3m3I8Y18ezeSaWB1wqLOEBWQ+xwKF
NzFWst/KxcW+nloikTybypAZUi+eS5cNkEELU7R03Fwup2pyb/b+rIJ100oxSWMFEXaX6Z7OAtXZ
+bPyyaLjIrc5FCxLotvoePSbiwR4im8c0pfEONZeOVWTd+0QLFD7qWSDznez9yvnbaR7l6V5Ucls
vmN7cDC7xg3mILs3YiXuVKkBrOKygY1TGYyrW312doWB77HHTOSkNBdaWwN04zT9Q1ZFsi9v4yD/
TaGjQ1HsYXqWMVKTJtgfaim0mESNOQXgDa9dQX7RvpLeo3cPod/+qsaJGi31QtdLNu2em1Mfxs91
miy0tSs+NKRFVNx6dMR3U9Nvg/A4qcFqMWQKn5XG+f8EuPq5ulJmaE/IVUgXd/3Ix9DRM0xrsqx4
+wW8QnvsuoNBfF/8DWmDf1z7/5cOnNFN44D5jnPI812w/M48ajVsbYfMZbyl52rHVcfWFKCOf+yf
mmyRWGN8O5snjp3h5B6SgEpNLosoc305pznw2W6ZyJu7FMb+7qCvfmEgF/i42P7HUGl8gcUI5+pB
TxlXoBX3NaepSiWl/tXGOywRB35LuEihmn39GqhYsjRKU8z3R++fysHGPX38AcX0B2QN62qjjNGX
TnWFsz57usH8HMJ4oLidMghCejJy2dQTv5uo5nOJGgFmiGngRBt9oAMMu0nqDjHS3/WIvxdYhHXc
UDPgAAzgH5N6yjpj9QxJ7ZlEJ2BiQoLN1dJH5+BjEkHmzgfst+j5N/6GweiUlOjcX8YlVxuS5niy
Y16enVcr7qEAcQocFsfduHcYnp0OGYjPEevf+H0AryH9j69uLQx2U9++C7duDCoMYXqbqWU0hU2K
4B+u1BGcQGkvnJAq76OKlUUzgs4GN2RGNiWthOKg5NL1VanYkVWvH1A2agwESg9vnFaWd+BcQwXh
wywvl+mmzCIH47O04r1FLJ413riQWsJjeUzujVkdSHqny9QH17fP2j6AKxDWuAajscum8ILdww9+
iXqm1LIUaCrSyamXxnSSRl0+VeZm3qgRlEsIX/kOZg82YEeZ8Y4GW+mlFJVBJyIRuAwtuETlnuMF
r015h0rfcxlzqndy9ADWdKeBX4VGOZTrrttSOF1ul1rrHbFcbD83OI4dc0EJmtLxlRWdCCaVIesM
V/PxJ/bqml3lMrU+P4kndpRiyhxcku7HcczQ/5EP5v6U2vByn2dWKzm8j6VxTwR+kb5k961zjWkr
xmWz5+4R0sCrP3hjyIzy3xyC97noo1I48dMj3uzuPdkNr+KLs3OBqvNsLbpxMioV80+gAEnwcNV1
Ps0Q+ONXDHVF6ON5Sq+1anI9dXg8UNFnZOHv3aXftt7C/X0hX2v1nBwMkE9WUsGFw0PAXtn3vga0
3fUWDPN4N1f2w69c4qYUMG/mKQhrEz/gUFIHuoaV+6RyC++znT/DZ3fs8VpAlIpj7XqCmKRELzNM
ovrdAXBugpLeerRykp98CbOZdXp3Ft1sbBA+C/Re0nCfAbPSuJROifL85lP2zWeqIUkMiBDcKJB9
MgpNs8EfFN1fUXQhTw13twLLuKwG6/n7tyfSUMrDZq2m2z2YX/Jwu7nHbsy/A6s5oxjGyTazcE8B
uljsjncuq5bLpwbPOQHxNpz1FrFytJIQyzP/30JlM9SnVDDwoiogXVxkYaDDryJU8KsRijBzQ3qe
2WlJ66/TMIFuL+iHPD0QxYo1sOZPo8occxofMONoQ+bWJmyFlC1eF6yXADXit+lzv+5BayK1UXa8
33keYsnbiOxBnagz5uHztEmrH9BappmHQIA+YBWDEX0ZCc0Y5HKzZnFhhPKnA5iRxplD/A4RbJt8
EtrqQDU7CWwRHnS5ilF6N/WWC1db6pYdIOmijYN4W1n709ktoP+2138ZQupxxjPnxwY4UUxTmxIo
y76jm6GxvC/HC5oKq8z9/NNtqcjvDG3zw8EReKzqx2AdiOqV4nv32D36QW9O4Afs0SoNrTcZo/55
CpEijj2wjqNo5SbmtxKPhfchfCVaHVgFTGXmOev2mXLvKu0IM6/xGyzk5kGlHrKMlyj7/n/t/7Em
GyIdsFlFwDI2qTIfMxoMMtWpnj7rbz3Y/PdWuuR8CTAieFlo198eSIo3i+97NUK/brehxwuzCG+z
S1nIYvO8xlo4xYHiE6xEFZLHN3cZaW/Qc/6rwUygXsAgKpL2HO5liPGALDfBxRfWVfQqiIkw/CvJ
IKJ2izuukxVWOUkvWT0TwTyPzRGpnMbVyf1drwgqqZf5+cg3hwhi0+JZnM78bSyZT93PF5xl9vyR
k9h2j4CjI+zN6vQid1L8YcWhfXVAseuoDjAnumlKJ84cQza22vmo+kcwdq6nlmxCfLEXWMghL9r5
l416yi4hhYQxmfqfrBULFPG1f6yZHxz4LkSof/ULrZhSsQ93bobcDoxj5fNJuWOyHwDTk4jkdtUO
4vHg0nSlIPX0VwZ6KPLIjacnlpdWsMbU/Nl8ZBAzeLp3o6itT8e7N15iJSU1JzWhK2YhWuEm3GG6
E68TOgO4X2l+35DloI076yc3835xb6kYFCTVsPa7RVJboRkrfZqEkDzzUIYnV+pJaNgOTwf3jU/s
rJPpLE1kR1IQKlnwZXa/L6y/uvwsyNrAfI2CcMYyMsN4CdXxixOT2I9BYYoZsFAAN3GLgJ13nzfc
g7Ra8k7jNsmEKwU0MseG0lW5jnfdrB0MMI+gaiDreOGvBj17wIX78bCHBiHR7SLi/uzGkkIRykcn
g8H8e9Vkv8XuR4JNVstFLy7+azHQlpcImqvCRDYf7dnyOSS19j3Vd1s+Wj62kmn33alm0QuDx2Rq
5NYkonv7Jy8/1MQo72nEpzbTeImIfM+ns33Xvi/O+alUp0WUYLEZOHU/nsrDKN6Zby6EmqXQo0fM
cfxzPtvWtDw3uo47Rk5ctW6mWdoaSIWZX71lO/l4vapMwKD7bP4G38bU62Llj6LzcT+9SWW6lyHS
3KFi4a4xVuxBL3bxAg9Quc0nPGlMYj7Xbn7LvUCuIJbBcTrPGbKBuPyFAFIa2aAc1k18cTJidd1L
RMsovCEkJbFwDGEMjkTez01UKSmJGn6bs40gTk/AUnaPiabcSW/tJOJjVJXBWB56On9Hjqcbo6p3
y+EttKrxXqY1DnR11Dece1cstGePQlVxct5ro805xELeQp3WGJpb/OkMvQHHA0sJIsfcC6WmpDQY
8IpO8azAcTRXE2HCgEKtPfYwDt7sXV1l1HQojgMH6cEvnOk3uRvKufnGmBMu+oIv3WnDkggq/4vL
8mW0cL7nORQEnJULDfXw3ElTlyAq/N9apWYxqm79PmGUYcg9TbfjvAhzJnXmLObKQMU/FNZOEeek
szBe5HW4T+iVr3Slra0GQnOhlBc4duMQfd4qGtCCn5vQwJWh7I0mdJP1o/RomDkeYCPsvh5e74AK
yw1l9KEkUQirlZMWFcQY4AyJV7b2SJ200ASU7w3LTRiVg1Td2FZMP5pviW4DpX1IiLdL/Q00EY/g
NUZsOg9DepmZnDoj1JIxDIGLxg7QCrX+4/PAUOpHk/nEcjBvwXUOF2m4pAd15r/aOYNe2DqOkuiR
tIeNglXdyMc3VFyxm9Wgk76wMJsth5BrYWMxndajl9/2hrbezSHvAOAfDqP9SF4EMzxqZKMfuyKU
mfrvAvvxMQBLT5gEkyxGv5e8kOnl0MBOkWh9p0ys9Swdmsd/X/mKPu6A6l0gpbEO2Z1H3tSOQDZG
m5Ugl0ovJm+glmd5WllhSuIDRX70rWOKoA8VuLG7YZRcXlX0SbjZepoCLU4sdSl6Ui/njmsAk6Sf
FWAqjCwhj+r554WS6DDJuYr76yqtVuULNIYIt65x9uX03y1AiEGuJ27qehFT5iiQ4NA8FN+HQ7ZS
17k5B9mooZZbsO4VmVPKlyPVe3KJ22L1X0n6rMFtbrvEPfItHrYgJ/eARbxafoJbDMYsTeLGnG0d
VL1PPB93dKPyx+G0bdXPZriFk+3Jq2on5ZXJBZB0XVVs5GM35gXRXkJVtaV2PVRfhLwEKnnYN6Hl
h35ehNfLbYPCO4v051pVDbcKetB0nzlfJLUvgyFbMZusL1edYlPk1Ey+nxzxSrFmOXuG6Eh9hP57
2rZNoX2qeP5B9k3sKmRZkhfPrHQSVlZZ9I+V93/JnA/d95I9obwOG0dINOI0zE3auUAYoGEOWQ9+
NOILVuF+5labGDOGveV2rWXTH2l7rroimO1ZFcy2UzSnTCrzWoN/p8WQghZE1nF0/YpAJ8aEAguM
m5/Agr4r3LyuhWmKjiS5D7PhnwC7+YCRmk+1T4QgDrmL5CTBh4aqAugiURc15xDL81nujtQmye+x
2Z4A3dH8EF5UuTFISEaWe9iAY5tlZTE8jSmRSAWSwQhQczwQuY4Be5p2vO3YXsX2lZ4SRIInMIsC
HVaCH5BhHtNFerrl4x8TrLUX2k/khy8SRzGucK5NXU7oKIHVk6sUj/DFtw/rRNXafPRFgQ1wyM/C
mM1mJc1svQVipc2llGOl99kkIhxCvff9u1ucxj+tNlbyE9Ufk8yRuyFzMqbKXvAvKUJG39BEeagw
Jzy2CyA0HR7fDMpWYLszvBPq2T9OXjbVkRl6W24KSj08dL3Ofnc/EEcybdboU85F9qFvrVL7WNHw
wekZNo58iTbVrPBuPFKIaJRgya+JEN8L3YDn+ws29Dunv19hYyW+gN6GbDh1Wq7W1tX+3o4u0qZ0
edUFr2Ho/4Y8lg4BLowqrbt/dvl8ZVu/PJ1DhjtUf9SWmUg8I9R77AGUQUfwTYvV6yuZiwAmJwyO
n/vp7agky6MGRbDdwGGQo6jLFsvBw0i2ex08Rttu0ZQeIwba0805V7e3E9/ZxQcxv62+0TefPBx4
Bi4QoDenPOdiBlsEA4iIXyynwX3NQr19tCrOQmSvVstUituyrIom+st+gqSWJCV/Hj5WqtxKy1SY
q3eIpJMQqcxh4A9Pspk/1fv09XEKEnY40Jj01LnXAcZGYBVlarzjFA7wo5S6HP/+PDpe+UvHF6le
xNE4YHDlWfuINuO3xrtYUIJQKhRtyP9Zm6BM6M+e3yJ+0HRdtX/7w3FYMOmsoKeassafsIH8aWrw
qEvNQhtEErvl4VEMB78DQlbZ+VIE0YY/kPaIQTWTkCAs7Qkelmysju4/69zW2sW2TtmEcYFVceTl
oqt5KCt39QvYfjoMHiSIIs9bc4JdDomPHJj9yJoVjSBnrhO3TvnGj8VuKP9DJ1Y5wApKWd1BlqY+
lfDZKXr4cw7HUgPXHq3k/FZcPqbxGbMakQPWF7Ko74sEWlpjpPBaYmo+04gTGnnS/yWbtx0QT7hN
H7NxChu411qus5YxfYF8jyTsiNZGGnk4JPpCjN+aBe+TkfxP6bh9TbpmJ1LsBpqfTs+RPBDx28dk
r6Z8dtMyIS/9NUKBBz82h+UJIQQJGWig0OK3q9WwxlVYW7VGNVnhsc9D/9pkxW6YogD3SEnsqvTd
HhdXu46hqL+XbKqEWNgPcLUGJfTxbPqkDhit2IMaWyqqnJ/jYx0S3m1Neiwf2yTG3W29PF9tKSZg
IQp8DUXvOklxVt8LQ579WcDE9cFhA9jS0/yZ77TxyUBJ6XmCHAQpfaw2orN4pktscz9/Qcz3PgPd
VTou2Ix6vCoHrXlWlCTUgptU2q39FeEngRu0w1GxCNrctaVUpMABbe8zlnXdl0TnlsU17jv55gAE
lXIR6aiIoqeWGQuMOyM+m6LFTp7lPyl7v1RsUUcKRnrtTbNh5QCfdBI0xALwR+TNL5/ULbKHZ/r0
CZLvFQau8uFK3nGPJK5JN/EGsE+yXJ5qiJHHgzIL86YJvzn5XX8lCpUKiABQ8U+9sJ6kzDpzifJI
5yeIosZqJ2CNFpJmdg7HuA0mtUvFsz3p9/x4QXW/dRZAp6JnEI9j1dQ05XJZHc+ESCMpxl7Nbc3b
3HlYpXzQIKM/F2okvGW7nbIhN/0LiuQacujsoqyhkxMhJ7R6y/E+XG6k3tzQgFnA4U5ZI/7DgyeD
4xd7NJYy0Agu+uIss2K0wIoouxmsDGYJN7pbOgkhDGF2aHzQT7p0vyEeQ7Wo6Biw7jkA3UFhfLdq
B60xRQvsG0CmIGEPeRxggvD41zJCBDEplxtUY8H742l/Tj35J7yRiUzFc/y/e2V/87xBtquaA35g
oPo31/4lUzb0S5oQ0ypP0wUJQETgL0EQ6WXoJDp6ESznFmIdn+Hgs7ai6LNmslYUuX5IcIW8Nf8k
F6vqFrM7jCTBh2pZ8F0RNsUQLEVmIoCkSOofrZxacbA0nahNNkKttDsPRpbH/kVpckUVAw4Et+5p
YCnXU6iAr3vVWx5HXW/ERy8t+gksYgkhIYPKQQrE7wA9zPqua5jlf2E6OPHxNJ9mA6d4iuWWV2xT
zPgF7fJOCnurRH5Yw13Bf5i6PSGqPw/u7FYXWf5URGoqCt2Qk/0V6J4FkmMbUORVZPfon3l0ZEET
4P08A5KBQsB1j4FI5hPuF9GTUVtTTj/B6SUi25eZPgGnpalU4ev8BQKvEhguCy29xEtdQr2erjl0
n8qHnVfvgqlVMVBrSIL/vDdlxOLrYCyyIkx1xeCZ5hmD6KT9w+gsKMTnEAlYJDtOFBtC+coBuaC7
yihq6UYvsaR1IIPbhVrB60dFLbkWRxPAbC7Ja3QBxRW1hSbD3EXPRJcXfGsLaU0iO1XkoceDmOP1
Cp8NkUM4dkqLZrSfYoF63Rae0c/96Ge/QDjMgr6rO2Fm5h3DU8GVBU638zLYI9zhpgbP8tQ+f0xO
DwNfKYj+wIfHDHMFuukVHGkl09LN/joMCj4IPG2SDf7dXldzHRCsBVtbhwUw7x34UQ3CiOvCqJb6
uOjuid3B6aay+bGg2t6t2WEsRDIMjWJ5HWEq/tVFyFEYhpWVaIAqxJUBAHlW6D4xQ3+v6CqnsqXz
FoNlgMbZY+97mlwcyqf+2rY5rKxAoW26WoGav9KcqkFfZpsYQ4NA6eZhdXN2ktnZsVa2gROEXEAh
Znw6D4DnBZxe7OgTsLeHeDk5RLC8IMgE5T9nXfX+inoWyvb57ei40A2d8mu2uzN+K3C1IqfbOUMq
tHV7R2AjpNUyTgaGz5q1/A84VwRBcfvv0DZnteCyQaudqHahLk5YADdObV40bW0V2hS3uAAZCnZo
iE4/5rJa11ZQ6x48UBGf4VfjoHd+/PwZunYmdndyTP/MSTc33r4DKT5T80HS6AihIZxbOJ+UBOYy
o97eLLLz2PexdCj/hRjTElG5PVnZmKulI5O7mmi0egqkBxrsUUj5PE9gWTg1PnxwVHT5l79BVZKS
Yit+vHaviQcPigcDK9cRxbNZFXNSFVKBRw1p8wg0ht6dL0MrI6HSJZF2nogXUfjIsvzbnvVVaHb9
m9QX3iOygr9PCA/SSunFSE1fLZMYKcob/3oNtDREFXt+il3dAJdqYVtY13V0ip/ANUyuAX5p/v8M
sE5gVzKdqU0Pj9BJ8XYYH6m439RO+XALqyLV39/0HVHDcb216sVHHSDH4brz9J+CQzAioqb2s+Ba
bCCW6laSGGdBs3ytDtYkZ+CZqcAhDY43Rmb6w3XkigC1+Vu7lc29/ZpZFx7kjgVzOlc50hCOQh8A
QY3fPOY2pr69OD18mUU9imu36R3G4TMlkbWic6DYZFrpjAeesuYMli/vHggDrJcZcdJAOOrP/GkL
OT5ZBZEF5GVXrTNQXpPj/ooLudHWzOc7SEt1GkGT5Vz+ir5XLppNDKQiyXGf0DnLoqalhySIvuuR
tW76Zyg1BVlTk2YfTqjzUHOg2+6C8oxDd9w07OJh7w0uQu2bP6LxHwfat5qrJtMaSNWELhijaH9e
SE3ZkTHpEl8XamBsn5FLysRbwMs8u9becEY8CBusPms/hqn/Q4vbejZEpjtNN9SiAB3imMo85QwQ
iWahXWTFttzGihbupH8fZ6K2/P5nQ8kyLf+q9fM+vqScRG+GHzUt6ub7+Axi98P/6V4MjoJdQLl8
i17e5K+tAk6jdWRv349F0g9Ctk1hob61g3xcyzQDaHtANh+5FXbeyVALhni6UmktU80REbWYe3nt
NiNrBbBxU8dC41+ij9wMixG6XLpEH+4C0WFX81JnUV0m7hpEEjNtRBCaA9pkKyjuZgWYKvJ6IZh5
uYc1YSH9Xn5zBecqAB6FqzJLZ7mKbXWgkJk5Bm1hrWMYNSc+uhlfEIBHQWNms4iBnUMVOMCICeZ5
V2r+aM5G39YLUFgmnZOp5acNnuOek3SQRkdI169PyoE9Qq1XYn9b9WOTuFJe1+42iLR5hxmXxh80
oz+HiRqFV0GqGUQwEAEOcy3DHt5ix8Hlz94kR7X5YpYqfpLWQJEc3z3FwqgF4FEUbLAuNhumbwBJ
LzQ7CvnZUDFEXUPv1N+kXhKUjPmaNxpqnm4rRcgmCcCNqV47jszB9uSEveDCkUIEwNVTSbuZzjJ4
fd5435VdL5y0iLBnQdtHpq1zGHvSr59qX06JqKhgW1deirhv8vchyTpRiy2CqcqLVoM8BnXXl7Au
g9dssXtmjbSrqaKTHYMFuaLfy9fHn1e8eDtacmKz9u6LnghxUwmXbIIGBIDo9zrR4DgVA6yxnTjg
k2cAxHLzaUyVQoGNy+mcJ+T/qDGwIEZBtD+CdhZ+4BEgqB4b7mWD0D0rI0/wSgBZlXTxug+gLWSI
zRR0rK6oYZSXjfaCYKDMEd5RIp0q8+TNCjPgF/YkrRXYVQOffS7qf5jtq/m4BpVdOPvojCrwdAvk
C+YL5j3b398JU5PnALsJGNvkMqNjDB0viuSsz3VZT3JcLYNCZETMdCNhyGh3A1aJixFcY6th12dx
HVz0A2ESM86kTa1WOXO1rSMF686H0lvhIp1STgN3dtdNC2C6VGJ8XJBQNIcbSojAr2NUSyvFA+ZU
3CWxPi/95UR0diTQUPQOifQBavuYuJvNnIWkr6nTqRUgNkBzKJc5iecnds7qAxP9z2OLQdmiLmUK
5pmijHQ5Cv2R+UUlU6kQPqgUXSn1DvIjWv4Zp9gCdHsnzRqjhGrD/J61U7lUOlgJJ77/i9BnK3Vl
EI6Hnzr7jjNW1ut60rbP1pFWW0zCzku8jVgFD7jbX0BJj5YC7GS/5ogSERRuA4nHykCF61JaWIQk
6JqMXOeCTEafl7rJREvShyE8MLxxuNyTfx6wCN4kF5lCBpJ+uex0C77T19rMVneht/45Yyci9Cg1
gEsccY4e/C1BRwCt+uNJzklxB7DHSEGhuTI2SXeDbDzOBat599W3Zpr8NjoUljnLhoFjXTJjZ1aA
91kxR5lKmkuJqsfyMox7fSEv99oc56v999FbPQbtAvimbWVc6+QgUYyfxSHr/zTw349/LSQz4nWX
O0Cbf3BDJRrI8jJBiFhcUjB7YHeUP9MbHtLWn1G7Hh0ukyZynposDKfgKxa2zt5kGc35f2lwJ26u
QmLYXqccO1W+vcZzLaOWFofZMURd0UubWQfnf/nTQd9je0o859tLXOV5tGMb0ocXbFUgPdv8ecBJ
JuCspZc6iIWZ2A1UwqpCZ6sDi06t8kiPj1/v6BWUJ0xbwmqtgdCTz0VYe2qaZNa8yj1izpT5Xflx
63SBjLmrO7J2nEMPU+13CoQXFAAQHkryOzGfpxQ5rkm1QZ2vx2hLarTtzNved1XwWDRIgFzWEIQZ
aMkhL4A49S7ShV8ABx/L0nH1BS8Pl/r5dVoSfnWeQZC/EugcyOVQ4tKxkQcXHqcmYrdJcP9dXOpE
eCLsBEMZGqO0fkMBxTzk4Z10wCNI7CEtyOLu0FPJa2rw2+ukJd+wIeaud0z6Ke2Ykj+6G2XVL8YN
44OyQjRTcGFGek2+OJ7F7l1I4XOcWptLJa+D55TOMpQkh5DPeUcFqTplZrtO3PaEyWQi/FUZsF92
YOXUN7fVhSpEF5t+0KKqCShV02Jy8z78a373z/KtXRrzzE3SMDjdIzhOVpy3TvMd9qUiZDoV5mKO
PApufMCVnJWz9CMckQOZh1kENOwnuMvCY3pwUJ3bDncm4aWNIG4QT2/r3IjiE1heButLpxspV+Jb
FWurSNGYQ/m8t+aHTBVHbppagif4iJno9Xc81l0V6PQLAVKetQe4SXfrOsl3plo9Pk+o6IHNhQDf
zglFfhUUj5J2vAPyrcOJzjXrWYDetUvKvfHno6Or83oHxTVzKuq+3U3LBXKsJpZthaHPoUT6D5s1
n3plBOColnTDsqcRYpxvUsmG+jNxFIBxJqQ0qZISNPfjktCB+WBkIlCejP7DMYlIEcqQ53zdn4Vn
9sVG+SaWuBb4+hTN3uGJ+2594P1P6gmYh8CST73JPzkoDK1RZQa0yjYv8WIqOogtcdEUxDEWpzhG
SWfPCCfSvDC5QjsZNiRX3h3Yp7otJpxw+pKZ+XJ02eRyJBXo7HpytcVtIHeXNK51YUPHzWKBUuxT
ddzwALln43IWMctcOtLxFNDwnOrhrJshobyAeFHuceNelbFm+j9ZM2yVNA4F8KNABppw/p99Kq6b
eL92Rk33qwY+HQwVmmFKcNtChB+eQFmIHbrx4YaPtYWd2kp8evxynQ7Ytl+nsP35HpgDxbYSOuhK
w+JEoebuTodGwbAeNDFGGTuqefFWF37OfXmcFnVyTUGdzOv+80MRS6ziEfSw0d4KySrBU3gp47SK
bfpxhpZwqPyoEo2t+oMPKNQznxjOLVlvrNBg9j0Ysryv1LOByCZwzzYhuGC666y/vet9GQxZmNkn
akTXhF7TpHvx9YVTO+GhB/nWBXB8S10O9AyQ/YK6L/286e8ZRkv0mW93mB87dGO1LZGEuAxeqlTm
KEBQCMfIgdWik7PVYQHkVUjn/jb6i4XmNWwuVBkVkqiDxukYi5wLUhHzIgJCy9hIKiPa/V++hHGU
XOgZFfnE9itdeyWPWzfS7gSxgS6knBQULPoJviTP96yacfqzjpjFK8vuDge8xI5WJIKOXR90KOP5
kyUOQDWkuWHf62UslolOHyWC/CpSHcPSgEXh7B5l5phrmU7FrWzZ6kMzYNcYI50OE+q6ExB9SnvQ
Hgnbl4QtrPWQmDmMzPJnKcEM0Rs+GHcGmObmrHt/OqeFuKYzfN/MjG0coY7UVdc2UbyBmlFSJMB8
RSbIQ8FlBDbnJ5lIVvKkG5yw+Zc1dSgHgoFQkn0pQw3E8GERcRLjGF3vsxpwMLRFjKT8qFZq0bzJ
U6WrQflrd7KN/XYJgMHQf4B2k0tqDvzrGgYzI3kkHbfQYb91V3OOmXqH1MPHRY3f8kx7KcEAsqrb
QVsv9QUkqBqUhkVk9fjBkTXIHlKXwiUusJ3Ya6iSbv1nAp9DxxRT4cGnrZQQeOKoTp1ARbxxuZSY
3XTIblEdTdLug5HUJPlBiBpvrjZy1IF8T91iFEAxdYe7FTTksfQJEvP8e6pDJiDcfl2uDVWLfPol
zAFp48omJrsFSBN110qNheRNQcO6DG45YVy/YzOMp93HFIUQL6E/0KKRWkUs2/oK9jwKmKyOWBAA
B48EhjRnx7FAbu/fE6GmFkjaXQl4HeVT+xRGAmFq82z1YuJdWnGw88ExggqSU48CagYWUm22lVS5
PTLh/HCvAgiE2Yn1RGa9k1Dx5sp/Qji8NlRFAQv8sbcwnz3ptRr3O1RYgSvQ0YN3Pum1B+zDPCGR
9eTVEKK+yQOmcbrxaK7Z8uV71XQe6a94RY4sjlKhX5Md3q5PxJ3EQ/TcUgql+yRzPPqv6iXnlgXP
6kXSg4TgK+AJhXjyycnqN+MlqDyWySL8bnELepkifrkjcH/SXnMPO/2hUEvM+akGmQouYz5TqbMP
iUkk3av/YoubF69s4maQe16Sppwu7W1hEAK0r4y8NKBIlw/nlyCNvvpH3Eeab6qDoFWgIZAYBbna
a50NGEUytUMT+BtUqwMw4rcSwfWTzbC4IYFEXSKX1eUubrPBG6hvV6nZc6+jZvrfRlcfvF1YY1gw
MGg1j0zQ7R4wv2YhxZHTfkbMlV5nZb5xsIsiC5cg4U3XVBmfz4LQlWPfZw4exGWXIZQ6trL4ptdk
PlSnQ7mn4T1NVAixtxz4uPCyHXzrl+Qr/+v1iELY4FSq5SeGTuwdeiLKOS9VcL242zQLISklCf+i
TR2WSwf2C0Ed0kK/f1fT3at0Af/Ft5AUFi4z7Hs+XQBwjs6YQFawX9Jrg6C+rrcA///Xcvzj5V11
/ZqfZpe7ZjyZ16SwrgMHu3/Fjut5weO08n+xSNxwBRI5bvaeXUL4QExc44p+Ic6lyjcgnPfz7jcp
S3nqsmr8fGit8/Ft7llHiy+VAIKml1SURY2i8RAZAnzmBdBB8q70HqIPRd0w1/kgZDXTblxTtV6L
bDglFVTxZyDdl8r8BZeOWPebVOPu18dzU8njpue2xXPqpT6miEhWowZyoDaBZpu7CPQqqzMWBwth
y5QO8DgAJXqhTT0WYw9u+j3z0QTapNnoxGyTmL7N1nuNeqRsOG9FqkMhPHKWhctgqwQDNVCJBmCy
zQFBA+R0zWc3nlpYbZKjo7dyCLsCwyV3rpHLDeZcy0E9xKrMLClQxSoW5CF2Sjc0X7UF+r1O67u5
3WKyrZH2w8mNwNH63OUKwslh2hkaqj4Ggsj94wJ1TdSmfF/SXuFfM1mFoGtjFsvQkKlK7KFqgkg9
tM8k4nheW8tL7CaLcA7kHuR7VRFryl1fAeNZlHfL7X8VJnlT/O0+GU17SKnLex3pXXKRa/NfxUa6
1QDFubI60FF8zYyxnbb6WOMDTK6rlld53xirS9sNk/6ujqbMBZJ6/d+n5m+oapuZZgigpB3XfnTP
jUjVgvTZ/9qeNRXgCZjB2wojqbPDV/IWTI9WHNnb5GUMqQUjMEOWHX0MkwJi4dAU4PcSYF7XUodL
aypp8IxO6PPUy61k37jv9Z94371l7dvbveGdhFrDrOnJD986MBvQTYpNZ1CBqs7EFGoekoU9CRYI
cNHvF0B1rhqnFqIJIiKB4TzQQN2A2nmZ/wqrtgVuq/utXCmDf32N5ID+fCAHQ6beZwLWPXmxQ3oC
tvCBFmRmFCU0K54gCTJT69ZIEaPqDe001mjLC8pSjhAY/1NLKV56ptoJ2VTaJyH/haxMYgpiMcFn
WdEQs4uqP8huV8ghD0C2I4lc7K4OHphYQA+sMXpmgKHE+l7wkfA3D56Aoq2UA5eoM8+fOp9MvLvA
0Udully27pBGgevvn1H1cSv9lJzOQRvIQAqsIsCzwK//8lt1TicGAGWnhbD0ez1NM/vH4rOW2Rqr
U8nqS1wYS3Di8BzFchmS1TG2cZ20urVOUPRnQcR2mDJykbvG1TbHAkAlog52yiDthy+5kHk8yJqv
mHk68vyFSd2KAtQMgYKTBV4i7f6qRB60BDAgb8XoabEPaGBpYdwcrpVgiFVCb8RDoh6EYBsMLZQN
dwTfchuq43a7rSucXDrirYvXQl97Z6scW7WYg2BeqGDdqxHuFasBZDqIpNukYqDqOPwk39EiZXS3
UsJKXcxN7Qft5uVmEJ9QBSSzn4avBmMOTK2LCW+vjoWM1xDqWbqR/8M2yVpqRjsCRaQImJIwt+NQ
bJIOpCiASnzLrlL4YqjzhCejwJBChh2GxVP4rn2UUua5s5VDgsHu78C2QS+SrmDQ3Uwh0jgsCutb
zM5ci8rz6dSRsRCCN8WNoAvNHaVkfQEBmHEDS//QOgFgEPex2PnV8yJT9rcc43z3Tlt0jDkUgQI7
DzONzMgtqj7TMvmw8fqJg54B07lo+I3E7R5kdz9O9hWLMV6g04p/xRzljEdaD7ntOyA3CNLhQHRd
PSISJIe9fNtBc0hOn1HXh1JwK/fDBKkH3l47T8rVIa92TRW93lkW2gV1LXTl3MT78wvRRSoiiIBv
kRgnJLKxe1E2qW3in5Ob+gvZhlCSs+bqgfK2QJEKtyOKvhfOAbMGihG9E5CJjOHOFxnAIrDEmgtL
imAIuHlbm2SOR/hyTP+E5EEu1upLmj7KCYCtv/ucHH+eUHAa3CZMBcSAVbc9myy2uVS/krPl/S4B
jAIXM5KIXFbZjJ9jZ20V+NN55GM7vyT2orlPc69zjyNRY6zDnBPZCAJFuEXm+msQLsBfrfzZrKGV
JxVXviIHUKYvnklB46V53CuOG9NjqPKN6Pb+nM+QJzhlUL1WeKfmKb6idxokIh07l9i7C0HtFoXN
ig/y9hSh1H6IzzraBRBGse08pqfKK12pkrPL0YyC6YKB/NBQEbX+7OmK8lcH94AF21rNL5RKY3Ly
sPSrZ1uT8kK+PJs8yxfKB44XHDmXsidBHynUfLvUmyKlRBvSiv1UcyiX+A36+RUtYOesOxQVEyEO
EewsR3x8DG1Gj2/ITdPyU1Oa1dHRsKQXkxXuMmvpArhT4FoJ4ictNFh7CmL2xkDtGK8p2yxE+ikE
CfYFXetdsi1EmYBcrcJod65HRsSugmUNzl2IGu3xEAJp7BkOWUkxmoxVgWfj8Nluf4DewoliUic9
zq9/Xi00O0IWEe2SY1Ij7lrf/yK9wL80teLRIovbKZ4gqTnUHcogNJ0+hsGlvwKEn4I8o3ccSYtI
lPPcw2Qw5lCNJCgjhlPhb+qr/7pgEnP0+V7byolFW+z9JKS0FhvmI4NCkU6AP+XPj4iaM7MZMxYU
2vpv5BeP+G6dX3qKusivsV8V1wWGvhFnjYKMHlx8Vlv2V2fKYIsddqxJy5L/zy28jddYtViUxcjT
s9OSOFvP8H+V326IHJZXehNw7jGCmIRCLJvNL3iS+lI3pxzkIa0VRh1LbgMflxE10ZUhQMCBq7JC
KCJTdCYtoHMhLoy9peIAEAkJvEYSiROe5TbpZPohkFy4maazIdBiohQdGbDBJTOlYzcbuwFi92Cp
emskwufgdW4VAZOIZ6DToAHg7x0AtvDAoDgqPF7a2KIMyqYk2W+Oa24SIz9n7fkQPBRKb/D4KV9L
fWdmtHH+80tLP1LzcOCY6KPHvD6IEMMRHNE1isl7hyXayiDd2dtpUAQRHywYNNA+yIRyYRrPPmSF
vsro6fvXxpUpB8/zfNFSlwJVl/nH0ooj6DfIz91J53gp2c+H1N+0IWsf34B6qZkqE3KfQdlZRnt+
HNpEJTlpmHgmAhlpIt+y7Auaa4SMslyFfqhHnSiCCoEr36i/b/fyrk192DjOlsJHq7zCZY5vhK5+
5KXqZ+sUB+fbeAYFojT/MzwdNCZ99Kd4bWVhQZvImuvNHuBZxN//x3FV6JyGUsMtDx/lWTZ+seBu
SDGSOnjmHhB+OSWDqSEhstXQvUGONOjXcrodrJLgI+fZqZFUdTXCleRkPPqw8VrSMytFCUuFqBjN
FbSuoGtFLAsRJx/cF17SK/LbxmtQxzlk1mL/M/0XnQApM2Hwe/p9a2NGBoHHrtiZyfS3HgtY14rR
QkXaMMbxdzD0xSIRj7byMKkhtHh1H5ZNobYSopRRUpIjYnZWgPNip9qW+ivFyc4tUncWZ72bsBny
4GpsIzeETMyLfSMw1susi5zIIEYfyBNveSCC+qNNBk7dWirs1kn9S9oowoFdnoSb8VnA75Cds+SU
rR7kwy0zeO6OVQ8xBtMG4mZAzy+VGpWybqMcsPsYdSo8Z4du5wUfE1SVpOmPmc7Ap8ce/dCHmfd9
nkGFSUESrmn1SnIBC3aLhs+jbEYVcK3ikyh8z4rNb1+LHpCFT0OQaPm6Gv5JGolXRTNCR5qhObQw
D/6tgxH76RXBp1mFq92NEeQpWOIZI5Nnh92Vi3ZbXsFZ1GW+X9pE4U1SdIWXKJP0+TIJcqgavZ1q
0pOwbdVzGH1fpmsmqPuI8lWMtKhQ8/Oh3kogQbni/8NAnZblZnaC0VdUCDSKhDuIK/k9q4kjsxto
AccA0GjaMwjtrTaKc2RrFH1l1pjD4PUuLlreU8AnUbpgjylouGO+GvQ7xzTVqFIpT43JyqbP51lY
IkWaylLyvRdW6EnYlRwMwRsqJbqSc/hQ4LOC+2QMp9e0DRpxaIhOdPFPBEUP3R72HOmpwGbPidyL
ZyzkJAui2Evio2/hmNbKeMSgnUUVHS2W2FBIoLOXjroYfL5crNbr0RPywgq4+sM/3NUplHNwQFYV
8T+VzQJCnLM8NypwQCCCVj/Dmib2Dsjf/4sykKyDndMGlv/p+A8/6fDSVinP2rr29XH6nGG8rvsL
tUWvRkgnI9jklYXsxZstQH+4MMl8cfnIJgCkMlXrRQS0wXk3pxcKB53L2h/tSAzwYDai6/WZz2k8
bCjMmVlUkhfcv4hDRWb4AuVo250fMh3RMXZ/tPC8nX5Lp3vRaT1teHdHVe21QOLGARapbHLgTIha
pDMzc+knEwt1ZTBpktYg9RCpmI92WKidMcx1LvXlkhQKPSQ2+zt+284ep+NxDHfISbFiWXnLvaOs
Ah5z/4KqutSTY/gU7q9zRn+HgWAMFOgjmy0TLtqpyjExJe8SzPQ+6rAgya5AcoJ65Wk/JUIcWwlL
P+UpwAdDvOMMZqr80AIdRZf0wC2VguT7gbRN5R4va7biI+x0hpxcTUwGXcwUCsYO9qDRK8+KUeVB
FX772YKDAom0m1sU7aNKdvOgF1ly+q5CUmhDoJdb63m4JjtHwQ48xjejocj5GO3i5ULP1FULItH8
yuNeyaOEM5SFLdQPN1mr0saADrapJQwR1Z+c6PrA4HOBXzUkO++nf24JhCstj9IeQxB5L70Z4Kzo
FUZGJ4z2M4JpeytE0K1GUbaqoNA1rd8hHYyAE0yVmycTmeDqKnw1G0X4MH6a/XiZEZzX8s2BT5qT
TM9mYky3IjnRK5RH8079RsT4+wivzgHIJlSpX//72XBV4WKfvOp6Irlaomx8Gfrssb7zT3244qLQ
LTWnPqCdN7TJhSQyGXTqt5aCGn84Hvsdc3G9F146/4VhnBpbSmRShrH8e96YIa7DPJDn7/yQu9aw
qM0tjqcmlVBavLNqAopR7/xDKiUKL6q4lRVn2KV1uilo/gmM5BY9NYeFS46BpzGm3xldgGsv8SF9
xhtGTYnPbOYLghs5pL7spYQyxzdwRdFm/FPnsev5xQREHKxs8jVNE+JhG+lssVmr1e6mwig2jWRv
shuiPbjPGziMQZ/CaI0a/LgZ9cQTO9YL49Dx2SddVOrhUUkv5xQwNRI1QZkkf7zkWq6I3Zsoedtx
n+vscdwb9qE35qg8uSk9Vj0R32Srnnd4jR4MYlTKh0DuzON/ovERIZCh52mwkjddc0GIrGeqwZIX
2RCQfyTF1SSsNAafAff5SIiJV9C3F3lrO+PwwCbg7gEd6mln45KIaOZzdinfGkmT8/52L0ZjwbJ+
KSK1MnBM5HBbl5g75MrTxXJqGgpiK/gVg8ntVRRT+gMeqLoPcyHu7IqXXeMmqDTH+ywF2guV3GyX
l6v3YMzGiBHOaT3DCN1xCdbAFTF6QZme0knvpqwcjXyY0ABmUs+bTNJaLXQxMFWGLAwomDKtGsQM
GjbA7ittHHHb4nSortQUQB1eqeO43Q7lE6UsAds1oTgHDBTwWm2Vu9ZMrmGUnu8E88AMP2PSOasv
0LSsuEXtAWQVOUpQicCBYcB3ng186xOkTXdgeDWSw4XEqTaWx9mPOJsmWEvF4zZk68RqsgZnyuQC
WAYFOBOdgVIGX34DT1jEHDdOWhutdQRwJcV271qXqiQYymXsgnK2A3X3TZRGZs40TEHnvUbVHsWy
ZOMqAFxAJkmGKOvCGHwz0c8DUrE4rNfGfyNb5bp9SobbRnydIvPbWFU6k6Z217gmwMAtH9E28pQx
ZLCsn6Tr3AOBSt5Mswv3ZTsUtfjmZmXb2KedwOA5mosk7NEGS/eBrt8zHRZzNALI8ioUOxvi5UiD
6bBC0uH4Rw+mSh/nFtC9z4CXR626urh/eERUWwt/pQvzjgnCnk3FdiFN0/Cv7+jbcJ7I3z5r2R/P
A3W89H46pMj+eh+c9WsRGMOf1V21FuUAGuu1exFR0Q5sx9+pfll2r9Kr+L5lf+U08NGE0MwvWZfW
yxdgzmiYemIuS6UXnkphFa3Kaei6N5sfF5YItXHWaLGtzUHqb/wgWmBSLy1+oIR4pzit0snZkVaT
q01v40s8Gp4Fhv71p8xeTBdFRz+aGbn3q1st3kRsYAyY4i5g9Do6ao7NFWkjGBXBkuGcbC6EvyAJ
2ipSYMnOVx1vTmZTjfVQ7XybeoNUTW7ShCvfermoICmazCBML3Rv3T1z74dtD2G5LEl1RgjZ6aGJ
NvqsRuqPumGx3Zqf6D5pe+/O1dgBwiNITkuXXBiMJOnvziXlP8HdNwcQhGWf4ofq1S/M46TZImnb
Eon8VrXAXwlUTYWg6YLUWMFwBMo3JZ5CwZh+aXj+VabgQh3vSSmyJNfbV4MxY0wte7RksxyuPKhx
6D8jxy3DFvSXriAj2modVyewQ+iIx7Ou3O8M74RIyRzZ8c+mStckAbiDeQtnY394N8tmgexvfWzT
1i75X/G8ppqsDtXPv+rreeGSt2ajUTlwV05XjaXgxj0APm91gYPY0Z3yX20Z3XWnw5QAu1Iy+EN5
+QtKER0JIh5QDGy3E0kzfyjpwec8pcLSw/RcLqUgggbW0jo/qOzIQxsGHwEOTkwsO4s1UQ8Qyivi
cJA2rql/+aLdZiWmI3/E8rEy8u5nJP1yty3S17kJSiL8rYQUhzit1DNiLUqBlryUyX0Xk2k+DSGa
ZWwpXE1Lpxt7j0F4mJdtHjJk1MYxthTsnUOnW5EkiDMPWj1LGPlE+gzr4tJsFkFv+ViR9P/CAHlf
dnEATkp0DRXlFmhF9jjBXr3ZNLRYO+caZlMfdOjrmLrLIPJ/kZSd8LxgUqAMpWDQIn9fS8o/smlg
H3NzPWVzLG2lKiXdflsdd7PzYff2cYT0ZEmSTLS9vNQtdtOJCKQLXCNbLeODrF8ISkwzfQAgl/N9
x4Kd3y+WxUNbQ3z1ca2u6xpyQHPGtMR8Oz1hgiKF+BAaLxgxeW5QlNe7p4i2DdSV6mmQnMQrEgBi
CYr9xKnWuThPmhHlkRgZxznw5GuC+hyPv1reoqispwczNBEH2QYsHBm+54ldNI26FTff/QT44Wu0
hzj2sVv7n1mbfbfJathUtRFk6hCBFJBQjd1IHX56OgUv83PTYfQlbVgpHxVVdHoD43l0yi19Qjiz
LPofM4o0HOCTfoCyxSL7wNZg8ZZ8E6S8hLZzXaEZOIj5NMPxt4gWT6AGOm85/GcrXQu8YWyP7Z5v
3+Z1OFFhx7Q8rzum7SYK1tT4ufc7e5qrBpcVO/a0QlGWy145Tjq2GzuU3S9Sazxb/lkcCuxprGBy
5rBV3mXmvyb40S7yLfNRvlC3mi2w4ZVuWnhGF1agFtvb5R2rOT8wMuFjeyECdh8elS0q2s1l2bTA
WRZFCf2UPCs84di/ojBvcEvnfu+07KDcxxAJtiCkIZwI2/u8OXKzHoVJBM0mlokgGv5/9PeSPVEg
mtsEpCMezJQeiuajqRqgSz5j55LhvTiTszhZCk7JxcXq/y98NsMjmnYZQ6DbhNyFTUGNY2JoBBrD
ak5fIHQCSquPzNjqh9afQ80WPtstPRWpIL7eXCv+xDLmqwA+aMnu2aQV1dOPHaBNs0A5F9L1QsuZ
H7LerVIXuI0nXUgIhyU9KJRNOfGf3OCAFYSCRe/e1rpDlUSm7942cn00s1x+bpXZVsGN69qIY4M4
HGA0CkYY82Fd72er86e2MjaIAqPoFQPqLFa4c8e/8P8hVFqWEC+vYzxr0+2ZCFOot67ItT32zy6Z
RQFXTYLeA8fVtZf08VMKPio37+/HdypzeacrNMSOI8tm17wQ6lqP8NhylQd22+bGraT4f5PUmj4r
z4wG8HQzh+xGJqF5dZjS8ueu8Ga8waKvDHHI8puEUAt/mYvs0s6JegRAa730YY22wyKsURRB6ycJ
wjR2F/hTAJEkuBvblf1OSbiR1XlOXLQSuqzL7GmhRAqj/O2dSDWlM2cxfYn2DHR/zNk/3erJQjki
7ztwppIqMz8DHGL4PsbzaFAlu8tMTOS9oV+6swRDBLOTTXfwJtTU+FEEcSRckFh3tUBs90Q6bq/b
4VivvLEowbUnVEMcRAVNELBUxjzudFS8AQOJzgaxu2f2s4G9A6KpEGLqgvXhI1Dhtdm1gnLd9DjS
rRcxTF90LAJjbCbwwlFZnrR/7RdvDyLYNZfKIp+24Vi6iEnCygSINeNnxmmHrKRSo66+EScLA/GU
y3hvugd3x+DyXwSh+z45CVxCutDg3m9eVuZk5xUaLCl0eGZTzVJKUpAGWFHyXpQJrCsnlLbtA1wY
cDBgKqZlBOTVyXuR9JzSIGExW0RhrnGuRJt8l2+Db3vOaYQw4PUvoNcXtbtOhUGGi6Yhjmji9NIp
yrMMhWZ+ekBQmxGZSo7SMqAjf04k7ROfsS7ghVRIrYDUGhkGFYC0XCUeOfW3UTjojPNJxD9q2mwK
krhfYJs5dPv8XPNBra/3tNLL+p0DWKu8jppxmx/rQU/VvL502SHlvFkSgCF55Pnux2n2p/eeSVrZ
xAHuzmXNlTGICfbqY66Y6gm2xIjPVCQmOuss4UCDxrQPQRnvXg5B5FMX+Dn025Aew7/X8Vx8M4TU
lbMxufIfSCy7FjYuIa56Z0epItYIIlj5hjd0K3o4JJ2uZ8MxMXKBRbnLdocEZSfgF0tyO05kcslw
kECeqlmM9Wi4XOVcPeBZ5gbzAhpkKR2PPCWRv7Q10ELUi5sv2fMMiXOUlw5f4Ga8mYYyT2q0VNjC
h3xzTqAdeSLDRTKu81huLT7bPrOTRiWhz1W+74eK4ifbixbbB7TfmQ5AiTZYYX+zgCP/FVKUKu5g
psb4aDj+yPj5Ysp3LBQrc66KVi7ti/PdPcCktnlM2fGtuNZ9z7zdfeJBkMY0RCVXT91v8Wy3LE9j
UU4dz2H755e4K/7aTkytdnW6ZYE2fyDgr5L0cmUAEt4F3jfdgas5GlMVdLBp5TrgAGBbDtYpHObk
AXEkJuyv46KZo9XIcefX3U0K3IBBrwC4MhHWLEZfany797JwSMnJ6bU4PqJJxwCXX5CMJizjYEkp
bG0KvB28mLDz14nC/W9M3fZyqhPi2LEl5k8yqZKjESP/G50xKYv0uELgfwnGFG3GxLDqYPkqIsj5
CFywEhnO6OdCaOwYmckGHQI98OwFmXICKO4jyLkOIu8Hc52mdMO/FEO8Wmvcx7fetra8Fg7P5QvM
DaAUxjNaG+GXs1Ik7v9Fp1yKYnIKauWNxuDunZMCAGjFfL9d1cPaSdPg7GMy/5Rlv0uqKdbyhnhs
vfXvxyfX7tUMoZ5B6iaSWrXPiakD9+IIDIEB/3Bc72tNVqsl14TqMFuRpKVj/dlLYGHcBm6jM77O
bFx+VsFt2XHueqSg713oYfEGb2VaSzokRDrz2QE4REZlmoF+sFYQwUccGwm2Y9fsyPJRlxyYj5W7
hLTQaK32/LJTi+WygvfpmK9NRaHoeZI7S/52rByHmnhGXPLVfoSRVRyIpk+6BCoFcicePZ9ATEH9
6qxdbwgYUlASZhi2uprKFiFX5OHx2tDJUPrcxBEVw0WLUx28HlhfyBPzayRPMH1yncCDgahxs5Fb
kEiQvaov2fwJW0NO/qfl+gjoyV2ocyEIu9dT+SZd4KfMLxHm7bNIjkVT7sR+qeodyf9nmVaiUDTW
TD/pO7BdIfEr0XxoyDuwM0GnSCeMhDsyuv3E8WyH6AdJKUP7xfcC/+IrAyTDNZ38gawwsPRLFqrE
jOdLD2YjvnJ8fEbGJwCa+0SBTKgny4MxrveaxJNkY+5bcZRtH01+o+4m/Tri4ArDm2xVREY8G33a
nONG6eWLRSectxqOtvTC/Kb/JLirWDpaz1Y7NDgi0F3eIvqmEsL3JoATYpUzcN//Ou/wLDf/EBsX
+xcT5I/Kk5sV3glpAf3snAdKO3D7rlID8/k8fZtVavgVDbG5w26lJhSRhiiFkshxS6VhStzaa739
mOZnJ+X8MhegMQE8smONvGrNRcZSVnmahSuMIFrES8M3u/I9KcQqyhQ4vuSZbl5RQ1W4rfTuIONH
M31JFdrI5ziLZx2lBAekPYaC69r37/+LNhDL9nc7kxrbFZQyUzkgdETzXoBC7pvOJbg97BodWR5g
q+IPXNZZl9IwIlzVNEOL1VvFpncrwuWq1Nx31fDM2+yO+Gd5gT2Ip9DksQW4RYKZVfHDaBaqE4Iv
qoVMEFy3ZcV1YXzuyVmNvy/zwNFqUgPje1INKGUYjDD7H2m5Sj0hV9jkItnojWeOjLWaWsPJImlf
qsSX4y61HS4pV3VLlhThk1Jjj2/mrIwnxmqf+wmlCJkGZqcL3KgnuUQCXHQctQgGeUnoPrvuxKBk
n4woIjrwRuOTAf6J8UjxETN1Xm8LHsZgxd99dYctdOMuhEE8bV9xeDXEA68p8F8Rn13DJQ+0iXYh
LdD01FfTpNaT8lM81M3GJ6m0hfKIMkDsdNHi3wkbkjBwxRYNiPRLtiO8WtHaRO0kQ/oygsmOqt5p
MkSW3SDgUhLTBlgZKUWVp7NiXiTLgHP5WoKIZYeBqnynHOPsnhv/pImuwn3adN947L4PD6BMX2gv
//uaXDgwAXbokf5Vnj+AFkUQNLaNSGxWqnTzznfa4XPZzV2KpAX/coD73OZYGHQNev15kFSgx1DB
vGod9otLqr6jz3telQLCqK42So38OY2l7ZLGQvWXZMClYmEnRrj+icRX8npPLbOGi33zY6Uh/5zo
TvwOT9/o1aWIIrZd2N0D38tjNFAQZEJscHLoaU+h+3CVxfBTY/wQ1TrEpgHx7hC4Ix+VSBQ+/Ouh
+6ijcpiLt3q2rz0CS3qYplxHhLCoSlMJQv7Jw5sKIH+9hFPlYVrokPeTIqv5ewv9r8kF+U4lu4a3
idN6GkXVp7bgvhY4CRa8AGsonY299rSeCGz2F2S3f0F7JA2UpgKGhwBymIt37MUU+nw9FigrRQOC
OPUMmCeTVocoFEDpx57ty1Jg/iBtz+UI1oOMig4FFB5qB7ePFgED8I9gYrQ3vlUGqsQIrl1gGl9V
mhSoxiDZM+qrKasxGMVhllpP10Se9Vualj7te4Xqy/fy546AJaO7UVelULEHt99qAWbKgok9jNtw
zVexIzYMbMybeRAG5Q0xTwTi46noBcos+pGA21Iv0Oo/5HDfjdBd5EeU7YFZXBUGy9QQRleRpwGw
cb/l3W46VYWOJ8pjAHo+Cj1VuJ+vBxrRo5xAFKTumIlB8QMIuTlnepqHvDHvcy323pAJ9yCvoYKV
sPq7pwx/CDHQGthDueZRynKpN57MglA29zFAfPQmKOlKvO7iWosvo7KJb4K4jW4cl8I8WQc8M/97
mGaHo8tXCoL/p0631G52PC3nEdJtewMDj/m4qgyQxKnawPZUUopifdTWbx+ffzBnNRDmt5sWMpqT
E4GaTaNZYu5rRyDNRaq3oZv6CGqXXrkLTkfVrkbSHnkBdoU3YaqN6MJIOOuQ64gkZ6LAUxm5Euh6
vJURf5omOY38Ot8UIsX7k7elRuiERJsiCW1Av9WgkXfkzP5FRv2nLExI2ko8c1g8AO68ql+fasGd
avh6bWzX2wOW94Qr8Xtlq5wzIE7w5j+6/0aNMCY1iCWsMr1alr99EAx3zK7ISRdNkoe1DvpkPZ8W
A+mMMK5K7khRA4PLzTz+GKmKdFbGkfQCk0xAj0uHBjmnBZ6gYnR1xBUS2y4d6g+mbNmA3tQ3az/L
QM4Ulfrn1ECNr8HF+v3pQcHIdUOuxzVMTcnpKfgtxKpVU8s6Tz838ubcAwbZLbLKqQuBthNDjNZQ
jXRU0k1HsKVZevh7hPBPKcI+dY5hsc36i9eaF1dOiGTWGD50pRqNl7uThODW3XQZ/op8j31u97/q
0Il7hyvdW56PvOSzgxnSvTTDkcxL5+FM15as9qcFMFIvLysjGYa35cz7y9oeCSxxwMiIf8yekgTD
GXNwCVedajrEjCt9GErkwTqAJCBq+TdUh4RBO9gYUkgAJNd1JayoYM/6zALP+Hf5uFe/VfYzaWQX
1T2zMAPK1YDFwHYeAzlhOhwoXQIiGHYiZmlVC8hswdvx4U7zBnZRDhHnYxDIepse+CxlV2IjkjmY
9DiI3GugVQT7ZLSI/fgnCqujfKDtjcIrh+yCvGiiUwVD8ZKjg2oq3aS+fhPsBSUmPUrPitm0eF+P
RP7lS1GONGOqblvYddWBxCJdRSFxECsH394V8KRWZcgN8zeBBdOl3fN0VF4Kg1BnE00hUed6svFS
il92OJU4Rdd5kARdv8AcA+fi1RIXu1BiAxpYIzm6aqJickQBdVMDlsDq5IxfzQubRsrWAAw0bcMC
11kJ16YPVpWsMoutLhSQnMUx61KINM0t+sveHzkxOuSpe6TCOlG0oBUOBwqbmyvs9ivGYCoqE6WR
nNRfp1j6Idiy4NOWKVilIRoDdgk2YVlBEMZyyP9zDFAbmCBYqeJ7ACiZK6bwm/UqOJeA3eI+NweR
37KbaAlz3M6jNgmSXR0vTg+5lPJ6iyo6TjLMgLAXKQgju9J2EDm06gBwBT03DwZbgC3zwzwgqhhC
3K+TVPsHvhxoMDazOHLD5Q01C+owolsbM4x+s+CoW07hGBGrxY7xwwR0gvm+GtVlv+Zs6O7upsYV
8BY8u/HcdpHhMa9+ddobHOaVcRqXQvvDEI/6dThuhujAqGvU6+cx2dMLkefA8FZPaK9wF6c9yRYH
rB98qCV+be+MX73Gh4TtwBGFV+AbTV5LSlmj9JEv8OwbGD2sRpcbS2roa3lUGgmiTSahMsyfwSRc
ynp9CnISxu8e+4e6W6dNZ/DeBLPip3M3i7LYFjJFVnAEbE7keDmE7BepHIhBIzPfebRyxbf0Uhr0
QTwL3czkC9qf5gdSB4+8sWsRJDomp/Q2rj4vL9cRJcqUU6XewciJY+uPpmqi2PnfFGMHtZxqqgdH
4EsZBZgQ7nsxgb5BNbblwjRSPq9GlWtSbkDnzjyKBKSYJOjXFcqeNjKFYAxhqk/3lYy/DcFhm7O7
gj3JYG4ot3p8EtsCYX20RBsF60MytWB34wo0Ndqz0023oBWYLgoJYDLk8tM5nzDg0afSADw3INgB
Aeq8Ibb1SquWeHW7AiZjxEBiSzCItbyfEfKMjV3zkEzJDIoAhwwWigJvnb43zW+gDb2B04iSke7L
UFrIdJAy65Miil2zrn54U0fCtuCpgpaNCqPPoBlkCJ9AnGPlECNoZU0V9ZrPlNZ5FqAbr0sAVPEQ
g86JxJhwA7njHRQYEJxfNqKrOyl+DThZwEvq9RHxi/kNkWJBd22SL4MXPZjm7TBHW4BabM8q68UD
cto8YS5jA5y0N1bWxH4RTZDmHSwJt7/5MnzmVQ65fDls7BY2AaqMndwCwQ5nprzsuWCTRiadqeka
etfXHXb+Q+L/oSPl1csEFk14KKnpzjLRns/3PHY8R60Wzu413IDGWJQKXaGE9lQYi8y7RnS/PQKg
A/ZO1WO10G3f/RDXQyZwezjDTOKfFtBoNMc0BfpwWeLdjBSMqoQf+2EfJ81A4OLu6xHSGDOSq1ON
lWmShxx5zgE3ookxtEs/hWQclSVH6L7P9zXVhR1I8WHlD8cTye45Zkn0g+4Ek9ZmMGYa3K3dqd7o
gUgr9Ldlqima6cywBO3dx0iMqFflfhGJV0ac9f1psimpx1ZWaOsvCXY2l0pI3GsxbTEWaAR85VTG
hw0wha0l4qoe1YBwzq/xaCScnJj8Rx2IzdV+5ZprHvn0zazf//DZttVVG2u7Hl0T8tsldh+OGrPK
HKK60osQbsaxyPCrQnsG78emRr1ebrEOC4eEoBJMUeBnzUkvYRb6FzbNHsKQYh2ZDg83WGwzTW6u
GMwtNDa63JwKNd38O1FJ0Y9T8cRpXYvSSSEVflKbsIIzvOWe8y2sXCMNrP4Fb+0xfTU1/CklR3nn
aYVl3EBwEs5MpAbFrxs1bxmELzjHz1ZByfkkjJauOZMI+2s4h9E3roIEaJa77zeGdA4vWQD1qod/
l1DBPS3iYREH0Wh7r5Q1URvx5lFD88Vg/+Tf4uTg9nefUGOZ7UYBfE+aMO0pOhLZsl5eeFIwckv+
s000mjSUbXK+2zF3PcPBfbwPFGxkPd1aovYhinjHJk1JqQ+PYjT0H8ltf0rD0oUgChxWTonvDx4v
kNfivG8OWpp5FfKCCBmUioyJ+a7AaVjJpcdmQBZSk2ry00ZKEV6Q5BdKMgHikK2n2Zl0W3OGKX8X
uE9n63r+R8J0LMGDEIWcoSbZ/ctwSXl2VdyzBCUisslX4neZSG5HXCiVdfZ/h+C0LlXi9DiEeiPL
oDrjR9hGmleZaNKi5WkmOE6xsGqtk41v4kKfIpivRTR8/syHdC/pN95MVloGINmEyVPjCA6ttLUr
5F+zC6bMVZgKQ5zjJzEm7m7zMP3v4wbwmNfDJ6C6zvBKDXLPwgsJdJh/weuayp3cPemf/JMhlB1D
qqDFoqIhv5hw/4JMfTgVkSsfVPu+ZudomvOD/iC8oMA43hdWPwsrIjucOLzSd+16qbIWfFxm7UOJ
kWHqNruWIYtFaI5BXLwhzpYqbQUwKGse6sTrvMUPmfJFhB0lkcPTgp32cp7uvL0bNL6vGgXtV4MF
l6eVmoXN6uwIRvIReS0mWPYQ+8QukEmnrriWbRXJzO8Rahxj5Tx3OUaCVtifph8SvZ9KIsu5kzcY
bZI9dJt9daBy6DUuar3l58SlD3GWr+K+081NFd51D2dafmv8CUw93XVqSnqSD2OTekKteTOafrQS
+pmvcz5uk/4LkjV683K4/YCYMFtrpHlBxdmN70obA53aRdiQBKgtqbKI4I7kZp65ysRu/uROSIT4
S0Hpg61KaRLja4+t4LkIX4GBjOAsxkD8fjafwR3qTBT+UTX0wbaPnp0+nHktcl020ske6bAcJQ4H
48ZHYgr/2QpxMqArPn4RY3EJr/4tLcG/dNL2kcdB9Ur2Ydg/8ZIt4xr5D4yny9YkwU2aEga7YRUz
iEfiqhNKaCldachs/sMg6NjpGzfuiX7Lx2dEGoL/V3f+9zV/XNUxyCMjta+Y+19RDUYJXh6edcMi
iddNNZeYPsH5EJWiy84IMsbbw26g8Oynwp0MPFnpyaOdY8CEBkCYN8WFnyy5CVOGSGW9rniY0R9o
tpAhfPcTa1FXCmmCBfyh3pedIeKo6JrQQ4lNdx3zffNr/TlycoAkp08EuwMeokjKRoA2gFDgQgUQ
V22t21hoaN6MyfNPZdsEjFZ0SdkC0ZD1VfLvETCxWQ638BbC2IMwZnlaYWUPiexRtDqdSrvquYSt
/jJZ5cQFkVHTCaRiRiUkMsg+yG52oKjLO7kWkAqScSYtPPMOIQKkr7OV+g++sa9/6EuLk0dexJxM
/mNDUXQieTxVtjbWhGW85IOMTwUlMD6DKCZZCQnB6vDgOR41GgIUwN+7QUgIs+Q0yLciWQ7rmS1k
Pu9uyqtKHqF0mdyBLrcfOd06qqjtotkcZomnYnb1h+1YxaOpFgDfMIqajDSdgj0CBZfXo+L4uIGB
X7E0wE79bKN3kKWFsDX/RjcEHmUZ6XENQ201WF6ms4w5FWTxNVUBo5eiKhzykMhEHmMv1T+5Qh1l
JZ1Ii5uCj1LojvbArZDmilFfGHjUmrCF/6z9chy++enNWQoNbbX3Ue2OW8TDSRekNxxmzKGG9O3w
S6/3O+dZWAMtc59fAs5hwIcDRbWhLnUwemwJLc61zfMqD78Fw/oLRr8NYq0rKfcS9wB3+VA0AGxt
h0hI/yFN7LrJZboT+7wjlG2U0eHrwNbhWmrhKw794ZC8kdkkvEj3jLBJqiwFM0bR3kFPRx5DtIvK
gKfXrkPWohCaXi5wxRbQIaZrYgy31ncVcAqr++vMxwRoSSDQQJg3ZU8qkMkoDLHVG6XKzdgNYXN7
A4sh7uJ2wjDh0YY6eA7UYd4z8D+UYDh8uqc4bHviRvOmIQuChGOCsdCzky5z7RbtBjS3BFXIW8GA
ag/f9PFYOVS2fSpB6s0EPzjFGAIkF8J3si0FphiVOhfJh/ZhiF1gjkBC3KhWxPwu5C1IgyPmNxls
EmwAeIiwp0imRufayNxFPWM+uC73UCgZ5dvKi5u5c16P68gu6lasG0kQhZ1BKx+Hu+PHAPlesW0V
E8WBDJGvMmVpfLB/qARGpJWht211++5fpj80wEDfYzsNg3QkUgTln80rpbD+76wjvGDkfFcJTRB4
AicWzgxLdfRAT4AIF5qzl3J8fgzE7J2stqJW1SM6c54jZAxYjZQOzxn0GPXxGbG0Pt5annWVZcjB
U2yKqgZmMvRS+pv0Dfm63+PC4zwOz6tXTpQbj9kAXw2c7gbFIIVl6jgK1i8/q2zNa2WWi/CEwoHC
6yMFHF5+9/iijOP4ZruI/oMKCs2ohaZg/hG4F/jf9ucM6EFxrWNZjK5aeVbIKCCtTF08ox263PzT
DIaD6edYtkz88Z+2XAn2Jj/DzHX1bM4U+QLHHMxiBlQ6LLYuCGMDKh7JXC5jQsv1qqYczlILwMqS
sku8QKwu4aq8Ge9rs9jrI09AUJ+Lqv7wGqTECRW1HFoEzC+qdRogpcLzSh8/NaEuby8zujPRsEhd
fd2D/hbj0dJ/Dqr9Oc8zAMhq2SQkXilR+ek/NXCpMXW+nq+sWHBXXypwQpANp9sY9mKE4+skj1h7
D3KqtVIegGh15oFVPlZQD65Rvi2WgAjCfaIpL+/q7WYD6psTPgWsqvdItiC3TspZZ0DGGTXipf2t
R6QehzCY+aciaA4mpx13EB3EWlvTzw40/SeVusk1/3b1C2ab9Np0p0VXl87XMaHIpQHATSeo0eZa
3ma3QgnphPcq1M3gk+U774c2DpfniCNVYqd1lfiev5nmD9rKag3Sg3GpBJpVg4E37EbXS8EMwcIk
dUe2ul1Kd1bjPexHCuiG+617i5U7lgQVGevYUc+m4sMEAotCAwgMxLGqPx88LXirm//YwBk6CwAG
i09HdNGkB2YgSiZMWY1G+8vCjMEa/0utxifAOAdmk56gO65nlsiI+hn5RrXXPDwulTgwpByd9JzI
scQXa86wVpbSES445D9twtLpgh1Ag3tHnA9eAf8U9XsYp1BVsMn1JqsLeh5xKFXsdpMe791nNd7S
VjstADZKs2nJduNPwjOJ9S1JpoEbMiQWcbIk0/eRy6+ojloNQhYrIp/eLIXhX9ZXFjjojt/mwn9L
U0OFgt9HbuLByzqXZKcOLlY6ul8nj8eGDonGOUeppoDUioRRHk1b5G+a7Gs0ZeesTg3Lo0voN0w+
X2t6XD/pMn6hjECxJ1aFXzUwvVg/h4pplYHDn0ekNTSFcOsJeIql8juq41+UMTfoz8Rm9ODl/TIo
CErcRHMbWEiLHC0f8Plh8U/tR2hAUm8cCjeG4qH1O1Lps9XSDbgvy4ZWNwa3IG7RR2ueUSgulg+5
j/qRbzFP56xuLCVwxbmAKQVqbUCDUZRnBjMRFADbmlmYQMEpgnHdpVMB1F5sKsop3+egIkNbSlTp
s5hDXJj7BasEg7sIu2NL22yfeDVTap9PjdSsOQvmOoDmTdD+Xc+81gzVP1rjgQdMw6cMoQAZf0sK
7o+Ng7FoNbZw4Paq9/RXxWH+ufgAmVEOZXv9Og956hx6liJX5WiLsz0sRKhJ5Lf69LJVCAXBV6YL
6jyvxd7FBg3mLsJTpgXlfx7nY8N9uGPaFv+pQCOqoA5goji+PlpchYne+4+i7mTmrd83AGMjfzM5
BMewgqOv75o4j1fbse8kYRKXOsO68qVemoOyQJeOR/PBOarTJWaPksQmHlo9ya/SMx7QN7gLfCsR
qCdf4kE4fG51JVeFYXzzAwl8QwfGlHvYThiPTfibRpj+4De/cyZqKIPabFcXQ02Du61O2/aHU9qZ
Gn6Pxrk88Dq1PkBHttMMlbUXzhgG+9BPEoLve13ai+KwHkP1r+JyvWqDV7qQWpiOOPhgU0oWirfN
pynq74mD6PyI2/+XsA0/bpinDsaipet2aU/3XcPYUZNwr+yTmQUi3jSgPqPkIiDKzDqNRAvir7LT
jvBfoHW5VR0p0WWZuWNf+Le3AAW0cknSSgVs1uyAjeOLEm79QnyFnlBR499pRR3AQku53C2lS6/M
BetvFwGhHDkf7EedAy9VnrQo4yjSKBs6sHjYVMKiFqOc5HNGLEy9q8K+XVHLeMX2XfopPA1/k71T
ur64vOTWPYWACVUxdm9QWQ5w1PpaeMyD7u4WUgwU4pfzCY6vauL9zmUNQc1MMnJ/CSlrC+g0HajE
8XcQS/TVkf/TzdR170+gYfss2AoKORhqsYQzRnPlY9rvSUegnkWZpz9BRGme5IUIi0JpjUiTuFXD
X+dPxrXKyCYotY2D1s8l34KfBjCAqB76ZUuCm8RuDi72g0zi1dzaETRA96DPL7eDGnQWLdNvz3po
UsCKyPEgJPxDQsvP/BJcrWVP870HLKi0N1Lyo86lb0SeXqN5kZGRvtRSDxl1mdbW4U25HMFbj4a+
jdyWBLAsyqXP6z6MjuqS7MV7durPSaXm8proZcyxaq5UxQh7nLdousUOqkpOkany9K0SDr7TjHN9
8aR7RmFKNgki90bjWxSQoI7rRKjPgjgqZUESJWwKxhMb2HyeGCqQKZQESeDNUZcSKIU5kARHWKuH
oYRFTznmtXHa6EtKT1Gl9T+8IIFO+ONF6itQTr17/lAXyrf9SuaSK1Q/OWnvjkBhJT6M7obNDGSb
Xyoa+thcXepQ/KSId1uQkAz7IuN9/nE39Rrty2ECCNXOR+buIU4e4nXkFufEu/ibtqP+PTZlNHYc
Zd+LRv8JcmspzNxmonfy2WLQWqwUzXpor6s1+CHQe4pY2yJE+TcDnShibazhp0b9591CueabuMuR
QolEwywNVLQMh7xS9jZOhSKTXfUMV73WF/KRUAd7fSbU8+AF3zEu8Bg0MwTcAg5uBnDGM+KPG8Od
cG7rYIM9QO7olZoDHivf3zGNRzRUGnoOtQaLAuqtl9RvsSSkOK42XUyXfCINa8mxXENN1DMUQFdr
yQkeov7LKN9G+pb6cOMjrxOOAVFP31CUxtr6ZcFsu2kHxnTnhLIKw12x6eDXR0+L1qNi50pHrdns
9Snr20/WYOe7vS6yuCvAbfiRRpzNRC05lKzIBNzgEYlNDiH22ZVQlfURw9bXBGUA36zq40CCgHvn
D/PfR4nzcA3AonXlg5rNfpB2/+toSKsDPade/xO5CIo2t0mzXwzB7P6M+xbVK+q5ytKyiYWhEDuu
ylRMT5Tm9S1VzDW5UwHLC6oVO82QnHytMt9Mk8RChu95G1wSteMMSVxyAywcGcnznjxjJUQn+Iqa
bPOOsSXvFnLJAqHCCo+JamLrQLNU49MEfY6z2Af6856Sz2RnF3lv2j3oih/ksbF8cZ+KXr345N4J
g1i7DwfyI7FP/yrsb0mreODEdszXQCnrjvecngRn7zcV0oVwAvrVxsRN9DJXq/bc6hI9TTjLJJvj
jxriYDf8XbvhXfnzsJbc7tudHxIc1EIQoN+9UOOwGLQK7jVpJXxSEhJ/Djs3yxw2xaxUjDfJtx1g
79uhVUm6K++8uMplyyO4NE0H3QdQvLukESsxf62B7PJFhuVOptIn3k/u+MQCQ/2QXdpcMbMjzwah
SzWMsxD38WCpLfYkfYMx6Wl8FycbjqRgnEEleX6Dqh8AgqrTuAXx2nutAFKOOd2Titazc61NSFln
q+xTtZXQfAFzZ4HcEQo5Oap2sVY5N0Bz6hobTkeJ55MYAmPWVMei/TtNtRduek5JJ/Bif8YqgvfP
A4GwQKaKdVKMtpKZMb5ZElhNt3CRA3UqgmnaFKspNI05tuC9pHaxJDtmNvDvAcj74f8BU835x+2r
fbJ3Prexv0F67AcGtOLilNAcmzHtjI17MkxrdoVS4LvxjSrb8T6P7kSp7i1Q7pZwOFunTPOX9XJ5
xv63W79b/fkN+5oGeyB2HJ1anjj9wT5WJFKx69m4cA5zGzQ2J+Enasv+jYjkn3kKNJyGCpzQ/RPQ
aeX3p2QMiIhRmh77adPQRYiP+MW0OmCmDmP/hs5ilJe5LQsk+0nOXVkjmSHMUn/h4U3wsVE9dEYn
fmO3boE7vbSVEtwwocB1nivKqFcbpAHo/ouEbusQWNwihRh4od7aUSfZN9PcWkeumXpcn7poodMp
y/d2rEAzHRYBoSrOam2rOSZhgKvxLgp3usDlRIK9vYZ3y4jWpSKyOr2ntSdFP+zLNqQC6W35mNaQ
8ng94E5g0Oivuo8569GOCOjvMqqlxVNqthUPw6FDsxSrRBPbtf9+/Wvh6sewFkbgGhh9IoDYAT5c
vWDkRs87x99AwZ5x1hzpz7JYkVQ+vMzMmyXUYCUopmcxkcI5pC2+iE6O+cZoOTCnWYehMHlcMBdL
8BAI38VgrTn74TxQqNgZbp8ENohSgefYx5mmq4g6uUwBv1xqaE4BQMB8MaHtLbe4cVNp9oZecjlV
NV6+yjKnu/ZhtOeEh7tcAq+a4MzWFVUVxv9AMOlDQpGL39DX7gLH4Gz7+weMSmGyGQsJpfLN6IRD
jv7LwXyEesk9f91yKvxPJKFh//VUNvRx4P+A1jwjQ8nftCxoltoyNjC3BaZJzD9cuSRcqu3fRWT4
3vHTOGgiD+A1lfRB3yMtsdCr5pP5LS5p09sP4qGKYxjeCyg9THZoLGPXyzSzJJdfQiFJvAbIR9cZ
8yrcpD579sxgsNvyGc4H0Lvb5g/uC2Rbdi+hNV0/Qf+uOh8K8M/icKb4CMZwMr1C00K4gSjB4o8w
a4h20XNKCrnHti2cpO3ujNS1En+MyGA28W/ggLhNJlfe5soyGKe0N9w9mJyUBlVie6Qdu7f6ikgZ
rNxx6IP8FjLN927DEHVUkFO9z3vCDAbcQ9lzLLtr0HsT4c/Y3o81NI76hUE3Z6Zh2EVmwPNfHzRU
WzS+HcujEP9NovXi5JcXOhYylEful0mOzeFYxuN46g21VgeMuGEj2iW3lvgaH0y5J8a7307rIylE
C5q6vU7fEkDr/g/40BOYxCCgRmehRyTxiBfQijdIV33MRANZEBnyXAivmcAq2g4K6URKjAjnfMOH
+uMB0KDoawLV+w1fyDbPf9YmLT8F51ycNDrPb74UiO4rFIb1Mx8tOs8Zqrl13PpjImyacN8SXbsl
SEASHeV5mMYmbpGKRd79ZL2q7I0anb55ERyDGcESA7Wc/yWuKT0KLgbLQvYyDAswfnbTH55/sFGd
VZfYdVsLmXOhbD9WYDV9V/S18jsKEcAuRpqZYM94SlHmERsDnMVxhYpS/3xSZyEHc3xabBsnWNuS
N6pChXprcRF0AZsrGTaA89Hy3guF1iuOwRTWw90h5FKZUON0OdLfg9w/RSieltuQSr08t0dmxufV
bqO/pmtgoEtUwfpy42IKKOJsa+y0Wnuz8diyBX2kOZYbDHe8+sIdOnE4Rj45SYutq36sVGYinii5
1Z0IJOb8FiMRPEaK02inEcqaJ+tLEqMlrYiekSpEPsjmexzZakJStca3KqwQXBEDEhlO/7XErMwL
y1WT9K1CufFnJE1Zcv2LAWdyq1CLsSW0m25iqXLS8MojnChnTrbewkp5YCwqnxMLktGJ4579z+YE
KJbRZLXjSEMZd7OMvmAtDyAGojKrz/0ZJ60LA9k7UhenzLGewWPjJD3qv0Wrq0qtqOS+LoPJ3JP7
nIRF5SVIKDwjJtXVhXMcxU8E4EnTxsCMOhHARLxVF9j/X+bW7LGfhP1JA9laWl97mSRn24xJXPDl
8TMHHbWNKoceskfvBUMQ+MyeTGE5CF0I8CNwbBVHJ8ugbX70NjioqmUB5QFM7G7ImylpOjbhmIp8
DQgqwqTmoirpSKjPn8oiLCSa2WL7E0XWvKjmxEMrk/ZE5FUZa2wVM573gbHhiEAZerb6LdLQ4YQD
vzbpyi210n/3Y0Iol9moXnmFYgXTO2Lk1Wfc9byp4v+3fdDdWn4Fg1jxe2r/3y5L83K6J447DDpU
66IqtHwxLjcNnKXbL5PxIqlpqFEoNDCNqPv2WEqnl6OsoDvgo8hdespCjcDm3DrwJuBGFoZ2+vWg
Snk7BcZ2us2dqTjqOGKrSLQt/ZYNNStMPA8U1ltUcfJW2EgCEWlfBUhpBL/JavOxkPe0L4RKV8Nv
oF0NqACKJmNzWXoAzWWQ4JO9OvSYe+SxKrkURJVsx+UOOddmiMqxp5HZ1Oq3ntS8irzkQ2tJbNti
BVYz3Nax7HAoUBQ6dOtVdnHDWVjGmPOW5bMOQZPdKLXVvSJlec4MSI/XAnJNV9tgNh3MedBFp8mw
IrZG5FbA0tp3drvOBsbry1uUrKBlZJy4Hc6PV+LqooJi/H808RUNt9zU5Ncu362uMmQavUTp/N8U
xznWMUHFtplEMo7OegMJz/OSC/AzszORYmoZSpXjBn+VcmSPrkzwsyjlH8E9km3XmL31Nrld2551
pQWribd/GYAHwWz5xFFLbQh7BsrZYWeu33HC2v5fTtCy1L4QjHEMpEHdJMBIu8EcVxKJZGH4Mj4G
vx/C+yTZLsL+o/CPIjWZrNlihgvIrRA4IZomsrrtSv7BX9tvLAaO2SWVPsum308ZH7cdR79EBtcX
owRNOK5LHEA9wgfNw/Fjpqa4we3eHrjRKZ2A0rSONePFBNHJHcogfnnNXK5vfzYKLeGd7zbbO2XG
3opWV+6RRXBMM8Nabri6sALT3a0I8WfpxsT+0YW84/sU8AqMh4SHZzgSGyHnebJUeVBbelN/Qjqs
ZkaKoaw9veiI1SdG6ze2eVWWOUiHcMQVXGldgO1quIyiwnXIWNJi3cXAG5jarLa45cZeyK6sYXyS
IonUU+Un8Glrkjy+H6ynvGxTPjYVIK/glOGqR6FN3CFmWupvfLixZZqC+cuazJNm1QEpoK6FSXZG
Ste0tG6+059RBBkYnCbnts6W1rTlv3DsND9vT1ELFWfK8wgNwx7Um4KGjnkyysKgs2pUvUeoV/EA
Tpy93yf1viNmZuFuc2UAo+8R6sqo+LuTDJYdu0YxUmrqjbvjal2soETuST7HV4f2jvuYRS2VBkkX
F+USt054PYW/CgNaJXguG/iqDpNIVRD0iRxKC74/LeJkrqVmhkcvIki6GFY4JOxNJIV+YWwzOAqq
DnBvUWF4XBWPPnf1CgfrVyLPpBjvDFSyfva69sE6zD9PMf7h4WheOPfxCiZAQfeuiz4zkb0zRjHM
yis/YaRkbCFPTbsuV81eN7hTEN9VOsi6hNrwYGUecdBm4yxrYz/nsjvowP5kV27krQptuepqvnoL
pp33MIFo/tF4f43GbFXKauTeK25i5nACK1hHef9Rz1pEPulrFwpA/oH6BHfuQsZkJuIufPn45l8R
M7bPWvSpdA+oFkn9w5cN7q9BvQh1oKj5nsJqlo/UJC+Yr0UsiuZb0+Z14PTIlOB/KOb4LfXo8Nab
xDpFHWSs+TfWm7EEP9AK346e9HbIhf6lVDAKlF8/5GyQvsx0dRGvT66MhPwr2Zv60Q+iu6MpZeIk
PB5dSlMgyeJ9pm5t5jeD4jX5VW/Mj3/EwR63brdNLqBscpLH0pdsnDrmexiEac6R1b32etckt3oj
GHeHvOWNucKzR/lBvYPfMABMGxuajX48SYcM+MqO3FUwqLK6V+UfCGb5OkitlP0pHyXPoNlTPb3f
eeo6jXINXLzVyazf8JD0Qpkn2hMWeUz8QsYpmKhxTwwGYpx+xSEp4euCo/Lhq6P55pbc/xSHtHzv
0SEUqT8pmcwS/uigJLjjA50JQc8GBHGOz3QOTCGlLTuUlRLe5NzbM22yVIyGlTuyqZNM7MzLjv1C
0x60XybZ2DdbQTtMNlAHuWbJ4BfL1r3VtvGpJfNMmIRmCII07qXdw+wjkITVM4ZTGIX7R23kK/rC
pAZq8B9pSiktH8175k3FMNU+cQ6ISv8MphmwFjJdcEKWE6jPTHv0gpJ13pGnUERc+qxVVdC/bcwQ
nKCfiBQYMsfVqOaFrGvwesO2LjAj7dqE6SuDy57oOHnEQKgaxD5hsavulqGmu9O5CO3ZPNghCjd3
ZmJleZdz7HG0OJXRlPwY/XhUm7rZNhVF9pXklw7vmCnGF2znEt0KUHwGTGjWpQiGTUnzglNrU6Bf
GiDOYnbBtNiTHvjkLRTer79H8Lizj3vMIL3ibcUBruZXa4IM0oWOTJ0xAXOxhY9VczMyPphrjUoi
C2wX5c1zP2EOcIm9TT8EG2uPFwxNoKopOLmZLr7ITQxOYcboMWrK6PbO1UlWtvrtdXKdD6O/mSre
+YpRUA/p7zinAKTbtl5bhdn89HoAnlv6HQEryZJmHN0/msrofCo1Vm1jdCbjhKHwbHx9UegNIksW
AsaGHeoff7Qf61LQaPZBBVpC4Zb9ejlas2NOK+vQe47GXLi8/OnhIhFcEeM4kY8c6dYGti8/0gko
w4kk5BDRelhSmGDHRbSpSsunXEJOaEd30S1ZsF0wowcv2kBbEm787BnbY1I2139gyL5dSuYG9Ku1
NQEFotCC3bVtJIHec9NP+8uLzVWOgXlM5Op7LycTSZ6n3V5ZlzhK0p7MeBoxQk9aLRyg/2cOrY4n
CszOKbsNvv3lYFze5bhe6+grRjeMgh2BM7mRHW1/Yw+a5lYzWWzou+JOhp661J7btRSi8YWkaAXR
HyETv7B2zCBJYoDD2tQ/mHe3OuIe1eMIbmoXeLev1YVkFNByE7jTNxoBhz6t9U2vUu8f3pQwuaJg
k/eFL6yECppKW4tLkSb+nryNUfFJ2PDku0HrE/g7a3xThEoqR4b+qvaB4HRs9l23dIdkuGGaVhss
Umf6ocAZPv51RDkYxChAdX1J1+te742djevmv/sdHsXOcP9mhcydLAesXG5V7PKn6XnV6EcBAyIC
D5277fe9mR6+VT9WYpb/q6t2jZ/r3XNayzrOHi6s20vrfFHtAokBoVcGTx4n9eNtY8ehPcxLZSt/
KP28QhVTgZ31QClhhRu+2kyrBmwOXn0XRi5nul2eR88ujN6U4pGFHrbtwTgRVWWQB5K+q6yvDbes
Kt4G4lvpfhro8AfUbQX6xRAxDC07cF2sbQ1tGHPye5QqPkOH10eiQyGQ/pjQhX8m3tiG3YJW7scI
lI3a7VDUPc7dzJY3T/FLBXxDMIEU7LrAyoBHj+aDUu1/vHbA6Bd917C5BPqDisC1+XZhgE+yvk5n
IQheVsnddc3XgPMOufBjwPATfEqcxwDTkNYGkLGQ5yzo7H42wmASkstEPxqTR7BkpnlBX/stWbM3
iEGg6AG2OLVuPatx3AUoHoCGWWzVk5j166xEKtaiSsz77LVJNJYJzYOVhRVvbN8Ql47IRTNTxzvO
4WwtLQELk0zNaf0he1ch8uzvoIP8f2pvojjeGTopRucRj/HLyaLYxcfL0XVPhSY32wBYUjbUK2NK
rH1H+xAs5kn+RCBCE5eBcqwPtGRUFtWVsF4jNs93bONLoTCr4fzcgdfQcg9Avbah2yesqNGtMETd
utVDck2Gn9vF7vXACeJWNUmxWk2dJDcVoFUMPurFUkI+84n0nKsCQ5ejtjkGWMTdUwk8vAHsoCWs
kUZngTz+XxrD+hW2WwLMa2v74EhETq61ZG809dLNCy9mlti2FnXpIG9djlL+3Lvhdqr49UFBOnkQ
FdVhJydFG8Rw9SfcGULDamfJmkdveqFlJfpvP9fDIgWBH60YWt1B8VG5Ndb3d3r61LjT1UNDX1jr
RyqVw6RHFN0MFjQ1OD8LRXxBLKe7hqpOzhVsGRqNwj1D+Ap1Z3WFfsI0yOOA7TNL6PMSRPcxpP5P
JmEIfdk1nZ4YZwZC21SXrw62ALcmjbymnMMO8lcogjdO3BYrgMDW8nI/Bp9qddw7NYt542IHYwqg
qOJDeyjr0OzXmmmQIX4OlspccJBvOaBG0kIdJ3D1OJ6abhLOOpUetW5DqCxtMb6n5RF+2M9Ne6AO
Jz7gw25lWDfetMtScnZxJnkcPQ+QlPtJf/Qh4GF1URuqEPG8jCYhagnh6gaPXDQdLlDT/4EVf1Nn
Ek4/HJDAwfupitOwLUF0FKdhWNzMz7Uwu2w7xQFRfxVV6739uzbA1pcznc2vdmKb5LNNx/hEkouX
N6VdpmPTWxrfEqg0iOoTVbYtUluHJGenv/q//FVKga/z5Q8nXbMtwmMAtVTkIWB6g39kMLBcfStr
odIRNaTgHxDCYkbqhcOCa7hBLq8/G0mNmL1SFCuShq/WnWmmoT4yIw0OrGsBeIAJJKdWImuugRWQ
Mlp9JK0b0v07OiALDRzrZoxD4zK7bc/VnvyjUIAtcTZzSKRkT5j8G0dhfdbB/rh+Ri0gf+u6ZxkH
kzmtM21J/4KvX36JU2Iho7bI2YZbrr7wu1lI4/JnBOBogUEWZhiGIdmlXInJL09bjYhJQ8+DAmtq
UkEM8ZSWGXi1brjSXTLMekCO3XvSXG0zG4iEJYSTMkTs/jwXFkzDddTOiMzlGP1g7CD1o57YZWQn
9OGTPTDNdvHN7wcZEf7EYF/gIGBUY0i2FM9aX9gitMT6tYUcsfK66kx3EtePbdjnKFmERFH3R2C0
XS7zwVQ1HKWY32Bqh5sBXTbYxAB7d4lDhzROb5ekqJW+0sxe5dCI5Ylcd0Q9W3598qCaq+keGAgl
Hls/8of6Vdm0yeeZbbbXVNqAzGFFC13SJD3NvG+lPBC0JIp3uRBRSrp19IKaU+t7mki5u/Yu1r1w
261cTJM4c7nPb+LVFTGPpXzLIrvcfu+na9ak2REcFcSAsC7YEENjzRke5NZQNPvQH08Mu6vbXfiX
ku8vsRu8vEuCqSahoVRJJxHaXbiceLjrTYJqrBueBzP7DY8kDtDZLO3vzHehz3vkwgRJm7p5Md8k
KjlJzh+wv4izpODec3ab03+PA+yA2x15ADeafIxeTyzkNeOQmZ+9s1C0KZf5Ntl2rVkeetvXcKgw
aO7mRDchufNjYwkP/5NQ+tFn7o4NGdKqOxEBXEOTZCsXMUU7hyjnqv13tMsKi7xu5pbNxZsdYglN
YPpYO2Btt9wJNcWToCKywsQ9a77dKLhyZ6b5EOx0FIofOXZ2ZWUQPbv1HT/p0pB+nQYWIcuKZS3A
g/vmplPhLVuFC5g3Ld0UfIAfmjRbOtE1ZygYONLb/6lHkmwazsQdPiDdQ7lzSWgQ+3Zv4RAxpQSM
8QF0jiRnN2BS/8kbHim2v4V92eTQUYSuMvzAOaDKA2moSKJGZ4VxK6jbWA91CxziRB75l8RUwX7v
j1AKgmBznry8rPgJvyI2oSwodeEp958WQb+DKH810T9mC/VbXy8sM32DVM29TAL6DjntZp/rXBbA
/AruT/MIaU6KYqYeoUKLLiAKVAP2YzExxkf9WWyDaFi+iE9f8Y/HJXIqQEvRhIB5oX81nfI5iv8b
peyNob8tH8ptz9mYxZfT/3HNCH2TVd3a23wp9V2BI45LojxfT9OdJIvVR6CJFhR3OCOvvnhn8goq
6IsqYYi5B64pH3ojEOHYIyGoxbOXL/VZ2lt5dYGRRB6jstUJAxuB9xmYPX8/+1aHVG+I7UHTf5rO
kBBM27S1vzs9yZcVOtIDcZc2XgSonSDPgKzGB1HE3Bt8m7EHsl1Jl22JqJrtD1QLhHK8pNccZ2eF
kxNxws5Bg6f+OJysJFPRKrEI+Tf3NriSmse6Mu39B8KL/06tgJtGaDwMjOoSKc0ODzpP++LtwTD4
VyviwMMyS6rKGl2JXOMF1phx4x8ukf2wRhNSY4xjIga6wflpCudxemnt5eVkL2VdSUnLCpoMfK9n
V9/cTaW0L/SRCnEMokxCZCInJ7gCvOWdhzFcnG02JwJ6Tl65vytUgiNUricUR+A3DWHo52IskVfj
lAZphcqRbOC9Dqrm1cThSuaFnv9Rix+V49m3EZBLDL//avAZxQwUs6eyDHJ17+tZqxIfzUEG79sY
OV+VYna4+EFD3FmQmWWxUHqbSRbWG4lgWF3oA+DzZnUU4qHhXGrj9eTaBiqKxhBbEnIFwNxYsMlV
qTcIbJf7y6/KD9kmxm/uhu5pfffAu85QE1y2KZczP1VlD2ZY0gs5+a6YTObAOpRUC3ICP+HGhwIE
Je6zSLZ+BhsdWiPjiwHGF1J9u73//JyDarSnX38T/nYbzg3i1xqiCd3Uy4HXbFkToorBa21ZdQaM
3ohD9Dg9tLp8ZLL5K4nVyQAp10rPugtl2osomTFxviWJ61yJRFvwIZrAQhNacVeC9dg5Yk2rhxy4
8p2IvpBxCFMocg0lItlYbvQiZuXn1NAL/7fUs2dYdpnzb77Iqv/EF0tgU9IJm0x6jcAVJA1Jwy44
h3CZKVfKVXHJTHfD6/kGvvHFRp5SCgdb9QCoPYdbuuqIuCmd/kJRRh2dUt5dq1QOk0bBLSwAe30p
k2iZzeiee3SqxyAbPhgd4hA15svcM4vPE2yS2n+rwxFVzmLnnTzr14Yj+e33cMNhttMC3Q9MU2ng
M5PK7GdGAiSN05XZ4ZPAMdCdiiQaLW8TPeLR8cMpyTW9jKCBb8gVOw6cJfiIvH6ixgFImcCGeHbV
H2P3pyPXnXSbcOzqd3JpDzXS22ozVCxPS9DSTdiLCTsVQ73Z7z3O8hIJFs7CtE0VnnIRPjPlMghK
MkLtA4VegyLr+Pidqn6HpqrQdSf6S68wjqkyQnXWGtNlcQLoiOhbJzEm0XWuMvhKZMUF6ksLTOB8
ykk+gyT1UMQ6bHOW9hYiYIcd0jAEpQ3Hp6jTzTvahvzpQuGbPF0wVaOYAjyF/aryuOAmr32j4TEk
5jza53+dnphMfXPt2ub7ZM8ni4WejkXF6gLDM/W9PKHKvy3ak1MlfDC0bn5io27Z+/oozaCB2gEz
X50OHJAALNe/2oUuIRqbcgobNkqyIrKISRQNIaxsrIO1+se8H3T73je1uXgx6m7gLKW9mWwxgSw4
Z+aXTJNgm0w4C2vFOrjMd7trztmkFVp0dBWZtCHMfxZtz8s7VLF2jlQNdzPeBCRbD8QmOKtRZVNA
6WosFtG5FL0S2Ic2vXh9hciW4RGV6++eQTk6welWyf447Sk4duZ3C9x5FTMns9FnLlZ5EITS7GMA
SJkKK/c0AuNi+B9Y+mIJr8mHvTsGTNb0b8hJzpkVM5IYpMEPencFZL7EpIS31Fe+EdS/jk7JJgxx
TsRIyCa6y2kWxTJgbYXFN9HJeCyfV63mHAY7lk8NomGmIgvWkp+eSEyjuHgQSQcsibC/DNo8lqTC
Ym6TIBjLQK+4rVbRoQ0EfueyquWRVskzp0V7woJ4RAigpkZ8Ln4CzmJuR0fkgA09h+WTkekgaeO5
zToS5qUMjd1fKr6SxIkwfn3qyzPKZWwJcCTFChUujESSqeqFu+TfdIWjWE5Ocn0dqNJTsFlfg4pQ
X76UludsmnCN/gnK2GDXnnobIeUwQM3UrXeOiq4+dipWfMW9I2kez6oHPmm1+vC3iwy5UzvmgbG0
vcN34dQPNPasWgb289Vat0QUZX/3EXK4BSPgsPohJm58HyL9zaFLc8AIojv91gpXTVogR5wx4LI9
CU8/rHzaNRLwhmoo4vVxKau1zwJSdA0xmjToaWjfZ6rPg1rDr4zlSMbW0YZt6NazMKMVdscnynk2
YduDqs5+asjDHIuZR4HJmhW2V+nmywIide3OR5nyX9Yjrmz1/8NjlOvTO+aESAC0WXZGnn+1NsZS
HJ7ei5umxeORem2F1kzsoJaWgiOifLOYQbKE/SEaEhxGaegdFOxn01lFyb2WLBTMVvzc3DHy34vK
k1Q3hEI2DiJ5lx/TdpoT3DhBgUQ2oo9JeV2Qu4D2KKlU88glrkmYfiWYMV3E5+JDPARmiKEBBOJ1
S6lZIBTO7+eUq9EswyMa6ziyVLmGkyeMtfuanjH7jgLYbHfEdjM1B1OBbpsqOJyE8bg6cv04q50L
7R6vXXlSnsGE8u3B6hGmrn6P+rgrk/ZSOKD9M6UDuPY0e/csTmg+Z3kckwGO125AxqNHJ+mEUuP3
3DnCrIs66yXi4ZV21bSDBfPu/w0FjDnpOdTPpEByDQiV7J++3Hzeu9o9dg4p+XWXsk9nxc4CzHyi
ut5J9uQIcBimgITNkOgBmX2Pp2Prn1NRHKMbRhFcitV9Zw9Jn/hBUDh2nDvEgI9fjzFPIQShR68j
2+nZrgfMC0/YaVv7OZUFlJXFLTWs28FbhXx4wjprEplt7JZHmqOF6lr8gAOtRTR62/xSrzgG+bR4
GM21+4l2XrYFuOU9MQF528/LQ5kv6dTSThSNfL33asokrGYBw2GQRF5zALMTdwZElw6xICYYfmpu
B7WZ3UHg8YILXsT6AK8h1VtVIae3BBzqJ6hXsP0qOg9Y+xXtjfOKse3fMCGwWMGjit6Cr8TqArMb
m//dHCYosaRPoMj/7KlPn9Pw6ziRVdnPvtlQoXf33LC3SH182etHbWhGeZsmkL+lRS7+rDcHPIAl
N3Cv+QpauAAQn3xXtvvcB6TrR9InG0RpqYQR+WQokAtYV4u3ME5t+mUn5SjLsu8RUvkVxv1FfedF
HvDSrrXZvksrtxsBYsBWejJ0MGDbzNDrTOlcfDgQSg+sqLQeNJQ4hg3TiqBmm/ubNUR+nW9kGXgF
ix1PI4maVcSqcImE7aW8QdRCWL2VcYTEwu6lYlSRMwdzz6KjiKBhmoDSTelKWxbCAgJYz9WJe7gM
a48DUDArmYsAT9hhitJn+N68QXIdjEgV3cKItQAtJJuiaf+FITvkH9fJKqF3qM9v1GzaFgY17Un0
BBJ4twzBvqz+g3QCmPDcw0MPlKUdSX9QG6BbJ3y1sP4riJuJ16qaAsxgGKOqjsYrCmve4EUavmYL
BCtdvrlQ5n2W/RTLoCdpDVnpCWDQ6lyJcwy71DLykLT+5mKY4uJn2+hNLIWoymZ1WzsxqBejLFIF
+1difAs7FHiZ4JMQ6lqYNZt5vCga0CGODc35dioz/DL3wVbmmN78LvqzWpFnsVY08f4KHqz+51se
FgxlQ8ox7qqv9zJWI18xwrBZC+yYE4yl4vkia8KFfYXhGYBEGyVnkyfebOslNQ+1kIHDVHY3pZ8f
bh0u1Zv5nAJXJ6rvPCCsHew16ILBl9yxJKOP1RfkS1YmOm4IVtArH64Bf5V3hPoWl9Sp3l4RVy6/
vAcYLg/ow1XbPSwr5k6b50jpIHnNKwa6la09x9K8Gs1/VH/66QhMQZnYsAIe/RQbvyJtwjfll80k
PCPoxwDppJi1DYbPPII+65TLRNs2bZleWZ8ISg0wccLw9XsPHUxZAkFQUkKGR2GBmIo7RQE0LA8P
bu95GI3bsfCupmJqffaw04NiB+0u/U51AIQ+JiQ3ACoVl0tyDRaCRSMV3IM5s50Arduv7BHUi1aN
p3SrKlbTnBGaMTo9NYyT77z7ycwHjfLpQ3Tlx/OYs3DvdrjLlhg71mhra2/BmUpMwXbnU86j8R9s
qEhxzWyoDpq7zCFpiX7rn9EU2fTp+CQdkYWb3c7xg6+/j3P+HezM7ZBSvpfIk7dyPhhcDRQgXpux
8wBy5oJVVsUnpzKJ9PjRs81GaxLpVfYlIXSKpBG1WK/9A5ZrVRb6dRR+Ip17hfr60ae+O3otzZht
2LTuRcWg+KAEQxJPbls6uMNj31nehty7CJZywkT3MuEl0BEnaONzdRnrvBmeOddH+fn1HCgl1LU3
GaHSvC7wxmw2iKo2iu9kC96+UzgUGNkGnwQFXVM7AlRJ83Z/zpARQ4j+uei5wmw2xhFCtodEt+41
K/ZwQTLzD7UusgPsXY5hiU5l8XoIgjYM3R/9zOBgl9Ed61pWbLOLP+fB3GNeqdBRsFExFyXEmJBn
recv5942Q/pNAcRtrPu8/F0VRA2CfyYJOGk5vbb/pvF2gm6jvCxs8R58K13KhiRP+NYkW3DgmgmE
R6hlAkW4NLh0Mb5j/7dJy3/OLrjG2vJ535dSAhxYJwpxeval3COjT+zvqkfQW78KjDbRZL+o3ynJ
1jp+zP+G3gHLq0cEYHDrT/AxC19rnXGGPEUjH2VhXKMNivBSCvIVKKtwGz40lEsfZQtLb8GH6cRd
HhYvjSMfCXJXYjVsuzyJChiinc8pjxedtosTeZ5BbHl8uxyWTxDjeDmehSaAaZXGgm7WtP5eSm7Z
heUkal4llbTKemLrApWowcuNHydzRDqZYQEJAEKczQtdDR/GoNgM6Oopa5k88KPeOd1c47mT/8T9
+qA/7FkTFVa8WV/PSQnVljWehDys2RIjuLhvjUBJC6MbPBmZx3SqMQxDXlGbbBYssZMr2ZE1KmgI
i4QWikDh4Ue7pU/RqGWcWn4ZJnM8YeaGhDYFOGf7CsbvAqdNsmPjYE22sO54ETGJuJTnLV9bLa0N
QjLy3UkXBo1ZnjEgRXdcn3C/rRPlxD5LSqy6HeO15/jaLnNVPUEdMRidUw161BQeYj6MuYGMrf2u
do5jk9TDdiiR2557BMk+r3ENw6z/rL6JuNIyCtrZOafXgK9x91bwXHOqD4xy4y54GaiMLP8i4sEI
7XeUxLXVe8HsDP+WTu6TiA4eDo0v74AyQ3eRnXfjR0ESnR//+oZWBrO5D4oqJD44UqjM5ilfFDrL
+wilYCI6HFdBWugbPXzmvrBsCTnxOVDvUa2S9nJKZyCYnMHTcsvtrBBj1IP7gShGAFn0kEezkdXc
yYOjrd0DKYnQJxl5RPffKpCWiXg5Fg4f1X1j58505jV8copEZfBwUIt071AZJQ1x8fnRxptn+4/G
b53n9rvxe+wrQQtaNoOsQQxlVKs6VKIMWGmQh3Ti8M6+lA49P0sk937zE5MmtSS52eCHqiLgiPX1
7d15BWv4IcY1YOlv794mVgOzGOBhf6eG5Ha5RLKetxQo/UmefKb3UXgZWPREs7CMNCs0qHb6NjwE
rGdLYWAi1nZ/wpPPhmvx4x83f8OzsKpjZOlH55anJPJ0dM2KSa/MlL+XAIQf0GR8g+w8uqWV5Frw
tpL7dd53FDhkAuCSB1Yg+SbVSfonT4Neqv02GyxhrvK3t5nr/6PWFZfWb5NsOfc2Z1I4WpozZxIa
bgXbKmJ/X2HD980kAUClHPrjOSQ1wmf+IGryCSX1MU5rX8CCNAXWHfyC1pgZOGt9Rnpd6pRCSO4K
6bND0/xV1Ei6mVCZvL4ThZe0ywfZ17LSEh9nLc+vl9lUmZ8agWuvNQi297VDfdQLoDIfO5qGGUNc
64OdOdn5Dsec8EltXTW2knypZ+XiOzoUEe/6rfesyz8qOKGRPGpFmPdD9C5E8NKcU+97K2tnmXhY
N4g4NDrHGHAQ+O3ahkN0LYV6s1uUguav+4jqZ29oAaQxLlMe95i85+nzT1Sw/x36riNV5gh9YfJo
RutoP+IP2ZzNyQVwsbTWczpG/LsKznW72JSv6DdIF0inOh0MW8Gg10lcZhuMDQnrna25Ak/wfh0N
uyNYafier228kJr0rkBbrSUsY8xCxfA/yaHT/pmRlRRpHosy3JkESoUFbpOKKvoF55uvkgomJcSf
eUIVZBNVIwCMdDjuBttU8iS8uOcWJV3hmfW7L1D11ivmlbZcHdVp+jdGGEZZge+NaJn8DR3GyvfZ
B2TKqmczx1c9XGVxns0MX2F9SKM5kcB1DlBQBFGydatw/Cxa6MS2RT/jXx6QIlrw6qLWBISw9uyU
7DvsiJyFkjtWAwDTIf8JltRGc6qNHMkLpbBjqkauV2GZWqqw80PIgTRnLttcoF7muP+c7S0iq99A
rIwGt0WzBx5yZfsRpcxvD8E0775czUcQWrDthsIifXRKITSNFoZzqv4/naekBWbfKiuBcQz05z2x
slug9qLPJth1J+UU69h8Z17gzpeDLJugb8XC12jRGv45uH/XEO/qSy9NfktEKlLw0YhYA7Rq8eZ6
nTUK5xiGF5DB/DJspzdxfOSeb4xyAB9SmDyvhUHPaAdcfMlQOnPIJVtLjuMBlyXVxVwC9r4bNpW2
fdJ2DofYFtNHuN7p2+03njsp6LeUCBU9+iRIftgKRdeFMe8B1zuv0O23i3U9Xw0hRq8hsEzZ45NF
ybdKY1gdu1H6rEHKSK8vQg0FegEyH1q6NxKcvTD0p/0FOhg6SatPHONFRMhuh6KmQiJVaOnkr2wm
4gZYlO9585NVFPEvvIHRSN+brgPPMSXyVjNFGmYlw94SRT3knQmNw7BaVfVXaF2RcRPbyGd/gl6R
I5JSmlyY80TmiQZridrNMTP8YF3v5cq2ae4jiDRxJrST4sFg/bPwm0j1GB2rV/4iR213ejhct8LW
3x5ozoVPaa4nv1AyFaypyd7sMxWZTjzz4ttod0q3LM3hHyucKzD6Ci0eFulUpVSz5lW/X66mc+fJ
G5LfS6C0li+XT6JyHEHOWDiKNCBH3Qo72S7NryoIGUmXV+QlMLkadwOurV8IFCvuVEHhrk8XDW5f
5CJwTddavoRPU6oZJxolqLuaDjvOmyJ7IU37NQiw5VjS2AEKg227LbOabqjjJ22jgwtzyE4/dLyv
amvbFem2XRa/RvOe1GLztAPmLEV2xBQljkkU//p7+p2VqQLCM/kTN2+hN05tpdN86M31Dpw5VS/u
GEcpXxI4g8vQSioVgp6ikEUaVKJzx+qD3B72caRZPFYEAd7MAiNp8pW2XS9dC2U+qQK3UnhBAua+
BS8vdxBhp3mENmmOkDc3jdyB7QYZwmesnUhIceq8nOMRG8F+lFiUCLtUfNUo40H3dloi/rmezLFV
xbCsPXCDZINjL/4ZELkvV+njPZBNrhdIZ7XECLVInt39i+wd1lSgNFrjM2c9vIXrSLI7G+FmeqC9
6jKFZGuldMLo4NejCLYcQe/7RgxNAcrLqJapes9Ret1Iml4OqCIDeUWbozLFD3H/6/UoZKZ1IHwC
up7HFW2zdpYf2ssoGfXO/c+Zs5NqmsHLR8h5X4af9fTIKFNGHa7Yl7SVu7ZuQsDf+GbnxEkwkwMJ
MvyGLkDGpYvYFpdcuhtOzmPmlbmJlyx/WzofBvoZFOS6ae0M2QmExbQIRP38HW2CKgC15J1Gpn8O
v/8qCWqgsyBANqB30CuEKTMeFjSv10DMYKeqGbgQ314E0IRERnCuUnByKDFVO+FgSJhIW58lBsms
76ZeyLGqbvPeKwZJjbU4iES70SNiJOkyG2DYZ8QsYboZU4rjMprnzZFk16xHumsQd4JsB84PRjRS
lH50y/zz/h8mDYD1j37KmKI5lTioSOXaMCc4eTeoRWFG8zWwgrz3lEOXxQ+anGeXuCfH2zq+0dG4
A9TQyAxvGWmILBMPxYAbhso9+LBugCrgPvvsAhmQyjf8xweU6J6ZlfEamTJTxAXGlC4fFgpHmreU
VLFt5t/Vg8ULsrwt1EMaYCbZzvuQFE1axb1uYxwTk94N8GLFJE/vVEnyacmQmQ1CSA5P9SMMNwtK
9NNYxstfbBad+PSupgdYZn6PtLQ8ZSDZU0Uh/VKuBQyOTR0AK0cmGcXjbdoQkSfUpg4Nzs3nnWxZ
YaJzTJ1aNENgVBrrSQUC0EFMfbTTRsn6l+30pgr9h/zqN5VuuKCTeJZC/uzii0Xzzz8Pho+ezWwV
DsJv8XMLFs5MhGtogHQX06GwfR018mhRT9gzIu9ZIDo7LGJyvXsF2IJAn79w2pyTQUIXlruzn5Om
zVO3HJwwxB1sqxz4tQ9a3lxgb0wYs3yXWUJsGXHWPnpdWuz0vuWaqZlquGKhK1bZYPxmZcEMl3R1
55vfszhFHSmKNqlUmKBdBw50aHkQbEPZ0VXaKhpOUPowegfqUdEmcplsn77iBc0pf/OciextdoyI
ZWaN1mj6VdDyCQK3wjavK7MEs3pulINpaLifU2T9KOnsXPNKE/mq5wh6SZZCu3qdFZaD/oHIzRWn
DKkGU9L+dxRfZZpgAfkYiQo1Xo+4TjMO/2XcizxWM/6rvMMpYfh1+y2TB6TxHpzeEFomcQ6Z251Q
Cp7+8e5bdbf8gmm1j2wIzGZ+XMP7MDBwNMfC0MCnMqCXcLWtB7a28/YrXB9/8JgP8sT6CJjvl/M4
8himaDDGqRLpk+QBgoxTStbmy4XfbGuL6v9ylA3lIID1db7Aqt+PwOm2mValMjz1UkOp4HGWAWWy
2MmIzEZPyKMB9EixOkQTimgKPSNtaIwTrKmaq2DJzaH0yb+P4JpLNmah905xdp2eKGZtN3qRB5/m
nRZSVVNOHCKPJCRPO0cXmImceBOs9kenZP6qI+1THt2Kc0I4l3GBYyYyfmGYI2tGVs1fZJVK1GoH
xD/8jY3GD9eMFTjr/7qSuO2a6XEcbzYie/nAbfDvhaTU8KjlTXNJzTs6VGXtkvaXUm/eN5+ZAc6E
MXDqXdLZUwLu3fbWL7krmPGKF6ELryvZU37Hw2yRlwozXqRRBSWDhT3BqIioCJfe3SBF/JOn9JPW
q8RwUFswUve7IkZp3IlyPvbeC0FZ1MBw2Ht2oeif350lQVqftRRX77zQbdw+82AYOGH8bDbxPxXQ
wJBhCeqU1JOvGLifL54EW6Dl3B6EGGpO3NRe4ZSTKRj7qS9Kp9SVKAF4RR6yfpspjU9BtV7Hux7Q
kSp99neNqhxLqjM3WKpRPEnCQOTwgzOTw/92GV3qG5g+gCnd4vxtDWrbF7waJsdYlPF7T1/pcvNo
PMf2pkXyS06Sq2RH04Xm1+33EnUQRdh8OkhqzqKGwD8T/vcYcNZ2jY7HlnU34X+RgeYIFQhbL6Nf
z82pVWwNmDM5Q7a3LAtCMaqqJL07HtIx9MjmwxXl7fYTTGPS5yvaPzFUhFg00h/Ts7U7tJJt16bI
/xDhWpDkQoDTiZWjdSQh3gUm0e1Syo1sd79Y7kcN6iN5rZq6vFOxP3p+fJNL/5iKNxNeLFkhrCpw
xzG0jz9iT8hnXuY9gLPbRpNxAZmL9sbND6+yetH0m6xQZZKMlqV0hotd9N7AV1gmMe2RA6YRUiDr
RvdF/1AFR7coJCw9/1wxT4ZMQBdK/H300LPEw5bJPWJnCjcV+cd7hCM56YJynkmSqkVc1idXgpjl
Ps2eyRYJuyaAT8Q6iMrv8i7mutgpjda9SE6e4sQzHc0tuhXPA+ejRUY8qe0qXOI5a/0t++E8mfJU
vNtLUFb0UfKelx/WSqUvwYFF3VJUWpivaGYgoR24ncbXq/KK/P5JUjE/sg8juDuk0lc8wSZ53zlK
nLFpTM/VUYyroWRgqjvQIsNPV2g0QRthQOHiLSqYVXsF6DaBWbDHzuT5bnquHvwAdUBkjCK5oGhM
P0OB/MklbajWmTbtk+ZNYaKiglgoRdr2t3keNJmQxs2OPGXvHd0RU/kbNtzB5DjMkpkB7wfVCRBm
XyXDa0N34W1+Lizhd4so+UmVcw578H1GCBMT/JiOuIst3muwISEAkHRKMFrIq2ano/eRYGXndwDW
Zq3z8MCnTRbrCMnwp0nftfT8F+rdCcivQ1FQGqQ/KWCdxJwmNOtISD4Z9V0Jcw3VifwdwWTRbHVn
7/a8MyYzO4xSXDkWtGc1hx1HqKyDHMVxtkCzBRdCVPbUlJ5CAfKiEbLCKvjP1Wkx2GZE5ygDEocA
aKC4Li65nVJ7ktATKfmXRgeQMmnPyUxuYAD64+E6+u7E28wi+nQx6cG+roL2iVl1bIE+TDpjXbde
JoIgzTu5Xe7qOUXAjNmkSDWv5UNhhud8StvZOLo/OOZW+5CtZfbrPKnUfodRTFurTQrYC2nWV9uB
ZmT6YvCb+glrWtnmIWlI7JtxJGIy5YpUFn77IyTq3OBtb6XLcc7X8ij1Ft9trMGzeXPrYzFQJ9vE
3bOBJEAXdqo2z5NHp3eBsBdDNe7EBcx2Z+D14OFaGBwkKIprYeMQxSgXz+9faxJSXKmWQdcEfBEu
NNtGDpmFpVsFz8sHeUyeXoaGkK49Uz7HaxFj59ql6XcnVW975KPnPAybFpNcpMAI86xhlQJZQmX1
QGmaVkW4yKmH4usLrs/m4zrcIrwXlHf6KJpb7RqAw1B8ocUj+GDpRavfWruQpBRADjvwhd+Gr+ea
uQBuTiUbPjI8ekvjEifjwONvED6ZZhGqyz/PBnxxxYc0X298ATkxhWQpP8ZEoAXK/NxzsFJHNOjy
JdyjdYx5oyK65gGqWwlk4Yk/2KpyctzYa0haBOwHLv6jb6HZzcxcwWPOKGLEYDjMBoFGNVn6SAXP
rJpagC1jjGh/f7O3hAzzS0B8KML1Ox99hvQCzAndgzKzIKpcrvBy9qzkK3UGYk72yfBDq5I/WnUR
uYW15LAzS9/wFsp2fsxKnH3FU+b+UuBFbcVF8eSXl3qU4P0fxdc7lVi9kvSk4J05YiikdX6GfZ1H
lwqz0AKcOXd+SGSThBgj7+FISOGw8SaJCJcYafAEhJKFCJxV/enYHc0X5dx4lCjpobtxBl1PXhdK
70pf7JStsbgT+RH4H7qtcojvosR6hugAGgUVEasSXU9xlwCfjpfMaDJRC6tYMqukv9+SnTSIAc30
lUllHP5A+CVr9py+mvr67HW6/cpfT1w3DzcEzfOa1LnctmTNl3K4o9MpbvUvxPrRJ1VRlaRO1u0f
1sr7DjvB1/p5pegKGtXkMFP05ZmlONxMCCTKS12Y+FVwMHQ2F+MX9eemyjOVqJZjVZlJe/zcxxkd
Lh80uW3MrBhhDHKxjJuMOVZ9Tw9NbWlyLCRd3wkK+rX7aONTCRbl9hfeVQ0UiBcLrzSr7BMmg5Gw
YFJpQkdMU3DVN/m70aSvhVW3deLqpQ3OhUIY+8A3M9ov5Be06TKc9lk3gmjG0eZvdTwdH0gfKrKu
9F5x/9G8WeVxNDUJbhO5q+ZA9iztPreCflgP2QQM0tvkLBvPfz19OLD7HGl3FFWzAEfs/l1QuqyG
+dWVaq/+GkttYuvGKU0k8NygJcgPxiayjCI1yVBFjL9C5/dCT2xBxwCzSYmfp1X6Cw+5VoA9Ai2y
m8Tke7XniZXs/dM2mMmKFs78jhlmXFFoUilUmswbeXHFDLtiuiSPzWPhRSH11DNI5iSomxBFu3mE
hR3ioypl8MrF5OvcyldnjN9QEs/7ECHyIqrqtNmG83n0uv3CPpXm+BxN5nNECgCckeCDIoBCPJeG
VNpnyjGX6cVXHbk5VXhVbKwmR2WQJBxZJf+WT7x781C/7cIybdpKJ9JahrXKavAOS/1dg0Y3jJQ0
uti4wCgVv4fT3AvePBogizPrsdxRNzhAGWmoP45rIFST7J6iFujZtEYmXXWYtnzRmQGlzIi7oEj5
TRhNGpGfkyAdcroucuE5kRAf9rb0VHm7FMuAyQA1vBk9OFvjTmVYPLFrru86ucxLwN9U/uaOJZz4
/+hUn7eVpP29knDVBIEWGQwEkLDSF7xRJsu5+RGkxpQ6gNP75dh844xsl/uD0RanjIFADzEYg7ne
L5xJwlqMxLnOBl3V8IfRJL0LbEBxaVpoTaORHgg2Out2/NbaPWjsR1vz8D87OTeat3ugP/r0D8HS
3ciRPcYWNPenFw8psuTk2OWMydl4hBR3l2givOvFGmH4nYQTzMToYRw1NSk7kVhwwoxBAWg4ZRZN
fSj7hrdiq3fwmZfoLsCjkZIxVMLORjAFWXcApqj2iOZRCNYqjzzxzdSJl6ca587K9Rz6daHjeCBM
RrWOuGiJCr51uMmqhcGWZyDNzWuCp19tkZctA2NdAraycKKFqe5XU57xKH4NdGsk2ddo8jDTCCZJ
lHpsJvYYLtO08tIo8TSKEDkTrDwDiRWdeSp4IKpXS3tfBSu22d5hluKTaPu+hZVeA8vczJ+sSn8/
UcMmCvduN33hDh/fBScsuD1coI6ARlJ3M2ZXJp6OHelmZ/Co6jZdtnoDGA+OYmFHOITYBPtT0e+g
iTTX2MSAyW5O7rTL6t3ByBxgNzHTX9VGijHlNFnfauEqV+BxguJlxiugGFBfZKr3iEFk+LNBhrHz
FHGShHErm2auW5PG/MEBsPT1JGYLb/mpIq8QSYNEte2V0Sa5jOl78dZUS/sk2ott07g751jw9Fzr
YXijdlyt5ux0oe/MdIGizW1WBzmzKNDihcu2DuCfqJeDl8b07tjqliE5p2/ylQQa6uGzn8nIPkX/
8TuQ6Wlx5/7yf9Bwn0gf7DeE+HJOHQNqqkAcVmBq/hqvbO3HSAW8gXUXdW33C09/Kox3UncZ7aEJ
ubYGb36XsuiU+fMA3z64tsfv8uOEqSsYbHuNhmTOPdwLKKAE2B88NgH1VOjWInNuuwp1h/B8cwpP
LFlZ0pKqF5aeqi/A8FEn2ZKny7tUjaF/l7LIa9akcJdFr+fh4iWjl3zyyRwbDSvUfz/acetAMLfM
6sRc0o6hjaF4RNdcGwOz6hZYJ8QIu92KMZms/DCySFJ143/dJI/9Pd922rclnGT1KUVzt43gQzyT
abaxqZqQOj2o59+MtOflpgCjdRvtoaA6M4NFzcdbcDengrymJ1mDpnL3quB+NXagEqlLyssxZAt+
xiomK4uWMciN8nkKsPxSLRChwYRUwI5ubimYj/OZyFnduE7sgGaMcbcSAsNaFRle8z6nA/cRwDBe
zj3fP1S0Jxcs2EMgo4ZwYj+3CZxQ744P/0Cq65u1lRDWrQn0IGtpaWUP7dVSnvPCKQG2ysb1VZT3
i3yP3VfHTYXdmFq/fTChHMVUlP1O/44NO3lYr8ZKXx/paY2WT6/xm+fMxuL3UTYDWXPUcSHLSOx2
fCxrIwf5apsrX8W8C4MV1VOpf/qfy72DHOONfAc9GFCLFb7hoeL2HlgDqcAve8UKPNv412FfGh6g
55mXcSkIFyv8vG8pdPLXN314fOMJKWxAC2LHU3ME+vTlyhJtylcapTLNBt+z8AFVzEIamsbLWd85
v0bC4kGJ98WSHInE8oSFW+byZ3X7VQjFe1XYne9nbvW0ZDhzjiFYHu3OXQIJ2Z5Mn4rZcik8QBuu
pdDtKxfJ8vyPjbr6f8eJ5edtxboRRsXpCBf3ihtW27S60ILuK/rtnjyGYl5WVr03I4L5ycS/5ELt
8NlQql4D3ORujzNLgPhpVYxNXNS+62pAGEUORr/bBsQ8+sNJGshj8eaniArRg1D/bG+0xsd2CvMU
6uuSY3jnoc0Gg5B6CVapdtv5ssI0bfwwAVRcmodkIjFaRzuawa7icXUhlKuhSkf93lYB8ym1H/zk
Vwe7NwHXi0QUl1w0D3peYO9Av3N2gHIFtG4A3Ynhy6SKhKDiTI0Zolg6Jg7ui+P/uDxwYfzI+gg+
DS4FFXCI/vT2TOODYswTT1TToXjAUPZBmvCHfO0npO1VjoZh2TXwxPV5g/cNt16cxmJaQa+nvjiT
8xg/DAAe0L2NKVDOTM1D+0T8Ly8hhWnvNZVHi3SNfAI8XbVLODwZ4+R3Wzagw34ttZMmL1LyMxGt
VvpG8IeqF4IJ0KGSC0zb2VQEnvoE5bKp3MyguldGSnyIYfUCrxuAolt9WpfTX7s42OZh59eicaK/
V7pzrZp5VgeN9NXWy/rbqnGKA2gsMErsIOjPu/x44Pg5iUHZ2lkGMfTmD6ncc6u1eHnrrbMY+Won
DkwiHZl1L3/dWPgJFiswQ+R+W1UbPY7NVuZ8pvIkrWU756ibd9c++fs8o6QbKGHLsSbRSFjBIxeV
BFPVU5V6rZBcHrLdkIPJaez/ow5t6mFHE6XmDZz3AJMWrfuCe4BefcFEQUXo5Ff/Hr35pstx1Of6
Yu/JwUGSQ0sAngXe9oyyK1kDtkC26KWRzXj9Qpwrzj8TOCdAL7kKTbMu2e1xGe+mFGv1iDu/GcA/
/1LJPS7RtriOqQ9uyHKIaU9MJ5/NOhGD7Vb+htoDUTgNK3khtDMvd3taLc4doMAhWyieG2TJ0EtK
cWGV/ho4BDau5anqbYrKa4cNj97nrZsS3b3VMOktKXUx/OjThuGqUlxRR/pfcD2HdQDbgC0EYe+3
bYBJZ9Q9jB10unBYPFoyTH5QIiZhjEKw1rHhWk7W5LLVfZQMQ4mIw5n5uFNEh8jF4G/54UXM/uHs
ctIflrpMulzlqAtyMX/IPdnCT6Pz/51FQ1FAAqSV/MLoHr9ZzSgFgsgHAHGKyanUTlDEnI6t0bBA
SSCDj5kkBXlcKFLw+XOs6/f0ZSx0UurKqQMMwDbvm5WGNoMU7P87uErcKooWlGZoIUpxEqnOSIWd
2EoDFAKEXjEBDWRn87eOOGXca9j++SlenkDmrBk+Al9bj6GP5Nof8siRPm65tlU3my4kzPjbJ+N/
CJAKTeK+CP/0xTyC0xy7/VVo8+QTqefj4g9pXC6Qbx4UfQMhkiQlGoWPPJb5lM/ZVp5dSn35t8EY
C2Q24qiAMMKCKClX8Thf5MdIqG30rFFJqmSnR7i1B2MIgUxqlFYxXeun0OqoOxtmbr4Mk1J5H/s8
9oEG7/HSGFHdlbvB/DCcIOCx9gmodV/t+Q7QMEKuYSm+fd/4aJWgebMDMi9IyUfxkwnJUcVStNdR
SgRDM+G41DpRA6FjtRyRt8ZeoU42hqaMJh+aLyr3mslSeY0C8R1i89oGOMWhTpaWJ8fySlXVtkBQ
pX9ebtS7rJhIrOn9gLiGnT5Mhnl5nlzDtjSinhnpa4uzrnNkzc3G1akpEgQ4muG8G3bAuSbXhxjJ
flr9erbJZ3RwiFA0JKF67QI4rtGGdaflFfO0NHzxfxtYI7EbAXtzXrjNNCG3NeyAsBrB0Efkd7sh
PkdC9feT1VpJ9jwLqOVDsboC3rcargbFMtEsQihxf+Uxpsk+q/c2kA5SYTwW4Ta7GcSh1EP1If77
bDX5Nm+SdbaM2M27FmWX/W+3rvLE5X1CragM9QjcUc4cLS3rdpMQ80SJzkz6Y3jJaVl0NqhjBGAm
MNf6NHGq+Tq0XFzqo1SHOXnMu244aJSe5vV5UiHeHI2lP2cd+t2/B45P7mcGphin/ygtvoEnXNn2
2ezJrMIG42HysrcjJDlU0gTVOKgse3K/3UMKmLIb5IeUE58olFxpEchyDyh/MVawU4hi4oTJS73G
zm8hGpTBCeVB1E2SoTD5RA3j7Z8oOgcGVuVXHyHLLuqAChXaBtOo4Yv5RoNcx0mb1ADY2weZLZQ3
xGvD3N486lva+z4CVsPBf3FQLHYvJMtA5qtISw8feOC+vFyvl/u/5meAK/92TC2OiC+51bMNlHhO
yfpjmREsYMHB9rD1RvD6Rl7qEu/F1TqG/yWZJC6CSGmxr7KyUcoNHQhghIlinLQt8xFlIS9l3hPi
+zX0/DLaZG2V/hOo+jEf5sgNT0q5bB4UU0XNTtqjV4yaseZXLFr6kTVh+9066lalwRbH1G2ldCwC
KjDYP4gX50JZ4i78rCplWcfGIxMxNTTTcDUaa1fgq2QpmmSBKgrM1dwt4vs+vSc3hTyFHwMdFOfJ
CCiXcTRjJgoyptyaNN8C7soF2HjD+x/uZAJ5kSpWl2ttaigotI0B9Wo48jcKgD6iE2bbr9BV/koD
Aks2X325pEZegkqnRSlGzsOmWCaB0eqAWd8N0crmjmRqX86EVOvObI7b/767CqLL6Bs0AtwmXQQH
Ny38JO9Fx3kbefbw3UA1ztYchBBsjKxQ917qB6SCf5dJhSJu/D5KBJmjQ2OWc5vbreTFaheEIBhQ
D/lmK3EwEkOwIrCIOBIZOjmMPZhWvTgU+zmH1SQMmGx/KnP4CmBr3qrwPiBzk8AW4QoMFtARNV/9
xlFTDj3nJlTlVN8766XzCzYa6N1+97OA253i0ccWYHj+bWs9WIqZjQQmjKDzNhz8vypeELcatZ7e
ZesBBXgIj6lKVt+F2uw3wOh9Tu4RBDHQrXH4hz1p5ZbisCdoBh6RMQdBSiZ8J/lggDd2XgRPW5Qj
4u1LU4qnOUDalSF4Ntj8gFfJ2xOaFdAlHGfvXYn0jxiHbHiijwoaxPMjtJN8PP+rAKqMJEzvdf0Z
1IrdNxiJtMrMD2ko53fKJP4QbAiNWAd6EoCso37AiKGQsNtiFrJE2ZnQIQZU/WfEImEaJl9NdtiQ
mtb0hFVdsmiwZmYDMgtuKO7x/zCxhFC24pti7z9xsElc3iUCsyXMNmRA9WW/TM+CPiFhaA1mkdbI
ZvH/l6XYzoLhcT82WB3s1qmn5yi3SoOSiYpqb8hTxKdQ4xc7eANGldcqSmY7eClk+IGx2xONrcE4
9G9PQ9G4AzPJl812KMDvP3aEAQuTDH9X/UqEIIP5nbIZTjVulne+9UZiERqxQ6sp98GRZkVXrdFr
ErdXb2JNCNz/U1kM2wrnokldPqxymkwL9RBZqgKiqj2PG1v18KtyP89XryXEjo27ocdwY6k5SeN3
yrdEOK27qgvUwr+SQp+EiyIXAAKoXilgZUtbcwu0++XeEGH+TUeGmhIl09DTz7pvPkdkiHcomXe+
BOhKpjVtSAZFQL1+6d+TgIN2It4FFRNCWfaeEN/849G/jvK04JPjNPTpQ+mKejODXEjzMWZIHjd0
dCVMERL32S63xsJNhX2loYqqM6T36Mk8is4uGCL10f5bqzqW08mnBFDpheI8TaY/yr++8WjgmCCv
D/fzA73afcpzpvNl+DcdYZ6/sYtUZPwy89DFPXJ19/9d39UTnE99kEY9DVfK6Ny+qFen7+rxgqGx
6PcavjY2Osw3HYTPOOc63GeSoaQcNSILgsrxVbODmtZfAw8l71tsjldYIJjiFrEjbMh/3VDeuWdN
wgFdjX2DsDMLjV7yhZ0MsJCkuH5HAnxTscpjtrTjn3jMOr0mplF+DeLXEDUP/oxny43oS+MAS/KW
P2KgPhncNZj+fqI1cur8fcdlQ9tVU6f9EXi2jj5OWUqWTHOUXin2M0tH4HVpmmiLMD09J64Fh9K5
XU56JkhTYVTdyKLvTzAowTigeOK2XsNjdAMAS5fzBjzil0e+U+9sVLUtSmHF8UY6GoJpKtNiYmei
xAu3uZO1UqwCtqC+ly9D2ooXzt29DMU8TjrD+4tHonO9vNUkEsxYqur09ZjpP3xaAW7JhMzb+5Qv
8foYmppFkO4TcxQZGAFZuDDAOdo2YAHwHLz1Kng6LhSfIW1d1imozBxJQ/nHKNX7KXEfTMWThvbq
x4lYp9OGpRz5M9Fxspsscfwe2+EHEGGWS2bpM3Kb71AmnPYSaMQzp+iTC2zl5fNZn1/WL5kORbqH
e0sIbI901XRxgaValvDz6CMlLCbZ+CPTq4SOIEudPgQghA+FewlGbk6v0fI7x+6JiaDYKVuUT9Ib
uVbvVZDDnpmKUNsXS+q1ivvTeWYU3SFdTXwqVyiTqXD1b7n0xOpnnHrKWmEmKqnBkP2hmIrSGzuw
jVPnsQDH0NeTySodEWSLCXIfC4/ar3y+RPknV9BcNumnIQi8zM8C3efsB4UYzNAVPILkoHfnBO0r
VGBhte0ZishrLXUhTa0WxbOlTwfk/M6iSeYMhvPC98miX2bQl9BKtR6SRCYUAH1cWtctUN+EREHe
1Rj/AFsDl3VVH61mscnzYYVQJnEgwH4d7+J6pFPjycRVqUuRRX4bCod2G8KmHvc0K0QgBu6YvCjH
txLSeqRsRoDL59nx9KcNzc5qJRL5mP29xjoc2J/3pqZrdK3UOKjbTYj1/VZPXD6eigvFPICxXMIz
1ykmQ3ocLfgmkZKV6jDMrc4Fe/ot/SM6fF1gfv6+PwYkQhG/LZn0oeO8JFF9nONy9Jms0YOTxxGS
KJNSb3Il606ObGBRquQ207oVDsq0TsiirF8V9xirxYEeTgi8IrdkUFYTnpgOBP2OAPmFDYRtHkRL
7RcCby1GA/KGzq85QZeX5JnoXJKPe3tC7GODuyMQ/thfgkcPGX6CZgRZ2zDRIZZAJhF4cnV2dvh2
NIpo7lsbXIPSEerkrWeJvl9PnMh6wzDgyCwJbaUp2MDKHhSBVyNIgYnYxVcrvnp/sDtNj7grqvV4
g7x38nBtsHnWcONCkHDao1BuJ9byphOftD56Ygb5mi1kS91FUmcxtiG6wXS374KxXYXHSKWGAmWo
HXKZgfdGv2uSrFyGJ127gXIwMRoEXWajfBI4yrNh/MbOnruqHuBz6fCcEYNE78VMVmAzEv51z0bu
SbXcv6BDsDZR0yLS/tKEuHMgRGuEkV7Dc5Cge72GvPRTVA9vyXxRavWvfnGLnXwDuGxyUFOZn3/p
meSO+GeyGMAiNYqpEZeorhsSfyHX4RC+DFXSO+vaahuzhyh7ZB8zsQB4gqyOtzbq/JfePSAUShJu
9o/grO7Dp0O9Yu4G/KEs8gwiZWQhGzfpJr307aDjlxGhrY05N36zdA2G2DyupRKz86CkeTkH0FnO
4UJ+rkePLSbcINCWejbbnC2B5/ZqaXeAB4z5Pf3qjN4F8ibBpmAJ8b0IJVU31oZChCrNAvnmmfZ0
omyXQD5soqG03wpD1PyTMWfTjdHQn62RLTuziBams8lSm+L1nZKmombOM1QXnAOCXIZgvUdrBpm0
ytxuYuVSflELb4p2HJPppQvIAdXoi6EUI19ikylw0iYpKSoIVpYkBHTFu4//GbUFLLhPgBg+d3m9
iyTc2U5ZQuLoDgPJSqOF5edm102cnUEj01wDncq3eNn9eOvRawG514rYcNiK4lOwT3Dwq79NXIWe
2QdqnZ+idjxTt4NpLa6v6CeT3Om9TBWSwPt7m8Tf0vr8iSbYz6mi822mA2aCCwVwOZpe1+UiQQ0P
Chag1UxsB8F11fG+2FJQbKT9aekrBjVbjDcjYa8oYbDNYUWsSpXjYCur3jnRvm2jl39XtGKJHyzl
5rzfMoZ9zr6Oh4gEjHZhNyzc6VBUimuzK3esUgESshd6gqN2Jvv0zxoYGsPyK5oZC+HFP2Hz9IGh
MVdIKaJe8eVu7bVUfxa1Z8jnf+29hJdS5R0hmKJ3hDzSsC/RCvLqnhjcwgfz90a/j5F+TC3cEVTW
2BolarEC31iqavKAOK8ECOenQxca8bLhmX0S7Tq4/j/Te8D58CXWn1sKPOw/Q2/cKPLul3O+pvbj
hydc4EAsQbmZ7MOQMepTYkYnqjskLLyQvqLyvGQS6hFygW8mFLd24Kz7tq01JyocHUSy1j+rfL/L
Qhi5LDqevPkwMcRMWbtH9Z6pDW/IZctfhY8E6yImhNGMdcUGfCdEm0DDqv/VlllbIGtDufWAsrkv
g/YUoB53VIhbBUGD+KLjPVR7M899Ho3hOnue9l6qO9wIQ6lipby2vqbCLhEwwqtFGkhQQLsd3Mhj
2w0UBPErmSLN/GIphbUpUxpFQft2GEZopTVnHjNeeQpotNcueg8gqFr52tgbCu5Fjm9BZ82Ov8Gg
9vGY0O1+52ROZ9657CboDr7SwjpXenCBOrxWN7vgum2+vZ35dn3cq4o8HyVHgeYHdgtTKJ8tjxpi
7VRqaK5F3RRHnXCCIi3ISz1BOtx9TtyKwZ4PHdXBCbnb3mcurEWwa9176RUNlB1Lu2tNQXYEx4ar
FZPYwnNg4at8K1rZH2f7ToAoOiiGZ56Wn5r14Dus1mQYwP/1Owqo3rf1CbbTtK2pDfo18dF82FLW
J95jmbCVRpmFFPZhsh5R39vj/EU26gyWIv1YcMAk5NsJ+CKo0Xjjb1fOENzDZtm9CrNgRD9eQQUW
t0HGvXazN7fLpPgv6zWON27Iw00UcvjzgFRqmhEJoj2EnDfMKofglC2ZM8x4s7H0JrRL5Moas2sb
GWHuO1pCCpu+aLjOYBV+XDfJak97euytyRrGU0oUSp9+xZrsbvzjkjkGpZ0FqmraXm9rJ2kCYlex
PH/VAYtz4rNuE0lNR/mZU7hTnQhurUPa8IDr6VWVRJbHkqwlC8ZJRFUPvLGSnYKrxqT2dxUuhEJv
Lyt9YEyy/ayuFl8CXM5YO92OwY6fArMUvmBhr92zik1XVeGElw0gnPr1tCRbZuDHw51NvyO9OBib
qjcBJlKr0cgR+prR5CaCUI9ZK1ga591uUZQwL7BwpUmGz+YsB72chZ87RqcZxc6YwG2bq3nXvDOS
ZDHcAIfqGxGRbWavC/xiL1S/XakXS10dKuE982PJBe6cdXT8bsdz8rJVsSUflOtTZAaBK0U3Jf1p
fjHXdnm4vpEdlapGg0ii/XI3rtQwRcPn/7PIf1Dq6Qa2/ZmlL0F0nhuT5kE3I5zE4hUflObfyVr8
wxygRp2vdUeA9OweMi7NDccsXOttuN5n3v3crLypmE2w8CWBrjA3FhGyAfK7PK6LErqViDrl4zmy
eTjtVd9qxbWkfIhdwPFLVNtcsDZNspV9aW6hCLRuiAry6qod5Mj0SyQkeszAJZWMDZ5rdehftpBJ
PobJ6eBueeaPfbdRjKVnTxOIXca07uFE15ORYXb3NCnHkGQmL7r0FK57pBDN+J8SGTkrPbQE6im+
l2qwYPCODyVG/gRo4YFYe1E4gUc9Y2IDjSDpRtET2YoqsBjaCrWFN7NaIb3vlsVhx1plUSi4AULW
X+kalsxfDr29Oc6N73G3vm2wq5mtfK2PeqFvVY0nXK1C1ML0HK2NUSCXwEQaU+lzcvM0JeAUrYWh
CAXcTX6LbJlpiSjO9O5X1yimb5vRJzCbpcycN0CKsKdIm13DS29lacD+x9v+oGf/XRTd1teJE5MB
o7E4ig4izNPk7wWwR9q8s+h8A0rV7DLGtWD8mbo+q2e+gfTOrmqMt2Io9RHMPyYfKCZHKJhfWcMi
fK3pDlEL963Y85MXJNCyeT115QO/xHDpQ2f7/V7+g19yJbZ38xDv2pW0LSSWsmJ94z+aTP63pRxQ
xYMQFgo/uy+cfQirQICwwncJ63RbY9QWPoK+VWbx377yp2Df/BfTlq44lXWkZ4DfR3venBzhKwKY
UuVEYk2vRjvTC1n4QE2QST/ztMT5LAdJrBjAdPx2hZx9MUKIQExlbwV6+480LxgaUlcKz5anPuvO
gQRPx3uUU2Lkip5Xblb/MmhwrCDGLGurLSoXjYcQlmkQygtMJhABzQRZE7BbkUzLpo1xmzt7+E2s
heThIZhs0HWfP3JLJoAtMQI+uUawD1aM3CJVqzAiV7pzkKo4DRa8oDS4UTPWRsFc79pjDhRhc8KH
gvj7auOJgoyzNecs10kmJzPLx+xl0qhcPzB3c0z8i2HDJv+ejXpoTG2fOIb6+v+WojRXhZobp94A
k4ARQb4+VLDfocaXiZE3SYkBjrm79OmLPWwQbCof65XvSs7u8FD4q3sLtv2YLhO268jCGVkXwRK1
jkLayJnzKJ3YhlNV/f83B4s1JtAA0oA1nngMcwV9iLxb73C43Q+EF7O7NYJZa5706ogZbCzqdbjn
BLfqFfkAkYuMRz5CStnG+HUQ4umVWeSsIZRDm9QApwVZNbIRqbyRIcPlK7VFrElvK6GcoRlHdDpO
C82STw87CXRK8GC3Fo8bEHO7I7xW0xWloaUPDTYAkgeDogRGlp7nLc1B8+/YJn5DKRgEZULOY9bg
yF6gV5pMphdF4cjamkUTvizIdjzAAuG3TupXpc/iwZ1uN9+AlMWejeMbNfQlCfFhR1DlvKg2iAqo
/GaoybuWjAkvNbf/2G+j0RsBEpJQcuqVOnqWrveP7YBqUwM4I6X1gqmWeXF74XKZdPqofgNklqTN
suX3ot4zkYwLOCFtlKLJfOglAzmTqKO2tqNwEWPW7gXKgrUDc58Po6YMLeIpQlusXlrSGK66zW6F
imUc1LEazMBxKJlcvFV8HlfaLdgcq/64obj6GQSKIuuvreGEAO0pS2kIJcKHamP9mmSZO6iNL6zL
HBtZUlff6Mdyg3DOBowSAZjTSydgS3H3MYCCW/dkgw9hLW4Jhur4NrMega5YVJTHloz3ZWG+K6Tr
4ytw18QlNYM3W6KY9V/ptC7cDXxnMwFh4ufdm06PWiNMLgmuhFQ9YWeOYvjN6cx/kMHm6vLNbyAx
ZZ6hTbTpFjYGXhJz+BNOaw9g3+JnAaPb/ZjpWvo60jEnopEGsFaOGuRgLijeUlS2gCKnl6uo7/SW
sjNXKQ9PKU+roAVvGkTILu1WmozYZqR5m6XtBjiCXJ3vbYxAepRsuTYd/INGOevxu5U6rfOGWDdn
YcGBIez704x+GpdxEligcdgYGWBmn3DjAf+lr8lAYg7UwgaCvvhzrK68QyM9fEM1UDFLMbPof1Oo
bhSXqN1tpqk3+YgJKxf0WPSM9V5qxkZS7nXshTmKsdnWgz2Vg18mkN/jcCP2sPLdzOoAy2ZOCnjf
fXB167rB/pmFWCs6UQqlZr4nWgDNWZhEe3K8pcWJ+I+AErqkF0gCIgG6AJgl2gI2ucQhpEvTKNiN
UIyleJcAGDP1x61eolOod6O+ffR4jhLxUiL3YdR/tStMT2TTu27zwIgrCv3nYvfJxu9VOQebsKoB
y4dWNGLdNb1l21Uh8PAEjW+nvZ0sXvSO6Cu5afIOqwNnh9ARf1Swe3byPpU+lHjZVL6DR6oQLPav
yI+PCFDY6fvgy/iW0eT9ENgMeZgIJ9knDPFA9/KsY5sH5PBS55fPumPA2HNRCo64gL6e3pOT8214
I+91IdLNfhNhBPcJXvxunFFM74YazKX17opejf3My9n7qCBBhUxL1nBULQGK0AC9ZW4hH8D1F26C
0AE7jdhTmdFrmtCuBuVPeNB+YS6SfvTzFbbrS1H2RCgkbgLhVQam9M6A1J6ilDQdWOWyyX0bPNm8
EyBdILIdIoJEao5XWzDuRjBaH/DiCpRenOUa9eOB6yx9PK6m4g6yzaY77scP2/PCrrFOUIqjq1XB
zOltojzQOpM4zVjfs4gAQ1mBaMikcBtaGMEE1aU3DshmKDpAd3h3sacYYv5d9edx+IC0PzFLL6BJ
Slv9Tqqc2cK6/RLApe2WlVvuxHPm6+yT87KlPcokDu8T8qWIq7FOdF1cQboX0tNh+WfR0Q6ihN/6
4a/YKjDv57mGA0x+xG0xxlnMAwAn9kgnkC7kGFGKYGRTNeSyaMUAUBlAJMzvr9fB0Be3tQKoKPrC
t/O73lEZRi3fzvquGXrUtqtb/OVuOK2ArOELNqsimzSQtM4O5l+R9DliYB5xwD8/S6D/ApCGBxmj
a3iK5PS0DKXFVQlyymf2dGKrgRRVByS+v6w+TCqsBQ23s0vhS+ICGQGSDJUsZII62nSR4vKLQmxS
2VJY1ZhjG99y4I+3TZf/vPFRbdpjloFFj9Kx/w/zwkXaMILABjyGBTv0MCwNhqKr+9OzUpdpNZQl
/SwTs0aLn1GNtMNT19wZ/zeXP0yxlQrJhCVI/DBcLBuBLRYyRux9QtYcLfM+tB0wVvXojnv2ucgP
1UuQmBvJGW87d/LhBjXXAIeXnB2czVJS0+VS0R95tYAPl4RJtQnwIopV46Yc0LS1scun+J4Qab88
SV55bcm9C+StY5UlUH/fuuWdazco/TMbavx0aPUulF5WklNtHm0BXz9s/pWSqRkS8AZkivDtcU30
A0DeARhzDRiTleI5qZFqfV/jc6/AZcvUZTgfIJzLWQyEGIipxCjUrAfgL18HPw0oEuWLY3fcssxt
NQ8Uxcnz71Dnk1ev3YMDpty0pbwC6U9BnBxBBsGYtZ3M3tYtQNwW5jwwLMB9gPOSHn2nih3C9oEz
oKN9DlMUFnRERzBTZawTnegn6FqqrDMHfGmCh+/OaQicK7oTxD7SDvxE90Z4dSrJt6T055k6GMYh
cc+5w8RbnyrQr6jRSZOnrqFwZoZItI3JzTqycSWjKIfEH37Y5ArJaUh6GfZZeW7hY6mQZyjwUtbw
klsTicd9uNKDY46TmwEL8zkDiV/CQcYnwOVDcBlPsbRiLU40+U0Df0i/vrfZvoCbGKh9+KKyCoFb
Y9AIWJ4MwkyW5s/mXHeC7o7F42VcPEqUyxoR7ufsc/ieVtDWYbtX51MdKVxrSrJmem0L4Z7GCRK2
25M9rnSH0VjsWsiDjJKDRRrocARnLs/NhlzAj5PWAYbsf+uSrMFt8uidQLyyz1lr/hT4z13ACN7n
XaEj4aesK72BBXKVbVAFARq3b3yeru0i8luH4/2UxKMjIWt6oFVYcYgK9Z0t6kBQg9wIoSdkgkJG
AFeGXm63qMj9udcYcav5ojEZArznPapXJoqiwepfiIzMLchekhimqVasqjb1ya+aZTZ3GPpM+Wqs
exKaSzwoTZjk7UhUFI9wnLEDfzIssZQXrxupmZiQ3hWo2P10Ye4WvlGpySoZ2mZcOSEimDb2PEeE
9FWadPLigLaFe2KYa7DqE5cgeWk2H3LX6sVmS65yT2748G54Rr+TRYoZvEol+4Fd9BjP/xdmTobG
AjSgK+HLFF6vo9DthIz9kFUh/E86lJppTHZ16IXfDQXFBPKJ2ReYYr0DHL/0LASXXLhfpcLXrPOM
phK5YFD/9BwU0e00xhzr0+EB/mndIkzBC9WXfjHZ838ZlKsxxcY9HDYhzTeHxESOLHJoq/FfhlT/
1gA+MviueAFZmye+FKhRrGVixDbEXeUzKwNQ66C2wIXFnIze5CI/d0VAetR5wI3lusZe5U7B5s/i
5Q4Q+FQkaPbroMMoOSZAORW7qeHarC/aO3i8kClK/G0d8UhfgXifAnT8BYcYuSRmM2SFsBYRdMeN
R85u2aWbOr2kIezHtMKyuoxaQC3q3/Y16h1Cc/LZpgIH7OhFVevaZpEzR+eiTFdQjDpqd6tAejjs
RzBg5hxc9B6T2sWfSdnSFqAVGOHKEwZ1W0o8OqH4A9mflekGJ3erAAz4e33eNYqW1Use4PKj5uoM
Gt/CYlEL+vHm0xRzh5n2LeZZ2KkBQCFjsc/4ZwHGEwj2ltRE4XPs76oURPbMmORxENoP5E+o8H7j
oBgTEZJlytG2tK7/eaP997a/0QXF84VwdC+ArgKdTD5TL5TGreokHk2/8U2C0h702eLBHnHdEMcz
qZ7r82tAnFGdq48pubzxtVI+k3O2gAaVqASU+71eqI4wKaNbA9xp8cOY7aXuc5bLCJCFA37DnOVD
JoUa6FiikTMZse9DHZTm6K8SqBiPqWYjdUpIR+EpG0MGdyuzocE8WJSQuuzINDB7ki8mq4AFdti2
OBwm5RV5sZZtzDLgjfvxOLAahoh2Ozz78cBpprcY8WTahGkKw6g0Y5ESReJD/cki3Go2NZOjdH5w
AnjNDZNPL/rXNMcCmNQTK5Aa0cPwniQTbVxAyMK7gAoJcNCl6Twqx2ZpT9G+0Z2sz22U3b4/w8QT
xpt3v3uCk27Eti/2/8DobgCpu4iG/Mwa3vBGKs7HCjpo0R0DIZ0afhUlt+XtURaIRPYmpYAJn+oy
vpIwog/6lZGG7RK4jjZ6wFUkfi+Zphr5k3KecXb799SUoxV3+0psqD6oc30xVjth9ZGjejtCmRUI
K4ixXYKo/Vos+zt+X4CsnXAydy9BbQ1Bl8y6eWUU+G/ue6LEASAWn176YMYxynA5fm6lI1V4ubei
BnPK5sFS8eddilPErrYafTny2/Kvy/k8r+WCQnWAgioc5Wy0b+c5M+wLFx1rA+/jZ9w9CHEXaCZh
gaEc+zpLOgg98kKPGVYa2VxgLyD1V6MlTaZUE3WDpagpDrg9h6Y9PAUIY+rFtq+fgA4xresj3GDL
grWcNdFTmuufXBWOgz1n/3sEM66PsC19bRL4ZXAeRBnZ62HsCp/YJ4Z/UiIF+Q1mbcVqZJA92I1z
R69fUHNXja6uyz2enkGqTtR96lGAheHp9NmawNiM4INuDs64EVap9ZQykY4OJDjG0idysZo8NCIS
a2Hizl8a2dgGJtFfYXY+aLrcsHTFy3s/Y13GA/FuylwV+ZpFzIfGUlf61UPkoDgUkNqnCpekpHDl
EVXDoLqwyY8x23nnpclKSrlRryITmfpalomghZBGLrNCq4s8PN5FEYdfOHxEFM4v8hARmQTcllnH
Lq0Pn3pd8QETSRM9ozxs+r4RJ/h5CfKJeb8NJEpzmJVJ81V4bDp4Iru6j+mejJGYnDjZg0UJR5RN
Vd76BrohD/cWZYaGIq5TOyC7ChKifSQOEi2bZUlTIUAvrgYvN/3WBFYFvTEk4NRcfCdb0m7mF90N
NyiF5MNDDYdr5mEWv6nvTFQ35faMWb3rmI6Wm1DEgFRftC+pvzNUmSN4z0OiHxRLkefWSj+LCuNm
nC67hXZYk+x01kF4ZiWZJ11H1oHWQl+opaC73v/wtKUMJt0yDId7F2OgR2ea+2lNd+TwywQhPOg2
yHJhMwERYErgJVWo5vBgzF1WfrOrABHBbKG7vEkRT8UDSpBQ1rFCuzt7WseBh7dQDFhtFSLFBB9z
B3dLV4ANaWIw7aQXR8dgCVW0pA1I3Pt27UrFdTX6XFqW5anVFj03f5RBPz0l/D3TeZWSHLGRixja
bwCgPJfxl1Uli531Ghx5Wn5s3q5fiYysdNGrFk/e/+YpOlp2bH6VxZqIzchsiru9nwn7w5yVb1qB
ReUWhWJJmBk9+XRiz8+46YzTK5syxSV7KflpB/M3QaSXvtts5OoSJ9JV/CaUylcQFGurEn24RSKn
UxoJ7wMALeCgYYhDPaGgQwsuCqNSMTsDy87xz452dkAKLfrwtWDzjuUt6wLOyLvMtLLQBCXmTdtO
9YTMfG7PZS/YqlGYVi9FhUx5QazuAaRGve31bpqhRxvRj43zxZLmBtpwtDtvtucVGAeDjQuK88C+
M6q1hKxuEBhhwkhaeYvyTmLKKnJSnQbXmGcTGNILhx+tog76VcKj7ioP2mFx9lPkpAdS02wEblyn
tFAHft3HGU4dHAF/j5xenBGPvgi83sojswRRrYRkDRonV6/M33Hr2oWurr07sJ1N3GzkeReIe7Lg
22Q9cJx0DlymaUGffgvB0D524JCCUHBwijzY9mztQ0dV+9IKIhGf7h1f5GBpWaAQEADBEbXocIAJ
yHppysdCkAflSRBR4JaTwiem1xoI2gvFsktU37Jg+n/kBgH+IwrXvhFKUziqlMgOhaijVru6yxO+
RroJbCYWpYqtSHKZlUnueUkb+fLw7/DIPyODBSpLPd0m+bXAjgWmdpOzX3eO2AY/dAXvSe6LwjOb
jnwZC93qsiOXAUVzMtdYyTtYsvXzh+IVtF/BRadoOFRuGHvaclrWuxt8A26assIxk3Cf1d+mRY0R
hC6euUXS756Acn6bQPiYqYVdsHWRT/JLcar38YcGOgMDxd/HZVovoO5XIWwHrB2UhaHy8htyV/8n
9jGHri1svks4T0U0EaWEijHD8Jvm4UWmmw4wMYLSM9hAmvzpmlgp0aUb6FwhtBP6IDQLxMR/GYoT
4SgFMUsydyZjFoIz4oWYGaXeJjFYUBXVWCEqHrySYY/hBRmrYGCzaUaZ7KBwyTKuTXZRs0xxkJxu
D8twIj6oRgIxFCslauHEutraumzNNcB9FLp+CloJVw2fRu0kZ+6AhCKyn8djBlNQ36rsK4aCUxHk
uuuOrYefXDX4xuT0MhUV5qIYAaxyz39DL5TUhuBgzlXlwCiCaYUosQFNSoB6TfDjTwXIKUPwIa4C
pwi6qqdWjJO/T5rnRmNDBfpFzCtKaGhU60c7FUVfIZzlNJIi/Yb3DFz6EiS5l0d39ZKp6L7I/UEP
I+u1ZefKpBSuvDh91qCkztyZn4mrgs3Mzg9XBhhyQsVXTbfIx6KMRsTY4H55YnJgiA+SSuKVNjLz
au/QPWkPy6ws31n+iKlfbbPRM4Y9K4vbYX3oGbZ0+Y8Wm0Ebw+CpZrzbrgHmGD5uJg96Bl9cK+b5
7ZOkNtNPoQWVbQS8GKNICu0EU77XxEK4Jf82S8034JIO4yHIqut4zzpxU0gVjcksFwS0ZKkMpIXV
hvMpoNBqwgnxvIFHbVQAmxpLYR/Xp6cTau4eKHuOsGPQDqqkDjjaA/BMFtgqbkzRhHTYZGWpgJMi
vUcxy6HwU6tdPkALzKfZN5E0MuuSiyrPLGqUtWGKn6y1jk5ookYCuBsqA/x+HEFG0R96LIis5X7X
EueQQ7rMFKa6FJZvJS+zSZde/z69wHJw1kSDrepHqFu4en5VL6tGokO9b/Lq2IlT7MIeaahh+gqp
S4fxKYI6R5C/zaV6p13EPS82dN+DscW2n1vmSOeql4FSwbGr5HHIv8uQ9tJL6rtG2BYWeaTWQ54W
oAuGIfZBMbzur+HwYR/1SQZ4/oc1gRxaIE2ITIKTITtyj1zsW0qwhYGbrZ/YprCO2ZdYQo4POXux
hy0z2iworUWcyjcKxy5MU5bLmSgRCVhE7ooAEAZflYag1S432n3kWi7JlMkdkuu/YNOMRS9h6jRz
A432tsOSJMwJyckBM57P19QxBC9hd4L+W13HlcOMHbPhn516wjthH46bVRhX2i7DNYqnaoRGCIRe
JTqnN0c9/Dpya00jO14IkrKx/5nziVkadFiJQtHfjev2srcHSFAxod30yZHxuBJ+NSHNq8VFQadb
CXRyZhyUQS5OUt9zKOuvHDKMR9xgoviN4ABDiwiY4WsWFSCJ+MYdXGs/TafwWiathtJGehfPEO97
mknmbdXe2Qbrcof+ENmgdGsXqeaMnH3kMA/ZqwEduO76H4Bjbe7xONh/Zy25YhZZTW8lqvS5Qij9
2AlYgUJ6eWfdRhDnIfD0nK1TrY2eKoHhz8qH3NSeLNTODaI0IAwvG8g9bcIYqhWQ9/nNGnk7ak8g
/I7CYmCIY/nil+RuarumVft8JkQj3WcYKNKrWzdiIvk7Hvk7HHIh6/rOEOFOcBMbQAksCk+WQXXp
iroeOzwsFubpHEze7wnXkCemwJHyVVpZwlXbQN4SL+j6yEchLONNdbZL4KTjtmW8S+iJXLqTD47c
m2AEIt335lfE73hspGzWpC6mzQRd3lkOwfiQ1b6p3vwp8OOV3uUgBxT4JDTAyJPqtjM6kfP6CjOi
0relCQE7NzdTA6E3gggLRj35ynU2IpaTFyBtm9L2n8enkobhUW9Y3zEbTrgr9/X5Xu0VS0CQnTBx
BKWSrJQp3CBlIF/14qJz8FZAQsAwvox7dOI8WAbAyu+hJK7SxKmXeIBjj5U97vTRe0iAljReTvaa
s0wny2HWWgjc5py6/VA610Hw5oqF15XI1kpOebR3CFGneY07/LX0V3tsJIUTbEHQ0KVPOlNazSBh
V0Tz6OdFbtJVVUIhpOpC0yWJkpUCPxe1sNoI2PByhSX+8p5oMXuhbzgwxfjcUfFStFw9AUzlV64X
I367QkNyxMaFQIDB0k3XWBjIqjcPYmgDvOGn0W5qjuAh1py01Pno8BSQml0aMXQMDyRCOjDMSM/4
l3pA5Nw8NJpPV+vLWbJC8FHtbYQPuxzBwJDeY+1YdcIuYssLVuy9LCbm9eNY6mvLD57qV8vXT+db
nRsGnC5PGVUbv+23hW/25CgfXd91034lWL/AsVi/TT/YLbr8ZK27dodZF5BZAtsH5pucgAWBW428
9lMbLQ1ZLFX4Y1j9I5wAIWd88F/UYwuZQpQFNI4J2Pxu8W/yo57Vrwt66scEQKIjfX0w7nRY/PUg
7LWvO0iEbjqnS7uxkqhdmDJOKvympeJ3MpoGPrHL9cR1PzlQ1IJnIRIJfrlzXhTAQk6s85xQSDt+
KqwZnM5yN+AXF+104BGwWendQLDr1nP7fvBE/eK4cwiT1L1F17BX0CgBiBfaaD+zBhCxvw4EYuVP
JCeKcEQ8GSXW1imu9chu5zEYdEUvg/5cfDUeVX48VByyW9k6ACWIjUIiyp0TVn6kNq2blgtllocU
X3vH90QpfW2xRW0JHohnzkYfnHR3s58Dm6D+katSkgk/kvjsh3KqeqVw0/q7Bhz8tFuraIk92pKr
18LytqZROqMG2BAy0JwBq65tSSw7qbABzjHOOat1tOsAlXBJE+bgmv0uWRoW+jTBMecIL4e+t14G
LIwnp1RpLKtn8FZndGfmhKmBNZyTrolhR7aiUK1tZ3xhxMS6b2/fZrloiNDHmcCyC3TIzyzdVztY
WIneKktAQAzUn/CD7K2pWETTsebrv5vd82f8i+CFMmiSZeHv4PaD7Xev42JfmtfDUMqyFGvDOe7+
nXTbJPnPiHnElU11V5c57M5bNytTgBnkFMTXfrrdEXh93Qhmf4BqNSNOoE7iyL4yIiI/AucsWm1U
uZgUlEvb9nh//yMDxVNLEgT5oIx9BTdkqgGGQjq42L7ESZyne4qQ/bpBtFowszncHou2WUY5qy/a
LeIr8nW+rm/zI1ShFnvUjZZ3/El2m008ovLmqXh/hSfUaz47mb1Yekel4wD/vbApCWGR45yaSK3B
PA6p4pL6wziupWzfVjQEq+t0AdZFx/0pQmxqVOZt+Co9xYi/eoyQihmNtW5jM4AWpGGR/WY8yIMU
rygZ9A+hy0V0Q5g985yeIsBN8vDc4Zgp4nIdWFO5GucMNi0re1rh+7V3BlSPoX5MQ9qWC/RPpeX/
tEbe7KO6RJpy0PdXfDsZV+2pEJa0JSx4A2aR9EvAFH7tiBgbnHoL9y/jb+5lUlcpAH7r/OGICQ49
GmPd9aQlvEuuywH+gzBgftmnmMqnkVP1U8UO4KalVwjg0tZpWXOomugGCpJEQD66fHB6XbSorxuP
5mW7V1Nfp4bffj4h/eljE+Sr4OgnuiZM2r3v4an1csjODt7WDOS6b0odPuoY4CRxdJb01XB0C/Ai
GRWhDpUpiPhq+5REqK5+ok+LR83Un8MXpkjh3PSISbMK8NvrPNrnWAcqWFfORyOIACQBmM+KYsQR
U6wlEqP3Fbb3r4DSmOCoNBAAhXEGmukJ5QkjV+WBakpnZz+Ny4xk33w9TiLBmpmS8A5OR3MopPKg
hPDXuX0z9D+vwCRRjh3shhCVjyPztmfibHe+ordnGmPXHrz7vTRLD3B9i/UptUCWhEj4xqCvdTcM
+jC/NpT8fct4ZrxxVdQdtztI5UVQTMUbuUbHGhsAcY5aDp3EKG/t6V3CeG+XiLrUwyAd+v7Z9UOl
bNDkcMheRR38ybqCQfQVWfA5juFX12lWYppeT65tY6A2u9PRJJ7COch7HUVo+w3MUiaa3yhoSYl3
QXeNaNbXrBHnA+8j5abOUUTp22GSlw/maVTgQyoOVc3GpQaXsrnWDrOxjMKhEkbwVre0Ipi0JHD7
Fc2dgGErUdEtf2pODV/gdgarO+ikHaRm2VzHdAQuP6gQbpamXjc3nnS+QLeLDSdTuh3OAgKsNtqh
R1yQpJbsOQCDJB1RCTePCiTAeL7LO0kicAgDXhL8oNDvIqoKjRlAYa4xY6iG8rqmQdztiZXIk4L6
9pfkew84GPQQIKIlfHc5rNDDUJmSt75ieIO5fug40JFDYO4wnIYbAirrNfTCnKCV6dhzrtv1E0Gc
jVkdpUoJ+rYPiRVl9Ruwj0x/9rsmgBcL2ssSovqLWr5UJb5Oc0FbPgmlfJ6Q9OzqS4y1XN75rTDH
aYZu4q3/SbzH7oG2LCXvxCaIa2ZCwClMzUoMYb/YY4LV7xzlTeXTwaEBmdL81+sRJypflygAN8BN
j+jYnt4kc7HMzwIquQKDVtD89EcTfdqQmsVvJdDFp8klJyTzjZz9XqzJEkI2foI45Q/b384RMhPI
ZdhhZA2NVX+ITn5ofhCepe18XFWmVIvHT401zZkTTFEazcq7Lg7ODd7fYMnTa8Yl7pL45D2beoxp
zLnCrCFD7yd9Up5Z3ICVUtDPi0MG+cpiEcdavNwuDm09nK9UXo+6zQquYnPPe0YPgrTSWBoN86qy
QZAsnD3qZqqCBRe4WfnhiE8igtm9LOPVVSh7aRyi/3ZrQ+HiVqUeyxHvRvLV+qA35g0fnPbsCeua
llx7bdEjEAwLdxJVqknAI6NAZwyJPi6whJeNSawMD2DEIS/25Z2JuC5IhPXpam+rfxOoWL0fS9kY
Z/VI6nn+O0jgKiZs/vYuhxdTlsSxpStERLxJ5zzgmB5Zu5S/ITCwgstm19wzth1UZ+7g75b5DZjO
6JnrS8jZyurrO5hVMp4FfMxNtrrjm93KeuEf81N+hIQVFBh3tr8A6iFEenIH3mzBgb6i2zCwsLZ5
blMRMnbxnT78eKK4y+Fv/j2gptEaXZ9Gz9O9RCZhtPCDJAL1fjEKCA+5xaNEpX92z01dVdgBCnyN
J00bRu+CKxZrV9hsfQFT93s7oZyw+o9x7hh1LtRhENU1wS0l/E3l3pKw2pJtS+24OD0MFq+ITvdX
Yz58wa95+obGDOe7DUQ6hTDCl5iAcV6eihFQCDURwa+A/ufbUxPiadusLWI1PXSw7JfL3WzSkj+h
36rE6gECpdsZsiVR6RBmhULOeuLNNtPJWBz0phDPFre3GXrxxxNKXFMWsp8OKXAAlO2RgJHO33Im
2zG9hIzn+sNsYMEat0tK1dVml4cLtT7qGY5osFDCQziCwviiUJwRzCgkMXjIP7TtZ5Z9Iyyq5JRB
p/MRFfmK3tXh6R3iu3hm3ziWYCqeRpvWisZsZhOWqMMwDPgY1tlKeKbE0bqfl9LzYryl3nuehOmg
BE40NjGiaQzL7K/Ip+qhn7/U4/QwocfMvsCm7hi8zJftIpFIzxpxqKTpU+AUuDJRRND/SWeh7v+f
2fK5ps2+8BhEH/0Ras61Mzx3Hx17SSilicolZ9E1Ph52Fiuh8xs9NckQQe/ke2ZuWnsknGMII2H2
aKslKt3azJQ4f0i1zOnacDOFHbbrw7qvrHdqynrgLWTSu4AAzPUqkP7AXnUEfZEwFWUSVixSmIcp
UPPJovf7DTL/VKDegu3l1v2elWh76KXkretvF+E5l5LJh9/cqjMu4lxn/5h0ddm8pSls0ryKmKSN
MtNslh8H0IB/oVXFupssk5hpihPCFJDWMAZFeCis9ou4uZYw0I2R20cxyEatusNMLqeeA6zv8VaB
oJijMNWS8esNhkcAy4y6apQ+NaCn9sj4EUPsNcD1MSTi9jtPhh6ksaN+uwMap7bIsdRY70M038dr
rLPRFHw5B05rlTxotrIapqP5f3TAqCSzXrRwLz8iqluB9MzrfSDPKfOvPWGAJrSFBF8WYulIbpkJ
A5G3XRvw/TlpFD99jC4n3YmnW83O8ur4OX4YdTmBs6fzl0dQRmTnqx2WXJDixixbETzPXew+NN86
WI1Uzo+ieqQG3DOPNgsbttgwdVj4geEt5NRRhAb/z1o5RfBaZwVib5MW7biB0yDjrfMPB+pBPWz+
VDBHdaDsiTCP8AkzBXiAlt+afYlcxZMUOigMrpxcn6pYH3aEoSjLC8LlmDFdJAcHkXwl8yjO9INN
lFDGadsdQepNt1IbWasQdSPcE41JRs/C+zqDo+ftMqIfj+mLBP0xZgACFMsS730E7qJAfu0AfkWm
1rsnQ4H6I3l4hXRycmnK4SvADQmqhfGI7jwHjaqDxINyUUFC2jj/C1ISVDe+DMUoOe8WrK80WfC0
8wmwJkcxioXfoFRhibgaHk3ltGo1c5huueE6YoI8OBBUCqeMhAdRV8vg5jnSEY+ufP/XKATX7w8H
fJcfUvfuyWTgQM66WEwemQxBqFY0BXqWp/dUHiAP0ijAILN+lFEDayZnNYTfvloPcGfrK6OKjEw6
0BFTHPXe7GU29MD3NETEb/sqZJVbhYswbxWt2wmfAmSaG1DgMxrsIgb8oIKxkNr2hRHIwPbGiMFA
hDyMlrbseJwc87Gj4Mn3VXeRotQ16iJqOHgM7c3Ixp9YrciMfrjGR0WOwXjrO6JngtVlmZnRMGuD
anR0itZ3P3traBydAijrxEZS+sD5AYWYzO4VRopcDNc7S369AS9UkX4/KLe392738T1ZXInTOy/w
6OeGUFM6Wb+KDE8bTzE+PoxMSDmPeezn6h67fcFp6qIlcxCQmHDyW9Fdk+wRIX4G6eyTmfODDu/8
T+hkK6TtXwqnIIVWJTcJpJGQxrk11mNFL57O46JOC++oeKMVZAzVH+xsok48l39COUCvonOCIfZ3
6+zd8TyG1fnqKTa5IrUC/AUhNjTKE3GV/fUFC36bYcDAN0xm35HswzJX2VcyEPtHu8k9A6JkrisQ
MaC2fY2LD1bXU6rA+HQk9WSCZbtgdqmbsg3tiNAenZUfDrGq6qNs5sup3s2tK+P2sUJr4pJwfyhD
Agqyxe/qLjCiyomN6BqL2XZlbK7Jyn1VgJcNqKFleSHD+Z6UCoH+htBLSfKrbTAy/rrDyuusYwz9
MoIz5T10X/1HjjKLdvO/pJ2vjk+n7HsqxQ5vesrXn5ivSfqQurFJukQ6P1A6oZJqECOExFhI7ErL
PaqiVhhVms85PafZybqE8/lL8ImYiReyRwTXVBOXRLK5KW70Lydt857Qwz7nzlb6542ylQ0qetWj
Tompyk0v/mSFQtgQNioglspQkvM9rsyXzJ529yqHGBapP1aKiUu8+G/8s4SDk9BbqJZfFXEPVmtl
FeVS8cosfeP39FuI0dtV8l1vUchc/19j5p6kQHwDis6QeQ8H91rw1nG13vZGB5By4PeGhgWiq9qk
aEkYbppUVuxhUzlTfteO8o3eb+8sQ4HBbNshAmNfMN6VgLKHiZ3NWY0K+rkoImsWf2pIBlAKAU8f
ckBI4rC0J+VFCovRjfXLsjPIoSyuruWZ9Yh9nbkgEy2Gb2t8p90i5lJXC0qvSqDwkaYL0NLkXmST
nLOwDbDrTMdyOk8KVNVsV96zC4WS7DPXUNZH5MdGpmGRey8YFWI+i2V59AroKTXgLwXOBkc3rmQQ
K/BLU7VZq4A/zFMhNPvA4ojhxw+/3gwqmkBRplTlguzmxPwgG7uY7BWQwZL5a9U5jNy11GGTvULI
20eIcsX6S+YAH1NSuaSG1iwKD+yCpkTouN4XuIRW40Yrnb2YDtslLlCODVn66/UlfFs2msvqpX52
5fpZLGxzRlX82lCjsyV08QUawElPBSR3PAKEJbVKIStDExdRLEkWubordVB35eDRDBx/sdoTnvIH
xJPn5/Qhdp9aTK6PiCR6z/bz6hBp35TqEM0I4UBfV3UAgRcju7Uqm1mX0DSjf/G16LMxEaNDuyIZ
VPyP1Cbsq+rn17c1yrG8uUw3NPr/u1siR1s03a7/aHE+A4whomupjQvoAQ3e/kW9nZFBmvh2ZLoT
z48RGoXHYXgdVD8nRxu+LQdI4f5/QIkutF+0/b0ivTsDCxEpoURam88o1JgPHxBBWuI8cJ7Fo9JX
ywJz5uMVhR3p56Ejk/GywASwFj3ZjilC9OhosDksS0tTgIQzb+k5Fq0AWW35lRIFbNCN163jjh3N
2CLWEUhsLuRAWAMS5ADLmKq0lY11VWD2MdEngUD3kjD4fdXVTAUoEOVhr2hJ8WwzTWXHYgtSYd3L
k6tM/vLNc6oPVVF1+rjfn9VPyObvnOO+uQfg2K2F6lJOq7N/cL9Y2YJr2vDEJpRqg94SHIMSd/Pb
sMa4XZZGoMl1r/B9EehF2PEWGJziIIF1Rg7R9AUbQYs4zQ80miQ5YHk8tzfysSLMxmrkZmEaEYNm
M6K0jINydi8nnrWZBrnA+/QUbDYsdW9roSNh7mEQOOJfeDBmwD/u0Vmcjr8NroWAbMWzG/VGPUPX
pQpdMY/Ouw4KJiQD1E8NBvgW4rDVkHTESgBQYnv++2kNWfZNc1AA5WmshEsSLm0hl1q3OfHpXCGN
TOjK6jh/UlUYBVNT8QNN8ajkflgWCcvF5REvoqhDge7YxUPlRhrMFvT/e2ZrHu0fUJP63+XL6xSI
JqBSKZfg4fS0UlIuqJEQltlVyrtHqO2p2xaWVntoZmhl9GQVpBrFbfU0HW47GMXqV+gWVzPioWYB
Umv2dc/RUFIcDs+ZvLTj6JvQCUU8cJ4k6aJrh+as4CKVA3R4hYxY/EzKJB3YzbOsWfNB7e2v2qtC
ZKYs3nMtCnW0MJWkggiwgA1+l4CkYkNx2B3ZDMPAiVRwXarhGFNiVbIh890CMyhqjGoosH/iqcgr
WvTbQiUPQhdZ8uBXWptIfW2R3es4yq1W3ZUdLLZsA2wbFRT3hvKp4sOpstBjJNSbk+ksu90CbUmX
u3kjscXfdogbfvwQv+4X4vplf6RDz4HWzigvWEuiu5zI4hy3/SVBa59Ufr62aLa089L+yJMw9A2b
SuRbNDcBZcWCEYiomHyAwUGSdnkvw7PYwp11RwwLvaFSqJ6rAtRBmiVPzBRXfJZ0WcQlJhWad6al
XlNOiu6nxbs6NLEDuQp63CGAG3e7yLwvBGGYlPTcYk48bmexKnvgZC6l34hzb6l8lZThW7GyD2IZ
wG6LVVdUuZnJhxqUZTrjTpxWDOH+IMXXd3TTvJ85XIPc5zPimegy0cYSCxkUNC72g3AMFDpOL8Vp
1e0aUwsqv6RquisRxT7jnvDbDRn7ldPxV0nXOFd8QMnazqNh/TIrwm7t+CTY6IV78WrMAL51I7Ji
9x4v/48fZT6vnCKef5Gm/JJhpOsxWgYTBi1V3w79S+0oUYzTXI60Sy/NX04fAZOPf1daPvVpDanK
U00dfI4DiCNYMXTjwb4D9aQxkC8SqI+fAsgOdg2I6BJnfpUbB7RMmzCnCV1RQQfeOApnmkTFnOUy
Kl+TYqq9K+jqt7NbFN0ak9svCLzGvzDtfHP9VGRh+4/A9jJre45OuZPwk9kJ5EZWj46tj2m7YaKo
b3wB82e4rYVPcj7eM+l3cm7hfM3OvXpR4QF5k/LgKjxA0EUEL2U0wGG3Gt8bFK5aH713/Ulhy96t
ejnadxK3bfrHVn2C5lwqjqbI0fXNyuS0AD1zedCgaXagxmSxw0/TOQaAdtrCHjCsfz6RbByrrK2h
QrPH/7oIzgMIeKilkgKTCGeFdrCvTEMV25q1+o56JZH+y95frM9RCntib2SLhmPMAYruX3AAqYiX
4PxwcZqPhuMkrqWon2fwsD6JCnG2RnsWBDfqPb9XK3aPuUOz4dd80XyfpCXyzn5s2V95+f6NthEk
BGGrRvIKvG5esNVBEY+pyBqm+br0OHkFRXjBHLxFwCso70qNdD+Rxgrj9frVXhHbB7mFtNCYNRhZ
CuCNsRJ/wY1rqI/hkcm9BPiQxFIui6IGr4VzQefCmVV0zDpkuWMTaPWSXcDaZMdN3SODSjCCjxsT
xIaGtwtiNivtSU4scyCTzZHyn7yrx+fDAVXlcpbaRgRWzt31tQ33+/VSPU1rQXasjPFI+x+MU3uM
NO+LqdR/2RxXuEhshQ0SaWG7vmroD8x6fGknWE/SwLE27X69GqmZ+dTRyBEC+7d+CnIhJN6GecbL
fotVFoW5wXN8csK0RzCBOAuVD7hx7bSUWPWPNHEcwmghW/lhvuIa/cWOJzVtUjpTBIlw/qhuYQ3i
rEg0/B3meTG/w7ylelxgR9YewtvU71GyQCgIlZ/eI4GB9yFprALiAaqQ2VrRLxPTrO4gpEcYxGRu
fkimkpJdMp/BgJBL+t624YPfoL2xH7g1efFBqbJyy+72oKa6mxQzIfh7UMHEwA/II2hrj6cc2Inm
o+LehhGMyOw6soaJhRD4QgpWb3ykjLJ258PLDbG/ju04nabfqjVF2ixyw4o8dfKt0u+2b5KDHgpB
cfYIrOsUxq1ZXurVRX5A9BpRyS/uvgxEPT4W3l5Cj/r2fgMOf7hEXivr8U4eDNrqnh7ZduD+gwE0
cd9g6+BeVNzQ92tgdQFyj7lV/jt7iccik2imCIabPF5jS8a4RIdk70d65s5kgoE0KREGMaRR2CUM
gHoKvZOawo7k8FQ0w7jIPSGMsSAyh8SMw/d3zmNo8NnXeVAOzMDU7hNQbl3uAhU8mNx2tSmCZ0K1
RCAO7QWpnEpcAjQQ5eqCW4/GgXecMWj5qYq9cUdOoE146u6MmzWV3dspWTmvkLX+108/wNdTHAwj
JDGdUTalGZLsIgviJmLB4Lv6ifXTjxlpL/mq1ZvJ1O5JSFMWdZny1pxFC/cOx5dOMjH3r/kg5NKX
Fprr7vaZbhgyFiwD2OankyfhBXNuAdJmYkiSUxBNXCKlnSwet2YvzGPipcF9kpUqsG2zDcFqlq85
+Lg+E+hBVjvU/rGPmJ8tzXmb+GqeyMbX2OF9HGoVE+cY+QbaTQ6T2m+AHSqiS6Sy4Xh/XT6m5OeF
oitVz9fItNwDGHqin6HMpNZjCelBl+P+M1yl/4zdxIZBHCec7AUsSozm4JTzcrJGa9CfM7XuYWIq
JPRR0xKgVlmVuI1EOaUOYsIotMInEvHI0EQmGJfDvREnxrC13A6lpxdTyW+GlTCQp4W8l73agFLH
/BtxqLwf/XABgDevzquimq/I71Ox8+F1FRFjdRgGA5nndfz5th3T07t3iYJCm9CpTuXVO++DxGzo
kygFl2JgORyd9OzPlbzIbbPGo/8C/WbcSjRihxq7YumDBQixE1HMfq7UGS2dcS65cR+hra6ghVzq
7BahoKRlpWYU1SgBDUg02jr7EYJacIBxc5MYvNtJYfRbQEfJ5hgK45Uq1ITv7cAZQEpCC2lI82ua
xYk7VTyMD9mN/6jJ5ZQmc9LeESVJN2BUecPlj6iYyBPSdeSJ4hC+mqkx5NwWm2drEENc2b67ZyMi
n7Ivlqcqg/X2NXtpaMOS38lz7dZeF8IuB+sPdwjQIAhGHffbNcgmOfZ4Y3urimwudznDNtRvmQ1b
eGg0O7Ft7UL4dKH09WS/HS/g4LaKkPoIjc3IQ2c7735eBXqiqzc8ieuahqnKuQg85VICXtAT5nTz
d8k3cFUjN5VJ5+YPrgGdcWnM+KoO/GQmrJIbaCB6vsLMYIr9+4v9YBm1vRNtkqcL1TI33j9vQoTr
h8Lj8tkys16OQLmtKJ/kDO5pGgBH38V4kZmBJbhySK9WI1AFOVyLGqhpxzklBQu/520bRLMD/8nz
1xQPdlTI2EIUHQpdNxMgRPteiYLjrGHfKQGriFPuR0sYzzFt7dh8BwaMt3v9331twz5tR5Kr5+Kq
oSU2yqzgFmXpA2oFvkEejtRvwLQ19ijYnBQsHnSofBZppnPG1FkebXxi3v0fOkuv06ojmL4kJm4d
kbZ5zgGY6dnBbEPEFplHlQWXIL3e0J28PK6rDMsLZenybiJPKci8FpsXWuJm/sa1sgzvrpJG3+Cn
Q3n4544gU6PN5ffQigXSP4vUx7D537QFtjiPONfjPraMn6+K0zgKyXAeWsr6L5zhIhwT+gxGYTEb
Ff6XeBwKrzTM7ZS/9VsAWiu7/bfIAO/Wo9HJa/FjZUDiNpxxGN5057jU9+xpcEUx8mgW4H3eO0jP
CILxC0Vle6UvDIFwxEinUpQy5zJgl2hL6t0FCPbQ2VaJhzPf2teB8quv4cnPYPhIKDwrBuenkzKs
jFOyI+5YHqUlcDA7QlE6oVEsQm4iWYc1+mOwGjgZyJxYTC0stsZJ98JGjckkcYxi9ycElBI1KGeG
VJHDqmen4iktFIiwAv3kznltPinsmI5gwgHTvU3DBftVazvqRGrDd6AMFrGBn+01AGLJ7uiRwVkv
iMACPvHkp4SV+ccyB4B2onpJ3//L30wn4Y9x5As18arn5/AWkgEoXTzD7kzSfbsdvojibZwnjwY7
iE48vsMK77qNDfMgha90i7zb9TJsmNLl7H4HZasHZNIQRWsYp+QIKQCXYej7OsRJlXTPuVH1m18g
Qh9dX6qlozAoqOYpmyKmoUoasq1+4euHvlsgyg3jQUCyMF4ly3OdYrdS7dw3GTTbFzgKLKrPDxGv
OixVERovzzLQ4UurKG7Dzqm2hoBXmdzIDYwlAmEVI496s+fzDdeA1vML1w/zksOsll0LfyGQMyQ0
0I5X4qCqkIR8dToxc/KfJnhclNItnoeKAJ1X5hTO505Y5wzj1UNliBafqeXIkntRG9jttBrHoZgh
FGO4k2/f9rjJkwnCQee9KCMf1jGO3qVbY3zXT2Tsuy2dDYztENMmYB1e3dWOtzthSxJuc6H5ByOJ
wgiGazGCCkp1KCJxVmhcYHPD5AodWNAuJDW07P9VvJ02aP1wAoicMl07NfjOLGR/XK42vVBNx9F4
eqzGloesPv6gWViIOCWgX6VpzN++M0amtR/N2mC5PAsZN88LDaPb0tNw6MvKJq/L0cu3TEPrANTQ
iJXPA9ngqIMFY+h8WG611U6CCBHWeEGh6BmgwksgzdpU4qYpZ0o+BjiUK2ChUF78ySt2aKzpyFjH
W86V6hX/MpfbG2uPDy3/qbwxMLWUhhlZ+PJ9yyjh15cr5ZBqUHliUOORnfqqfX1IMZkK61+fxxSr
jKYldHLit9AIsxMkYJRkiIJ6/kK8VorNHF1TAHrCrzJJOVg7cHVImGvmvnPlqJiuxa9c1p3CmfNl
S74G7sbtxlZVq4e54a27ovRDQLLlDFSMGZSDLGpZJhE1uqJp9ryNKjxPkiO47BxKZtuNtkOfqQBb
XCKW8yJiSPyVQHhJheyLN5qsDieRHONcihdAMS2QmTP9cExC6niNMqQYGvW9hju0cxosW0jCj+Re
ujY1qV2QtdZqEiPuRsfyRM2/hSdP+IzrdB4tfAgkgL127LEmyBrKo07DgoP0s4YZAgelO4eDPdFO
8nfFINtCxZ8eeA0LBb66xSHmz0v6sa8UxZhhFifgXzPZPT4pxycPrzH+SU2m5PJ3QBGUJ71rD5z7
551WEjFUlXMkdcnjAcV9KJCw4hrg44VzhbiJMl2aSH6dKghVF7ty3b5bHrq9DqYk5tQAjXp7ifUh
pt/2CJj2CG5yZ8T8SmQ95UnCU0aYw+5nauruDReJZGD4Omq3pH5fWjTCG9Y78y957L80OtXs4j71
XZYBQn2/vphOnamc4qJBnsU2VhHa7UWpyaFKEN3Uevnt8Pm4m1UzzkSayYGJnFSDgpx0x9m7oAas
iz6eyIQHVyL+MYpdDDnXWxNZp48sem4g+pmrQW17djPgySsktOhXH+ur8mppIBH0iPFSD5oiCqGF
ptFYvzqJXLeQfXJc71xTVwHJsnH5WdL0DZsIfPbAebyj7N6AMUmPiqCda88gRuONtap64kl0ABDL
kNgOYjswb1Efl8xSsWaHhhDQepFDuBw7OJzli05Ow8hgSPdvRFl+bnfGu5Tlh1uuHIh8r7T/28QW
r4tzDOFAEBeOGfIPnrRJMJoNwfqZzVxTqDZn5tovEXGpFu+YZ5wVKThZF8hLNFxMiTmp8QaruNBT
Ma/yeILq1x0cnlEwsla7bsGhTBFGRS8B8Zk2G2dC0hNJXjND5AJZnFmba7XgOsXL8SYR0qk4k2kb
b4h3sDl/SZzXQqiJwE2ysb6ljMPduCfcZJ6FUW2UyBd4bVMRj3xkWCWeMbUQCMaenLB7H2kjmhtp
lwaIOlHAi8ZbD8ghZ+vzaObvsoXHwh/8FEk8fH5QhDOnqE5AkYTCO3yySurbUTYCqDd3zx4rNXGH
UKnznoMLlwMwC9hohCLp0YaCK/dheTHMS+LIOaPdTCbmnbIHZSNlJiAtlhIqqapvL+xgTYyR8j1n
Q5NdMzz9fhZ5LRtDJDuhKwa270PoCbkuBso+/gn1i3P4ipfy6LfVJEDr4RxNTyfFt9tUSINirbKD
OV8j1izH5AmRPWrhBnv1upzC7oMIpvqGuVSQqjZi/S5zD8nljVbAysQXPia198VYO2seqhEP9q/0
yteyVSjvqOow+13MEfgnL6Af6oAJbYukWBwPqZwu4vd5bsHnELWDwVV7PodQLemSpKrcD28KqgNI
g4MTL0y0YwX0QYw8ZwJLIVvq6RtHdkAb9rWLb6aDHvDAzsxsI3Hy9ByXLnciG+u7z1DtRlWzgoEU
G31g+keWjxtQnPcsbauZ+syijUo/a4wT3LqpwNBSYc9pBnYwR2fl9cZIaZOdW4tOj2I1/E+TcNPt
ciNe8RDz3hJacp6k5ypc63iR1fzHgWUmXO3qmNHFpk/niYl6e5bXLE+evsUsgoMeCUheVWmzIfCC
MKLMqLPXNj6Lr/d0jf1/r05HDhmY/P+ssjOXHcqMwuisiaLci3Bh9wJ1rVB2/2KYYSwIM3uYzbQH
6xNyaNxOl/0kNhCCm+eTXpsKmrRC4xn0yf6Nkj/iUvqwTaUjLZOOpZGsBIJiE8WOeW0YUW0T54eM
D/VZE+Rv1XCkaQPWe72aYUsVKTYZWGBFcPRRY8KlzZL5oER2+KoPKg1ujSqEhS0ubEiEeLatI258
/bDvFEAVqRyowAvKC8daqtr/QikcqvULHbLKTfrUW4E+yd23myKq18fRopLYDGMJe6o+dcxNMAE/
m7p0y/RIMm1rDleQN4SnZ2UYmid+JI/Oqp0d5tiTsis1ijZbi7Gy+UI6Rcoc4KZ9RPuOh9JYZKxe
yt1iJacX+HaizaVyF/TWONKkBwt2r8UZM9EnSwNGQjP2KSvOSPF6pvm2epsEUxmj73bYp+fqqrZE
As5ygRra8pF3Yrll55TNgeGUWqQhlruOAjs0/37gWsvTMhhcJFtpqPF29PwOLNqAg5DSy6Rs003Y
1x7oOLXI/Af8dgTnf5Jh/wZIWJAqfuYEdEqawzULxA8+QHAkN5tGTlauEzFZcgmwonCYiPvBtx0S
NPPSQ+bqUNMZmRYVOJRfa7+qHWSbTWjnK2BniD1kHTiGWznKcQ3pkHlPqvNYHNlg7SFSwCkAoWcX
kZtJHtPRRTRThCrzygYQ209fqt705DjAYLu+AAyjyTr+1hzfomAXaipNR++WG1JLKVUG+YemHnDf
UAFagClLBjz9/4y70eXklJd1gZ3c2NDKOzBeUpS0e8KIBY9Eftkr9tSSPeWT6O0tB88mZIHU8Zo/
RnXqeE6TJJRzvRFAyKVeym+4XFz8zpqmXgBVlxJtC/Y3JDFcEKUsH8gO2XLYAm8SScCUdaBqJOXH
MWjEpl4vOGetWrrmn86IXi6JnS3pLgZQhpeDEREmrLQsrAbskX0kzx1vwFn4SusSBqYUMeSDK1i0
ZPK4/YDU2HbKEt2G3K4x6EPg65Z/LPMCDbfdJ58+U2WgM10vVuQDtvppgstvxJ+BNtg8TLlOa2lw
8A1kaGneJ7Z4GXF8n6LE8CmSepxHighgDPz5SOLI6isNQLYAG+YsmMjLmKQD0xrPQIC9OIeLu+h7
YvNRhVxQFFnJnmiJDa/c2ridzp2jzhl7jjJo93OmOnbnusApCbIKo81/8v/1n/mhqETLbfsl2p4R
08U+eOyiScg0R4lEF14orENDo5/KSJUewaefeAhHaS5X9XIZQWrxcr0822lL+bCMQYPaaJW/BEJL
p2ZLlo6MCZyhwxIjXshCINnzmvq3DoYMmP2V+iLeppEA8Dq2vIMHk7FIy3v7/N4w0c4ldcMf/U94
lTkupFaozOy4u6x8G3GCZ3u0veRmq6ENZJdZydPPaXwAbxE+Ydat8bIfIGlelz3wnk5hOLxuhfqp
dmQaTHmbFQnnv/SI/n4g1wX29bjCvSwwW9cjtvLpWa0AmqBzCyOl8vQCFeUC0yVAt0JW6maSXFuS
b2LwBNpYLUQRITWWuppKZcRsF6va8zOvkfcsTJc2af/KqeowyIYdE8iyZcXCi6GMfmSFpIVYaziR
2CaT190S64vuR4Su3bQJJEkIFq17QWzIODIa5VKJb8qE1zpe/Vpu01TpGDcxbpVpV91C4PVry6Jz
1CCGrnBBX3lOStW0MN/XOK7B7rz6ZjBkVeXfPAIxDolm6pET9O5TZ7kyJWNWIJdlBpS797mYusH4
xKbPMLn8ZAoW2S3MH2p1fFmK29DZCYFLL54zo0UPCFZfLf1KbsGag38MzG6bmih8YJ5FpAurk6AE
K1I1aaL02URyO9W538KPKNEASveCsEJr1BaagZtVTYUh+PVbpCIRDlG16cyDU0xtXztUWYF1cpoH
aVMjoM40Qjse4eupnKcmoduO4f7M3NwHw25IfSYKWXfsPlLjVb/LAOwJ3gMlHXbKczRURltN8dwL
q4PcrMfxxHBxGzNjM1uYGMRVrXuG7MN0ddcpsFsgkY/CKiy9a5M/JnDQvoFWrwdz8wZlP+muvAtx
kK482L6MYPiYZ3dL6FMekpETywqqb+Z0bpb2EXf5VxTroni0oakgIJlKx1BuKyN//bMhHcWS3UoC
SHQYx34jGJSAv+ke4M4d32bFm4hkHkMCXP7TniHijlzJYFI2ngmXo2+QBo+MwBFGFf4vKzHCJy+P
vPTUTQHTPCETeWpuvZx8AxSZNv5bj85yh7qGhjvEwTINvgDEONaJqpkQDzBj00KnnSMBHbrAR/cs
ytreOlF1jquhUagYgbA0vKYt+eKItETYXyABiwUxZge0cXUaW6Uz2mW1qS5YSPW2keuMdnrbbMem
Cf7qCIZIxhZib39Gi3f/UWyt4jgi0RelktmVL5P+OXuiO9QoPw2nUwjI94GAHo2vm7zbRsRi+Oor
cqyledasHG/pMdY7Zp5VwtWujq629IoDV1SgP8Z8TEz0JRU8zOeCbILnostH1QIrbcERvqPb+4AS
oFK2Kj6x7T/40ddKEyTnwaN5pED3iR7LQY41UOPop+cyzEoOGNREGVh1vhRJNUiLleI+6uTZBjPH
2bT37ly0DjFvmI+oC8Vh44QXyA4vr+hN4fMmaR3vfkb5H/wwxUMU8reQavv/WZpD9dgXSGGsCA0E
7+77Eoc0wSn6i+ifVl/SYf+5hiy2S7DSup9lBRUSdiEThNF4jW6RTv1zxoMoPp7tdCTgwUH3pEXF
/z1ye3KB4DbCb9yH7jYoenNzBqXfPSzeEq/JwdO4LxQ4jfp2tF+aNzPpxx1Q9QUMH16eRiLErJt7
ZZ8y9zMdVsKn9wVcuVULM76KBILwRWQrXfTJopDw1VtOWslQouv6fkWfTvFUrVUB+eDWvhX4cNKG
52NSqtajkeFAHy+bghHZNWx6dyuEU1OX45CSIG20xF6w0gPjJt2w1q94u0Q9Yz9u2qUBBkPaa5VX
xHjSOO5SHkeSXVWkx8DbYyrHyhqwm+j0iLr3CrGECsHHPoBc3oeX+x6WC7k5bjXPv8oY0INo7lzM
MScQ0EzBCwn2Qmr4+Mku8OkwjWp4SGITeIj8oHz6ggwvfV+7hm1R/frw1h2ZyoPpgevmxsuUl0mD
eBi8Fvedy2ucPIchJCHTpOF6jXGgj2ua4bhwa9Z9CxYCXRBU55XIY/90g2UPxcs1ck1QcbE3Hux/
AWqJk406otM6iFYuwr0rvibBv6abMV0WN3gH0dW2XCV6004MulH9eXRiZJBJLin7sDQb6iJa1ucY
ajRqpoZtSPvfYwSncaWh19u8D20Qcc3mL/28yRTb5CodbJY8PeL18XbYDzrEu1eK7xRlm1FgkgCl
N/1T2+sJBhx14i//7MSU5Q/XAA9stodSVc24JTWAQPxy+o6ZuQM7eBhxWPwCv5qMYBDKsgtmG7VS
HW8yTKCVC/G4e4MueCFLJv9RLJrrxET+gAz26Y1M7TYzbgABCj+Pq2qESTri2r85O3Ip7CBP4mjO
jh/bZuC9cMmRyrNiJPuOH5Ep6xr2ISOAEvGBntDiRMIzL9Hzb1WXXgZD6e+zUC0k/Xznb5i+srh8
Kv5CLRyH2rE2CGSzYvRk2MkZrsKjeyYnMFaQxsJ9pZVoEKSw7ef9Axk6tnepMNBmyvX0qSSgZJPF
aSFPFfseisyMckWH2+Lf+6dxfB+s5lpmL7s4d+Bt5uugbPSdcUf5hntVFuVeuzGlzo6QprqJ3EXa
QmI4b54veigumjlJhUyl2cB/4FgiKLWrXkG8b1mch59XB9HG2+tBn8aGoKoPB4VSi+rr/+NAOkOd
wrXN44opZIfJi3e5E+i20cx1uWvPwwoQS/IUocAm3Vnhi25J7njInCCDyrn/uZlevntbQeowLtEW
1jf43xGOAaIXWF4OHj9OEqP/mrc+H8AEfLIECXKmi2GD7FNYquTaGDaFUVhU3LQrmkxS5AkhegbV
2VGitbvSI8YoMjlPsdB0QbSNyqFUEqQMGbEZHxigXj/S8yQehNR+oFNNZ1jygLTsTl1Tc1RZegZ0
jLcFFpSDM0G9Xx4GAxNjQr66CbEaaNuoFkVto8Lb6Vuu8Kht7o1VzxTVdt9GMUA+f7CjnHCvWXQi
0XaZOd6gPA09GdMk7z5A7XeKt3iQnzSDbQTPyMbzIfzUdPvRIFTbWfP5m4Z49HRx0C0W+3jvkb31
vyhmMoCD8FExPzyXrrhyIhitpk7Exn0vhSa+T4x+Tfa+DAKRPu7XVffJBKxuVzBiKe2S2a3xYERV
AiQaYmqOK+wzLG5V+iwPsRJFTaI22JPa0CIsBwqfocE9BlJfSdK1YRQfGkdtqsPWEeoqojVnQ98e
Y3ujyQXlpQPtXMwTA5hytevdsAIMVMWi/AcmWI9Ga8mI4xhAl6Fkc7xkr/EZhzJ53M/i6nlPKLoI
gM0+6tIkWhxwM4NRPv0a/bFr/ctQaZ7rysWYWPAw6Xdn60J+lXZ3dQXSo2XvlZb3/Yw7OytN5Gbx
722yOeciuoX/LocFqO9sF/V6EOK7afGW5NgoPKk9W2Dw+EA5qN3T6ZWDjHHkFiYBu5JzIq+HLU+N
JgRItV1EWkPilSZMbR8TcjmmJB54F8uYeDrEaq7Huvr9jZHj/v+b9olMVqXtXa21ToEEnlAwCxed
dJCbQanguMq0m8t4aOXcZnb9R9vfzXKE1Qy35XgLjcJbIyPLbs1qANGQC9DGbx0dpCdmygh2Rs0O
oS/MpME3+/Fxf2rccj4dFVOWeyh/WLjh6wuGD1edy8NNktNbO73mSO22ZFnwr3MibqN3zoUa10J2
oIhd5R6YcAYvYdIR4PTsBMl5TQHrfhQ4DaNoT3vPTgAM4QqDSlUECyp5pjTqQZuDv1TvIHF8F8la
tYLXb/4JJ/rDxgdTeaV45Q6z1X53TGAkLYcNu4oZbjD9o4xa277WnEezXv9Dtm+3dm8NChIhr16u
O5VFhL6bjB2CZfvYC3qkepJEYcp6bQrHaDk/fiaaUoNvWlQdcNBV3QDZAQAvAqsJPRpT7sR0rV9F
d46F/yO7z975wUVQx8+46X7rMXd73wdxt+VrYBu4xaGrPTPL4A0B5oSzdSJtscfQUCKZU2ikkzIi
z1JLNYm8EeJgb/4x9hGMG8NL3/0CkTHEPPsVdxUwte0qQAoXuB5AsyC/r4QLH2PHRZd1uOgFxuJ8
bdva6SPYpE4jmALHLCYrgzBRMU9wPUuwO0Togi0tGgj70uIaWVwEmG714Az/E19BVG9y2pEaF2JR
HPR0/9Vy6gkmogncWwMO2GnBj1YnSuXZ+XJe/fhQcvNqpJQKye4Olb7QgIii5Gwq72k4jF2GJa9K
UWPWdRj+l0YVr4h4XTOlRwSsOQASxHxjDDl3vVnkdPcYgIyCbTK5YBksu9d/AlzodnKRzFkj6cMJ
zlQF4KBNY0endfK7Nr9hAkgQKPkZOHDwqRXskH5ExcWa+3+V/QvvWKr264MCfkwXFFFYRbfaKFy9
yNxcEkNujDCZgZXOkK2TM0t3za3xxSvBzn3oPzLXgmnmRnrcJqtHXShPHmF0TwMh0Lv7+IcIsNPq
DfEVURssq0/g8hWJkRDcf7rl/9CxpLXkuSSNw1jxjADXnbEnlGE+ESGjc/AuJnipg+DrhObHgapb
Wc+aRnAywYScGDIf3x8hSuIQGEaEMOpoUYi8rpI3oEtlLtynsCaKAH2MNeD/wvwPB5z8YBOSXsuP
YiNv19zuHrxU77tQwTo7h7dTHWo9DjPw0XTDKTGkmsWIHSPUkpdnOxLpJQwarABnj3s+3Vp3Q4/g
E5+0v4Q33yrfmEJ+SNhyy65I1w+uyV7g4cFW8pL/HjhVVPU/6xk/BqvPQ6FRGcTRPqdmEax0d0RQ
2E5PmBkiPsj4czizdHyd4PjPmlURDuh2fQFA0rFGZ94ziR9r+cyhFv2Yxc+OyHyLD6ExXc6yHlbQ
vvz/pgGfYDHmYi3vfwd3/ov/tdYV7Se0zcS3AUobp/OnvHHd6GEmvgTFzh6de06RwHwmJfpSGiTG
Y7UrQRflPu9nneQ4Xsf0eMhYJ6OJhoPNKPVnC2aEbUp8IzvucYqbxLXecES2fZVPDgGrCp2pKTAz
sih5PylM7aCZFTEtjhZShXhd8/Bu69FbYArMbyu+Z8mnctqj2W+PFx3HqNqTrAuc8AE6Hn8Uc3yO
0Cd0LaMEZ+vhJVXAS0wQUrBDiB6wErwEDZwFJEaEtbb22jFXz7BwNRykPtIs2wnixkdWbtVCw31y
qzac8pzSMqTaFkIOEzLyln4Qk+pLcIwB20sd9Gw+pFdQaB2Z/JXr9OO6noFwAiSn2PNeQ2VOXpiM
OSKxDJSdHYYlxj3K/l7exBBP58qTpRZpApZSQsbI5ieVlId1iONiHsc1q/vfPkK4HAY4y7ofaWi9
Nmi/HkVZktrQSVINviZz34AydhtJjpRIL/CoJI8P1zYUOto0GEqqQjiJF/zllzKd4WQpCWUl+P0K
/a7nQ7f5lg6BwtLE4t7BC75lfI2TrhG5jX0+yg/ITk8dtipMCw0sYgG+Md5r5xymKVLU6CtUg6cV
BPoCf6FAQyPnFLX6dq5Y6zNyF2akcCGFsc58ft3bj0VlDq9sm5t2lXvv+DshYBATbEpeViXh0CrQ
7mrtwmPaGmqB64pjW5SCfo1TvQl6wLg/VrIhCIPrrlrGwrylCvbV75tqhNlArIIS0bHf66nSWfcn
SG6pM9x6nywmlgBVSSGTVodeP9gXM9GHY7x/EBuvIfBpkuQFkT/Pu9Tyo6bDCVX7M38h7Imdt+Qj
CIUA4ZWHp371FJF672qvqBkBS/krY005upSlpo4t6rcQGdQ5IlnBkyXu0SlySbmWyACEkbbqv2Il
6noSCOCw7lVpjmJyJMQffvskBvdqBcFE9J+lhaQX7eFOopatNy2HqXx7fb1xfUL5V5xkO+voOi3r
P/mM4AbOBUU/rpKK0WAdMPEPk9bcJOElgqGYdNFEkl4eztJEiErGeme7bxqF7EzWFSblVyzov+xr
5oBREvpraX0+o29RNFvP8eA0MF2xLAPNssH8RI23ehK89xlr9NgSoP0tswuVlxDU7XB7p/8sycHG
/PYPPYB9SWA1XlUytWC/a/mKIDqBZEIBGgPIC6pI/2GOFDn/zojbN/Q9qRJnOdTpyjSrvrlUq8kt
G8cSggazgTc8o7YlMfBPTi1bZ+KQCCAd+UicFlI4D1MOKZ3DOP3tJUTcEO5F0qa9cJa07Kjh9F9Z
gDKTGHier1XNjx96dH2QGpExDSDooBOQYbg2dWdttmQmfRajo4WrojoqZ8UH+O8FkpbWGyz7k7Qw
L+jx0/feR9+SetVGcIRgFAfZmxgiqcftWPFTCg+WdZ8O2KzBGau6R03LWhfTAD9evEdClVr/yWDN
6X+XtnWENuYaVHLxlB+VrwHDbKv36ZtY1Zpdjsmj7gSXyM89yDK/bb7tnQ53z2LMIbm/klkYshrR
4YucnKhmGbAnDDpjMFg+nDe9cLc8AVx6/wxl0kUsUyxwj3WRPaLm6yv21sGZ1JN6fP/U/yEy070H
0Fu+ZQBawP0QUaZSVaSuGqd/YsrgOdlqRKm1lFXtVDq8Quct3kNB9Hu5RFbP4BLXadRiwsZJHva/
rUE3CTe0dUdUmxqKke1sMAHrv7rUer+FJ7gRCO5V0ujiUCLYNPJgSjX1A9E1ayZYxxvkUYlA8XYv
D+7GuhlyjBJGlps/LIG/w4dLtp+3Mm6gkE3rCs9SlVpZkSiQeoWVSLirbr7WnCsSgl6ChV89XPoH
H7XAILbpzy5Kc9U8/eONx8DlJCDew8lYlHMIciJHoqIouCTWAtqv5kaWpJdF57efTV/3eAWKF4HU
Kn0RifbdR6NxjYTGwqE4gbHi1mFVYVFUoWH7JN9GjQeLyyeyoZ/2PKGoCT4oTFFI+VcVsgOftI8l
hfnclBpCMEKjhznfjpkT8vstvSIfdrUubyyhop349Jy5uKWs/etATkFqj56XpFTqIG/n1c3pg+Uv
xPLQiEpqP9VSOc42log7fC7f44bTqtyxj3OZQjiRCha2uVfeRkfmHuxYwZGQ4dMtr+nPYwe5HZgf
QNXy0J8tsDFuLStYuzUYFKw+tYNNVWJvNd7OgCSjCyUooTVLTWcMhfQTfrc9hqiZwpbDOhPOxjC5
2l8bK77RLTaKq8aSz2Xl0iKCPoEZp27NR30ASf4OEv0n/Gk5XylcNh6u/4uoFjF2DZxwqHV9kF/x
Y1GP5KxhCzpXK/DfWRzCPtvILlSp8CHDmEPExWo3AirU4u03g6Djw/vCRCSjnmxQIIhkHxAWhnRJ
TUn7Bw9ny8vU4DntqkcJnlsLHkWNGen4KjWr9TB/swh3zArxvzxw3m13bvP22YEmqxEvNFQTnMud
lH9HUXa3MPLJbsBitX/Os9zfm9op9uYDz+Ei/Br+JWkRxPKsE8gVFqSchFRxfqkjEtsQnQUKlrgo
6xeHfFWTSJyATdatNUGpKOLqMT11+0fyiZ87KBZvhKFN9tbcwzmOR8X+ZQwA/LpPjvw4Q0Wq/9mn
1G6qdwjrGTSO86k4FlTzJpEHNvTd0dejmcW1D452hrUS5AHH6K3sBB+R/iW7mYFJ/0Pefnr11zB2
2mUeVuIZcwA44FL7y95HBBYMAN1cchGgfOtXukfpM5TFb5cyBETCf0EfZ2iX0If/hKG1jUlonAUB
AAhJKZ09iGCkIDbSuqdaSFl6LB4WLAFTXv8+dxJaRC/H8XKqXPsV/eS8TJapH8ZjTyMvW5/4NWjy
WCu1T1jLA/Ris53E3b+4pgLz5+IFELWN5ibvKSlS6fAkjBDw5wiKDL1s3ylMDj2AnYVcIh7zhTOZ
2xTzU4qqKRrhyonGFd1VrrxkHzkrW/dpYNaXcQHgRr1Gyr1NYpFH0zzb7TeIjpkKDYerNyY42nIe
nND7xzrl/2tZpcdg0fMnnkBgSD5Tb72E3SPz0d7NtqNGkbQ/BwAT44nErIFMUn2y0Jky4erxqkvM
BbB+1ib8dTIZWChzkPoNeOCSeAuBEtOFvQWTkL7kxRCQLjNZOZqdMPlhBJJC0FkRuWkbCe5xA9MG
KRiAKf3WSoX0BPELE4S8HaXSCH9Jy9Zo5BkaENMZAe1a8/AcTD7+YiV+zgRd9qyKwjX+tZGh0yW3
hXSLr3RHv0pkRswgsP/KDfpRZkDw32QNNwl/wHrhHgGf04ZadQu/FmykflMD4zasLoBQT9FqL+jJ
J1qExoTFTNzNcMNSgNWXVvlIwYQifDds6kwveVKyCezIkgLNQ5b6UZ1StR6vSuE9NoVBF3cHuFZR
RMkcCRy25xiTbd1wv2uFMGLdMg6tZxHv3KFfouCUDxLRUHJVAV8rLjrnZfyVY8R+cBJpt0fj3Xgm
Snj/BjK7hIPdo9zgo4GP8PAH2Mh44bOrU18O2B4nQuI6dyoZKFXCRB36VCG8EumzZ0eRT+tP5Bdq
EYGZk/LgWwbPMNNIbrpJK3EYC7/nX8KPi7S9PVnLa7hPCMrkJUdEPSghw0yBX2NcXatdPcta4EUL
1elmHnJscA+/titJMWIXbkoc+Ff1i0cBM91pDhbGB+aq5YMvH/YLDREdMK2cwe3cc2wKVeHqn0XS
un2sdgvJGad4SwhrS1iQoqA1aNqqc3qYg3kc3owEKCdHDskqPV6fKBcSRBZrY9naLJXPVFLUtfD5
gaQs4IJjjNjScMgyr7vLYiat9rX3y+AIwLupG6+xPbBE8HH/UBAZq/XKzlHSapEYX9WgiUd8g+0k
CMsA5RU5w3CtTZRXGafSJ6gJr8/3iGelz7t5uqz28GrWueTBHKoVUxhX0H/sXChH9Gtx9uh1B8ID
kD1BBMaus85R6kUA+zbqudlD2yV3iXAn0NRXjMP0bYkXlTgvDJgLLfUnBrrGbo4InC7zMm0He6ta
GzvWCgxuURvJjV2LhfmEEZ4LdoLPkIBiEieo0J6aIqtKHG5uXlC82Id7UC8bP+och5/okd1+McxK
nsi7/BrA+2yNQb821mG3CduaVwGTYXH9BZFyjFYrZXag2QHn5tQhMKpf3I2cqg+wW0dvhCme/fbX
L6SfPSCq94nPi2GzB/szzFPE4g0KCIvRnoXXjvVTdvqgRG2AAz6hsiowhm+ZOW2F9vUHbePvjica
YJJwWzwSIjoVWINQb3L52CUyyMiEHwe6d+0p7B6dB+WG3CWiBqUz/lbocQ5tfQ3sGz88xE0x/NNi
PDp4pufZc+q0nwE46NfXMra/HibFYsLf/auJr70vX5qKJKuPe+9ovGZPwJ4rGNGo3EnVzV5NVfRR
thMbGAWl3qHeTbyTtsmFIU4STKHTTHnsahzuaVz+HR9CSU99rE3lrq9bkdikuf7MHewRti9wqbcR
lDHj5WfW+4HexxtJ4EPEmVqLF4KBIgWnNpCrNdcbcNlbQ65/ZqunH6HZ5v5ny6+frEwffGt4N3Jr
6GgKup2TjNu3UTWT54L4jXcfUtgqcUCYuB8EEg414bSVdNBNh8mMo0hBFJyBA2az1DmO2fhxbQTD
SUU+oFRsQ10b+p4zzSWRKGbWjGA5b850OpFu+LqPiIVqvn1nx9dkEd7L/CtiSU6M0RAqLV18lTIo
0FQZKFZTAU8KH+6GEq7btgHNLGifhWMBC9faQ++pcdgrhgJtsMmoDr5ccuuGsC+dJnOUqFe8N88s
G1SDuK29K/qhlwPglI3yB9z554Hf0Ykfa9U2v6fU3G4zu6ABlbbiBVDZapqqODvJXQ98UN9JpN2D
ybaj+7pjSBQxplk8a6nHI3NZ1o9do6Z57Bt6yVWrc9RvMUlItdck6PskWpjMpvNDbRMZgL5CXd92
0ZApK5WGAPVXl0KUg8zGKEcsyGPbnOnBJmEKslUe5BFwqFp5WVGET7XiocuHsUz09SMNhCQd1G6x
14HgaKYCpEu/4Sfn+rJ5UHOzZocIiv1hLhsK+0ONquOvpCCo6ItqxoiBV+QNYiXH2x9A4feWUJ8j
No3mI7Jop7vo+ZuEcUtBG7fNMfpblF17c/7E8Kgrgxgf0OCm9QMZ0SddgmdMIF1eerRUPl9Ihcnt
m+kjq6zkeTfxJ/b8wyEbcn0i/Ozg/+iwxsGsYEd0jAtj10UGAjEizpCYuWAek1X75kVbTkworrNj
nPrhSiC/zKx+azNcFzawfweducjrx2P0+64PFDhayz6XZIfCGTkUctC+iKVI6ME8aoAcGrbd/fbV
icBblCl1Ae+6cQQtEdblVtMeyE5u1/TClTh4KbPK57cP/9jAyWAIdOeuvn38gXMvis69dxZ31IRg
dxXiEW9bpf23Wcb/nEgDlkuYIOm459BViFY9yF1yjhT3lPjrtsmAUY8mhsMpbIwNX6d+27+uqsOO
tEXmpniBhQr4emhSG7jWTdIYWEl1yaThWFXz0G4PTx6fqQBVC0/T9n0hNdtDdmJg6Rc5e2jRJcLS
s517Zll3YZhTpJwMVxClHD1QUf8znQHp41LPS+VFyicjbfRoUo9vjz/wfxTfXqmN/EXoZ1dqDPgL
GdZIkVpVOQWDP9iSgojlvwb4KoIk+QZtQF82+4v1WzmGhHRfNN9xLU0KWxi0VFtVluDTRUY6os4h
WoTAfB5ukJ/f5yg6oxwmOIyhEO+mw51mkXiYJvtk9twL72CzvdWn4Utoj5wrXJkDh8Kqui84NYiI
OWfnvwBsbMn0iEOo5Bgm+ZnRX8KS0711XGHAsZbOwOi/RO44aReIJPnHJSQ1iPA+SkaoT8vRSJI9
AZSKJduD1GK9+BlM+CA+x3njVo3SLLfNWCphb9/giPdhYgJ2H7pegPQeAGdqY+/Ac5Rvg3f66fsd
/7TEJuhYrhswJQ9J26NQIJjs7hu+TAcNhZsQH8IE9W/P9YmE8taLQZ4lewdwvH04ktGYGDOgG1da
IKVCjqqI1IwKoNd68rlPOl9UBNN2GVp6A5np2x+kSrXHAsAYQwBp/5mtChxUtmZHZH8blVRfEf8f
ZwpR8MnIGHLZ3JTrTg85Qsk9i+rE4Yd0ZuK6Axluy7ciah/Q6BMod9xrqFlPoz/LZvylAu8XbIgk
dveF/y56A+wAafBW2+IRB6uMgWOyUCTzp52C3BVls5Kio/cy1RO1wellmtvW+oeRo+2bqZRd6GWY
IOXQBawWTJTz6/HVHi6qf01FUIfXMkSFj2L/FYfG+DwFieWnUS58aZw7bzdg3wcGgZF5TOb6dJka
hPDuFsKA/rVPvA1BF5UnhfcIf3Ye9bm3vepk12GKvvmNriqWF6CMSs8Qky1VNr1HMkjoSXHmd2Ha
bkltao8A8i8SRXAnaYlrA2XSKZb+WsGxHSl0SyJyQ5y79fL76CpaL2AAFUCuV9cgonqMDexelXSH
XdYgu1aSrcO0l41c2y5NZ1uNIJ5W0ie3opSydtKWXavnW7L+4ljxZF9y1Yz87HYe3+OZBEJnQlI8
4O9xfLJcHR4eo38Em/hLMWuY0HvSJX4UmE6d7a7GPgBWXGz93+VFwa0ovjxuHIGvDvszRUEWjo+e
XSF7oBtuR96b2EKO0nTzbwB537bGCgGvbpXds3Bv7t29VuSAUBj+mbruaH1RvhOx9poMdjRkxfLh
JA+Nan84nRpyLmwbKQt6g+aqfmJYwHLziy7GTQBjxOzmZ7N2DA9WdfuD2ZS+XHNdk0laBSwdQ5sH
hf+2WuC37jx8NNbY01Bvf5HTX9wtjaurvOEvNdGvWuPVpv5tQB/2LO5gbJBVCtmTqzyxfNb5v7y0
wU7NttI0ZYjkFulaaIgQrVcutez9OarFMsoxoe0VjSUa6FPm1iP3mvS4jRNso0X22w8p7j9M7zux
oOrtMUGNKUzI3dPfeNI0m2+++7CZXvD0wLDVSN8WzEm26m7P67jVOcHHERmNFNSINehXMneCj9yL
1BJtbcXVsoyksAdo8IsiBSgYhkY576Sod7Hkc0+uzDk1EiZ2eGZbIjp6TtqbS6F6b8qZcKgfeNpN
DJbIeTwEOUv6fZoI4po+Pkb4OhCRG4El9PkOIeOOBxBmmOWA95Yg457n8R7YCrkweVBpQ79zmBSs
EzbMeA2dGSNGvmmgjy31i+N4jKFcD+3CwNBDnSp0IT77Gv/US1EZxAECXpdsgHEL9qW9AYy4Depx
yhDw7kKkuTxjL/1gDa0xjIKVmnI6dhRBo1QOGJTMPkKkVp4EUS68S57PNX4UbUYj8lzSlMbMEugd
Pib9mdGtEDCf91ziNdICgU6Nip8xJBYxL+OVd3yVkySf4SPje+f5w/s6H8vpV/PYdQoGaq/8Zb45
8P92KtPpgaxiiglZwvtqvcjUg5kc2Q1l/eXQOZ5e3XO5anzkbRddlGAsDCVfSQn2wGwhtODzbGoI
v1z+lLaquvCbkCc3/LqdQ7W0dgt7I79inATOru2JdtHa1un2LTY0iZfz77pE1ot7jK9XvdeT10gd
KpmEkiSh98cy0oemdt7YS2yYz7RR2EVL+yWsewORtXi8HeXO0F3APRsjLC66r4OdYR5foANrLuog
DOPiVqKr9XFvNjAhfbfYyuEnDmuqBp7m3o99LD7E0WkjoSeVNd6+7j9C9Zp1UzTgJUFfUZ29YVHw
EGlfKoNfz+HrSOo0wBLiCPWTy4iQdFfCr81jS9nrKvcZLna91yMN71nRLhaQoGEN8oCpRsJr5VnA
mhTmbQ7bHIhCSYgFhoAYudqnWSPEFdgFLEkgggbaHPfvKdtE8imcmZKIxzK0Vp8RKy7uP6QzGb2T
XxgA00YLBCdGx6G60Orotm2+vVI8YyXL8LgZOgyKmve2DxJxDI9ntVCMrFOFfe6y6cQwRtlde4g7
yCp+V2rQUdujW/I2RpGzxCQQo3Ca4rUJTO7YdwE5FRMaV1pa5OwiDyoidRxjZhsTo3YU5702uzi9
Si2IuwV2vg8HRVkhaLGX5f8x7Y9Ju9fbTqnQk/I2FJSz+o2HVcgu2U8KWMrHPCcDCJBq/Rqm0j37
Lf70AGX2f23KMZ5bR0lu8Ydp0u/LV2cYMaPNRhrxHJKLjhE3MOU/NptCzc3UkyZv/2THcE1XPDtA
Ths74aw9KScrHPzjzRY6ZfuR4HeMPLEPwhtk6Vaw7XMwrRFNz+CnNkelNSA6iCJLCDjoQ+/tTylo
ePg514DcfIdThtcK12ZukiYlUOnwnSS/FMQLzRubkriNtIyiRDSyFb2W9mR9M45mtj0KF3xafgn4
jTXjjkYOd01d78roS9e50DaxGPEIwqRuZV1AiWsRvghJgCQiUbDW5uowREPOGWxisdc2lqIAZq8Q
Srb3Tya5z7hog3bobZB2m7vuhTfK85PcMNTqO+LjMLndwqI6BveFF7+dIBC2vMp32ll3p/XzltHM
i09wnhMncfEBrwNq40o9CKukD3sIt1P3w4g3RAhe9nQTFFT3lJ0NUCxxEhmNGuPyevfPughx0Rl8
AXgLQPYN6CdW0o5w/BoCiyiheLRmgVlNuZvvu0IiIJaEhY1Fk6rYf6d9MB0VxIULCVguQZF+LxW5
Xax1Vq/pkz1gC5+VL0INEtRBt22vU0V+IrU2/rWpaOtv2bE5xkdKxBZVOjonBGqL2j2zjbg6GIBx
+qtOl5Fk5dDE0vsjNBIwicqk7vnmlkhKk0q+LpXp4Ghpa3GiQHNMUng+SxQFmnJ3T8vQJKyKgFds
oevQR5njj8lzRXHqrgO6yPNNQ/fGRIb2g4G/nbYHkrqUuRUUDnanrrZlsH/4IJmd4QKFqgH5V/kH
JTdAF2rteGpYQ+HWD78IO9+J2s9aEnC21sFnPVgNm9Ov+N2Oh6TPFKZpIvsKCtrJmRFpm7jY71a+
/mJTmIKbwrUlW/U813YQP+L/hDw+4o9J5klt/Vt1H7JnQRc7g0Qy0g4AIxCKeNxCPFsnBlxNxZbQ
+h43ENeP8fugbw40GtZSfGUs8FHKkW5mLm2dlwoVxMMUO4BvTwsFgKSN1JzQhRvUtyayKD66D5Ee
/eDl8uXE05v8S6e3QRP4R5YXQbcU68ZA+vR4hjUkopztuBZAY585r8ZS7kfOCwFJREShW/flSaE9
nlA8Y1L/iMlcVDw1/tE2Tm/Ffjk7E77RRxrbs/X3l2t/6n19fYLfAEX301ygqwv9kA8YGr/dl/Db
BeF2mDo0ffQnxKPwgzRGh2mAAe8spbKqM46yFMJejXSNQM9KJBQf+u/KU30Yo7d9TBsfE+sD+ZG/
RrKWjPKIXEZTo6rKa9ExdCUA20gEfnhoomeGF6u1g6h9LLcH1hcwm38sPz0aSKQ8eH2z99UQb4zK
xjxp/oeBcpkwnESvx+8cwGiUaoR93P3jXtCbbixC26YuL29bGr1GPtx5s/Pi10900G7vpykXtj93
i12zhGyecwc6gK99YuYp5Ii+T5XEhbvKJlL3L60SZIpAXZvJ1yUdSwj2f5oJqwy/2YMXiTuI16YI
T3H9AzWK/PgbRQiH7qMF9EZXH9aXqZQLW44BnCdSBzBXeFRGW22C3IoRLEss/mXxdLouQPcdhlpm
wrcUUnoiW+vvc2qEKqXT2xb+TEOxfxJ+vxFnMlUKw8G0ofmHuhHMkx+HkEgwrSGFWM3D6+EA0Xh3
TGPFTTyTcYN51KSCzxakEtPpOq5raeN8n+9JWkrqWnFW8Dweoie4Qwb+Cua+oJik9MUBvV0rruPU
ktFIGbILQ/sXtOaX3jeCi3jcYHKo0uvzjy72uEerGs6IeoXBAHdgNRdHa1NHDIrXrKAfw/0efSLK
L6hxCS2MhllgCwCeeOtfG4wP3nhaZRXKy4VHtcRT76mdHoyYp9XsuzlMaj2lrNgQc2JJVjr+HmLN
p5z+SkEiFbH3SWPoOlwuAuMRCf7ye2mJ1zHPX2BRFcvTsU2YhZ37C5IKWHW8x49BEGu7d4jXyhSK
uReifkPw5AwQW8CKleO+C6xKO0T4s8ANdumdN/tBHleu2CgvNs46oNdQbnjwneb2JRJIpEqbVqYr
FyGjhgWPlhohxI/QApQ1ecSrk3JBoPUVecTh5AsAE9jT87WG70o06OMzyZvo+stNpGjXa8+NiORb
dh96oAxZzDC/E2/6U80j2FC+NTxS2YpFtuGQsI+59JpCTzaCE6cyO062VLFxL687kEck1Spy+EbV
ZirtVp8r6uNvH0uDa+LuIa4XU71kxZn3VJnM3ppQMQAkMkTlde80XEe12pdmUgGEDkj6Ij7ZUsBg
Unp6vzTDoAznuou1VCjPETqNFs0LZNzeWaczyK81suqmVTqkUtnIe8xGGyr8KJxTpnC9F0rxg2ok
7ngW+etbw/DoBzZU1ntOlE/XiCyCVmFFKoBOkksGiQK6H6R5pdz+etfjcJj/D7G90kReuhdezlTl
5xCn6TPbAbmJ+yZ9E6Il3KlGZ0Z4HV437VGZKSv7u5a3sgDU7nh1jPOrWIR0DWD6t2LRPwU5sYeR
mE58uph0ELzctEc/j7y9wdT1NHVl01UYNnyBZ5zg+OEwfPS3/Cil/ffzDfAvLbSZLtak02HYi3eb
we7f4TE06UYEk11bqABE18DJzflveI1v6lVc/199OfEcviJ6UCJmlT+f9vklpyqar/myWtqX1PPj
AxvqPI1F6xuNJo66EQegl2EWOpd7KnpnsccQWu+JgnQIn+e0zP1oqSTQjTisYNGE9JB7oZslciZl
vJT2WuFa7qaOi3snuT99WeQbAh1/NBMX73/AvNNwokGDc92cPjM4hWlQ6MDJewxEfr/S6DH4x3RA
PHBPsbfG01CMbm1aFWvleAJ521KUtCZ1oucB655lg5IwPrNXb1NQVhFddba3K+p8gSI8P/780Kmx
Et4rlylbpP0IhnawCOVn4Bi60FgUxN+A76RMMQHuKDTNvL7KDfz5go4aLKkr6GR0dIhuxLhu9gCe
D8kELNwh2rs2yAfi0eXcJWvgfOtCLksGeMc2PgB2uOqJtlxTkbGBZ177vd2N1rqhFm0tLQ4swb0B
nJTf11ADj2v85U6fKoAS3QkoYA4cIfYz+UeFkN+dGyotlH6/YxAIkqFMyayoGRURamQrHNZdb+AK
iqJkrVEgoc/dYtNGlyfB6X4CxGVK3JG4IgE82K18eZRxAoOwTezr1ePIz1WIgevWDq5GnFtyZNdb
IOB0PvRApAo5WdVzU4/X3aqsQWyXi8lx99nMmW44bVpuuhv+WC1MtjG+1pFzO0XVHzXgRmRQB0bw
iHxes7WA3Vy74YG9oNSFa+fipQncsJqgz+QTeNef50MgkF/an1UJrKqfkKzIxQ4CsIddxTjcJhVM
uCDwL7BY63he+uC6BgkF596ELK7hnv4j8M+1FBlwRpG3WBG/zzvzVWllLdJ/QpeqhPvy0czWTUgF
XTH8R+XJEy8gsAB30Rw1Tk2asX18QIV73O3Xs9uVUyAsWC4Jzh46rT1hFr9x9IzTla8a83x1k4c/
B4hEbicg6pOu/aycaieEgg0svgDUn9JQ55yOu22PogTXUEvxAe0iV9adNd+20MBbumxqtKS4jaw9
uA1daemcHCZPG3aCunn0PbLO1EibL5VU+ceYvvqG8upwLFYJRjpxatMfp7kn920ckYQR07pzR5RC
aYfWtxOcWnvMKGQRnQb3qjJ4DVA2msfyOE2UhdGMJubquiVKIQkrL5IQOWAau48aKjr++/lcwaNt
XJ5UHaqTnzuLwqrN5E25nsiwNmQx6y4zUPIKe8cOgakelsU61+ZKvPNg1Vk3SxDrb/HP9oM0uWYU
n99hpl2kT+hKyPragn0N1NgFIoSQGRDd+TQ9bskdQ/r9uKGRWK9YvmQGuN4Bg4ySFUgxIGt153Lf
Wu6SvWorfvsXATo/2oztHhcXx66+uluYd8l63FZXT4lnCiyyBTWbR1z1rIbhAVtFxUoVgjLBPtiW
yAoRqVIAbYbaQoCevItav92pI8NIHpkj2e3TrmvkfzOONdTlAh/kHdd6i5ktODBo3B9R7msN4xY0
v7l00Cmy2lPjc32gmqVGk2yW2dKp0cw6mnS1kpt9BujJTrbOvzT55KB0FHqYium1PiNyKEjm7gdt
B/TuNQT/sKiyJOgrraq+drI3eYL1XqLZQA80eJuEQfC0Q556TNkd0lO346jGEvZFwJOGgL+qCP1S
B79aDMHYNDwYOe4lXMK5wyaOIee4ZMF9I/oIVSvZe9rZDb+8Shehif3lkt3MyY0WHDhKVEVX/Xvw
IRGOLpriBGtKBKVIPhup6FStrrW0+A7sJ6UFTc+V8kY6TnOAqL/Uhezix8CXi4vXz7P88mKw6TTy
vJAjhmn0uv4IYHe7pm1PJo15uOmIyOXneoplqg56lrqbsUcc9C10tlESy9FTCZ5nyDfrbTaEH23I
l+rFm/XU9lR5XIwS0JHUZqBBtUay5aT58YsZHQd0YfRn7MDqA0pi/Jx0XU63MmmfQAQcV79UjjeR
FS2yAJJ0K7BFIaulov1T1NP+BlDALwihTNf974/G8zS+H9pmpv7PDwY0ix37wIXDzOutBJkC+wM2
oB2F+cPsGvHEOakT3b1QGMQgyCWK7Yb9LENeoO72aFi40QoKdCeid2OzbofzfYXR5Z6ruTLiCKoi
NCwROxiHAGO9NtKzJ59n1tiB9immW6R5kUaOPE62WMYWgozksvskj1mSNiDD3smlZ3xoSUNI3M6b
iexgmXQWoxcYs4wTTxBvfZ0T0q6pE7reEJNKUW6AamHPLqZHmFWQEAMg6IcgJ7hdYDRISmYgZOkP
d4VzxZTrVKiFrnHstOkztPkRjxcpfKFvt0tmANQuMFs4IhOeblnsSyRK/i+KvJBGVx3dfSOnFFDg
lwhCRttE6jIRWV2w3kgSDiENwj+dOHc9svrUTXrG9npvB+yVfYVdpYlhX/8+BZD1DWFCm/l1Si7J
4DKopZ+FrgXDrftVg4STuDRmn7OBpvCY5MJIMBuX+RYLOk3mHH6qix/T1cHidKwOm726sR4SJIaA
MqBgmb+pTU54/s3QTu92pKdxAOmgKuK85rJqU9ktivRXCAMBeZMzns5RQLGKw1UHMKa3xtWS5zNj
MYQRDO1uB6PWin7DLk87XnQTibmKIwLpWqF+isExO+pnuZJ4TssmYJpKu46L8hVoe08xF4XNVSCM
oITLweq99aPspbFdUPDensiHScTuIEEjavRhgsMftkxuhtJnWlrCtt9fH/hLMCGXJmXom4yao5hp
Fq452LA9lnVYpySS5XFoupw7cZr0jGgfw6QY3ZPwIAL1YLpa0EDhnh8YbPJQ0xeriy16wXEE0oXE
d059/Ebx6AON2u7XRbXCEIuHaxU1XJ5BEkP0PUEv+YOSYAVYrmSQNXklph0cNXWPyScFKupASqAj
kkHABployWneYUpFFL3xCXMvlC7IxPmwSNrf2cmgurWLpY6R5WG6NQLaPqf+/LaWbNoqUiISrC2+
eTj+yRuth7nu5kiqdrKTC1epIES3bJ8JD5gZNzv9SeZuDYxBu2afBXyKYllwL1DV919imY/iDtdo
Rc0Niq1dNMOQKLqAythbhEugg4v6DuBjAzOsLmYD5yFsYyehEcG8dlcq5TdAuHhmB+Ng7gxtvNw9
jLxVibnhmU58dgAnX/5VpiqYKpWEAtwf94AAJOmGekoAv8cZ4ojGTeGMZj+PzOXUnmn5zhTVatDq
dI++dQxLXdo2TXaf8iZX+4nFwo829B/jtB7+h1tUIpQPOsNfr2Kf9Tdx6FZtTsS69WjZ6hXRKxxg
T28VgwMFXdagHJH/b1hXBSXd010aObfcwQK2k18D1Y/jDt8CBLa4kU7iQllwgnjTXui8WkxNEA98
xhzsr/fKFFWVyHVUhXxUfHMQ8EpLbEm2gHQztrrtHPG+PRh9NHP9zeqP03G2Xc1UhFUgZmi5RM30
wkLKz2opA0Qh9BcLuI70W8pycP3yJqh0WCWFyZj3Cl/3mS5QyzWad/Bw8dYOmdJmIfBttoqUfuJZ
yVt779PQJTmT2ir/qoYtLvnPmXkGNqzeFIr1+V4MYZzF/6pAlsww5Eg2sUQ0QRusiXpV0s+g7kSM
N9YXDsqEZaq24m3wpKRww+GDD3+xNkf502r9CLEeYtpWXlAjBDicFYw8l+VDxJjWx1FOFyI0gjDH
/P1zerOIapRWMVCWEw3NB7kCkxGM6EVHwbq9tFSXZDGQt0Lk0UIpZDiipSWQ8zFFgksXjB6q1sRb
Xm1HrWV2qY1juxZSNQ8dllOrdkicppB13KIN97S4TYz3E4wHkEMxvlvgWxyPnupgHLUMJwSovJDr
tHIZMdTiFlvAT0OF9DJL+mSRIVd/PnM2noNxGQs5R+G7xC/kv5ZBO2jAhYYdjJwrbhnldM96HZVS
mnVl5BXOTeuAcT4q2bIYjI8ezTAsh2Vmrz1uPmyis9CRlj5f7f12me9wJx1o2S7DEDv4VzMdKRhM
w3i3jhzEBjwh9yohrz9bibKmubMdyMR4AhR+NV342gJEMn1/SZdxH+L2EBD7QhAbIW9IF0vAS6uM
D/eryk4EmlBbgYcdM8dpqAXoAgymBSiBdvUJq0DZDXjxfQeqntkg8/1WcxcIs/Q09zTvNuw79Jak
9aonpXSajFHZxf83LcvpYep1lvrC479eCLQ+yvLXBxqWblBgIgoHp+HFk4yDE5IlZYioyqtre8UH
n82b1IIPyKijDwww3KX+u33nrGdpeZHoll5ah/yvTn3c7LYi5wZuxZFwwrLQ1KfUPoERe3EuHdwb
GSDSxdvMlSawaRSMyrlHX7dxJz4uYfS1sare4QilkcOWps8BFC4qnAj4o1uSHUyEXISNHQwGdu7j
nxUi3dDjBaPsE9am7iLM4xS59FMcPqOMB6eb31/P28JURJvqrdL26lpDduW2RDUiOkThktJ2T2c6
AXVus+SlTM7tjvGeXYqSl/cKb8R3A42lCf8f+3BGRz11kgNQob101w/4jt45zymkOmioSEd7BJYL
FP9cSU8ZD2eePE/gpNtEoK5Mr9tteF+DF6bCHmrzfYru2+TNXPhZbORZ9d0hO7APIaHdczOeqFMQ
tPPage9WlJYBVieVZyqRkttZ0Peof6HspOIZy5/HB5YlLMpiJrqjeDHUMr2BW1v/LHetYOafZhOX
ahqQk6bwLZNKkhHx15ykyDmm2xJbKDCxFiilZ706rF/+ktYyTLj2lhL7d5UCs+sjCrTifDTynNUI
gS92RCPCkx+XvRmB7FDGgefIXmssbQN6X1Y8HoqaFdC+cA15SUoJFnjkiYX6Rmu3celrfexfobih
i8E2DTS4B35wDt1HeeaLEcIb585+9DYIiigOyv2VwQuO1mWMAYLtrfYSblE378hvsLL0KpVw00yS
4YmtrpwIghuuAAozA3988wrzFZLuN429XAKfSQh6dLaOXIcaFw8rqaNiel0vHcxR30QeKfojhTYw
zAHxWa6ppBScgpJpIOsn4c67j9Ygq2qvkfPRIQwlqPcuTypXmKBGA/F318adHc9mCwJkNPuSFzP5
SCmY53sR3beF90Iy6p7Y77Ztq1mtNU9eCDPRfsAsD0oTtjltfNnptxM/MBvDDff/9IytBeuvxONa
r3hzlMnyeZRZyYqPr7nlQ/WXGPDknSU2py37tYICEQTVPp3SA6LUXFfuRo+LopuB5LtwRiEL70NH
0izFZ1nh3x4ZC180X7PGfC1JiSYZo1B7nFnEMsQQdmM354UbCzhlg5at2OkpMwzFbRl8ey4B72jS
0ZKOIz/AM0cXTK+jKlcy67K/Y1guz3trVJmqEAFrNnyufPFOnP60LyVOcdJk48oJDZ7EBk/oet+5
pAremUNZ2aYCD/lESubG9+ZIC6y7AgxtwLlqYcyee+mhUiH5P9FF9zBunaH6r51wZH76apZkQUAb
qF7X2U8aa6C9sQ/1NtzcA2AA2+0X0pkmoJioCIs4kv9bNTMJ3v9nD59n9jZXVAj28uXNPtX4Irkd
3GBic/IY/4jCIXSXflcAspWZyM/h1AFsFSxNBJLvwn3OrUheJXccEaO84jA1JSXTtcpcF6ZQ6/W5
8O5JqEPgp0R5OFuHhowgHlp+C1bEGtDTotyf2CTeZVWmqWLbx7YAaaCK36qfRQVXGxQqGenZsikj
qautww4XR4Nm5TlSQayZiV+iJAYcH7oq/nZDIUpNV009RyEtXsuz12liUIRe9hY3pHxAc1WfzSP6
z9akQZidNmcM3QUfBhAor5ff4tcd9fHkUpjzK+5P7I8OZ/ztBQkQVTwX48CbxXDhfs5oSZVOiC0z
noGDu6yafnEHeBXDRCMi3g3Cq0lG8B1ivhp4ACR5cw/J3+dmEkUjR0SNCYz4MK7vLoHVBNRAxfEv
s8kK2jui528iLVIO8w74Zc8RxkmfJOZ99rn3qKyw5uY12PyiSd9hZnC3NlqR7QWyKuDDIDhMiwSY
ECJIVjNK+p53YW16rNL2idm61io9sYFAk15+ch+ATIHxM9QooHS90hqevbv5+A5ACzc7NfGommvl
9p3MP2XtuSfN2WGtdLa9gGFlhZCzMnBVvZXWlAqwWyPrUCJU83f5K9nrWcL9xh4IqJukX0hiqb1l
3n2x9bGv9cIAI4hud/eoXrRGppmJl4UQi7ZmNvdGIT5EkuO2muUGkPMZYBYb6JDC2G8j29HpNIRe
iWCkZgzNhYPGeTmEHED66UOPIltlW9By5izOjBlUgQTwZ15p9nezv4tmDmGq+Uvglcxr18gd3vAz
ZprsjwwQ7XyXW0RYBNP3dAJ1a5CvALk1yWUlmW/h1Fs0nVxd/rIbbLwIA5uLC3NEhIuth/IbHPPV
JWYwqJNTzTqS215/4jJb7RdZQQUv7g+dYQ5G2hTIicGLFa8GOzUKP72Fwmse4AezzzWf/qzhaRvq
wm3RT0v7g3ZJdgkoF7S/hBDQvzzTuT8ADYRMiJujlgjoLF+X+xqUk4aa0xPYBE2EMhrV+m+Zo904
HbUetOz5XLWDVmm+GMZQ9rkLBlcHLOMDQppfPdim69EFc/uHwRnsd9E3SdTucycGQwvBr+MZLzmc
EY6Zkfw+QDwXLjNoYzH/JNWWZB5lNi3RfSnoY3ObL1VZbNR1zDP7oJvs3OVXehNnK4azf3KitJys
rJ8MV2sOXR9IL2J7UVlurj8ApOqYB/6YhH8nTJsqM8ajYHFNnjB5MV2CoRtW5/iIWgp5VKIQ0fWb
e2Rb32sNXVxFJstWH/2M2Rf9qcdAdhgCqdGtcpUbT77PNI8fm8ryNrfZA0bBF5lzsVJgxFcpuD7k
jLViObZypTgkJkt2gOWOUCDOPNtLbqRwVtR0bXKfZEmhv7z4lhaRVV8hxOtZzlU4h8FS60bmtdn0
sb5AmHET8BjQjcDLNiwdfmN4nufoVzYegc/hgugAzqLJ31QAFa6iOL9S92IDLXm+dSpSyVNzCsXv
BqnL97t4C3Zu8WQo8uXh8owNeJIQ/B72XGDKjoPSyQztlzArz+BIeHr8MMnKR+GVDfnNFLVzcyxS
t20Ukkti4Fy05Xo6iGNEneVR2cb8tcr7+7Rr1zQZgQy4xfcrOLvF/Ygh9M5LADk04T4AJ9Cn9BYX
2j/aT1bLWxlIn931X9Xwj40Qk/jXQm4AfGJmbHhw484g3sa23sKam9tlq8oOafTVBLmqrfKtIESO
Vn4mxK/iLgtl3ZnzZ95HQFPUcSMsy2RZTcijZQhBfhGoEXWCpHnhe+VQsFdVJz0QK6d2h0gPxwsD
KWBbh8rpo4TKcU6syvp3EcfihgTsqHqlAdBAWZSNSdB3VvkRUg87CxA/tA+jCgZELDVn5hXs5dpl
6jIHVBIk4F4Cz62I7ml/+XK6oqDm+l05O7Xkab4B52oKEfvO5aUd16VFQBkVRM8Jb94oW7KRPmuM
2tQDUbXyVUOViQUsCZ7r7lxlqb2qu4XsVCX3yCMyAqfEXK7ebwZOxZ8SkaGJ/Qh+peijtOByf66S
UMxEF1SsvFR2qown+2k3Y9An1wUVYPXWao7oYCxp2Cs/l0rrcdguqLG89z6GeOF2p0Bgltutt+ki
II7xj6Ozb6djZnBtn/c/zBcDphToO8rn0sE5nZPCMFOi+h/6159A21+m0k/49JTI9tZ6p3CMuSpS
DXhCAGHfMQ+8DK1xXVcvWH+zzaiGzNDo7B3qKz+Oc8ff0ZeRiVVGFrN0cIeIgPBA3oI3ZWHLixDP
QbC6Y2rZO+schH1Kprd+RItzQgim/4a2UgDn3xtdyvd4upFegpChJWR/oepVvKMXDMxpyRKIb3+U
+EjJGVJq4AphHCUouiWFbvXuKCpG8cVdZ2lrPlnG0LeZ8CDslYcSaeTFOqcnh1r7ygU2jhi9Rv8B
qoYv5vDb4UncQ9hX62RhradKE5c5eL0fBF4GUv9+LSXVfhjW4knUapMD6K0U/67+vrcOfoQOD7Qm
On1vNpro+i/ZM4xQdN8WGyoviCmTLZ2zJyEIjl6cz7gd/zqS3W/YmKH1CJalpTAz4sCJ62rAEA9Q
sCDiZUtKxydgkNLiPt0oWhHZ3yb6CdUHXJMoo3ytBRrtiSp/XXFqhqDxDZmJj/IjpX7fMBC92MwV
w1yjkLcAQhkt3jO3MHY2s17x+1Pj3WXgUF80b6nGQ8eQjLJhuJUSTcxztMz4PUA7/uKR9ua2fyS7
nfVL0tY34KNTVAdP0lzHKY6iYA5MJ2NglxyZ7YUujUP0AJJMe5DZIkJKCykbnjW7ByAqBnA1Pho5
DgAuj96+MsGPv4lzVE95hsxmYGlTUBJJ4eMcEp9kR2tclzIXoiLEv/BEifrLs26xN6C2aBD6SFC0
Q1OkhI1g7Pgkb2aI049ee4ABYhfubZPkeIqBkGM8aF8RZ84XM3RriJ8bXa7if3ep6dM6ETHu0mog
9llh0OjR/9lEGWTk7XoRDCganOolP1lAPoqq4GmD5Kr+RMzgtkbZcUAoFzwmsAtA6Vsq1hO+EO81
Ji8OBkDlNWsGXwSwDYKkWtJUsxZJv5iw8hGAami2QX/LbiMhyJOTiSXmemEw5VWrUoCwWA3EjWEe
ATf13yeT8Av+fN8C1lTummg+GK/ZLthe94JpgmjnRHQWA7Co+K/eYeQDPQVIwsJ7vJHdY4XYQFSv
w0y1lZc9hV4lsPXIGTHshVsO9fSZoJd0a/akCdf7xnlxJ4vScn4msFSy4lcer8QodrQdd0b9LJoQ
Vv39gjA1LYHouKZElIZheSx4HbZsjoSw87vON+2zo5WGZxW02QrayZfYiRPWKR1Md9H0VVQ2/erk
CqhNrufDEGdSMXvnVD2q4hNJ4hnEXKwywgUTXPOmteMMCwpY0wcVZzjGUHCRH1F86qSClGUDcDIl
RDwS2VXdBCitVhmOc4dFneoPApxgBZWQu/WsBo8PqVN3xqiT+R5kTTALCQ0Zy4jGuapwpN4Lp7H8
5o0tXerakKhfH23t5N14caHrqpI7ojBfz0QQxuFM2G2PC6ZRBe05dzYcyEcJkzIqsbnU4kSMsfZy
wndAEENO1fRy26AS9BNnOu05vf0G4PxsK4NcfX4fkzXZ4QgptVG/8+5cxT4tED4BuS+464gLAPX5
4VskuDwpBK0f7zfGkq2lNNLU1N8QVuSeb3JdosPJxgEqLxngyN385ByhKR9HdqUZKkgq1HyvoZsZ
XceN+uaxShHXqY6lPl/GgO0j5b4Q1anWtXtmM8VivSXa2+iHrsghzRSzD9zvA9ZA5u+CRqoZUQdr
4ljB4h71OQ60KCmtFyHbx9jSt6WzirLUcCfr21m7VS/sw/2J61OViPLJQuYxr/gUu6+CfjDo3lok
PRstF/f9U6r/Y4zaBHQSp9bxvE/ZppC0lhUKdj+JcnoA15j3a3aQ4QuvDoNth3apOygw92vMiapN
1ChdjQexG9kxOt0UzsOsmYIaVH0H/PDANIF/WEdbfU408YQj7jy9dvsItWW0RrvVkKHfC2jxU9Au
gGBb7ybQ3zYvj9jYc3FazgrLkdGOk80T2lFdpTAmP5vA3GiJX13Gy1Rc6FN+WuSmznlgnRPGOD8S
hev6c8TbCD3SDfpG/k1TdynsXmKmffSyH7uNz6hspdT8ujmMcRSBRGlPZiNfHjG91+dpA7WKEXZh
XUdMOYnjbTUmVJ7e/zYHVFFldpVG94cij1zWtyZFHvfmExWN43ycQ+zYzLn+UUO4m8Ysx+2U8IkS
VPx9kGTkcxoiam8iTIxwZ+2nGKLxNVqxPgyAFCOK6+GpmK0kDVftU38+NM/s/4dKsWCCWWls0suv
eDNK4+79a30BOekgZ7s6wEwk5i3AX0Sg4RQ2J0ZNkDtROE0vKqWwbOFN38mt5ensQXDZm9gBdpxA
jBdRAJ1s2WSrcpIyLpZXePBwkQZBXuhYFag3wi0li0fvZRXLz9j6fjUt/6YbGpht3xsNbOdXK/Yx
jzn9VxBEzKV+gG4+699QR2EwVSKHwBV4scZBZFkmxd7tSmXOrqzuh5T0rjmg+QEjVfVjjKjuu9MS
NDsc+Xlx728+n/wy7QgOYYF/EFe56wYzw99Sl1aIw13U2IiilWVkvK9TVAVsQccqMeDUuwx09XUu
DhWtB3m170DhSWx7qGyuIYJ/agYqGMuB5ovrrUX3t7h2F4OfUDInXDFyoI9oi/knuAq5B1j9MteK
9b6shsLA9QiMBI86M6QVHRxOKgooPmyg2PtRviZ4Ebx4mLAcH26WxAkv2t6kYMmpTcSy0gJXIyAi
ugt+hZ3potdirCp4nyzr3kd/PS5GnyF/7/duR0jBJOj7w1B47EUkUjK/R9zU9yENUBN1Vn+MCB2h
rUCWgCMrF4ET4Cu6nxnbpxiKkzlcLqdTDI+W/Z1NEBzYU1ay1DA+fvcV75r8DcxvUe/H6y91/mCf
X2DOgDPwGWglt1zN28siMbABgj4Jpnd4CehGpqkkQNl5gBfNkK9/BCKRUN1V0rkou/BeDd3KIf05
oGzrb2xM26umOf+Ow/Lierv/AlpASGzONor+aqZyVMQZ+pInmpJ0e1jPxgYOcbInUb1qjZb5YChz
V5Eitqhx1rV+d2zA9y38lyuO0QjXJSC9wLcuNXEqKZjxtg14nyP29bpNpTS5PaYfMwFzl386U43Q
yUlmyG/czb26BlAtCfEJAio0zWCxy62UZuF53SfznpHRRWgykiHeys+2E0PnjKiXCvihJ4HSXvmT
ZYddhBhVppH9856wHhcyVk3HQobDcW7JNvdZnc3rQDfB7LFvT5B1lrS+SqB9D/stuv5E9jGDPB6b
qIC/BHtYmNQFPdgw4z7hMO2gBF+G94blHBeCHXwvk4hxlMWoh1HGRw8X+SZBkHJsjihpxTpVFcJW
TcogCeIIqZ2fs7iWA1iV9i/YdECKq9YHtgClrdd80SLaNR/A3w+ttNYZb7pnJU3yEbFaFQxvQnPU
AMOAO2O0vk6PXG4p6CwUbKMNUkHn//f9IfBJJfeE/2KwsN81HBD49Dz+Lz7ymoku6pR/aVceWwwO
FKKSIUxpiFUXch++5MozMnhL7ukLsOejjdG7aGmBqp/13C5nqbljn2k37g4vSylc1B16RMVPU3iO
7hwcmxfXK7nAm202QDS/vYi203rwxlmma2xgJsaDFnefGR3Ey2FPzprIqXdQb0dkjEWZeCJTKjy4
tzdeFyd+6VsWRChk9xEIg/VdoAt4CL5YmrBs8Iwv8j7C6NeQf0zzEaU3tgdtEQiaDbS0l389YaZa
ndmSsWyvWftp7MeFpTaxKy8u3ztCUU+LFb6eDCYI0AO4cyzAZjr5bepdRGgaywf6PmGdqvvFuhql
Xlb15GQWlQkEdqorllnFeTeqOoACrgE/v4gF2sG+IqBIeorfKn6g6hbZjPjRl8uyg4d/f7ioBRpy
3Zc9MyCw5qmFTuAg6kiqtoGC+lhP5TCI6W1BHnLlt431SVOK4XKpL33H13pShWgvHQ25nFgn3Vt1
peK5mFcrkcBX89JOSvfD+1cAw5kiO7ErxfgV+dYHM0z5b1eJssqFK4IfXKSxPisLGkZFTIkXRMEK
QnxGx8jRfYNDPp8+FrPVLkzX4VEWNv1Lz3vsDmz7Mwfr+x/61E1v4Fd/y4Xncmkqaf1eZmU/ExE6
9obBmpue0YVo+eNLbzH69MjLXdR5Dza84EMUrCqqu0ogfU8x3newgK9mDrOhhkzWpqW/2iK2PG2t
bT/iMXuaOYRyf/11+i2XD6qpRA0KdfGPxx+rWmb17wwqVnswoTtnEu4CAunoKdjeKzvcGu1rCD8E
X5pLn7qNoajL2nk7QY6apHKdNBZWNpTksxtpiq0tU4A+Gt4yULFhW4qYpTBVL+ZIXHIpzrXXlV6e
XOG+J4VHqXDHZYNLzHsiT9twEM1l3TmWDet5tedE/liz8DlSA7GQXJKcAQ77ZbmGvkMUhEq66GWw
AfByJPYqtKwN1+H/mjwUNLeWn0bLuyFunTJIs24j8iLa8+R8gQOce2ZmG9iu2TaHpSxQdcm2vtD6
0XOEseet+DUPowvyFdpSQiNdWYAWYBts4bdpYMM0UIxsvnw3idxXoxw1EIfZ4p8ZCiPZLPfLmjRL
L0GXToP2hzMx1ZHlVjqiuYU99yex3t8vr1Jet+QIQQCehFsBnAedNDVtOzYZSy6jzF7dAW/0XHvc
1s46fn1zIU3ADGXTpbFPmm55vEx0ytcJF7pibPAVEGCZGZ8lG9Y91cBCmb1x9JkthFrAKFEoEpYj
L9jmg3C4gVruucZrmFyX6ATJZcP4MIMJkePTg38YuX7BUsdfxF3TuPWjE304xUegttuQGtqisNYX
tUvPz314PernydCTN4Lk64kOorWdBm6SC1WvxWTr0/PS6O7P7wwhXTZxsu/6lPqANblYJTyuNcOx
0LOEOULKsEE1lR0N5CE4HUQBCQjQh2x//UW/5nTsBD6bVokNk+5spiOX1WorLnY/RM4oIfxZofY/
5DImV7/g1WR0AUJDPE/bmu/UVqNr4A7k3TIx3VOdUJn0FyfheDgy2qdmko4dSBzE62+jluj/ydXw
clG886Zk6Q52JyGoOHCkhAtR8AKeVN8cMfmCwvNdK22LSXFeuw8Jzqt+0BMfyNOOo6M3GFqshJRu
teCpNZR30DLTglTXZaWlVoxlCyYQkv/TmLm3S2Lol9kGNhaaYM6gj/shw3KFyM6y3vJvGH76Ikp1
2t1K8y0AS8NQLGeqeG3hbmcGRMzQN37xNKUgs5MTrWeI9f+JKaBKV5rB+5wvxN3WpUwdvJWOyRIB
Wsw9oWP2ca1ydA8/zEBmy7CG+nUadujGjdN8kiJzVitVkil5Isp2v/C7k5De6ogxCIX+Yi7vgkID
hmFcf5Z+iPwwcjueuHKOCDjqcIPq8R996owOd4iedthVnXup9G7VKnqjJ++TWrk9SR9QYL66Ef6O
/kuIPJkR0hthi+7V3pNv8TmvLRX3wnPY1ME54Tziytiu6ra+2z1dkiukNsXkHSYyFs7/LfuMw9dX
8R87yL5/YvH/aNNuVr6kCn5fQauZN7jUTHxCdPBT5ZYPRdRjxMU+9UnlHBEWgA2OYWK/JNQhzzae
bPLOQ77bQaTf2wOE+33nmz/mYbiGH+FA7S29GqBX3xhQv/AhBd9G41WWkXmGtnV8eoiWJmGEaKDc
7ZfLshRRye0Cph51ALOskxqdty5qvwG76u/oMIbgJJ8YS8HHZ6RwfMeAAXPRPapysHWENYV1iJoh
5ZDaVO0YR7b7RBz6aIrDgPtbwWn899fKIOIj3uG3Gqegj7HDyh8FybaspEvDm21JhB/KrUwM780o
M8WRu53mfvt/KYoqBPlsTg1h0J/60D8IpBzhjI88Y432DV/ON0jTp3WBa6rdaJAoX924S2zDTX1C
N/P77vhg9VHzedbHUbEQjaPVOga12cqKiH04AI8frUg+QKxluRusCSUXPWJjS4fr0ZpqhIcOp1Mk
pdMBzRZtFTYZ/ZdZn5YiByQI2blspS4debJISM7F+l0I8QaLkdw7WL3FzJmjnm/ItfHY3fEgCnwH
6HiMHRMY080B3L512Racqf14TfI0D/AN6guL0XjsEa7qTDNC3I3jkBAuxz4BHletqlZek8QQCZVd
x1HpgaImV6GwmNTLc1w4oMtYxQwf0AwcpT6AR6VrUMz7MAOg+ATpUjKQPELChWhqvhoYL1CeirTt
PVaGBYXdlxuVD5WY1i8uOeTS+e5cmbtQbey5JmBhE8w3fx/Zburb8HUqplYYy+42xOd+endLtXMS
l1n2jZ4JeKLkRZEGqwyq1ZYLcQIvvfddMzcfTZQVnwCpCQDLh1g0Zpqfys9wpOAbqM23iKzdoL3G
ZQ11K9f23C3BBCtbD0wy7/6FMp6MM4aLtiSL3p585vZxYCpB/nSkoLOHDuDaOvp46fXyQAqYxzAa
rL826yrUP36LyUW8JvG/gGVZZ5Rxp9tXmU1xS9BJWHBLn6BulosJq5Rz/0WNJPMcDfUSQJGgO5O0
Oe7HU9XiNqKRFg+2dEL5+bUaiAkYtFFV9j/Jum8swVq04SPSy8Bg2QjoSDgC/EoXXJQLP9KZjx/I
GZJLR7aGOxk7uJnNNrJn1B4vxKOJu51TOlM8gpTrFbkANm5WWUF7sqE20dRHSB6RWzReP32C1F+Y
4N3rNxCkJnvkvIqyw89t0Mosm27NzYjAnklL2svX/vVoffZEOquhOcLG+pVyb9z8Zh5yXvrifFdt
M29UiyS1R+zfy4KuJ5yQ8rY4q5A5XAcywGLs8+BVB3C83pIAwklvf5QNq94LGzpl+PFG8Rey995K
+kvZgNB0Q8Vi0aAktTxN8W+zFT6x3zlfGqT5DRDUHKgWf4eY/S7PK8YE6VrdMoj6pMUqB3zxzHxt
ilMir4khaZbTelH9ZvZWEsCtS/vkSJb9IkRNbVfhhrA21DniXgH/bszHPABFYz90McExxCHPP0Gb
9XQLgKTUeCZmRK1/lrepAr2is12lUJfgYEMJRHfXw8CPRYGNqfIOPpi/GBkgd/mSo12izRXggE15
IMrCMOYOl4oRPs9l589kFApPWvpVfMYkxDgdBKCSAcQNIb/3kq3hQUCqieaYX/xAuc13GlpQDsP4
Z6bsEH06zBJrp3gV4gkhWp+bYM1d0kFfoZCne/0xo542Wyf/tk7qw3hsa2SA63s5oGxKfJsTrIWC
X5QKhEGg9XhJTewMat2oRn4M/aROYRY/mQVDjtjkr9zBFjqiq47Ld0JQUtm7RrG7H3rRdP5+qz1x
furVgEtioO/Hi40fHxif8nDmEUWIg0iwNGJwcvVDT5ddljAx/ohvOeEdECUUSTUq497b49H8jtG8
zoEZ6RzIQ83EOL8C3UpfkSL+plSv2JZ/ek6ofMJ3EA46xfWjJ9jQ6u5Dt52GI+J5fryuiVvGcED3
dQOsIytI3nv4RJVWZjUrv7eMXxV+BRSfuw7B5xRgyEDs78a3KtrLq9dpcWh8fiQBpJ9Z4insg11d
oj+2kVIP1iB5XqX6dlyXWTuslAtpUUiCsjqM/ZILZZJmcd+6GEjI3DlmLnxiplFpwtpUNI8AviWH
aYuk7lNQY+Edams5rAi3j9f2yB4FI8Mw75w6hABr6b/wNBhfSDiEUqMSvhImTYXbuqfF1BSLOVu2
NItQCA/UPdpEQ9WL5XXdo63/e6HpREfDa3jvfSOYKDvufbub/sDiw3+k4cbWPoccKCKysOUrfkEo
+KMyYaSk9rfwKpzFG9mc/Lw5WcS5Tvuo+yMVrUnIMLixOSdvjvFTWra/tMQrQROdE8ieGB0bYbl2
cmyEz0LfiHSKV4gjndMD/+eoXN33x1yPY1v3htGhafUXsJ7VhKZPgjaRnlhNIyVBcXShk3Uy0lP3
t4op9JiWADkjMFl1YUqrPcSu5jDgtEuFmmvZWTVkq9peLo5WGrdSFUeyWtSg5Mhg4MQODIVWuhv+
n74F9xCSwt/FUjkSZBti7J/gCvXcX2jS5CLOkwqcrJOqPHt1eDBBljw8qGTknkdHYBaFRUnGbgZ6
aZzAzWF8gogXbY0WlaQvitQxnb+r2Hrffy0TkqIhHhnGfw7uyXljwn+acF7v6xLrD431lmPV9nLn
+/wqwO3K1nJHJj+q2WzP2mgP0lCowj+y/FxmBwTVRmjz+FeJZLuEraFtEJ2E6YaDFxGg+aGr8Zu8
YCqWUhNkk4rudQ5H5DFYcQkJOPNsczS77aywZuwdu3y8F74hfaCipCrmTv6gz0XGozX7ql6yqvtH
RJ4Bej+okuEO9O12ALjclmChTl5PEFrQTJZGvtZNFWVdbu4W1QJftefw1qyK+bbGFYo8wvcvRA+g
DFZOPBJ9cvaLRYrJGucdz8d4R9KcPMcqv6W3oWZBSZcFpqp5KEli02IUGqID/oUQwCo8yB8x6vjf
wAhee+brHdxGc+Mp2ZxhkvdhBtVz9ya8q5LCAOLBZFrpLkHbrIL1ENwabpecllvdUUZtY/Unj5O6
2RSftAVEg1xFtk7d5SiId6Q/O4pY4uHki+hIIxFZy4V7mNzs6N8OfU+wNWCQoPpr0L+y9/V6IqsS
FcNyvZuAhkY3L3JZjgHn5YUL6/w1VxxAsXzS9QW0nUwScioWi9PCCzTGXKpBeURCwdW+NWatrE69
RISPLWxLfgOFFRAv45eK+zqj12UVo1ZwR3j99mQV7Arur4CQM236GtI3QJUfcXQQNUXEK52JWcz/
1y1Pg0Ui8GJ0iZCjJrYw6zOYC6o8e5Rj0xX30Rqskck3/72rxn2b5pF7KZQMNuJwrdeAHdhbvw7U
ppvZg5Czgnq1x5V0HKPj5z9ylA6+W0gjy54F6Pb+d5dT3aG2CO+qkWfVpjk+/X1CgHo+LqrM58PV
7dJDnvFlM0qwAD3bj6z/kF50dgE8cf7NyPtiv4RBT6UAOOr/5aAhHDoN903TOTZ71l0/0ijt8XAr
PZkZf9P9QYjCH3NL14RS6UbQ+zEJavgi7k5Z0Je7fs0Hi0svrDuGbC8eCSseufHpiUS9rCZdKPLq
rAvcIcOtyjr5jHDf5TxSgw5zxOrc4oL3rin5YjVNfAXtxtaXk7LCzp8aMQuSLqKGt/hjcLKP3Vj0
QqlEc3avUhzrINkxYkcTUNQj7ngMdGKgBVnY1lAUeCIK2Je+LZvZ4sGMmKKU5Ic7iBk3+3aA5Y4e
Mg5TaZf92DsGk2wbCCW78AX1mmPjutL4O8YiXaxoqu9xaP8f4A5KY+Itgalf5estDjFamvKN4geh
95CpQFyNlmX6LwnP0ENFCy1f0WnPZ0z74aBwomYa5DaOz8ew+pCBuqY4EbWUXEq/zcqfrAmRBWfB
BV1S6g2Q03HI4AP5XjT8YuzmqtnPEfgDhmWjzAXlnb4LTBOEDQTa5p8I0dbpHHzOrOoVNlGy66dh
IlNKwT2IaLZERpu47fHuaUrYqgGRQ9SWDXwVZgpRzbybtj3vkhkiC56mBv6fIgvu7/bbxE4+eFf7
5dTIeJARbwQ0reacXFlg+bAuOJ3amXZvaEoqF30GRh/qfMgoAmfvXW0Rhuounm+7+gzEafoczYbO
E2f3I+ssh2sFRTxhaJZJOG9/jqxacOSDqE7dtJ2+UGNkwGQA1EP5ulHTPmYle2Wc3GJ7PNWrni7+
oD8dsi1lIn3GUJLt3DVSFlvUoovL8zIsnheqEPJfxD8Y/NV6111/I1ZN6U2vCZwZ46b4vsu7KJUZ
wumAWPbw310qWRM2XebO3M86iIGcx8zlZtFH/VtIbbIlFJSUjangW4baSaNZCfS4MNdD4snzyCAP
AuZr2v5FNuU9mMVYdm5IDLzV9hb+sbVlDq2b5aTYM6TmhRxrwL5mS4YZN1FWUmlELsMayQrKIdLe
bnC+YdeKrdrZifeapVMFybA87FLrPWZg/+9v1P1B4biYSRCvv4TsCQsZ1i280J73clGLZ5WmnqEi
UR2chcXdS8Bq9CvjwvMGh5LC38u0ge71/IGoGXEuUT6B2Mi/0yx3ush3IrDdBzC7RV284LkpiTEZ
z6deNerp2AwmFmhVegV2gZzVyyz0/v1wHMWrCe3R7vP3T0VL/5VSt9TNaRs8AK/axYEb3RsrmAvl
RJsQdx5zP9g+DPTKMhX1dD69Z+Tv+AAlojpYhIuN0jax0rjDOtdM45q0o3R2YKqKZY15SiQdSZlk
WYgfMfmBE3GvTfsHQUYXdl0aA8vptPsmtY8jFBuL/0z/vweRuJJEEW4acvEpL40i7wS+g49owr5H
eM+s7ZuB69ImoLx70vVzBL2MbDWp/H063Ozb2WOdI6nMOawR14/9odA7xE9IY1v1zPSlvJpa439m
iZpi14fNa2QNl4oEVv5XG5IEfSo1fjo6IzLGes//wR8oxAIwCP+/hQi0nn67N/RDL3LfG2vK+IVz
DcHDhQ7JGDghtbP3nolaWcxfdqQokHl4pbVY3AOzzpaSiPp/kq5F6WfN7cX8yrmyioyXq64SO45+
FYVbaScyzaQXoUqsYzT9udYrhuJTmnU/HEg6/BgmL7fwjFXMFuMgkV6IJAF3cN1Fu5PTKveMT0c2
RBQSfhdaazodEcGzp+eojJLScyFzhJR9xCwpbFrFT0WjKFV2DrZ79U0BL1z7FcHxBMZ6K2/3sYmm
CUP3PrUIly3C8ObJ0LTc5/15WsmBZ0b2bV9hjTvFc9tWoHQoeKj8PolOTa2XE2b9j1GZjAmcvQc/
FzjOj2wq8ZCeb+8tMO3eCAJYih4gV9Q+32BIHcISBRXeMOyZ6K+a7nomR7/feVMYaarGDjieE3CK
KkG3DPTjGaQf5sxnZMrdQCjdg5ZK7Gm+4HZneLEFAY+JC+S6uGiTZG8wp3kVaUY5EbhCHCsRofYS
GVrUFF1EOo67iiajlBSZEJyDgm+l0j95CngYEb8VQv6HEXxT68L3nnqp4JnKN0hHQAxgVAWc4MHU
Ecb9VCCKx3xRMN+28EOh1PbEJP60CB9Gz0oFJWD5ZwWhx4GO1QchdWXZdpgkZN2Mm/9OeXDf8mYc
2CR1o7ZctZqKhpVp3tny8r72EFS+SIIbxB/PeNoTV2q1JoJPWXnYcJNXmOCJl/XT64AGGcSCL5yY
AAwhP0pT+7LhvuPaAahsAE86zJs5cJGK8XTryFPbeebyk0jtkA3K4s53ioUqdeZ98wZDY4YYfRiZ
wSU1ZipUz4dI5N9TLpHOGbJpAXuNiUclDB3KG7rNOAr3M12gx0Fxur7UJ27ZTmIX+frzRQvTmXAl
NtUyNQI5TwhneTFSlI34WyJRAxdcMPb9OWs2DjdKDUo/iKPKoKm7J5SxeUpYrSrlNwYKSJ6NPXAc
co1yVMOw1ZVHmSXK8vD8kA2QpCzZ2NCZFsJIy/xn0Nlh3XlnOLPOs3qDVivqR0DYIHBb/iFGov60
P4Sq7/Ee1D9f4s4luIT96VO3be4zLiEnkBF1BSAepsslVFEXoVmwZ/bp9SSXu+seCdQLjUb1yChI
etHLvyr9mrzHh6kr24qJjcc8gtUWRaa3+umAtQEg17o+vZzpgrV97x0WZTL7blBhPWnzQrQ7mlJf
WXywMBQG6XegJPJ/Ng7T7Q4f2iooHQrXAa3j75OWt4a1tV997DmyCqN3vOmlC3ZJkxLWkE1CzB/i
0UT2sU44eupklmuD4HJEAmvI+OcS+TczxOAkhLf7y8g8EwlhrVyTLZDUPiDhHUaImtt1Ckain5I+
9iwwcwJWwOZ71QxDBpRmc2nV+Y/Sw9RUmsZIP5asPgg50dG0k59RSBrnf+L4bgoZJwDOpAEQzuWI
zGuPFUvmY6PqdX/+jbRoTzWyZ8sz4KBp9hEgMVPGIoDfRTGit5SWTbiJ3VDBi29u7M6aZ/CXN1pm
buNpv+Wdz6XsdoPXHlN/kZ67oXZClva4lFlP9Be8240x6AVoMbCVTzmwzpQ7kdaOV7HNpCK+OUpC
uEiQfngoJARpcAwNIE33OBTCHLx99Ymb+6mZJyKf0ea1ylSYpXV0pk3JyZ1u6YHRRSKZGnYZf9xV
NSbPM2gZgABwSKeV7CmxO3koKdOCovkamjGCtXBiGZBtIkY8rWtoQZluyqaR0Iz9su7XNi0meRdT
1ScR59do9LtShRB27cW1lWYVesv4YvURqgyFyFzEO884wytnEkDTF7D+f24nGZb1Z+ZZvNGUI4gG
GUvz7chJztBVJJRTwBFrQMNHCp4oHp2M3XPElW7Huj0ZBkgx/DKZ3GsDpGWW0XdjVJosaMRijYJe
NhsojgSxIgbpVk1+u7dDvGBE7g+5WMt3MvC9VjIeb0DRX3y0UjS26E5fHbPeSKghk+tbGvqmIuWX
qdh2OoebVPSsb/ks5iAKSDfyNvDqjedQohqx/mmR6bP/hhelMdnveGMkB9PeE+EdtlPC+bidqHZh
1s1TyjTRXMnHGGL1q4j30DqkkPLXaOs3AHG5FbfhF7GfGcA+swqBXki0X4uPEnkm3PcoXN0xzJj6
tJnz70HMB5KzSfQIEGeI5WYvoUbHlrq2b4qyy4d/f59TxFNTfozIDUa4A6sYhco+Uma2Ng5fYRug
8E/ae4bbsoYQmFeFvySmblDaC+jr92dOKQlG1qCm+cz24jjnigGq/x/HtgzAikuH126A+BjT+LkM
Gc9ip3WVbcdWZZ1Yq0xqFBAos+CnhEjNzAmkKFhwE1B9T2xK4wYtGbG3WXtFSWyZr7G5OraqEF2G
y6ugpvwkxvk8pRUxtCTYQiAIL9xB613vEChTj3vbGiVV07XHdXKMTQgt5/XNf+9KW+xUfeKpKjMY
DwQ2UIGRuCXWKL0/bUsOfao0RozSJ/Jjm+DBBIqM44PSmlohuAvy/V/rvV7+r77dWyaJgVGO4zCx
p3hQtMHaMomtPo0AnE8MmxO4FTOlZKjYaszS2lnKlCwpksQ/yjTCacU44LEBPWP3cPRwREUceebP
euoiJjRl6KQPk3jI2jGczt/+9ByctWUx4k03D6+/wfjLCOL0RyfPQUoGeQXlcLe8U3t+PfXSkEqA
wTJnnk6JiULbXfQiYF3iH5aY5K2YeQBD27D6BPNKQ7JQIgtD8A+JIK30x9eSf4vPosJWYDSGGYZE
LH3MUohRN+WxB7e0YibYVjFowuskAM+CAjdISsh2clziTVSF1XuvZeUvaD+nBJNrYFvJlVk2QyM4
6ivGCWcQ02ARe0D9WdEMOfhg3iSk+X2nN0/XmJkrYDWmG6kWEK7AZon4uhUEyQRksT5St3YsIrhT
c7epGPxFG4lXktpjChrFpMUfO+hMScxiKa1dv8LdGn4I8KFd7cNH4lhIhxVAiFI71gToVjaOZP3l
kzZugpby+SIduHubqYTd6uNtNDXdO9FSMSC/bKE0uIHaVpKGd6a0WeCipcxorfvKji2FrAjx3wtf
VKnWceuvDpMkGIU7DBFv7fOHl4ImQddeVIKcQitfiBzO5dUZsJvc8FVIL6eEDvnDUn5XOvr95na9
bRIN8ywqRJdInKFRsYY1blDA5rwNRkRUx6ozLjU44oc7TmEIyloPlrLFgK8Z+fDkB6k4oB9Tjy06
YEic83Z02dANpPmMCQU2mI0Rc4O1bEf9TVBD9jCujE/D5KBvzGZUaCXaowp430WZMYLYyYhG7/od
7GswpDRINg2fRVh7je6RtFv3fTXCEc4j8xrqGzVFewu5HxHoNCuVL1MNFkUBpXb3Kqsf7fgszuTC
COsX+EuE/mV7OOf78iNbrUA/rMpfgTVHWL/AQ5nWpxTUhuhAjQTx0wh2tDm7V30/FPzOE8AEbgBd
kErxdH39lHwfhEJeabRf8GNd8JR3JbLfB2ib2AW4mGM8dJevC/6ut5++DgJvDY+g17E/ceHlA8dx
4SWrmiUP16lPFP1sX0EMMUdvCNxu8cZ23FT8YDLuV4FIDwhUjRKMSlvXy+S1UfXN1/CmNcY9MoAt
wTQDqWqAU5y6beabDvPhk0hfHf/FMEIt2sbfhzhdC1I+0CLSzD0nzXiW6zL5+FevV888kC+d98S/
grLFhLr5UP2LvKLRcQKJASigQsIwQ6gHYtbR3HADgW7P/MpZVDiNw6fDzC1NtVNs9I5Tuixe3RdL
FjN580MTJQVf5HiA5uoCrBPlqWEgX2v5vQdRj6MklzijoEFziC+e7k+/n/E1bpQRDPDHkug/tfXj
8U2bHG9bOxs+KIqAnluMXk3+eJJYkSfl0dQuGP0fETkYsivjIo4o4rwv9C9f4TP7H/RcM9jFFxWm
KRhJbKTmLtj6h0jv6rGzmeRP1A0Lh8lq7RdzHgWCuKUkjkIVCJYmWOeGzbJ/MdeLZ0GKx7FIohXY
rvzBF8qkLVNY2gjCHuwAsidosRsVuyRpFT/Me4bp40ohuwYaf7aIBl3Md6sfEj5FZuZMJwLKNEVL
3hKyBQzMomF4THkMK6EKVk4RE71sUqkrmU11JfvPNj0vjjKym3o7qDCCmZWyy9nrlsBXVf2OU8CX
UsEs3z8mAk6h9oCyyr0zl4KTtq8qYvx1oPXA6LODHlJFAVGagmXbuJSGnm9tolIjnSdULxwiEKBb
ie8WrUh6bM49yVCGvh8ElMT8BDUQRsMS+y4y0gDCfQqz5ImD7QltxZrGGJEP7fu5vVmojFsU3Odf
bHaptyoIoZFt40zuFQlsgPkjv70x3knPhUvE5nKGk3zYVYrAxtStmXP2cA7drCmF5hKQSgMazOS7
EZPH7vYOIxh/iEw92nWUjEwCfvzIyVDXQGxEX9hZVYD5HxrfvKJNh2YiBPbD63SNUvrynKB1fPhN
5FfUq6YECeQTWGrHwacoyfZQG+TTa2mbr8liJKy4NOu+wytScjWjd2DgJ5lD3mIkn/63PlAbM15F
OTVtfWBVe5nk1IU5YeJDJPxxrBgn2zrWED4XgRaniUlP1eGq21HCKKGoveEONT7bGM/55piqsq+K
I6guHO+aN/L2UMaP7GUgEhnvljzLJHIdUynB/tVNO1rnU8TwPIoxLBo7/xBfc6VCJwNrQ4sK06yr
PNfTcPZL5g2NYSrQHvKYp2SdWxiDrgMd0vkn6M/vfBPZiYFD+MqPSDoPRokIx8Ei2JJmsJ0ySukh
qDwfIFL1EFKbrWXCS/5NXgfk0Sk+3vtIbfus9sVFR7Ma4JVFyEYwJyOuupWIcMHuk7kAdzcI2hnS
S/rEK+GIUTsxLPriFHlJbFsfpOGcoiLXKdeA+OuQNphfvEw993AbHWcxEyKlsGlLdytC1+Vr3zSg
MANK/y77jD9aerSCOE58lXnnuQmHcKE53bE76IvyerzQyyPV6NcK2zS0uc7VGObo8se5v99iyp4l
ZtKGw4AYNuEQGTsV443PeVc33avZhpvBQuUI9hz6b6/FwIiMAPBn+LM1m133HB1VAJWBgwBepOZr
VDOTXN2pCtS66/szb6Fc7pVAbHsUzgwVdLzD4+3qre6oyBIEjVykBVgev/KJbtGXBkg4pEZD70OG
fuQe/NoBH6UOykW/UmRCjnEMwHBAlgDtmwbP9uOC7cntFl5Jx5W8EmMQm7pcGB9ODR28ddCEPApu
g8OccmVLgBvxmoqVIt0KFsYcSN4pbvaiBBq+N7cvYsWiZXjewuAFjgzjgR8N9TsPDUjy46BYwOGV
gxVSnrPrZUTqHdvW7lt/tCHtqnNL8vcCn1L/AZqUuAEZ8GwgwgssRiWo/t0/RBEn8BOlBAX9fLAJ
aKVQn/awiydmg7DrC97UP2qIMxAmGirlBa/FBu6B1zsGtBEcJNhzfzd5fWgEMPWuIkzd/USHfSSP
ePfBkP63bl0TabZya5GuCFVrbL1BKh/cTvxGQ4G+b3GJbsRHA0tBgEWHs8xWZhsUMuTK/37p3swX
dMy4Z5WFAVQaTY8NrYQzfRJkDb/4o1ZpV1DnSQ87+dJVAnoUSXHSzk3JQLtbyCsrdaGiCNV7pZ8y
I5aKrlLsZNWTiPZHrl4I5iB72AW/3ullSq4x5fxOtCcrXOlFzCfkIB7RN75KOfTXbuKCo1Ux6iIt
/fpR0glaCvdSF8vfX/V4qAbUEx+l6F3/sy5eS5rXufZvdR9a8MBu/JKUgDeQCB+wmDg8DzrRMocb
9WND82Xl45wpatT4FaxP+k+SjGPgTLg/GItKC3dGSNnrSIDw3m2t2GuLIf1ttMqtSF0tjKq7dP1n
MhvjXu2YeZYQqfVnRqQBvkNK7ZIn46Oijz5+jeykEFKWcwBeWT9gtnW9P6BfmbbXZQwg6zKM0tTa
RDX789b1L2Gg2LeqO7a29ye1ghKKHoOY1OYAWGq3zYWLByHnZ8Vz1zFpDPJp7DzQpnNuBLByapry
TWT2Wg4A/pvtgw93OMtvJ64fu/v8XHU0HrgrWrsUNo6rnM3MGmHYGlpSyd7T9HepECuYxwB/yaYw
1ULNQml0HJ7ZUg99+R/dVEQ66VMYywTgc80UgqI6Z6utB2uRn52PBGzJTUfd7VI/c7kCF/vZ+uea
R3GLx3TygJ/2BmGjl+bAbowuwN1w7/kc/v+7Xddk7ThP3ILgH5/YbfOuMlPGHk9Gwl/ZvE05Vfoq
I5EEI3vV8OBi235Fej6wR0Cq5LlqAMVJo7UWt9oq8rT5vdI3bw0kp4aH2U3smGZhFmR9ZZLNVTCs
tIITaHINXHfVnaTwgXhO5ZaY3RsQQo8223Yg4v5jPMb5jk8qWY5uXxX1I4RQQZ7ZL+XS9FAHFsQ3
hdVIRsXDCzQapZiam2akm6ZW8rI9T+iM9cia/bKRdY5D9oHYCXD/3fI0X5bG7yOmIvNBI8XlmCkI
pMQwNCHv1aFNeBV/CVhIzsQHH9p1i7+UBZg/wET3yxpGPVj+HO3/gRLCJ2KnhM17bYb8HhTe88WY
BG8zgZOhkxGC8AefSd2yjY0uvJhDw/HgKjFUHXPlci/m8ScB5Xs+J0HdyJAV16sFJxXKD4g5Jozv
vmI5B78e82VicNLS2RomXc7bcqgGjyUiUojeXh/Ex1hEhAOBoERsHzEOMJQwMw+S7hs6iEdstrDg
6HN27wzfHSVXqaJc7bDbUy0sv6Ys5WOWoyQBdQtyiQwKZhPkyrFnPmxuRJ6MxtL1NFvGFjwPEUUr
MZRQsKO7vqjS38k38+mjYhHcXzsxtUL30cVVwCb9byD3zb4PZ44lhLnpamDm1eJz88cOJ6QVAOnU
H2bPUUS/BScONd7GNXzvvMEpKfkk097syYCOb6xtff64uU6PJ4+hv4hgHoqAEcaMRpxmR2r8JX3H
xjM+wiMo8w7NYor3F1VDFXCZfVBEvuddpd7Fbc7E/Yv7zgzZGqax96B4y6D35HW6eKCrHJVy9zGk
vkBmQVhqE5KxMaFsbfQ0mhFPkZIUAVZnS5FINboJxKFC8ePbNyAjm1QreP11UDxEutjvbG7Mf5pR
m4xt9Z+8HcTYpVFFZckiLYuDU53OkA0Ze1apPsLsqsxmYT0ROWS74uMEVnGXAOXgUkp/kOYuwYbv
lr4zCkLFAxKz5eqqhLlY5HYWMifq7C5jLI8kJ0koF0AE3v3ORWGx3mObIa/rC65tKByAhU1r8PjJ
8v6KCJhM8P4WjTywhggvY4nyL/LjMYXbv045Puh/Zd0mzMTqNHqT0pNvxiWMYaastX3JTZoU8oyg
cM5mgX/i3umTW3gkGlDcpFDva59xXvfv8YEctR+ch0eQLSWuuek1O/kX+DHB0Xl5SVahw6LGUUdb
F4h9z75sa3j8kKs9bv96/YsLtz3whMI76cKS+FWwefmmal8VjlYDCKjV2ap14Pn22NLf2M9CgRZv
hDQgZU6uK81EYfti8yyxsEQfWhQ/ILyL2KWRS1oq+Jo2LngyuT8xkJNBedDoIt5AlOZQTKDTZOL+
N1/AbXeXWk5nrRsCADLye3uGooQucwycLgrYSJbpQHFjrtjD7/aOU+Ey6USn/dPw+ifDtiddycDL
nztnZ9HlfnrTaLDAchW7LN/MIM0a2YIDFmWZ37OgAI+PtKxWbS5TQ2g6Iv11fQe68Ti8DtvHlan+
GsXM8lxDrq/ZfV1HMnlHeX5RTTLxwySAXmycDHdYxARwdhmwJuICQ5sDq43IHAva/iEX3aaekeJn
e3htSTP4Ms49PtBCklxSrPtBFfK8JLR8+Vv/ONkXyGXsCj0XEjEcysq1tKrHU27Yx8ljh+UBB56G
rpG+9AI/ghL+tUOAJz/odLVC8E3bv1D2lHh4XlzzsmPcltbZak1srqKxJfI/AvLnekCOvkPF+ijk
9EPwuJ86/m0PZT5qBk9DUJQIgFMWzo88P0Dfi2/TXowrxWnZeH0LzzOqEranm1qWFQLXPAaGz57j
uiV7KBssgxbL133K4FnQ8ghqxkvVPm6ERM69xph5aegARHKET55gwq559eQk5N/ysWIhTxZr/FwI
d+p1NIkuWEM5N30LXtyRjuvjX9PFoIXx+KGH4ZnkvaCSdn7yR4wAFlVu0E8wug5TiuVTt+pil8yS
VBx0LG+3ECmOi910OHo9JBXJbqxTiW6xWoWAYTaPBsB7CQZaS7ArWpxYoIcb5OsqlshM1nd24YWz
7k0GI3raVLYtmLHUXhPjPohiDd1kZRJVLM00RCdhtDFbSTOqt3+eR8ExynRibM6UIzLGFbjmhjzD
uGmWQkMdTws+aTDkqEAnd2Te/Kf2y8xGDw5FOAYqNIhWQyLzKrYS7/sD2eTiYYtWnvj+IpctkCKz
mM0e5xGstajPXLzox8Sw+TNxpwbwbopnmmHD3SMg6Ql56Hyy95s32KOAUZKQVTLtHE6uioaP6Ub8
2NT+0ZZZWOTlGy0heQ6B+KnArCvPhS8cQhFTRzjE8M0ln9RXzvcomgPDMBph5gYPoCWxqmFiYeCj
PXiGSOeLOE5ZHCOJrvSQcSEaJ1u/Zj741diFrOS0PMfj5xtcj+monKNQVX4LSup34k4p1XH0Ytvo
bSKmsVVsGadYYRaLoFZwsf3YaMofthO1Q94AQaFvWIkI6AYe7T+QsyBzXQSKnEaXFmatRdPnWg5b
jLdzqYZtYS7JQ1wSiop6XXVkeE9ZoLUXWwNIJnKj1u2r1YMCkvcHOMT82FoCEU7wDx8/GD83LrIv
rKNYkAftynK/WhhUdc5wYOSpAEb8nzJGdNZ/uaiNFpc4qv0wVT2JiJ3Tq72oj1eOufn8d/EX5iH6
+a4Ol7kOL/FgaTgXj3rwrzINp4CYfKMyINITbhb3Qp+ZEhXemFkiaQcLp5BOtaQtlfkuNkcrSr7U
uWAmr5bB6ZMEw4Qr2tmWgZcHpaR35LFe8lvT9eAozbyKWlyr/MKVnEN/bty5fBi6wTqBsmpMvjsr
YprEwi7UmowBa3VToKCyJetbAGDodTrXHsPjcLv47Rj1AIbiu8BMLYkPu73WsB3g0pQmpv0Ubplr
dn9T0m+Eh8TjSj4wOvCGRoDUg5Wta6bk0Mc3Gvi5jqBhRYl6GHaEqdc37+YA3s/NRt6Bs2PfFXer
V+HRy0f0+B9gbUh39kWDtSAsNT0IPqM+VhpW4CPrqyygUaRb6ak3NDjJmI9ZtB6IEmdu0mS6XvM1
w2x6eOyREjyskCXm9xQcmgmPjU6eGWo8Xbr2GIANQG0G8FqWzmH/9SkofYCRVN6IkGDV3QWnO8tP
Yf6mQOzNNgFo6RRIh6TUELLjxLefuDSwxVi2ILbRnzFMYn0wa7Z5YCYM1jxw/CwoxPZwQgCkX515
1x0/95LFdKBaqNENzTeLuV1RL8bCXBgmoYZBfQX2ojMcnHog1KCn7XRH3WSEP1bSU/+HyTZKozRT
wNx/h+rDuDsmXInvsvDkCNDADtlT0xoGCxj17kbJQ0si+I4N96IHh7R0jWgK1aofnjQkYOnw0EpD
bkw2K6tU/3hrCL+cdDMOfLJ1n9kRaKwFhhF5bH8oPJg0ySkpmFNqDw65LyXqotiqZbkAu9IHbvfj
FYR3nq/F2mO6htz4ckU4uSChYVt05RJK8158JpRg4Kux8xlicDK93jRYDv/gEkT+KhhySE9DnQaJ
j7plJsLgRgTSVcuAZGyezG0W4RNjobVG5g/x+d5MhsINfH1N089iea2z1af0r+be6RxvE/bboWFE
vbxtO/4Ad3wPGzNoaJbRmDNs0f48f3eRL1wBGxiwlRDfAnG1yW/AlsPcjk9UywrGyhmbJj9Xw9+g
rOHNzlKVhvjP4ugva1pdiqj/NW/1H6C6tVzvhwwCS+iz8NhlKIK/QJD/8pTPhdXp28M4fHZdfpds
dLIfR2y3tbi+aICZmnWGVFNta18CkVaH6w4KN96F9+flAHJlSi46JB3cKpupyb6E7deZmME00Ef4
q8cA5h9FI8dGMkWn1ZhW96bHmmDykWa5HuGMhJf2pjvSZnz42E9+wioSq4O4bDrif+TT6gyeAyPo
iY78Gcw1lh93cNqWO5EdtSeYac58Oy1URIqeczk94gYUG5vt4RAhonfzeopE9rXaL5Wcuq8GEa42
+pi3BzvgYYuePm0M1uH+2ue7sekjP3suFoOm7WKQpnACPOlfGDsz62g9mQzqoOrRmmB8yuSGnB+/
WfwmNTxGIyPCCIbJ1bazf7NywSbgeEelQ3Ne+Lwu1pZeP5pI3fmxb3YIAWOk7ftQFQCKhPbfLi4y
BnVw5i2NSaX9Cks+aC+znYwWmLKOcYEGYBzOswiniItQJ8wZxqM6hi+7VWJz4vyz9tBw0Ae1WQZV
EHjR5u2tqnLqNpJZJjrr9ioJ5wIOUl5jMqB4W8bvispIhoHgHgwqaxKM6XpORXTko0iJJQX+tog1
3S5j9DVnUYUhlKAM+zRQ0yJLZXbPrOtja6h/oC4Olb0tPpQU6fy2VF+Pbk+Pl/hpFS1akQny2c68
eAr0lVLqJC0WYXb8WD37yDdVHJv1rYiSZ5TI2X3rEd5pqbISsMnDEvEhgGUEIoAVKnah/OdTH1j+
87zJvgbWag38We647loiIbDCcSbBZJjoQwwmeHX2QnmIMd7iDPzbsOg6w6flsS2uL5TlT47oemDD
GSSkaqiNedxKgNp68CezR2vXzIJJwIxzPY+nBxe+NRRo2e5aeT9iivFDX/oenpdQ5RmzuiRagwgy
5iANL918JcS/tdHkjGXRXs23JC24BXT8s0e/bSAwuBcPNuI0s/0zT9lo25dNo6kSesVQ3cNgNClp
puLhuRalbaZ333OMKhz+1I7KY+FS2Het1JacwPNyjF0e41Hs+G2TqpVKHbTs+mKA8TeLJioLR9C/
k064hQ5a3tA2G0STqFN1nUGAZGctxIJSQEdwoauoP32e1ZoyaPb/oxDg4ZOIr5Qcaayr7GRthiX8
916RmeNM/7HD7wWDj5JHdhyjiDnAWUv8N15VXL43Wna44YtRSM9FD3Iwfny8edKcxkR0wODHLLpd
ix/McWTbylFqVwwCsz4w18nmkkSPOq4Gw7Cx7iQXaOn+JxkHfDmupSAIxDhsPKb5BNToHPnFIHfG
Gjeib+P3J2TSqF7O/gnjTqZvBL5cSvQJprNeW/gjLx1BvRyES7Y7ZtcK2rN6mGoaY9vr6o/zyr6N
WvSexCZxhcot5rL0W1Di/pTkNpt0G5nOwwDVu2mlhaFXlgJnHsO06mHzLlrleu539EZFO7R22QXR
LasFpZM0qAE2K04OKHiTyUtTD24A0tXeB6w8rIyvujTcS8rLU9fed3hTM02y0WIN53oYd1i8xmq+
ndJrc5rkiY0c6otmLRiCN5wBT8FWH8k73kyIRhuZ1waqB/onOYO++I6bU/Ysm0mJXZP6d4kD7z2q
ffSPcBJZ0vsNt7DBgYvNmLp641MXKrxdeYTdTa4mmRxBw3V/vf19A7+LYTz/+x/8bKMkW+rEoKNW
cmc/120qti7SDAo3JVr0+l25SqXEO0m1HHhfZ5rwedn3J3h3GuNPOk3LjBRpesBz/JjFroaiv0qY
JcSPhaCnttpPeujIW8Jxx/hQGLu9oKApdy02LTj1QaROHVcCRmcFo866MnqlvSsi/rkqnusaHe0T
ww2awOEsfmLWofQD94iOs0iUApkqWoOX3t9xarCPt9kS5OZGNxiQ3hRZYU6t6Syd2jDMUMrN900S
AuZ6qA2NtEFrRFMZtXdipbAeJikNbWvYfGQcWA8WvIzPeJKUvj8vNrO+OT+uYJsc3lI2sNvdumpz
vkrcDCZhHzvK2Egu4eadd5T1S0fvDsYSJBXKR62Vq6cYCavr7F7N9HZC3/hMA9r7gT6CN4eW3tsc
YrkG+jp6MCwhx/NAiVbpN5bUa5LR5EBtGAH7JrjOq00M6ROBHhkJD/21ZxLnEcpDeRjmh1csSyGq
qAA/iAcTDHumxIaBaJhr8nqygiojC/Yx8nMaAwek7Tm7ui8hh1CGCbx0v35Ky237mWs5TxNEQfAr
iZY/pDwVZ2PfuNqaRgnjLLO6cPo3CzDC5erbkJvkCTL54Uf1y4bEeGgyf1x/FkcSajmszPh09kcm
5n7vAR6Fj71zknDVmXqSL5tNr0X+mBHQzjLIP0ezP0nV0nvSzjL3pQnbVOJPQ8o0dC7IvDF+221Y
Q9cTcmEHOCGbykntAVQ6l6zmWLKF/ziC07XoMQU3IN8w/OP7jNCciKUggRcx4v3jnMw1JWH1woyK
XUmLCjTSUME6sCmwUxvj/Ij/e34Fd/9D3N3tgKILH2cuKw50q5Eu3b54U0FdCsBHJnjVv4jmtGoY
wOFMVcWE6cb/J0MQ7aAfK5WaKMrIvx1Vv+jUa4XrUFlLAvgkF6qayEzRBTWRAQjRDYQ5DLmNQ+HT
frESacbDDuU7FXTsyqwKeFr5K+zKt9xFsy5EijBxjL+41g/M+rs6C5zSebES1YV58m7+Mbbd+3XG
S7JAErqms/vtY6ckfX4NV5RW9y96s5E+OYtfbyvr81vcNJ1tzoYjCKmlnogwWMDqpMbUpUi5RJlb
twxdwY1gJ1LD1jfIRYwX7bcaeh2Cc4WmNKN7mu0mbB71YGyU4D68htNWr404bLb67zTrbc2svt/2
NBSsWcVwu7WPZPcLgPlDfkgGM62jgabCGFc4XNkOiveYH1vSaj3g9MzbnY9PoWoSrL9dqaQffuU7
BYgju81zr9aoCm+K4fExRa4+qYFvAOLSNOvQU3/n9TO6dEKAfKaxvWLAkD50jPTv5BT92vqZyAJE
HgTxOcnY13iKTFT8tXj0a1b7SjW3owrOEOZ0SHuzs5AQbeEjzZ3nAMwIocZTFcjOv8TM9a59XI8t
nhkZaPWmpduUtk12BTKYr+MPDA9Umd1aYsB2aVz1QFN46zPGlnJgiQtc3PpM9i2VMEdG5vH9OtOi
z0CWVbqXxMgy2O9NNqn7KEI6qn8Q9xPIxsFa9CYqa847zVN889w6iBNqFsRVa+KJsIVJhUqs71Ip
IFoB9QSmuC7yHy5/oixsEDhd9N7K2LrYvEgrT1G6N9k4LXeG1F0KyGBQJq/QgnrKvaLv1PBD2dxq
3vNOhICqmBaY/mevsdUx1zgiF5vitP2JQp6CrFITByVJmi2Y20dQkgbASZWSeKKpVXtryQ7xl0Qz
EyQ7YaGgn/gR5RxRK9Wf5Ea7QhzikXyl7K6q5Sspf7P6gYowVkxfEswxj7ptH9S5soma3kcGEByf
qq8pjruFHiLcwqLABNc9PR7VqOrYg0n9rmwTxwWQiXU7427dzkjo4i4xca2TuC6s5D/sh+oARGbR
KCjiUQ0+//qt1IJesv/AYQJMspF0NS+kmd4B7dZJVlU0zXA4YZ4rOeaah/IRasvU3NEct0OjvYGg
OOpi+HjulCbZfCYqCuJW2iVoBfanmIJOdyAyORyh6i+Sau+K4+yJgOZVQQi7HRcpmtQVqlsr8i2W
TXKDFcc589y6+4OIiV0EgB3UP3m30W67ptsLSu00LDUPJsARgBtNok9UTBXek0uXnM8u/5OTmeJe
NdWkj9I8LQbYCjm+P6UIbybYyAvJbuWyTLYlYfi0K/7KjT5XWhcwPmukq4LUYiuiLTzoQwFW2cCE
4FzMYq90OoZno/Aqg41i/OYdIuObAxTxWKiDQWg7cPPiUqcrGKK2f69v+vdWhGb+pBp1yJPXw6SJ
BrHRIzxyP5WnwVmDT93WMzeqWQST9rDd9Niharmq7u5WCfLjDbQDj6ZWS5nfVlZDecM2wtDVPc/L
QjTEzdju02ab34dLnZrkegiXbBnnR6Xy4UQxEzeKPOh5iL2pC+2nYKwkU3UTI97EuFHNqz+MV57x
Vuwo1CwbwHJGSkVlYXrBoaTh4z8C4IMfc5LzN5gG8OK9Aa9StxFJWdOurUsdHt3qq/WgCFrQ31J8
SyDxYdX32aCBBlvSzREwczJiNA8NRM81arAUZjCpisfbVEWBwbr5ZC/G+lWEeImSIzYA4Zr6Wypu
VDkRsY+qP5v5vSD5VOCIzc3MPQ4MbEN+ZnxAREyoEOGReUw/JKgqS4MVutrzhvJiqyVYouslDmFI
W3y0B2D2qhR9zm/KhEe8LyIkmJRdXLLNEXLOyZHUFpu3TePXx7jG8ZiDTxAJQWVZDN45g1x++c43
QDORmYhpSUI5aHeKUtid8wfZeGvD8r2mC8OxsjKVGoHkWDLZVYxfyWSoe6Wv5ny+nXtAPf+k+KqI
+wnVpe4Og/XVjUA52XMF9CSe6ntAVoTefvssxKUFtBNtjs0XnuzWBUOz7f3psZa7Yo+xZPpkglER
M1NnQG7smPVYe4yRY+NFUJ4hky1Rn4nr6wclBqKhx7AdQbq1Kc+LzB6MhxVEB5ApGBrLZnl33M1K
NjxXmeYNBD8nl/5JJecXe1XeF3CixkJnbB9nAVdigXr9u4H/c53xfLEfm7d720PGgpGxqGuoW9LN
qU9h6QNiNDYrZaTRtH4FMU1GSpJyy/t8rUfflZxDatpwnA0ugWk1y6nK3gNNdEuvX1FjcHxxxnFG
IBezyIKZLu8XckbcMUe7msDbhVioFGwZrhq+pmtogFjvgQA1A3vrLYTtxvShFDH0Hvz/VpJTKpiO
qU1z4rDmG6fBBrhirSiKC3GpAMIeBImiErvY7RHdtsk0FKCg56Z3tz61agVlWOJkSYCWBjL0K94R
kIDkV+m1N1XL38hrAafS+rMT2gVTK7iIJPC9Ppxhd/Tvtm2vuKc/Ggz8YdGoOlAcE+a8Bk9bAPU8
yiEQu0kGIYeXvl37ZORb3wV//6NQANoEe17AWVsVKsp1IJqsv+3TmoN2OjTwwy0Pq2qWE8DvrxFk
cASwg8OakgUfI4utGUjP3hPe5tkCzxjcwAwF18W9uMvh74dzHvw7dI4cpmCu/tt64rduXhUAOlMh
nl0S8y9Tg7d+M3wj89ED60KoFLD+6u0EzImEdKsNz0LodlxMgXChaMT9xDhwtvW4L9WbqNkWeies
vW+VOZtwtK339tjkFX+gTuPOKNkCVwYoyEzWucIYl1wgv+pVXeZDxXzctOGjAcGneHAIDXlkqcpa
rzVinCUbxH5ELCTygTcSsS9dY7IQRYluScj7qTS6l7i7RoBRKJ1OZ0iYXh/ldbHFnYYunP4S1cPC
U+1tp1qTDmcvjuv1vPKa2sNQyGfxyN1f3dvYQSJyHw5pE4cLPAEjREuJCPn/NtheThbwRnpIr947
OD8mj3N1KTgoAtuLLL9cRn0AHqsUoSbiL7ItJ436vDBHHLdBiXwY5GvFETelnmHH9FS/lJ+/I/AG
XOSXRwmNS26zbA43iNqN9uIdRhR82htSqlVLfkoXThC8o+AH9hP6O9DdSYOsEKD9xHIC79+13u4g
dTAY8/O8YQyu0igASTkeOR6/0IKh5YpUrdyEgkIkGqLrBkCJddekGjBVot6gFQRvSfxb27RJCBsQ
cpHuvpEpG+Vl1JYqCRi/52A3uhal1kZ9VnweJ0fipOvt+ff7XVCpqo+iughd/U6nk306m8uFMzOa
IJXplRI9D4F7T/NVAhPIo/BliYgOM3HB3uENidLvUM9Bm2btX+Jqv24PluOfX7vZjOBdoG0rluUF
OsGt4X+9JNqCZKvhKgloq0gn3snK4eoCBj8izcJ4+s3x3WKIIVJ5f/eGr2PtLbMd9raO5RuJCc0G
L15JuDC1x98nT/75RBim3dXcSFT51ch2Llp1Wr9dpy3fGuX6K0hvbqPcaPy6BJmtkk+nrCyMGhce
pMDT0ioLpV9AU6pXdFYlcaiwwxBJ7Novo7FD3OE3zx01F2VOJdWRlCWQW7+gqdMIvwEztJ3cyVqO
I2toUEth5voPmwCb5+Z7+hKTrvGv+VY5rWiBysgw7bRyDzJQb/JG2tBL/SQvDGr0ba7drF9eIIig
pUKD8THKSu5OQYVqT8lCtwRfPnVSRKm3vVg9wfu2WfxfkJ4VjRLSBHn8AkRGIitxW94QASwRI5ib
gB+xWRn5N1je6PfzfGSCDDFEtfdNuiAJe0K0Zla0YcBESJ4it3Ty8vhj4zzvtvku7QuHYOKMin7x
rwsDd/yfPn8Hn7cwHeQu2BzoJIhnydzk9m9L8MeqlajNxPGp3gm4CTNrQp8geXzGapybHgVKm7Ez
wFEcgYvkgFBqXrYFHGqexnvdAZtY2xaMr8dW7ZoQtuxTiMmEc6dkTLJhrZ+wCz5oO34NAVe8ujVC
R2nVPtl7DGd3jMtuHXgRx3q3/ipyrwsuFZddRejx7JgIHi4aZhFVJDvWCkFpQjupgSHN44Kr6AG9
qY4DktxmCtupTb+TgS3plHx31p5ybaMyFsciSu8hku1yYAu5N/haZ+MFUm0rXFNmwZO7WdevHIc4
XBmqJ1IdFUSosOqDnF8np0Ow5bGhNNi2hOLG+kdOQTJ7VjOzUMOyHLJ98WdwipLXu/n8XCrH0HH2
nvCLu/UsyTczi7X6gD2nPwSZ0Xx8FWgZGVl43A059xVYlC6SApsBoa7xnZkwNN9/YeaQPTrkP4zT
QpiBGi9j9UPDGB5ed7yUKlMNdV/INwOQELc3dFSejag9Bz+z4O1WYxk24fDVDCguwR/dzzvzQl4h
zatd3SgtgbfA4gFNzp/Ku+6brxLhkwGHxdmGdBdccwnbfZJmu7PhtKEih86phLEB2MlZs/MZjEAY
KbNgJHktK1zEj7a/wA+38kbH4dR8K930BmcqDajEE0FlgVZqNjOZ/jSF5k1dzCWcgIU4nlxmKhWw
ceS483fQNDeTdxAssT5YERttNfrpmLzyDQnfBkW8D7JGXd5r2uHCvelDHP05rWy1LnJDOLFo3A00
mNxVuNeHlqSA0tDODcuQhSqwUJS05hz2ZYqOzI1Q15nzzZL0TZb1sCk1kC5CQx9o05PLZrtHRBBl
WMRz5UFMgQwfa7sI2CU0cxW+jooPpsUnACaEnyCN+PJCkPLORDwdqGnZvMrJaFBslQ6VhB0jAgm4
qGeWqAL5oAQftAL5B3/CplagUSSnZyco7wyllQ6QNEDExbWH8Vf5HjYfSn9sXC2zIndEyUtZ2IfI
LCuMiTDnGtl8CbtTVQaGl1/9WcTQ2BM4xVOkFuV4LjN0cpTf8zvxGuL6P0JRu+fj6L6fJZMWcTp8
DLwTfCoLXL/KmGuOO7n6Tea0l8OJhie3gHrFVVfTOmHZbJNtHiQUZCSdq8ducw7k2yW7kf0Je8to
Uu1yRfVpheQn4Spjzn8EVUbAPR5X0ElYzkcTFpS6qJAGhBHxku9dtIqhZpeAZYIZH9MK8AbSqrw2
nKJV7yaZD2Slr1CbtrRujb/Srl1kC95UrMqSKOuaUZOCeft/lq53mmwfgUjKb9oq3n4z3hZAkIeS
Nb7TvJRWRZL6arOLuOCJl5M5z0fFO4W3KuewQaEaplnvySpmzpRqVEIFcr1vx3D/L9Vr39J/w+Er
a1bPgGIcM+i+DTzbM5NRBkCg7lVNBk5qlkkPNFlNnUt3sGc6x769GxYVOCIyJRhXDPf4WETmnk5K
+d9S0AL/irPerg9dQO5TLbL2S15627K6qXZu/F0lLCIXk/ocmjHXiTE21jMgSApaBU7iS58JBcPB
+aagJsE2WOXyt63cHj1Pdr+38r+C3jdlBDwekm795dQK3ZVKlgOZU6upGs7nEmKECtKkbdFOcux0
CV76qIopgv4qSauBbpPgubVyeFoW9etwrcjdHTuRXiFV4h83ta7Q/1acfU+HTtX5/IUSQeLiYrLl
myDCILsm2XvGGTatc+7ge2iXv0on9k+ImcbHT5cGhFT+qe2QHSitdyNxxSg/lRrqC6z8KkYQEe/w
NEbT8rZblJjm3/2Wqn+W+PMqlCNKlFiklm/8u0FCbBxHDdamxdqI6orB+iiBByiRY8oB/q8nCNmu
9GGqL2CNrO6rkny23HQRHzFJWMSnnz1Jxg6s2L5kLV3KK2v6oXETGFyi5jguGiHCLQ7GItFBIy8q
HZBHGZSPgLbn+oRWTZcfCDaoTj9t3SP4pXJWsAXqCe+YP9gOM0u3LtmXX2Qy7p/rFdCIbm/mahx4
jUhYEmUS/2A+xpHA0CY9jInWK2GDJKk6re7miygVv2fGlsVd3P9zZrt/y0c8h1h+2UeYD9GKjF4r
s66QjEvxcVmzvuHPpUdHVDupMVVP2f6OPFchf3Dpnaapq0fvSEx8PBxiWT4qLp+Dzcc2GkyxmXgU
1rpUrRERTIQU9RWNFrpA5wggbGqgsGN75w2rpmFZFq9B7JUm/JdwBj76jycnmL7p3geRp8WRAa00
vcDC0zTjt/SLfamUdVhkClowZ2UmEMbGWStkeQMxSD9eNqvavTwVCohPdtT6MYYg0eDVEd6+fb/b
ILgfAk6xuad85vlcxzy3eC5m759KAeNtNotkn8hDJqiDASaXupGaO9XXqrL8jGfcD3ksW6sRVm/H
wtxc+4+taLiXgjehrbAzhjXPCjDz4CqQEGLsSh0krIEuUFPzmjTMU9IRu48EvTEu5ap6UIBSVZvP
5/AzEI+qrKDvC4+5dpgvHHBiXxn08/E4gkHNNRwPAyrWs8HjU/QAVHefKQBNCwrhnmxnJoRIOu8+
5pNkiRaYxLKuFBrxH+O9/KjW1v43DEA/Dxb1FWzKhpiGKDtdKol2EhwBY0kBIhg1fJNzoEJnWwku
apZsN+dlaQDUUIIyu49qZ2Hi4ykRh4MdfLqr66DM58+/FQxUdW/8bkjYN1HS6V3O5M7dh0nuNo0x
zFIYEFbdckj9T0Pe5pl2sNefP97UIlXeDoD5CdXPC4quuwYjVegLYDWz1IfdlvY/UbqkSZ3EtMnu
rNVAqL72Ytq7Qg8uywAP1Ji+LLwTJyMhLnEnBDXSxEg/V5ME/nr50kYMGIf0Qmso3qYDvSI8xObT
iizlR8THaqykOnkv9zFL6MNrvt1V8SfhS+nPAYQP5ASux1YxmYD6fXhK5koS/y2p4FpKEIZCIUZ4
5GNO/aTkSedpBKJP445LMEqALDF6Oabrii7iDGKQepiGTVm9uwTb5Ux43Fop8LM7Cw74xQ34XSde
7XN9EMyq7g9CzydOGW/xjdNQT0dvEA6o45sx9pPodoEa9MjuwzFDNwhSfF6XWHBI5n4hWQ4Wm7sc
VHSer/F2qBJAs7mLxEXnHaOcCfucB/NrJRcxR3PufCdB1v//dK+vwdFesBRCqIXcE9m5xFfiQY8B
XsN2jqI61KbC+dnzc9zqQjwVACDxpOM35vnIfjnGrOlu4a9/h7pgA7/K5RcXC3VBrDNbOjO9h+X/
RKrWB5cZZqFCM9e7AvJxBxBz3qjAUtjVDvaE+VQUhZGE9ohGx4mJyQfEpAmQnZLsiTuRrPg5QgK6
nfHKUvHNBcFEVh9ZA+GR//pw+zd3JhZ/Jvv7IJ3zXNUDo8nB4D7QQPMxgolelLTNwcu4vz0q4L4K
B4Rdr90evcopYV2aH4nKBVF13j2BFstFANB9lq093NgAHNFf6GWB4ykhKkbKIayKqhfGLeYPIlOQ
JnEjc9A/qg9umFkEx9aRLlwsQUW6O8m6dI9TjTuz1BtZhjUFNIuyxgJC18uvX9DEmWj7fzAeixDJ
/4GF0ABQxtO956lbiiQKi1/Xrl4HUmMoEvp+9QJBJlnIbxfINdw+z6eTeSeTXB8wpUNL8KHpf4qL
g4C/vRga84yKdKDMJw4XiEY+Vf554xFQNDGZDSiIwrDnIcYSIDkoP8U77v02+k37LsXU0AjmEusE
4ZDQsxqAlictZZXm5J3yrc1QzHvEqq4i3SqyqVphPWoqgQqLu6IKbn/Jsb9feG94iVE2W13UbgVG
OmSnlGK9Pdt92sxqSZy81Dz0+ukSnvF3MWMsGWhi0iaHJ3iLYHH2BbhnO4/SjLC3oTrZXYm4xqI6
fZ1mW4MVK9oPWtHALHmrclu671NSeu0VRW9U6yE6GvG0MS8bcvB0V3dwYw8yV3ofaHvn73pyHyz/
2E6t8GMLSSv+l77ti+sJHQcGyY7iaxHEqRuQ6WyX7LUkfoCjBz08LSF4ll0USgmwxm9vqLUZ4T+F
0LxAZ+MnSSa9X8xpOJPgMTGoh+hsyVEj2SO59Z/WB2He60UQXd7BGbGv18tUEJlWUV/n3nAeyQtI
7fdca2GcOaQit7Lvr7S/qD5tlvs5X+tzpeX8W1HbLDfkdVd4GiAlSkecTzECY7SQJTbPbsTSBD6x
RwwD+eVdK3H9iu+0xMtXoDT/eRm7oAG+2/cJ0zFA9dnwaM7Bns2ttn0iTX5T96+l4OiSuS/azp4E
Ee0P2kBAq1CwV2m8YdtDK2BM9LsutnrDQzthitPHkSlykURfsryk2lFqAOP+HPpU4LGe+gaAZQ3D
wbXQRT26cYIRagS9dvHlMuCWNlYAzy5c6cFQcIH6cVJ+KJd6y4/4SlIbV8ubdZuU28ZN9gIT+BbU
82tEVmWnxA/JOY914Dw837g45rKVnQ0d6Xyv0R5srZdwl0jVQuENroUTFHvKoYCdyP6dori+cUyr
eKotl0DGSnyUswpaHl3iBe7tGKk+rWJ+SOf9gUKGp4TgPK45BbjDlNlvXqgBRQaZ5DSEeqPpXDRU
fRR9j5VshGSU5QV8mBxvcXWg/ND7W8YVu/cIN9nkQyZyLGMgzBaBdQ5De9zZakLWEpS85S9Y2xu/
Jvcv47VIi01xMqdm4fk+h6WdRNvKBwhQydM3eHW7hIq5uTFejmaSlWiRCO4NsNIJBgdv2XrwxA9d
bP4JSZitqTmKVJR1QZDaVaFhJyI4V/M29N1dj4D4pLM7momftZqGoy7NEzARkYZySNgyptu31nhy
Hovt6czRHPmV68y6iunq8sA/F7H0GTNpXlwyEK4ZsMVWz4wcje3Grt+Ker1u3ieFg3Ww4WvX3Vpa
wX6Xxj+F78STHyBBxyoeWsLuWoYkJTiku8/82BkBRgMkrlH5cWnPjVpcLLVM9h+pnlFVNM2E2U0r
IxOvrZ5ryCfVsJzqGQKA9dpsdtJmVsXxD6a/lYZgD5tqy5yZSx7D7CoEbqwUpbbnnvfubgMXLVZO
juRat6Z3EAETHaPl9r+Kt8/J87SxsBNVfxHfFdz/Rhbkzarszp1Ey5tAPM5CGsMccG+F2LONFCvg
MhcrLiNkWfo/WGliSS52xHOiMwK51xkkDscbFRcFIxBrwstHGZiw+qBZNRPWpQ8q7stNMIksBix5
qoHUPgOtliuTQ5GQ530SccjP79T/H17x2JqEN60w1BZ7T+Sr16L/pNZdWPSN2LxKPhiFqVkfAAoH
ocJc4RReN0b94CumpHwc6qVIlHgFjzMgep9ecfsa6cQyMRgIY5olkvC/p6QRV/9hDIHtXVrQ/0i+
Uw9OQWbElFCMqMCRToDkn99wzYFW8cR1clJ71KtmJQPmyGTwS9SIBALjWvuIVtcTY1p6YUJgFtJf
e8Y5rmo1fjTRTlT6RcPMmPxYL67FgmSRcerfA7R12WkXA65qu8g26rKwk2KjGAYs/8nCDQjJs6nn
U2hAJIkfz0DBn8BgPlJFZaKae3y6ZeKSHY6t4AZHOoLEsxC928U/YKsl8/KKHa/nFjB0Q2uZWyGO
ndsf7Nf2bGLW9zR7Fe/dLejkUDrmih0/7PN9T/Nes/euAjtJ4eMDrW9d4WQEZl3X1ESalPVAfN1V
Z/UiBa5eVD+DZLdbczcQCOITPwp1Q7DyyaO+NxD3smJU+WwACcSh51pc1iDPY1wKXS69pwSHF9Pz
Q0QDJK/Esv9ktuddQMCo1uYDQqcXia4ORvrQEALgc668+dH3ouc9QryMkiMgNIpVCpCULJvSoJ2B
LXsjT4gPSZY4aO0GSvoNd8nBG9wLSC3t8P0EbqxRaGHhf7YUZBCWvuoR7M6Qtn8JphCHT/S5qmiz
zXQuC4O9Z20cwcPE305892B/Ze87w63BEguRau4ozcQ6+wYm4rCsa6DUlwuHIg5qjU1z2SP+FHAz
8tENjCVK4PhKsVFrCukHLoYHCqutwUQXbx2NT0PNvho/FCnna4QHSlV4We9qMqvb8TKV+8odxv2H
WIZo7iEdUgkMJNLJaR+Qzo9XKr/qFDl6+0FIYeMNGMivhDnF9RsHExv5yaI4zNeuZ5dgms2CVh7d
cVpZDIwelp6XvQLNFyauIpOrFf6OHPdjjeJuTklp1BAcLh9BUb6kiqcXn3hRBSzpLaeJQPeWVaiE
Db3eBdBTgixx74GQQJMn1v5DogOX7LkGjoZKNY2HHL3RF5k4ernO4WB2bqm3Ii8MvgqWY+IyqJBo
HND31QqRBdRSOljq+HC57US0p2Oa8/bPo96UTLbrntopUOSEywM2SjNsEdrBODpwv1q1PfSrgJf3
of2hdiViEWi4+EqIjB3Sllprg6WT339xLwLgPg7iRpF50EY8CcVOp6GAO7TN6qBqR0ylFDPPGfOK
95HccczjhDQ+wso9Zlmtu/mQnEm6mKow+fGgtt8J/Ylga9OKyW7/22+G+7WKAghb3s1215B6aPqh
ocRu/+w+CGluy2xrf2gvlHNsiunJRdGz5sWuO97Pd4gmLslnFMdX81TkUgn2myqaMg7plI9yXXsy
cdygl00P4rl6e/PFpor0aBnWAj60SGKdhgK78QKdD01WuhXYxaLZtOMUY3Myuh/Ju+wW28seYyB9
Sw3TgZSw/6F2g+BOnzrAOAkrnvn8MaNmm0NK/iUOlALA1XTKPeD0FWchoKJQBmEbD15LeMssoGtc
+tVZ2cHgWEoo+SO7IZqGbhbgvHb2rbGojHbrfgW3b2bP+Yk5MGLn0ldbdqACSWsw83S+qnFG1QiI
kepHXgWCxjPOd9ZYreoTeS6uNXHXvoRK8N+uL+HrXk3G+3WZNhEXU5/bghD/DVCwTCdUrsRgXvwu
urfxAm4Cx7xKya5YTiF3Djj1oI2VrdpzpTEkPEiGVrlJfWOjSjFexuT85gYGUuip0uhQhSP7T+Sr
N7FrRypk5cItBsj0k0fL3bnPd9ZNqpiiOkqRegajyFjl1LrkFfHqvRvGcvvIVMz89s0eU4VE5hur
yAmXa3NOjNxyliHMDUW8PN8QtwM6UWYHzFsloVrk6EL23iY2ghmKhsPM4Bee42el1CTIG7b1nqgb
QNRtrmL/CXimiOo5/S2ltrnvVeg8zg4VY7cUlE6LaUIm6IKlhF0VdHnjTgrnpTbvm4J+ypxXTbu3
+tWkEvLuLyKgmmMARQO+IDuLEztsnexlO93BnIsUiNxdm3MR6IoKknlzUnsi6B7KDIE3+i22rOHU
7vALVqArlXlGJIfFC1nI/qCN4Artm+aV5A77895nJhamU4I/1iDxt1N/5/8YWGAmN5R0nys3yPdT
2gbNnFXjjeBE1EXe2pf+QJeepIO93gS0IX2dSM3k6Wti7zkctMxdMT4z+CF15BxoKIadRrfzhks6
WiTPOyOx0ueCGObZEN7hblUQqqvnUlXyH/fwoyN2hFwgfBBsrj1BP3oZAyWVj8BCPCly3X242bOW
fmIJZhyamDUbHo4f/oVtsHabmEguOVvM/VFuzbwbqi8vn9DOMifp/4taI/hbljjHn0KiGjLwzgnN
ckOCAzyeAHuYpJpWGsFPKdp3/d8Qas3+dP+1R9L9J2yF0VWRTUKbFgVSMRfLHSpKx35o/Wlk3LDT
x9BU7hqko2r/K9F8yq3X737FkGnH3oTUd1ZoHNgG2WZjyQjrEUyqnB0nENpV5OPlvw/1Cl73Fzvv
0s+niGZJiyN3zI3q4FK5hWuM5KpbW4X9fuuiH3bp8iYkanC0JDdUuA3gcFBK8DU85f4EqW5U/yUM
rHiXEFtFO5ckwaKUDbXZWcbyIG6QbFMLcjWmvOT0/0Q/kRTNkKoQ3rYtiI4v8KrBpemf6LUqMrRM
S/CXfwciMQxplDbxl4vWjJ7Nbmti+xFzDtgUGZIkNdvbIxBnoNkogjrcB5fBJFtc/XcD+syGvCdP
bo7vrxixdnE4q4ATAXE+VKxHvpGK61Q/ohiq1FApQF3Dfi1xmjGFErWZIlKViL7q8XIkAmA3sdBu
WBHKeR/O9YYnpoZXZh8v5Vh7JVTwwfCffoVPJkjp1Vdn/rgVnBvF8WwsFjuUrUL8PhMKeVgpWDRj
T+ZwCniHkVbm1QO82DGOSjF4Nzy6I8yQnkTOaLP+X5ElzTh+vzsCKCVnmi715xkLX4HJ2fpPoETm
lCCPNKxmw0taX5+KpBu10W0OsLp+gqR5uEGy5QBR9O5RjLfI7MtMA7sNNMb6bC3AxJvZxhAnWFIU
Re8BtbUhFlcFhndQyfWQfSAc7OxgNsM5J7FNpawNt6D++YbjmkExxBTWWzuqGYL8EhCcwm0NNtgv
+cBo2EKOdKuKNMOPiV9bzK9kI5nPQmg1c/z8U5v1BvynTyXE6qVB0OuGRkjUWLDFw9wUfLFmJg5o
L1X29WHroS2nH6M+7ksbLxLKyJI0O8CB0iv1eYiqSgf6mDJxAPLcPPrb2nnEmXEkKP9mQNEbGey3
UG7EbFLzDOsrBw5LgWwZCM+R1NiBJ+Xcq04IFSerNvjBNkePTtqajz5B3O6oUFGPTUmLvDIS2YLO
8mYZ4I9Bpf0x3ZRPlczuicQrFAnJV8NBjedExicnVMnkezFYR85QP/YnGA/RWJ9SXaZJ4BFlMARU
UoT5aBsYzDuOHnzaydh5nZ8Q/g7FRl9mb6lK+h12hX7RnFr4x3Ck8IenFvYRAannS7BVI6E9kvCB
e3QYLPIGVSjHg6Q7ZY+QfhIdwl50g3Vu0YjAq4Urtyp5yGp6uGixGTYIglj7s9WaaCO4QZc1d+Ej
VWNJr7240nOOT/R3Cy7UN0ZWIWIzDXk9U1LhdzFNsReB27sjdd0XpKFGkvgulQka0ILD4ZoC/Jy5
MH/2S1QpFa2EV9pNnyJadXPvBaCyX4nQPHhRhaNcQn+T2YoVyV8qHKetVc/R1ieGG5KLuHBMJ4Q8
JXysBFqJZC2peXQsoylyG5bq3y3kQD4mKPOorknLMYOPBqawZ8Zu+NVdQTrdHTFRXIU00xC1nscK
6Ypd51gCTj6YDbHn74NadrHB9a3jH7rafG3ERmabxVYvxx86uH8KYknZ93BMSyK55pOwhy1vWSXY
mpE0Z9ph3VETMGE7Fi2nDha0OEQXRD/jXlA+YGDTLMj1/5tJ2CiYQAWTgVCMG9X/5OIzGVXzjdW9
UhRJ4cosGb1X0qyFzcj8OLKbA+9Gtvn7HBapyGQnzZDS5woUGysB8dJ8sR/FbK4azswaW/t8sBYa
ZenS6IgbaWQRTRIPfLxEwk/xBlxT/IYBSICqpP6+74bsert7OgJCSAdrZFfNYyq9B6Dht9QeNAyC
IFEFNCH4PU7axetxv2aRtq4t/NeeRHYHEOt8yfdscwmfxcPI4c4RLoIlixHLTR9kjkjlsRWmfq+M
ONJ6Xj7KlTjqyn39fRikdYSkaIlgM7ENt6SuCCrrAeeYXuGcIlRryatDlOxDKounT+OaAqFo/5G7
YtL7RwuaW6syBVu6u5q3dtbnbic0+1QTRAivy9P+FRd5kMtrhoOkY5h6JShh+A3WdBSuKxHRKyD2
As/2MW/AvLFdZDlLryVqtszlc4T4n+RnQDjnGY8vOrd7yEMG303e1Uz6BjaFRwr/Yzs7D2ij+2u2
Z1j9QI4/Ph4m42O8hlTBfTmzm9Q/hUg4a7B0ILCZukjnH8QGqn+ldDbgiOiOz7wJ97/KXRS3KcME
hA1iffzFl13XvWThYNMQbPSzg4KB8bf+407r2QbTAFuuHfsfqUP+9hoDPc7RFLWtpyFHLKnZ0G+3
k0BdHqQrHS8z1bd4q45TlbTlngOolPxWDCz2o/IF0xCo/lKc+VQ7TeJB3PlmmXlmR3tCXctTqCIG
80fFvMbENEmAxFygSRCzmW5MN9CHW4buSTl3TnJERIPxFpVKq8GrniLX98z7XGjLBQPCZAMglscZ
k19W7q8zhxY30WGLIJs84B5UH8sZIa1QR97wo2GipCgJSuAd4BwK9A+Yz6KPN0S3F4eaPfScbRtg
sZni5nuRCPdXW8HBo5WHZtUCbvHJotvTceC33Oh05a9ddXNfazkDO4Obeh/k6xy8gOFY+I9UmiTh
I/CXVFgh7ndwek8v8KkBSvsXAcMQ06n6ggXOX6kAfqOSo75zwPMr6Zheg1r28NsUZlscT+8U3uuj
awf3O+3Yq5WzFZtRA+cAqPE0MetGqqSr5Vi+p5Vu1clxqdq+ZimJPJiQCl6Mi+iXqGXzVJOF4YPu
aunQIANfF7sK4eZSQ5bzYxy/VVGsTw3mYR9Vvx8rbgdGzt2dUTi9FeHph1f0RCLCucc1CnNj+9k+
2XazYPex22XqdmtxPz3w0C7tlE3MB7U/qe/vYYxjbkTPt17+07s9jB8gt1rCm9SfrIrHk8zfyYOJ
66IcyY+9GJ3hPijIGlhsrKAFdbdCNaoAmlsPXfko1afqLP9KBxAQ5MMiDAlbc1Z6Iv8d+uOyxsfP
vbq27Zd3KsByF2XTBw2yaPNWtrHKxluIKRnosvZIgoKlQYIOJgYNhtdJ6p4Hs+rozjt8Pqv4cmdH
41BuWtzVpEC+srBmvzciHgPfsc736KuEyebabylObbcWItllIulIhaOcsCMYK0+hVhQJYRusE+zo
OLeJ8z+0EmZnh5dNdMrL30NMBm3tNEv1Fnkc1HrZukfD9FAAZXM1g9DiXVd9Dl/Ow/iV0fN8U6dT
Nh1qHXs6LqVTdUfSYKrAifFKKV0Uopc0a5U3SeBCmoB/sXQcbdVZeCjCKklMWLc+hJn2nXTNm5OE
2Dx2mxqqcPMWDDWOZFx1/gMwUP1qld4O+MUHKhQjTFV7HxQkxO7iLbceIyo7VocIGpLFX1jwW5GZ
QStl/gez+Jaj/ODPld5zuxUiRF4hOKTlZisQhA4Hele0WBIkOkZP71RzdMZUdFTSZUb3JKNfITQa
N9UbcazfIzCH5NRPbOZgvkFAdl6h0JK3a7XeotvgLN9QNUxLYjKv1oY235M4X+lEFsecO+KUOqxL
8hK7ojo1W6UAG4ro+7PRqIb7yXpb4l/1vZxgY5mMqtCqRXnUrQDGkJlUk6IxZx/OCBpvHX9kUYd1
Pq3icY/H1f6/awJVL+T87BWnfFhyILPUPnFEHLZozSfMbXpYgmoNR/ADabSlnw45Sw9XeHmgEkid
jbfLTVmYSH+BEystfhJ5YCrqA8y3w7NodFTLfF9y7+CzpytaYtk5hfpfjnBVdNkV4VKouZ0i2k/J
dOrjFhQEJ298xLoFYiGfqrtjLoDToM8+9OJ3tqrf1hLt5j4NGb1i52cWrdcxz7WS1JWXzW6pbvAe
/ReeLHjuuXsiB4e2TqUXdFDXce5xQgDYFwLaE5VKYiVGvgm/mOlZBx0nsV8294a5vAhC8gg93Rgf
TebQa35Qv2hXZRfpPWWKuymIGOjoQaD1bnqvf9OsJi3tXnfYLl30fHlop6bFEI7fHkMdjo9x1rJx
wB6XphTFf9QZd30zhwbebKuIZ5fPW9squ373J9wu2jnxsOJCK8QuyRQPxChbVswbvL5t4VNoaX9U
uYYNT3s9fHu4LmqIjjxqt1smziNxicsuc42+H5wRGlWYMSZ5H3Kwx6G8RhUyn9u1XxT8MBX5wVUs
P6vvVUvfXQI3uczakM7ZYw3v3Z6GAQmIPPnDVzDy8aPZuZO/WMUm4pups3sUggxJMvlMXpY5YIJk
aWSr/mGNHIsAMgCImXk2gDT0emNtgsTCF3ljIDGoNqmcQapGoqX3KNdO787BbHpj6xo6wsjF8zlx
985VdX+nNsSatxc/8CDzSWfWfymq3VzpZqXVTOqMtBsDfiJjGSbVUaxFHJLGdtuX8wMVM+Qgy7n2
jyf0gnoK2bg/vQhvYajPvUpKbbIMRtc0WaD5aeIBAhZPi8/4YHe5xwTVltCiDH3d4AQfaZQczjjI
FIrxAFw+KMkb2WGK4H6V5QM2Ypx04ulQdnuA6/4NtCwEruq9Fkc90BjTRk8hFf75oJxt88swVv8x
8n7F1JA2TCWrlYbuj5LRpbb6PqnfbWX/NQubZc/e43uqIcgNmOW/VnFhUyAjPbF0bbdGKnPr/ypp
uU+/adYsyDcQXWJO9dT0Ge+Tvd0Gen2Idsc4Zy2Mc+XewUPSi7OZMegqAEaUJvuMhF9yfSLl/x6C
ds28uv7CHzJtpLJPjNmHj0naPHX2akc78n/ggXLB+90OwjZalmSp93acAUtjUTNADu3i85mc3tu5
ZU3/qUfajZF/lFsu0LvmGQhUhVrxDvpaN6ycJad0+wS4YSyWnlHuPEF8W5Bvr8djm6ByoIg5s3mR
twPkxIEWpWsF6x8610CSsHv/SzlyxsrErtHon1X0KDODR3QlvtR0ZboA1SlLUu1dwmuGPuMvI4eT
sBP/MjypD5mN/QInafd2LhGLXyTTsxsmGZeVbwZaOiUfPRVoh0XIAMpPXFBRX8gu8BfDidtb7rCM
IbAPc9GOyQzUwByBjJjhcoktdtEzVcKGXeOow35Ki5cFGahD9OavBL8C6e0B6o201WUWAyaa1QoB
nWxT6M9luYWiMvxpplZQTzOgid6eQaEYejKszEmX/CmX0zmkmPFz8FmAwA43bcdhOTZIBJcD6x08
6NY8hDnJ4Yf5tLZXgnLVTQ3ZD+WD/3ME6K/k04f4tmi0GDakWuRLfu8Uhi+BfJi856k7HWkwnhGA
uq/YPqTuiKgEMRRobtGPCVqpMulRHhYhnTnRGGHkcygMtMU6QfbnxFauHbXVrGZwB8YmLBySwOAw
yyNBIYiPaAOF7w73N5KIVCLildm3oDEleBBBJRsjIWKbX6vkoh0YnV3W1gnXeD8ToGKOttUlJ3f7
ePoujcqzkZPSwU4C2NrsVVC8FsQ20u/mSo2lHc6XIJZfS47lPgSsx2t2fabjOsapyBl/RWmiQi7o
P2HzpGG3+ujfJoX1HX3reDbQOiHeA38U99t7pKHoPCi1EGvuwUMiulIE4Cga6VrnB3eFIqfiGAzD
pv/jhYdMxvtyp1YGE6S/Oe4s3C1pudEx8wzBtDufq/AuxyQASu8v/WUBbWg8zeDhiZcuf4q7sI7a
kmOIW395gMtLdbj63Ng+rUTzcq2LE1DcEq5TwCPwGhGnplyMrRDz5YQRNKgTzWRTgtxF+DhImkIB
+xFkK9f9GzYJKY7kBSBJghgx5UtjTZ3Xb+w95rrNU0wFHmueuKmrjAOPpwcArKM+wGW3GTiu88dA
mmPwJVHPy3K9b80X+R4ntbYgrJ5k0jSUdMWHs1Pn9vkZBe6tzs12qrLj0yVC/w31I1WdoJ4A6GZl
aMfXC/nAxaNNA+diTQSuzadytc2dJRO/E8Y+iVbtzgfL5QDntD2NRyyebiJnQDwW7fW82nCtSIy4
Mcx90t38naWribH6TOJ//87D+t+AJIRsY1d3NiMxt7W9ImJ86ZuAthjysRu4vxKLX+gUgJd+0OgV
SRBeTPDFync2QzEe5ReVXj8Jyz4bILhBqhxFEmxdEnkThLEqg7D1xasy3xFohSI//NcRF18G4rUg
9Vhu0yKp3mDNGgziusjlXEY9tsZ/FVac5YGj8sEC7MgTT9/gZPXZkj+3w1q21xTI2T+5wCcChD7y
ml0+KT/qGLTKE/BDV4KpZ79wcEv+gz2XzJ4IPZQ68Q8+gWxZPLMfze/EdPEr4Tw0Xr/wGE3/4NHf
NuhouByRDxJeA2lfDMbt4lvh/lg0SmEsZYNLrxs4LUf+7ggoCq9GfHjybluHMa/j7ZAt8Bcs/aa5
HLDH6/sNBVmKJfNZviWCAFMXYgfzvWjeGU2CnTulP8aDTR+xoH0UEkhpWV/tIFSkghr+A8tHB7ZO
jS4Bo6ncDPdA52MOLDtumwhwQ4oRfQLN9396szerclgxsnH5ER0SA2IYX1fftzvMN8u2G8kQqQwL
1eFFcP4vpRB4v0yMVyyHFPDVMeSG+N7F8tYE3CeVaIMYiyduUO81YRz+yMJTtEj4tf7C50EwZgeG
8UxSYsTX6nuw3pTLSgaunOwDkfZxwZDFKiC/S+Q038atmDn50j2aSL2iZmZGuuY88WPchrpBMb0F
7okLgewPFCGLU27n5qC8mzAER4eoUWisoOuXdJ0yLCoLCteIIHajo2cATFnSZdSOoGgCyYJvZzKj
0NfKlDcZfTepz5nQyg5fhQn4jstfCaZm4CW63jOW/WWIqSjl44EC9hlVxMuQ2eh70JFUyDPjCFcp
4ofXRpYh6DbX8ESlzXT/WD1a5kDSW6gHi3T7lJmJvlp791QNbzvcvvHCEFgJH+kXXH6x/f8HzIh4
4tcgJe7exgekbaJYLRYuD4arcxatDTiCGbxGM6GuoSdQsc2SbmUD0i2btZjfdixl7aFlJDLgde3d
0AiZmo/MafroUenX9SKGthpCg/bMoOXMBdD06gogUl3a5Mbo3zdRXk124CsRdK11NEuEqxAdOsQG
HRuFiYZuhAPVeOOFm0lr35O4KbjEPUgPihb3s8UBvQl1jlwL3enCzIFlpkfWUJNO6TpB3K3aXNE9
un7PD2/orx8mzYigeWoWzCGCz9frY1pBRt1Wesua+/iM1bUnDNkigHvCo1cg0SIqd5A5rCrbO5oe
5IRNyeydIaRfUNWpSG/RDjxxevlLoMERN6ail3JienAwEyhMm+8yuiN3wYKL6G2p0UGecz25tF8A
eCMemL0/LuqO208W/kGZ6V0gdvaFBCnEkxiLlJeA6cD5yzfkV5xRMMc5PArR2ffpFm585sMkgrII
cAHgogRdK7H9JMojvavtOC+o4xve6iYf9FFsA4jhHYBraykCvZREpxP+xYWU84h+JUuqJxcJ+oDG
musXxitz+KWU+QIshFItkC9JOgageSrKi4CPsRnmzNFAlqo8XMD2HxdHefQtlo7H36FIf2eCXJ0q
k/0Cgm4isJb9GtggtoMSo2La0ODcu3JQIMb8TQy2Ts7ofJLxP9XbCyLDdvdi6AwwzoM97+p2Giz/
6snMcvolUwyW6Ifv26f5EGY7YyxaZGXqI54PZJEy70QK15mAQ7DOCA9IBg39kCAK5fUldQseBMwz
8qL2XcnA9NVKufLyhO4YwJIEt0GNhcYCGIseRobdj4K82U0ltVDcG7TzchZxBOPxDF7R4rHyzek1
kSzLv9fnUqUxWOVutDKnBVQ8n3JgSEagK6hFmmZ/6blL3/TjzhVxj/A+/dLRiDoy+DdGRATQgchQ
ILs7KRabvCIPTxckfxkEzi8Eh2AjuyBNEwlEDdBZQVTte+Zsbn1eqbSGgQXxk6ZFI1UIptYlie1b
FD8mGSjDp/P34diGUj+w7sdKHvs6OifhVzIH/wY0187qxLXpwrBVMXd6X0LruCmfPYzZ3+CzpNg3
uHKE3AYtJ9LA64n1uSZuPIhzWqXur1kttmX/xP91k15lJ6lb/fSji8vu5bdTmYI9FAAcOFo2dCEK
iehgJ/21zjB4SHUkWULFgyJ6FZ/TJqt6q25stkAvmp2L+/a6jyf040fu+xTtTumNPRZagzFOMzw0
khPhtwl3we4uA/fq4MFEITv4KnEmBP8+RN25y5LEQBxoRW/Pm6oHxv5e0bybAxFB1Aqik6Px3AG0
NWwjzzs8u9pI/HceEpXbkBvapxCnsA/0NGN2oSyMmVvE940ET6gMOFRLSnDVQldG7CO0fvEyWX8K
O58D7c8NYaXI1sMEvVF1XkZqz8/a95aTxZ0gSciHmhG4Vkw+CQLlsySItjiI6vqDXl3SSkeFPBop
F72N8/I3++mkL3TtXRPtnqh3gbTXWGPDkJ2w6vCR+0BLqfF3pXb35CyTOAha/CagU8F2thxomS7m
Ls09G2I5jMP4HREgkccuhnX0scUO9W6IqNzm/b2cocF+JV1j1rIKS4Q62Q4vXs8BzV/OZummSdSP
J39YFUqAXTrZRsACQ8iWOX8pTuJeTVPS76Z4H9x56G6NhoybZkIJnU9vpbM7SlrNZLn0A4PKaEM4
gouxY8+KdNDHp2ca9FgrbXP+KIMyIORpPVgPmSR6+7Oyi60lZU+4an1StGaBSLeiphnbox9Ide0S
mbKY4/8g/g06KT+l9WvC0WH5BlKW0SC5RuqZmfjdT8vE4V8PMqu4EOUV5hlFpSgTmrI2Lkm4NtlL
DsDP8xeJ9EcAnDXP9iCdgqbPWLS8N72sX+/W5YbhMBLZiBpskRPqSvuviiB2YvJch+FIJnYllVA+
2PJ0GWVHL4LLcwD95SHekN/xFsjkq7Asoh64dsf1PzpwvmbskabDoL2gJrhbu3FGGH80zzQsUrbj
1QKLItS36LKN7CHLndjMQHG4WKc7K+bJ5o+vu2D8YzgQm4H2olFPnXLBa19UlAC/qRBYJsoDAauR
oZwiVSTUL0bKKZn02cdYyZf+JwDWGhzOtclp8icC5NM+iJjYURUyjT5pBMSwkg/L+2K+gSjPqceA
W5PvlnW+elO5P9qlRMoCzSyLzj3xpCaHBWvQLKsZ7vzswR2hKpOSSMvOdaYB6y+lWgu1YB8kB7Jf
8lh5yuiKOS/0F82zPVD64WAF29qLZlZ7R8/RxfQgqhbM8lVUKUJCk8vtk2flHm21Mnjf4Vyorho3
nUiAR1E9/QPGMQfz0Xi4O0rLREYMI8qsZAMoHxIDc7lgc+TGdeA/AMhXFbNsHx6fhqw4HrgLN/WC
xIRj6LR5znPWZJIQJcyaQZ71n9BC1/fJJfr701uM1MMyNRPRRh0PqBryiPGj6DmfhcWfCutpnxyW
EBb/E38kFSS14mzy9R4Msg2OKxxvb+udJZBQRmYortrdz4Mfulf/rGCZ/tbas7aCgNw4mxhuskMr
cfza49oLfJ8566HSz55ZQAhzPNljjBt1GxdSWZfL5IntHMxNsi0Ku/XwLZbp3puRmohuKGUI7W9d
ZdN4yYwlDc30fFJIyXn6Ap5gTuaAGLPlmiJas5Kv//C/Uh+0lUEhHjHy6WP8VOBATn5oPvVyFPnI
danGG2fhAfGyWcWkYxFu4cep/CCN5x0JixgWgQjpd7wf2gmx7FYEbZHoDtYWViVC1f1N01XncaLl
llFGftVMro9pisWagKCW/IVWceZRxBUafp9jaHxrbrANIjtQzV5j5QYsLWsgQPBk5CNZ311shUtE
7lFI2Zo5jchL9rZw2FSxDjmzigI4viUzCoLA9xx+FnNx8mYjs6fTTW5BZ1PIsDomWArgVoGlROKI
T2AglXKJOlm7HxSfSVVY/pca1ZDvDk4PYeWNhHw4PRX1g4zlt8chlozrIIP0z/SkM2Be2JQ/cP7/
+XzObTlkJWrM0tPhExhyLzJNafpkxKQCZdNYvhbWwHjPCN6ZeY5FvSaW8wCKfg9bAsPWrv+hY9g2
g0hb0Et52fcHq72jdJUlGL45xRLHFzWuesbFBlF5DAMcNsSX8Vb7B0yoB7fKoBNnemVeTcwbOSLP
+e442KEhK0yN1udLtPk2zXmY4T/ZeaAb9woSJOwtVeHb8pHm0c9hGsJspHI19m37NlmnPwwdtdhi
rgxr+8rOlxK/PpgyE9SB62xgax19iB3FC6JuIPjemCHf+jK3HHnIqvWjR+LHBXmQ8tRGMYsvALm1
2efVYwIWxjnRUKGWpNJgZuehrugtnnwmrFiYTCqmUkkh0VBfumqV7sbt5T2Io/Qqj60w8O4W8M3m
CM8Ne3pI5qN7IB2NPo8tPsRHGHyPHOi6LMoew2nLnqdZpgKZ9kju7/TrhYI/Ak0MWxRVVu/0Hibo
ppwsoec/FSJVj92tbK0tQX77jv03eJLW5PQSKXZ8JZx4h6aBsGy7cHgIq5oAIJ0FXme32dxbblZs
lnGK7Gzx2QWLP6qm30IoyIJejaZ5nPDzsQTqIVeNKLP6vI3ziWLdD830DZYn+6Hiaz2MlvvERzPW
uPo25HSGzsytFkpPUl90XPUMAI/MXJEJiz1WAMlwhE/Pe/B5r52yN/Skeu2hbUB5HxHeQiezzsX9
JcNGLap0w5kKc3uhHIiU1strdmfHDQLv590VhdoC656/tzCKRFklfva4Uz+z3lcb9D837N3AIoJW
hbMQTJJSNDRJ5wDKn37pUFPelFnxKsb/B5iEouT2ATEpKUKjuhm1HZW1HwDeR6vrC3VDC+fp4iqY
WsqqW7XtxAVv+stx7IPARBaCyw0CO0oQ8U/DQkcECQjtbLo7PguT/oWmaRlxT5e0wvVR2L/z0aso
MMW1o4JY6BsxmR3LOzXzv83YozAwHfzp85UAgDO8RiCc13eU7zhZicCCi8QNUzgGDArOe9F1jnTs
FA9GcZtQHLELLrETUGf247SUWi8xV8Q0A1OoXFa9srnmNbZl2zT31enM4Hs19gqVobWMhalOrI+h
MW5UUk+Fu+qquzrJMrw3khEHuflSOu7nHRkyfNXs4HgLh1CEG7wxgcpQc93Oo/r+COy7WVZk87Nd
xbiqktFPR/5A4XVvDbkcQYzKUr/7nrKx+9nFTrJis1fl5Qfk/4hFPisbhU8vc0/TWLAD5JIjSLo6
407USweqwJCy/QlB1nTU1RhD7oos5CJDpiQlEhgr6TexnNPt9OdfHesG+1K3THMEyn1MgekVq7wO
E5LtgCidiKGokEekjI86tJ7imP9NV9h1X68LLwEOLwM7lg25p/VWo5JkyVR8aOuuf5qmb04HnlF8
vLzSQdnzg0B/HegGJ2VNEEmLq15+niuZohBxhzCkTrqbOQ2tcUohPP7MQdHcMULxaupS/MZpkHXD
lsBYSw4QMpTCE+PNYtMgua7yQUWUcQnoHInR7/VUqZApCSOSaFMl5x9AyjhzcRx7WfasKzd+P7DC
c0XUkwKU2I3Ugo43gbHMCwihR4lWY0zKq70/YHJJErsNz4VNpwO+vP7hh9U0Zc19fgQGiIGvhK5x
bj5WRtNLCKCRRFbn0UGhsopANoeMmJdPdf198WIAz9q7bLyouJill84OcDIcc1UCGBFpCRLERWRC
sWttnbFw9oe8s4wQjITHqHzrkDWjMEIeajeL2LZFjmr5gOZJpb0ZzmP1Q859Cmh1tujhZO2JozaH
AiqCXqBsPr8aySWH8lqS0vxrtAecS25KIDs2iP0BmJafZh0iGX9Iig0RqBLcsFbv/up9bTg1HC/L
qRFqHPOuuxW4edSiRjjGSqMiTCZqIZzl0boht2U7NFwMYfg0tUU6uq3GSaXULTUmokTR9MYLPoT0
z9PrhFCDUp1qYOWCwG2VefWOR+241m17LQxlWmv/81zRu61FFRjNl9FYZZvXz83LSwdiPz7nBmKk
vlOR+dFVKC2pKxNdCI75XnP4npiNWRKxZalX9+RN7nZC3NFObW2skFIcw7oQD+GIcB1w3wy0s0Jc
K2so3cqIJj3Ea750Df+2CK925E7ug6n8CwZ5ARqZevYssAMDyuwsKfBwHZn03SXJmgxrcvChJmm2
lTZMnok0SlbzCXWWzYgHtID/djjRgB8qvR2GtRdrNBpJi/vSdwyV4oFudR6SI14fbnJ0eZTW4HRI
NHTZks5SuxLsNN9bO15xYitR4kAEPL3F6y2dlbyEHZPnxQ3JoKqq8KavaSWFCe+K0u6l4bpGrqY2
xuV/F0+QdpOgqIbgel5iQ9J1mAW06oWg4lV0g0aOUT3PtXKvi4JnMUTa/ld69ft7wr6k7Yf4O2lZ
2iu3trJM49r/9KmQn82w8L9ZAghB9bE56i1It91lkelyTFiqSkT7czZka7xtGWhxASkqTGZl6ibs
nojW4QFs5mUSoHkwjyLvb0jjsVu5CYUvV3jSkGY8ecBGECxFTqvbflWnm/LTIAKkHiBBhsHFJlfZ
zRDCPg/5A5ccvfRgFaxwcgPvCymGGouvpLBBevLwbj5ntV/jyZhA+90v/20hoj9oy6Y1WmjgJ3FG
DE/VIx7mRUNqCpYIIdgEcvhjAlTg+VkvLb/R2ch1ZthqsmevsGhxcWYSzvvEqGXF/lVlfy4sHAvf
k2SX+EDYimK6Td1ag6pLQ7bOu5v6VHY2iU/UYy4XLB7/RKijLZJTFni8dTWV2fGm5g11kXP3o0HH
XBJ3Scd+FYmxqrD3ic2j+kw0cs2wuzAHhyki/x1BrtJ2+T0JHJ8p7v8UZfDemMec144eem3xFQGC
aObLRj9DogdKHBT1rsVXjvrU5rltk7wAO1jUTm1K84tHZKbh4CbUiBe2n1miZqXTfbuMvfTSNl27
mfnrotivJrk4aYG1qxPxaLWTSLbZTqOqkpzxonqdeNGSkt4+cjNL272UFsLSMg8OgReOq6e5f5c5
oxWo5M8gkU16MuQtojpQZsofKxI4KPD/Cf34lSki6X1cF/nRYU9TMGTIs0qO6eJL/S/g5UBwf3+R
4jjhT4wls2aJrmVqQd8oNJUFDde0y3+ZCzO5aH2Ln4+UMctaVSDCYQHD8bafMD+WH2AD0FSquHI8
BJX7NR+NG4kt3EIFanGXNOvDBXT+WiYIARgQLROM1Yp0bBtZnblzmwIL0VkCgZHUx/BoU39DunGF
BRH2+4OjW52sEwlncqDohWcSZrwJ9i1r4lFrnYGU7qcXzrYQPDRtRgR2Fg6SAhBnc9wdaU07WxBK
gT6P3rumLrwQZsA/KRzdEQRmg4pN1+Mfw0mddcfCr9ndXGo69UYbKSrnc8UUvMJEYqILq0n/vlHf
yHNWDLl6KAoKlWIq9hgHwpsb1DwbBMdI0/A2jjNsgWLltJNceOxrM0S8QwRu6jC2BgAWFmI6Zdob
cxHhfHmjDIjQJ1RUHwu6PGVqj/tepMdViayb+tF0bMsvpXvPA34Mu6uiJxWZPHG9GeBrqWYy9FdO
yy88eBB3opIylYdsqj+dyFOKP5zF5DS7j6hIrbJwxcDmDsksRjes606X2BvK0kBhWws4XU+dKOap
CAVCuWEQqONRDQ+ZisLKhAjTrCR9f/Ye0P8MzXOONH7jin53knrG7doC3QWOBkMsoHZc9R8FYSma
EtU11LJqFKDqf9OyJJG4gq4bt7kcwoUCBhnAfKjCoH8pX3e6gqOdEv2/4rqne1WwbWiH8D7+/G/h
5jidcx/wo77wyrus+oUWtKXprlymKOsj/scefZkPcl3MQu3meFYVD2TsgqU/OWiVgrUA32VVRMi/
ZykfDp4NG0ya998vVJUpPsxcstO015aqAQWjioC1wo2CXGYI4o7+kR16E/6rsIAoFYxRExKR78O2
4rioMlkTAsPzIK1udGhADwjymDWPj0Yt/ON1Hn0iXO3yQIonPh65vCETs+ED19cT+nvnTQdBZsu/
KUt4FGtZS/xjA7w4FC+SGhGCCIprI+480GxfrNp2oE/ovJCeJ5JZwZFJqc3E33/bB0RCs79/Z1xE
g/S9JCrhxF8fDXoqxTVEKyxUpl0WKFAPpdA9OQIu2uTKIdhFfSiVWQ5ihw3KyAFTjr5fmZMHPq6Y
go17iVvKw7hJ11NTagXOobCpNWXvVDu/gEW1QsM/XyGN/Gb975E1KUSPhV20l2sMMuZNg3/lMJED
xVtAr6HiqsMPBpah6QKonsMI1+aL9oEYzjHDkeTK3ScTgLlcE0IAw4zXQl903AicXm4FPT4nTaYs
5dovws+Fz2bgBbngAvLx2YAhRHQS33ATbelIPAAdjLcE24gdHlxSoM14tF/aET4VzGb+6ZUXN5nz
GnfsLii5oWuNXLHdLCAXs+dSjIr/NHjgB47HLHbIntTVp7awN7clwSd9yFh4W87bAabccEvie7zc
QBbaBOHwFwb1No90CKiNK/dgHJmYt3u1PsucJe0yuVKJhDoNR90t4XaK20akcc5u7eY+2xvnoOLK
KP3cbl6fkAWmdVh9gE11B2uAyrKgSS2i4BE/Or/WYRK9+h37vyCc+HSr+pV12YNH5Ms2gFprlOWq
IGskN84IgeQfC658P4b3nHImO6sFN5t8zUmd2PGqly/GD6LpXpCFQdA602EKDhL8uPGZb0locJo3
AI14AnI9ky1FBQBajkOYrDj2+HouDTOlozL3nhvy9bzfwjyVzmo2PjtOR7yBuI1kzmBiGrguhw4l
1GDulMi3xTIZb19alRPgbzi5VPejB5SkOirmvsOp+kifDtsH1SLzdpRJ6uoF3EyzXTvQ9wuxVmju
xpUrzsT6h/+iIcqCdoMSQCT2hC9zCg6CDLy0bGNZd54FHP/jbwVV28je/m9kM77Ag//6FudOjIsD
DJUmFjq9CT/YXl3/J27b0EEEctqGXu1OespGsLkfZPb25iZfiNIcEQyLJC5Y7t/YgxzcqiJgqGkW
8HHa2YLngmW+9xSO808gamc0A6g77tkSaIN7IY5M082Yv7W5fPFLX8BbIK12DyxALHXuWHhIanM6
bsgqdXqLYHdSzrOCHtjw9nmtYdYtCq+USsi9QGOBpHs+TYS9EuWrbu25PwF6V/4I2e+SbqcSVFC/
OKGmz4dc0unajGrOtp+8GjRKhc5lruJvkZpfwDMQ16/Ydo8rqJakh7EOYjXiaZJIdFEDOf9SPGIe
S8tzwK79cVtxMEcsyF/nNMh7+3HwO9OJy4W9fHqcmqqsQUe3Fx+M9d5AFcLMh1KOGN0znLqwpM5d
e777lRk63pGzU0SrHQodL5Toy0mCpctux0oG4p7xSwsblrOeBds6ZGuSP7wOe3h9HE+2jpn7Vyt0
fpCb77eeynzfKFzrFZ9bzxQvWp3nc4BM/5QoAo9rPQ/mZ+MDFI7x/wYsEbBZCJIXe2pmDLwulVd7
qcKxeS60fhLu30tiN0//MTcWjUMBTjEi5KCdLW7Pgpyzm2IxlmLc9Od+pmN21rsbAR9ExuMXBq+T
Mxqo11qKtD6YB27aFddIBiKFCakY3b9zJUR87GdowUa9lR8l8BG4tnh1EQHpbjsMkpM7LxcyBW/J
VJBZItLaLKmfvOG4yTVMFYMf7sci12evfhr0Ym/hHruq82mVKftnGGHXCUrn4XoG0x6WQSGBqIlx
2HVC9C6Xq43QyXzs/LiRBvatFiQKqny+3hPgPz8hBeRF+mMC8lyVDVGBTdttAuXHbhKMUyfU1cvA
6U2n6GAdvLWzAGs9EZwX9w+EaXUdKUowPyUgHTOb2yZscec26Jx7ofTvL07ez8SdIWwnav7jCmTs
LmhOGkjT1jXLVk9257SAkQSpNA8TxYE4+rbVMY/xC41EUpTIrfdyIwHEfWegb7xrG8WQ/IKzPMpw
8NBQryrCm6BNPJ+MZ1H4OaPGOZifpVCiylxjWi1v0oX25a60ejbeFV35ug1SQ6keq/Cju/WHzRuw
uTgmCXQtfakh6DFAcp+ctnroZPAFpVcxc79hoXZiUQ9TYzDgmuVhhhShdmkpY8Dv6vDVjtEYhl/f
QShiDeEB0TJCz+HFMuI+9bikVKifvPZNIvGaOZSdI6EfPPGrk1xgqweUaShEiGmzcfQGpA2iX1cT
hWpZ18i/6H3J6ncgCcMa57HzpCdoxPxpeFgEEN7LdVQImxQ/7zzYNGTH1LMx0xjVK+DxX7pADBx5
RHkD1ZIVPzyQuQUuzbjrobArdLZMs9bFDdWKhx6/SNJfQjeKj63BsBJCh9qjx8XyiJEZTc5YUq5s
fASMQvo+u1eXitvdPpQNiGHHTLKAL5/p7M7ZWKp9i4HhwAPldec7BqjWltCEEZwDrHoT7NCFSp0x
AleugGnGQ+zmIEYw1iJMC4WX+w8AO5DFJKaVKIduLCiNXBnSVbrc0luccqk8P6rwN11CcuaGjlnc
mi7As9HOy3fcZe3klUbYoaID8tQQWVBHKieHURvH04gIco/bLhPaqmuAjESy1NickuAPn8AHHqOD
wSut8VVlEaZVji2E4jbKcPa7kGorX4/tR7K0tY68qo08Zf1E/XEl9+ld9JY3LXNVKcFLosR6iKhs
lZ6uA6eLQJHYiSuJGUnLcfHKY/YCeniFC8kJpE5EXSkccICIJE3rP2oAYtsth4dMxFZnU1hnN82w
oePgYQc8TLg/43p2fIfJHGFcrlA1PbcTJ2qM65Opr+CK4PpimYuIv5sCMLmcDJDL8EkIZtEZ/KMa
XxITA+lQ/w/GYm8u0gvpsuHGMlIucAZjvBBt/Ye2rP5BxRyLz3GqrLNWJ4C5OQOJEMMLfB7CUusm
UOyqJZ2db0ySl3he8I4TYwp6illzX2dOCWPWjYIGY97P+p2Ace4hEV1cF6CU78imfMBBIekrlNYo
yjGEM9jLhX8BDZFaABEI7kU+aIcjOIu7NQzyzkmzC77B0kmvrGYAlkGuePkg/jc3sOPhQKyhPGNY
VwU8mTAi4f4lStHbP/hKTcNc3jXD92OJbph9tAollg1JsBZEz29VNprUnvsO3h2XJCvoGB0eD9kM
UZS9Ca7KQMOwAIYUedLhyIbkNdxe7cNJTtoIx15joUkGGqZJ+iUDSYrm9QXT2z0A/NYEq9l6FwN7
Q9wrARsRlZj5dq3RIrI6BBq78lG0lEuugw0+RiN5MWjE2UI2ZJMox3qjWeMxNOs0UJ4fPVhmt5YU
x42VMm3hifTm+JxLOeQuruQz0sSD9GJVwf3ERNp5ezwUpnIht7gE3mflLBlqNdT+eHloyFbR04qE
T4icpqzFheMJqc8xBpb8r093jWSIn45rRQuArr+iLRdE245L0bjfQV49lkOf+3BHl0s4DAl5Zmrs
xd3uDJtBgzTz8WUQ7B2rEJqWLemrImAM03B7wtDbH4q3YTi5Jwch+l5hy1rKLmMQm7xnDeFil1q3
hakFgLVnDd6wq5eRrrPiocZURLzRlm8VPr9VuwLADfAp4sSNIbfpK94/9g9gvk1u5F2ktyHTVSnO
EtMNJ42bKxs3BRgg8Ohc49MGia4mcW1NGKqtg0zRLtgOCyhITAIAgM63t6kT7zo2VSC1dUvd8LdX
DBGT9gEZaHYkwNcjR6OdLonzxR7FBLZ8mjJk1Oh/hsgnuamghptAtDKiISHLU4x3fxitW/PjTz1Q
FHI8LiNmWO8jvpJaHRRSHY5pWWl6G3N7rCY0xIhqfUdCQu0YmWefIEKfIxS0TR818h44mF6aF/aA
l1q1aTA0/jsA8rP4ZoGcGEVVPkgZVboym3GasgkMjEf9MWuDY905p4baRTROPLFg3RK4eMTOIiPy
hnJzGrEWBFRoEWp8SJWCUe0t9fySSiR5VK3A4C4+hBwLeAnvKQxo4c0NmAjSoyyZ+xes2oc9ULqB
+FgSZ7By1Ednzv5SeWhq1zlGr4kKmW2mhnSXsQlPH92orBJlUmFr0C7S7/v+tRDOhriYuYKGCx0j
5c2SNdeE29napgTboCnWzquxyLEq8K9FYl2BzgrkXcX+uXuRejLuOKcymyzXLb4848YpF1BM67xe
bUdL2iQWfaqXZfH8GUgV05eT6UVUMP/fyqy3LWZoisbjbqZccvnYgjdr93/tz+Apw7urASOVHcme
BGcpDZrsI45/IckhpKv5zyHTjUjSPQAz/dxdWbo7lzRIQXoQnIbt6ZEUhcvLG4ta+6vpwSZrJZvQ
ocK7OJPNuFx468QoJ0Ffoc/lxTE/ZlttVEwvgsoqHgbuodns85tXIUveAWWmJdbuYfPHCCkMb2/L
M4LpKc2IH7SrCEBnQ2S7/MTvNUlhgHl7SPAGeKzdEnbEEFh9ItaCWcfsIoscC3I548hT+AAPhmdh
kP9BLpdjiKls+8obwKvenNZ4GXK3SKMmMvZlVB0Btj8GMQ8DkyJ20RoO5l60laClqm8nIVxqTLNn
BxmkU7XHNkRA5e3EYRV9FX4J+Naf9bvYyH/z8ZeqFpRITmU25Bk7bPmVO/tQtYjTXgRApC2UGoL7
KjXQULiYYt1IJ4MLZzS6InztU3PCzO5/FRbPXskCA+fgqOivmuB1C6v5k6BHYlIPTi1FofRMoACA
v7YSxsHYPEvIxpYrC1s/vHfygih4n0lBefb435k7LrvNwT8FGURslSIxJPob1kGVW149KZneQm6B
Tbcf8op77lLfWyXB+a2sSOztZStiKIAehg6XZUBxg71eIxldxHn2O1JpTJceFt7TnhTk5+tkXovN
cznSfv9reouNebp8PCqaaqc/l047hqk8V2vuS2TVE48g/BBqqIPpm++1jsFf+w2xDGA+2/OXblg5
X4OOw1vEJm0WjEBtHEUQoXTrDheIH7PiMCdB4ueK5G6LJXZrbaWkuxl/kod3ocPH/3iUqSFYkSC+
6+pEMutYET8olk0DPQOjV09Ik51yj9Iebn8U0Fp/MRWfOtHe/qusdwA310CgJkHPC92DTvderFrQ
nSn+rnxZ2/G/aVAoKyEO55SlpLcadNUA6qFI+bEfT+Kb5ablfP2pDeoTp9S00BUGikKbmavMlyFM
NiPzy2LoFbAacOINax2e4WI2OXMnWDR+0TGEpogyCaeUoAg8bq5hVzG7yh+4rjEvoTJcHVUAvWKu
9mTCHbD+Ef8Kkvhd4JtAeAgSmLJKR01NbSkVpZdvFDGkSysLSTtxeOmlG0f2F5mClnX8ETR0jjUD
jhNjwZZI4yWjlWHvuhtsdQm+47LzcP2KK1rEapLrHfwrOEfWqtCUIs7wFhDB2YEfL1fcVow84elF
Asidurd3oTl1muiAfNKjf5MUvJoTK6KDDZhnTAHUPVyqJeLmsRlKU6Vh5rKcEX7AJQ4q0NFV7O6P
hyNIQ0OWLQfsKSwinTvLuUA5CMv9h1BibWCeE5UHyKwSmps3GCdaX4WSn4yM45NBEAJxnrWEaCHF
U3eaqnH+AIxV5aWMkzc6vwG1eIh5UoRPDpNVXnhGqsQe8bYvJcLw+jnsBJdnI889V20RQkKBtjeN
sbaPAQbdW7uvr8Bd9W5vBTnlQMyCZToGXSjcP2JkHtH4Huz2dF3IzrkWnLhfm4EAIQs01PvwmwIy
KbJ/nsy+8bB5mtTTuazIrg7qLElJonpAjHf/zI3+Mzzd/MJqx2y4FJEvR1cwNDdx6Qp8PKagIRub
bBrtTkz1I7MqjR4p0QwwePezWwYa3f4/8DrpexYknmtKPHifHbxmDZ0+ozbWH5R+3+6CboFDDfNF
wAmV/a3M8YLacByQocucfsAuW0Pvdrw7FkPH1zb+eOVE3rAeEl3R5leiJr64XVLCv5TAqzDl8528
QdSfkbry1AByBzEZBl4nGtYlNko7BOLyrAMEh1rg2yG6nPoXilaz+zTZmus/TFZGE/0OehnRlmzf
iPhjdb259neUpfXGSMlvePXPp1NQTSY+k3Gqp+zLfFWXpgytvxskuDnOd9o0VDLlPlHHpWiinGBo
f+oc0ldEVzG0qZz4aCst00nP6FiS0t28Lp4uZPhxGLyQmzuwFEFLX4JtuElZAaxAANyQ+EOsTySx
Vc0PFk9ldk6SbrMmyo6sKw/UdLqbFW+s4SQRbRE7sWY1OPw02YtE3C3QXKzmT39/o4+K6MjcU15y
t6liXmNji0xjWxphGvMQ1zW+kUehexFPK/QliydTEReH6LQ18ddfAquA4SyYxwt/CxvqhzpExq1t
dYo9lNUxxhDVzDAk6uFvyty49LzWCP/PDcevNv2v5UECCR46M2XwLpjS70VfV2h2g+0wEtqaUm+r
G91nB7onfpaz1dBP019lL+fYaIbNbLO9PSm/aS7ehLuIJfwNFdquIdkxlsYhWCKr+LegyToxsYWY
dSbb7SGSdaUrZ7D1ZYCkkYgiaHjBTaaZarif8Ziu49FjefoHMwartcQHypabj0iO7K8XGk7Sanhj
2p0pt39sn+NRbyt78AtqrIRgSeT8qVemzkp8nlBDH6cLXryMee/tIGZaXgWhOm6OnuwyvWtBebia
xEAQVLBT654lt/Dmm5ebds2qaeCyuCsVG0rIzjxjKUq7kvnhffMsWosH/vEx3Y0ClBSIT9yS7s6v
L3lQKOHlXyprmHATJ7/bB1+8iG4Wveakj/cg8ySHFJrcFC4zUsfwOoVbSIQ78gW3U5Ly5TeltDcw
G+L1f+0+i2rrI1t14gPsqEMHHMoy+8PRPHCGtapSyPaBEHKJH3xMoNHFVUZTSKKUd7fYc0R+dk4P
53wKLD/jkgpVvBsbuUWzYtr5QL8HYF+yQ5OpvjOcRwcI031+0VekLYAM+f9YvsPIQI1Gn4OqWcAx
x7DbqYtAsilqzBWipjpRlYvqEef+4a/+rk0D1qY1j2DAufFToia9tDAVOXoak/HQhTIFPbGZi8uv
gnFLGHMH34yfZIKPdnLsVRGApLlnf64oU+JcFcdSt4eqepq+qimhE76PqeP2/dDZPVS2S+C5XFxm
Bbv31YMrYvk9t/Cq9Ucohxidyans/j0XHsuYIDF84eoxV4NR3yeoimw0yH7fU6aYRX6NokLfrb2B
1xX45pcLv1dr55B0FHLG6nqR/MrcK0T6flRSXJw+4y656Iu1+GWDiLwWMke90Vw7AxPYKumXu6uX
OtkZ4p91WzU3rHV2G/huBuIyR+HYtFyK8YWHuFO/4c2j+Pq8LqyYC1D5TMztkcKn2kiil391U0zJ
nnQI6CZ4SBty+eIrGVgSztZsKITPiTdKWM5yfQ/ehJf8S1OQfa3StuN/fwhRb60eDFU5WXAOB2Dx
FbcxVFVEWnDGxdVEwqVWCO9AoheLrV+UicptwGtJ3UpuvnZkx/wcnJ4kOH57/N0zJQ4UlfZTqejq
IpU4Xe4Q7wQiS2YVtE58kS8jLqciv/oJdzUSqU2al2vArbKuwtBRvQ9YG5f8aNbbhswinYTr672z
wYWrU1k1BXyUHNWtNrTKunRR+H0Jt5ITnKVopIaGURHwmE4IuwQRPPolcafriQlVFQE9a1uzFo++
5S/X8wGZUppoWRkHdevxnukpIT0Ajdq4uDjI5F+n5gjumR49NvFZRoUNTqms0bzQfe0Vx61Esn7z
yVPPzmaZiPDsIxl+9eIXzn3tN9j7QdHg3IeOTZa2Ij77lVzHlRLSAEXc9tVibBYYAsav1PlTo6Pj
fisWu3+LDm/1lGSUC9jM4LGOuSFRLHhFAmA1dIgg4cwX4zTjHX7onpw5SAKH4zD0mBpn2AlYgslu
QWDNnKXZvEwdA0E3itTq91OaHRUMKjFuZ0AE+vBi4gpLn+dkfibZdB+sii5xYEhbb/e3fdTn5fz5
GqgUEEdn2M78IZnH7cRSvRfYTDgDUKB4Xr7zdqoq8fYqT/hgUyPJMxuYWNGJwUVJs+GEPzRA4LqG
2bvr3Beoq+xAqvezC62RLLoEc8T1hfoBTTCApKW2ZyEJSvzchllNvbvNCE7io1hldbXJENzAl0zR
RfvA49qFd3HR5XmJvs+EptgFRsmM6qHoVcRV/okVQo7MOH7bEjnZdw5TY7Eik4auFX3cSr7BQln+
/UOZ9T3VSJSoCQaAxJTecLENT9YnSWzj1nJK9inmgvpZd0LnqEUV7LXktJrtdb6joEo38o6hs0bS
kwDUbaCTdPB8C31YWhP8T/FnG8VQTFWSGm1YjDkMnOCFhwLMpBieYlNHnk5fZc0xjfit0vDYgR3+
hTlpWY1kKgg02rrsgNCA0eQQyr0JJzObANo8BrLtOXYdCDDZhmkj0l8b45dOhzp4XT45bpUFA/f6
KKij4f3Sv2cepG2+OSaPs+tZnsr3d9NoUA7I3LPa+PLVmdhnAvopod3qoes8xiyxCx69uSFd3QJA
TfZK/09eFPig1P3+dWiuMwyjMyJhFCVOP5ErxRklSppA+bttcJ1x5iedkdydGNxEpnEIubsoWbLt
MEyEpLB01ppAtzYXGt6z00agmmSVT7IYP20yDRT6sGt4tdS7wIBN6J/P748ADzVgeYPSWZqqDHKv
OQWecqY5qVb5TrbBVDK1WKltf41ksQdEEDE7hlnRB8jp7PNwxmND6or1Wv01YFjmPzNo8DGcTlD9
igG4EyfHBxeqGLfwaw36wPRehNlxkaVSCgXnZJCoAipn+M819Jb4Osvg2qYZQFdRS51s964JtKDo
5Gsy10kAuBMr2kCLdf9RU4cn7c/HGdbzWzigBhtpMehsA98UEJKiZuKrTkL8+sbUj/yqx9z1jISp
AoVSJMbzMETw3rW88l4h+5AQF0t2lSlAooDHLCVAfb33mw3WaKR7zckO/Sx6qOZdGdshRPh9tpZr
0WZWdTwGeC7bD7l7SHARGXYFmZfdi0MyTh9qshGSa2SWkJNy0Jt5vXXW14e19m9Y2VknMbojwvg1
/it7fvRw+Fhi9uXPj7oZ6dExLFpxwYlj4yPWNVHTpq+aH19DMQq6n/xtmVq//K2IGAjAPmsy7s9S
iYyrNZZIec/u5RLCCxN+AvvOt035ZqgvTW9qFxWVsGZoxKrZJ1llr2YUDWKuay3/8m7f6S31Jx5S
9bcrEmUx3LIfZhhCcPkSuIxVF11wHbcm3XA1Iq/UuEuxJFK9VbPz2s28XmullpCDXlVnx69LAQm9
Eg0OqHNs1VAUJLzQ1OkYbVZu7xXVitKDqXc8m1JhWAWep96BhJ3pOz5WEdzRSTTUFGyzUaWV9Q54
mxePWNstroI/U5ouue1cMFOYXq/uMCjqTDa7gorB+TWKRihupKBAGNhAvxdjYJXDxNYytlY9ujxh
Qu6/pFsyq94pIGczIuu8aI6fs0qjteiYs5A3PGneSlBrmDvlBi0r/jB+38DTHXemuBa6yaZrjXUx
h+63irM8y1VdQ+zn02fDpybJcvBbqfPUpe28IIGYqpHAeroD1SHXlXNHtlUi5E2/7YoCenelmjFa
vgF9hshZS+X2jMDCqylO/WDF6YBUM21mDu6V+HRrE4RavP9bs6Eb2BaS4Wpw2G6GIbPNie6xmGuE
NAxXB9WkNU9TZtgJWtUSPhdUtbZO4r4rh3jcNVlFynyzjtgCJ6bIZ4+vSLXFtdcH4dmWHc5raUtw
SoDlXRl13DVd2zXeHXFaj0PWlFmA2NkGJmue2oaEr+JQp3WHKNu1l56/QloOmOkvfPI0kR0lUsqh
L9+N5Ko7cB2LppNViTCr5bAz4zhnKiuxM52JL1TBE+8LEBJfyQ7T5GGg91P4ucYfyJSqqjr7swDa
FNZWRKePYj5S7atKFB9Mr+PM7bOQ697U01Hylwx/7lbzjH6DT/TUAV7hJmMbaMkHXqHaROnfbLZU
gPGDzIb9vX7mbZKbz046+ygL1p9bgCwq8Os4OgfNeUstqjVrlDLYTMT8bfcX2g0XobQUw0pYkzV1
/i34UuXm4Bxl5caIA0WBXqAcI4ah4u9/wkKrPXetkbzwRq9zIMzzjo+5iEp4zjRtguq2wkiM+jG5
JezwOiOndJuw6dCs7VzApV6ciIjUFpBBVRjLhQcMpkQydnh7WXTFCVWy7q23h3cXCD974LN1SybY
ZApRnVJEWH6xHjg0iOXZ11pJ/bBb83KAerhBjI+Jj75Hba8zrj32J5LjjZMRiAFASpS/pUheM+uA
uvTWgRj5XLng/brtPU3V0IB4rJx6kKAEJ0OuDJUIDFjPVHjdKhmActpo6XYajhMTtQyDY0NXUY6D
ZISZABFdh2h3PVv/dVpSM82iOk0sXWFtYsPf43gf2K53IP0+Hi5zK5nkp5PvrpJ13cwCWKqRsnoX
1+JUdKw9vaE9liQuh1vauWa8VLA4seFcICqqQE0qP4f7jZCi6+DjCxPLQScigRiIDDte6IY8D2hV
w5OzyiYI2r/WChNYiiak3ATTnF+3uwEbo/LUCyXFMZq4rIPXnzjPOsxxFVcNDtOfpyEbXl42bI66
S0DGhNa2j0J5iIUsKDUbASQxD8pqOA0cNFmdk0rMMKHFYJMShJgkJdXvksYlkw9cQcq+puMLpHje
CRH8IzXOgHpk7XQF7lVL5oN6Jx6hNMV7wBuImbR6M7H9GXWzYaSBrgDjwmFZi/Cs+UUE3/3/+0xW
1q46/x02eOdOZDALJKqfiV6A6pjFqeZmfG0Nfc0lBaaUYCdf/HrXd72wu+CEXH6hcduPm2ApA90X
eWSv+nHHxfeXBBqcdI94nrJRpgfk1ovgQ2p9fOpZe2LCNsBZjBszmFG13WTAcafO1szw+OCi75WZ
8/T2dcVF8Sf0cES/BMphLfeGTXfavAC0Bk13Iatpw+M436K7DoSB6FHbiUS3uGakGGdyVOO2JZEW
Kg8zFAAGuJcZMWbS/8DJg4fM6eOcFNFukVwyPf2C7s7BLVl7oqHpTxChfuZUsjwfIyXobBrzFQTg
M8K/W6hKbt7T6Jq1jscMXDdYRCugCLOPBh5POW//boO2GIr1b8hWJFSmManBubqjMxtFlRKkHnb3
/RI1T1lTr2TCoc45ZHW3HA530EMbOJWPenM6TWmjWTg8IVwdr3Sc46i6/qLb0+dq7Pakrn5EHo80
fMYM6TfxOsyRDwdrMyR0OllrGx8l3ZkdbaT/gtebVEGgZCjKjK5ERm9g9HEm7r7/WRrR4SvbQtn4
EtbIzyY9CUIIC5zpNQbNIH3pehX3QPHB99WDR78GW5BlP+pcNvLEYJKU8ZCN/uWWrS9TVhORL9TR
2UrxPUBAQAACJTIuzdLP6t+dIdIkCXO77Cz3ZJ3ehPJtstMuoSfQ9REDgpbLjSqTSQ1dIPvH0CDD
b6NDB/qOmMuajP83POx7DurLstbsVFSdC3BlgCK9IGcdO3SpoX6imcADTrBIdYpqFiKUWFRL+prN
pkdiSTVAM+aARMEfBXHIFCNHk33BqzOGO22iixrFjgIxIGkcgf3IoGHBqBmHX5fPHxJPIkKoNSV6
IpxyBeWutGBf8JxyQFivtToNlonjTnVZomrvnqd73dEHRUSyuZnsgPSSIxgHAW8mVtzyrO3KTYDf
1j56P70FOEkWDdB/3w/vtPC31XJc8Xir4uawIyg5oTW/UJR58ZZu+tC9g0YOiYeZshdDJAWFt16I
yT48CmZM0+sf2bzfHnYIzoVaFD7kIOjnLjAydRSyX1UDmgUBZjuB+3KNHr1DTNU17YtaGzMdj6va
Yq84ub5Tsc9CQTmn7LH5X7t4+CT0wJkZv+vtrzGp64HTQW+HD8er4TzfqsUGiZ1sIkzcSKMFMnjB
b6PMY87qEDk8IMvxHfEhr86UhZxC1czGVtSxYtjWCqjV2r7cWiqNsVBAjMZtK7yNWu+ndbt+UOUk
RPmQnZodce2gGiQHBVY8jIsYEITQPnk8zcyJOhtCa4ME7iuWdcK1JUblknd/tC/yJiaFQmixMgRH
ZR35TEZ7iBxSaqRUFIAHpIYKRNPQDnnZHzfsyAvtGUtEMqnimpInqsk8uY98jezYyawon+JJW4AH
5P0TpPKNT8NKs7wGEYG++2c16Igc8iCxqWtz84WK0kygpa8PPhTR9KTmXFQ9ILebOVbMiHXHIQRG
a4P/t+QBJ/udsMVRc0LHyI9qst6ZFyjJD997wH+eYyjW8nsdOlfo80QNocsTpH5G+chcbD5PEfgK
e8GHO4HhW2HlkZEgdT/gbY5cUd6rGu0PyQOlceIwasZxug+Pzm3kkTj/5rm7bzc0Xp0rpFIlk+RD
zCk8DGMnmgiCQMiUi3QdCXPmRcXxTnUnwrchHy2XLlvte21EidAO3B1x4oz78TJ860bNajE8WA3Y
g8JXcPS+vC49qADFU9wUrZSfiGXjA1uNESzaV/awZvVLmGuY8VJiI0z1W0/g2uwGXHJQHJoxTBp4
Kj2aQkvHfilfS5XT1AAuPtehhGhbC/L1hXx+DGZ4hdeCgfuLzHgFUDqS3cRVewVw7QLoyD5EWQa7
Wmenj7F3fSnMhRHX4I8abEJ15nuwA6mYPpqeg1e79y6IGd84SoM4ijLd1VyDIsOjZZ/utClrbabn
yNiIkX3zit28o6g8Vw49NcnPHIKj+bJiNYTZjyEsQ3NGQAsmzHG6Ty2obVxa7GF/lmrhKfidcslo
6JNofrm0Yo6MTW2UVKIPzx/TDiPazlCGnqy4rwgKufEgpjwOTs0XOwPDWnQw2ym9qmNhQjIYylU/
nrFRN0mlXUCmvT25zRdzYgIQGYwufDAm5xZf5uO/3UkZBFoPwoHB71kYreYY1mN1A3ois/nCpCvO
XFQmBDt6nM6J2pRbwet9qLH7PaBDXKe/i76IczGOokMLRk3FfhuCJTsQNgGN1R2wWamgghRK5vyr
1ZfBmgDbN5/mf1Bens3Zd3nzRS+5w7A+MlQ402zMYOx389y/lh+ByvlnbTNG+r/Ck/yVJ0/06DIb
eh9/4yAMbBMm03RyTRqK4SNrwg6AfxkeehOD4sydEKTJ7HZuEzlCxX7r4HTCmnmDMu/QOskFO0LT
DHKUSj71uu0MoLquDpHVxRoA7lqSMUEts0zMptgMIX3mItZ+i9D643BXdI9mP3zXz3rXqOabiUVN
70R99KY9NUzmbFKmr9Mqs0KtCDyclxTicD32Vx2wk5GIUMymePcLYsYHDSHSudgXciLRqXKAayyc
V1kyxS4ruFVv//VWjXEVsg0r9Hz3y6IKTCjF2i77VsYy1zNMlWa8+kn+wF/sIFp6vcQLKYOUpss9
YF9p21U/RuPshOatwWdaF6iMzapmOdiZ67x7ak2HfEKUqn+6PidT/BZz9iY/DytoApDZUUd7USAo
WWiwucsyBeBZVpQ5psYSC2Q6JGbesS9kMUru81vLOjt+r4+2x2MZBrpiG0iELqemUNP7+IeP3Hv1
ma5Ax5UOvWC8N844bX11Jbl0Ys1fc5N/WxKnyQdgLkiFCFanxlf0PvHhXKbqvgm7IPdymxraCWAp
2mEsN+OnduQ/w6Y4VD321j5nGrvi8TA0M7wn5wh4hAf/+LWGuCwy01aw6QoAuJUsPpO8gOyYXXdo
5lQGdMWb2YHHGHvlKVOD2bCA+quwGCmwfa6d+QJNDQPU2qP4WMiu211orOYgRK2z+r6Vs9oCSXL4
lR19kK3TaHQTZpZkpMT6tXa5x2WmzjMZKrgBKSwqd0V6a3ojoMbDrWEIU8LrIHaoik/zmeKwiRGG
njNkNNv2aQJO6ZzgHztzhKpueiGtcYjrFoS9XfrnRxq1Uw+Xt1Lcyu5ghtwqxKJhCp8oDMLf4plL
WT1Qu4si+9yP4tVpL9yFG++xL1y+j6moN77sK0IHhArFrpkg4FHxBYjFQvbiN/Rtq09yfG12+dmn
fDcmtIk/Efwa3Q2SEu97lps4/yNZe24b7pphrrpzEp7tqWp5R0JFSnJu1cKWqQuxuoq9KvHYdP9q
p7BznRg8lo/Pz7JnpWuKSruiRjcKPR++HlqtDEWK82AB2Q1KqbGqmtiuxBDyrxxLOhoTSYZQaTGt
owns1RSAyGbzouib3V9+XPN3J28bQ53qeQm/qL0nt48yobK40Ef5ZnmF9Ox3TL2XDJA1xXMqLyzL
0YMfl77+BMJy1czVKoHDvsQPbAMdyxOvRSXPwcg/3SRhwQbmPmRVUEdibAmpondJffp6v+8Wiua8
7dOIjhqcSLAz+Lr/eC9ryS1HfS0XK7ax97uNKsljHv5xe9MOCZFHEAm01SwNWUCIryVfD3PGSf+8
ImbLZ3RTE3GecKdN1JyhGZKDjJ9HQ78gYxJcY0pwSqujci4AyVMal7cqanP9Z0JJ+nvT8vWbW7Vy
Lfr7llGpKMFWuI2T0nClJFKWhfJBzryAB1XyMJutK9U2PzqUwR3nqXASzJ2yDkXsVceCJcT3ROpS
gQN9IAucsbeDvqVCZ8nLllw7J6KU6Q1r93as73bMy9MYyRkFSsOfYWW6FGHUWA/v7Nu+BWrd//jD
VDC3PtGNJoqBJJLCut+fAgwA5mNrlL5T+EmsOvsdtQMJksFg8qYkaLecvm1Xj1waeAb4KQbsDfuN
HipgnLrlviFBuMkGyI6bkcrPx0esG1GJT37RCsYTvPuHJTudzvCoTQEb3+4Z59G8G7ALb25L/jEM
519RINjQAGymQ8Sw4CpID0WcoRFRnE2LddUwavGfsHoc4vGRcIiIpRxQbV53yxQfc/JVhJ4kl3Pv
O0S7TK8RpPhnwNBBKh0R4xzz2GVY1Gnua2Iw9Vz0Z47LPZn+aKlMbkAUvNOdxVlfgq/LabLtPALr
Es79N6FZUMTxGUMbHEi8SwPIcGhFitB4trtLmP8/t0U9sZkVZnYSAnNgMa/lz8nvpi/W7UZH0dgj
hlp4SQ+fT8jqoPPpGewOxGW3JgM2lpqHOlHgyGE8ULYLvSMerXdN2oVGPifKCXbyridVHZ/5rHNO
JF0ee4aexgCzSHjJ+N0w+KGxZ6n/c0y6EcEMeVZSC8Hyh6MLxuFmVDgN4Z+OKo9yaBsEhCV73xAw
YDW2AwSkPOdR2to+wQloC0dSr539Eec8V71TzaW+RhE6G8ZLLs6sZl1cZnvhz8I2uDgLl92hOz8J
CJ+vGucmAUx+yXz2zpkLswlEQldgbypvZYCddcxKlSPhACc+QN6LPgbIHKakQi7dcq5sV3HYLX+i
uJTbqc70j4/8b1JgNTeZ0UJIJKWnvzq7uJFPNI+zZxuAR+lz4sL0+vqLZo6rjbO8jInvbaDQ4rtG
d2CKaTT2lEemD1lepyXKmrKHt/OuX7kBD0xp4pO6W9yZDmcPrR6yeNa7cIjjY5W23OrFprBtkp1t
xw5SgozS+A9PrrZeveMtML5wReUNbM2K892He7MpIEYuWzJhv7T/v9BmLc0z/HbiMDBLlc5FrRPL
NNUDN1DJZBTskIf7n+oLxM/V0m42UTfM/vGmrdHXrV/SIdcbhxRJfJttmkhoRb1ksEDnJSqLsW+n
HT4THhb2gieaz1NYn1EGpPY0Bp249Se/bX1QhP9f1f0aRSwZG0Hf04G9cBiBmf4Jy37KtkvX8r3M
phuOfxQAjNLzUkR8QtsjLfofkXn/bUuybNTfXvGSNcGcf4sdg4hRzq5MnNYLRD4ub/S7T30HcXO/
F4uTGE2gOj1C6RBO7H0OuBPcCs4RB8DCAeawCN1wnImRZN2+so1bN+dtEV8xW2UhprKIxMuNbSOh
mCThC91kQRmPFYsZNrZBT6WkVJV7ovPAeewP5QCBH+/WDh6uE6VIOxHvff37ghX0GN88qDe6UptH
3NyI23YJ5274Q21DwF88vVFC9oV5kP/wrheGgyySVK5J79xgKRV2buMAiODf8esSK2vP0XvazlXz
Pxdi+dWdZG5o1n1+JiUtanYYnXf8B+6knsqGyeQkHG9cyl2qvSVwHfODdwIuy07ciu4eJ33h4XV7
2HQoFVFQ9c18seK0op/0fV9MLIbl6vUOWywkofkaw7HhvDh7GHqYbi3p0UhAClElZuiJCuH5MW09
Ayz2JnSkv+pB9aLRh1ylKNsDUMrXUG77SLPFyvj6aoBssWmxKDJA+47yGLoe58+k6+mtIpv3y/hW
bAzgzMMf8yzgofz1loR6BzcAWtfbRfkvzQbxe8xfwPCNVtBNnV6YpbWNviKGNRKvkV6j/maZTYXm
aWEsZQyVoyrBracdwUOv/83OOnH14SZfzBJs3hkS0LPTJ9Bky0LENn/RkQtlKTtxx/LAVsOscgos
6/MU5hT79jR8S7MORsQ7tm28t3r2aPt5hsCF5/yp2N82oSKgJuXUGulgDeoAaWH8XhR/QcCDYZaQ
+42Zw/BpCTY4JNAmNxyXdNQHqBJwx/kRhdemdEv7dKAvB43DPJeVi8uSywfV6J5k2+tjl5nnXskX
9YLmQMJiv3mViZ/IrR2bCWt3eWze7aEhYzfuf7T+tHxfxiouf3JRmZdFV0msH6rN1tziuP4DPJrH
/Rg8xVxF9cYjt6eQlZe3Qdu0Wh5eh0DN57A+OBkPzotD499lxMGxNu2AAMeuQBRhzNOUf7IuRKCx
b8iAUm8PWAVroDdlRF9BrCS/eBZ4g/HAL8cUgIVETLuLV+SFLQT31W+BiCNBpSpqOB0XzdayD9ax
6v/h2IJQht2Qrb3uwnOCvuxXLLPC4lbac6hLorX0mr5P0M2rByUFNCgNwLdfVuu9mEX+7X8evcS9
Ub2NYcYGKxPbrCKet2arz2pz5xW6RpAatmrErIoEZbQ/q1OGNDyuYrQPHAXdzHC/u72cxznmxOEm
NNqLhOe2TVGT9e88qd/lamASHW20CdCYP8+1YkN6zhvh+2L5Jl4FhVdTAWqk7fCg+fZhHGEFIdg5
ZTRSyhOBPpVLEgvuZ8iv9IACZY3l8qjmVdXqRlXOCMbRFRI5pIawWbOtJ17u4cUGChpzVcNHR5bG
iYiPvV+biUF+g1Rn4J0qw7sLlXUqmDZW3ILqTtYycBGl3o3n59N9FRlO5c/kaR8Z9sOxbrwpZJAG
rsEV4fCMPgvLoU2YQJbjrs90yol0nFjdFpLdIOz3fmxUbmtFFVLv9/l/y3P1sqdv7DwVi2t2lTWV
oLfF7XWn4XEgNgcsDnEnyu6JErln39vhJYfwQaOuE7RwVf2zD8shiZ2EJIaPn8OzN52OVh0QnMoD
2tcxSu0Zr+KziG0/w/w3DDA05dxrnfwXBWEbbrIt73uzuY7QZwzbjq0RGXhViuE/UvotsGo+D99t
e1ziMUsUxPHAWx29rTtbFyAq+ccimX3Z8BjbCelZaY/Vz+BDXbYLGxmyY1qSr9mSqpE20VCTkbEa
AnOLA0WFGG20cC6cwBX2M1YDiZawcCfi6nE6P4qQYWhYf9rUX2T2eQ21um48i5geHi5dthSTW3t0
CHN9FcFtBdVMP8EnVueY5gtU3hqpuF70SpDWCg1rnYj9hmnTXQGptb/ZEKirkgcU3Bqf9VHA1/aR
++pM/foUxf3O7cZmq4xNULGFSQ06T+s7W4xwsPH/MyO4/xFDJTxP4oIc1hNuXkyIJW2v+ab5ufDB
gXwIDP6hDS/aiQ38IXQ/MwLTYsKHPZRweFRifyzK64DJbK1cgH2bIwWkD/kZZ82UwdbBWzMURuXN
EC77/yW2HBeSYytzfvkUWhjJBe7/ZEAywBe5DCH5sO2/SyMjY0CwhEx9oRNiwLvafm03X6PQy2XN
7zep7GIAvSR9xJ4tzos8PSg5K281tyrV2Rit4stsMzXGZvuRaMq2G+lJxbU+tMHP6uBaeyjuKWS2
/4kn4cXGfPmhAdg4rVlkBwJgPWawlCaJW/BIWQsdPbOrwNM9T2OnH6UJ0zBSF/9i/YsRGz26VySr
23yGcDHLCozCSQZbK2svGfXStDCELJbS00Kkh/8Qa6gSRos4jgvod7g9acfuaNTyTOpM4czzUeKo
7D5Q6qsN27eFw3xKUdowsJ0TYppLVubzw+km8ZUEWwtr6ojz4Ki5NNNWrNzL2bT8336/g1LcGSFN
e/kQi/BgQEOB++lFDd/Ht110ufS+RXo2xQgIK0BXXBQm+cWOZcfpRlM08vq3i9Z1GN2GoLg7ss5M
PGZS9aGvck/gw2hpAQ34meXMMa99gnkjKjJ0GjRaVlDvcKGsntLQh/6e3SQJJRc/UKgPsHfWqWVY
1090BrOsWTh9VpzqhtlDHnf6GurpxrI7uaG63XRIY/2SqZ5h/ptOQxLKLzAMjFXc/JuMxfuNGZ3r
yBLHnz3meEjPJE09C45Zig7/aNe389IGvvn4R4sX7Cw8rX6iaTr4oBJ17E5nZq5hoaqOWj7PtIlH
2X3pbRV1CsoguB1ttK1i16kiTEImyVd2b+LvJOa/oTu3AHnFVwFsb/89r3CSJ1gOP+06JO7ASi10
+WtepvWkg0vejwIyxhKgsJIFRAcYr+b7HvrhAYdQ0xnYFTMVtvoaRm1xrXZrVHu/QJy6CtCOI3EP
6fPFNrDIa3qgq0uhFtshGVZnsdu22OcEw1GsdmwLm3/nqVxTaabJaM0E4EK0dOSWbgl4N2qVFJb6
MYqiri0l99qa6r5DdUE82cjYyjx0TZJicv92eUej4IPQQLZKGhbux4+olFXWRYbacW3D16XriT60
2mXDdBQ7ALZAdc7in/DrcU623cyv/7y5fXyC8faWNC4aeMskiQNMa9FWYHCgRmMm/XP0UnnqwrAb
TX+qJhw62dRd3Qn5c3UaAVi+DFwzgyY24pph7xii4OR6vE2+ZJxrQTWrOPCZasyfF4Mrp/DNXLXe
AWiO7cOn3SOh5iunp+0MtQ3NjfYfrqqnsapbjtdyNvJ6KSDJ4v748SoVP1KYIdacLuW1sgPDLqrk
AfaMu/hyrUWHgIG7KEBr4GJGqHIeRzhE/rPLAUxupaUXWHMkqVnDLN9LlFFlZvPpNKbheUwQWP5u
dyhZWe4U5PjHTEp+i1p/qBayVZhUWEHRKCGzedpppsubJFZi2JVoUsNCrNNaOqXA0FhcHOnG/SwK
l8fJl73J35bQjZ1qYkB1bgAZeSX2tOQMaIEC3AeU7w3vHCzXLKoYe/987D90gVKO/9Odwjru7Zik
NfsH94yTnPCVdz77bSBRN77K/HlT5xfKks0zfllPx3NfxUgZOGOxJ6Grhw92/qpP9u0mg/L9qGYB
Vg1SEnhsdSl4DlfLQFGUNKiVOAM66Y0GBfKHDD3uGHjtkUAvNbgoaT5Cg2sCkrU6fJmURlqk0ueo
40n1QMACYixGtg3VOCDAToToGvWVcl8AMht7f9aUg4Dkih/CTO5xqDLzM0WtsDThwjN9yBYizG1/
GDI1RUzfKxEgmNIr+vfadY/1qBzuKst4hD1eWcmOWwN6u9q/n+9xIeW517HyLKImH/eSxlewvjIG
kDxxCQ33jJ6vL7jkUoTwWJ1mUbVMhGTRBfPuneEfxbikEn+5dI1ceqt5pwsf77FrZxi/JZCIgKNR
kLXUzSjTZtppE3zFoofYU78z4evJwbGsxceJHRLMvvkNd0rl6801HVa75mSDL32Qtn0viDvzuscO
WIjZBcXkNPBTUhkZJ3fqaMbZBJmfoJeRCz/UIB4GK45P+OvJZYLq9gWYqmxfpfxbzEeXdbznnsNp
9hP9qttq5mLVShRL0zi28yn631lb4k5KJKV2PuwCEiOSDqJRDRZjHZKkKFP0cxvVKkb3saPNLov9
PTtdKwrdvUXGSFRbLhh1MtlQmNDkz1OoZC8Vs9sa0da2U++BLygBFW5ZHEsq41jbE9zijniV3mTQ
yxJ28r/j3B35CQgRVZ+2QqjK05zo8snvDHQqV6x1NtQd9xe2RMrk6I4alq/qocBGNH+yTWPJak2m
LRZpLUTFwlWRkccAbC+EoAlno75SCPQnBkuNS/a4EFFd9PpLo1gkpV5JjByrSnfje28qOWQ7X4HB
sFQWumh8KhnAw4EwUw3VISEvCINRlNfllBPC4h35zGbje4Q/n77qsBTlEmZ5Q2VEzZdpZ1wegHBz
Uv7M8z2bM4hYz2CubPp5RhlNrDYTilSOxJ91dUNImaqsuSdrM0W26W1n8CqbMds+5JMEzbpkzlQc
m9agmLpf1GWWrjIjgp45KKfomJSXa3FcXQI2+OjWhS3MMqkwUcTdW3Q1oYFBxNS+ofbkG5GlfNIn
bPR3p110VQubfOvb70m2LkWnDZyEkmhEFytpspzA8Tzk4xpth4VBTS3RnHe5MZssFPJgArx0zZot
gl+euBA8sQzHwKqcGyh8mS3wUYNf8gYMPn9+52dGYFIIVCbuN5tu88PdeYttPnUM6gBn5RJShJhS
7XF7tnoabm0e6W/9fkEdT82JJmuB5vbMlUR88aoSR4F2sfZAoxncCvbZ7wSyc8ErWX8dRN8PC7Zu
gF0bY9Q0UfLzTP23XP9/+OLX7t4T9hFBWxCjHXlWb89aT9qQf6BbkH1xNsxg1DZuye0lk1VuSwDV
TvdIDaRqJGCN7GZ9EIOmwgDhUcqIulTGmTzfDAXt5sduh+iqXlL9F0MnlY9OGKwmOzxu1MBiuNFb
GWbem8ekIeG+Bh4FSCjJsiHcMYJouOKM5ECFtGMXfoQS9b6LNsuJiuM6MHwMgBs4Q+bdrP4PvYpo
F5gNfq9ceq83zt4t+C3dmI8EloJKN00aGiIfhhkl3gbOlyp4qSTIvRnauaSWKmLkYlRTcKeK+UrE
+A5GX4rtpXeeyDxd82xzelBbO33dh74DvHmzZRv9aDBwQ5m4BP80/npHU5alucr3ZSdzWdYhS9mb
PeV3E/2PyL2AJDIuShp06QoeIQ8Rba+5+lo8UYE7eFleYnQI+xVO5X4pN45dvfIVrl1PnmmMhrjz
wU3vHNWm07IM7jwBpxbUuxfY6Do81ippVjJ3XeT5YGKe+XPYGYH4TvcuAC9HB06Zg0nrKmzh5Zyy
8P30Ljd6uT3mjwdVNOt6WOQCwfs88BJ4EgGBpBVzyKZjMWDnB1b0j9uDNCxNtFGw25pfQ8A0VAiL
aR5I9rcGDUVlcOJQEJ6JaE5OJyZcuWl1yuQ63Ju5ySz4I0Pw24OZSqCG4BAklxULvo8nmsixWd1p
2isdQ2OM+r1zgDv0geX71NM84VrXjJKaX5tiU9BR7PLsUAqwV5mDIdrIeSj/d/NHXLFjWVI+cUkD
Uy4xnBQ1DmipfFpd1tl47v2XHhMZTxwnRsxpPmNlxswDwObta6DFopl8zVLcDIAAQQPlmgG0p3fK
N/gRrOXaMt+RW7/Q0wu0SKVKfus/1ulhISjOYWvAI2aFxGhnz8TdE7xGJ5NrSy+Il4WCiCz+BjLj
l2deWhf16OWavHol+83tLYfPxuNLh6N/FFhQcLkgrAiSIfAqULxlOrr/wIs98jY15UBRmTcXnLB5
U8IWWOtNgt9Uqxxb0r7TZI2d+iZI4AOrHSsfb6BLZYQW/0pScZgwbGhkYXyEVbx+mX/GfB4OJ2Uu
eIH+CZCv2ioc14HcoFmEie5uUZfWdfCQsxERRunxL0QKM/JggURowVFOeaQq3jYk52nG1BJZ7uBU
tL831ImGazW2uKwvKVHBtbOwg/7mmIVVAgKlc9JR2rie7BdCVhrhIxsdhe+3wZ7pkv1Hh7xQTH8w
RPPogwQi+OE16d7HWe4Ug8iAcFUvPmf4EsALQA4P8NWHI1FnhbSn+BuUUkZf+Co7NMLSeNovJLYt
MRdGOX/QIGjywznedEo9gYGU62hNuONJcmPxCEvH1Ij6MVM1mOputDY5NZoaaJ1xstvh0lOcDAum
Nmcwk233j4Eo2ft05Xn0462WriJKfldjUk59bmZ6/YBqHdYVst0X7ildtvKgwL4DDPN2Z7BTV1FF
XJs4i3vaDby0temEfexrdo/2T49djB3+uTAS0cm1rKMmd77Q9JtrHiWjbaRp5tytJbSwzbsCve/j
QcDdY7K+7+OArupchd2MUnFzhWdKnAswIM5lU5LbfpqVVo6o2ey3Ryf2QwYDxeGTx2LeJvEHOadG
6wuuYsrwj7wkOBQ2ONcRmmLjgGh6vWXSWV13iagfhENen4CLX5W/8f0gGlqUkV2vVWaX8SqwJzWh
hsu10Y6tSnbGHCozQPHFAbnhm5bM4n18aXfBWjTU/oor1mO0XgfBjlsBmG9APEpOwVgOrFiLOQe9
7Dow9i1d+Z+hXGprofdatd6cwKWS4xn18UcjNRkPUH7jj/s7x2/rrSV5khHbnv60f3a0Km0r41rJ
cCzrQX8HGOFw3R/iBDivioxHR+3vjan6PffBD3qhILwp3MrwVUxj7FCQClP8cJc/W+mVogGZnqfi
A4DgRqwGWVDCf0c13843YFgQCierySXnVtgYHl12ZT35a74fXMt9QZs7f1GRJYoB1gYhRDrPF2xr
HI8ouyH/mn3ipfqRN0xUZ9V99OqwfPp9iSbZyNOY4gucEn++vFFs4nJviJ2GpqZQyj/2vXkBWr6X
OocTvSUxZ+QRZkhE/y16SxmqBOFnhL5rrWidUJiPgTRfthhTqo2zL7S33itmiSFTZHKhkTpEHh02
ufl33u0PK8Bw23Aq+wYxnFY+0Ulj9srRp7CNdohWx4BSrDYcEeucUL+A63JeaD7Q3ed0vGSDMxYs
dk6tgH3jDEh42e6yCFk5ax/JBhwX2r68dKeJMaaM65qKWFum0WCPkWf35y0F/fQz1iDiLQcAgMsE
eDshrAbkkiUXlpgvkwnVgfhAQFEaFIDyC8qOhDe8U/VjwuP8L8P2c0bO39rxjQ4q8F1QNR0rTNaf
nS4UaIQMUk00AjhJ+dKmjXhPowHOsWs8QoT/1NPNTgmoXccWcfgO4OcC6d1jR4RNjOu63kNjiAfQ
kYGCVijjNoNMNZVCFpXQOSXyMSr0rw4GMahWrMpiLSrhjg+Tn5o+Ov2I1p9JsK/yj8RYENafTmgx
U68q31vmSWXumekT0tVTEgYQ6O97wEcHAPArcymXMti5dzZVyU5f8ejJhGFLUkzh3G8wyK/SFZCQ
eBRxG6d/wzTnqJd8cmnlJgLZk45lLIa//CPPXSl8C7B9kTB9T5eoGpBhV6kecg7EIJlReU3SAL0c
qv4i5wmGz8fbGRqqH3emSiW6xz7uUrnWoyLR+K4benEkLGkb2F2Xt+eo5+ZOpwqudaq5xkb2i1YM
ehKkPJbkG6cCl902Y9r1qVUl0sRkKtOPKYPVVMmKYsd4o6BgDNsb2kAozw3PRt23C4RPtRdNALyx
VXyWA7t7ouE3+65PmKYJtOsoakG8EuzKPc7eO9EgbFX0CmWn9I/L5pRVgwyK2xYDUA8AIOu5TXw6
N7+Bam9q74j1a4aVSltSL8ihvasHPgg1sSzUoberwyglNdlKRLZQv07O2cgIKKnLOKnCDNE/z4Ef
HXtzgToeB1KV/eCLlL9jBWoeHF+ND4r97t2Jqjn2Y+7VpS+mzff0rvWpbewl2Z/uHcANExfL8yL7
E4AhTVEFxNKqqvsWNovs0WxaRuJRi2Rbk1bW7HcMbJSn+IgX9mvf/01rFhd0y2W0tdZoPdEh9K23
XrAX7Z3mBTMzgo4q/jMUWzp/tvdGuZVetJA4FWnN9Q5XPtfR2pM7j8Dy9XrOOa+q52lASvTiR3xh
tl15B3QSPnWkXnXPglmCDhlv8fg1atvbvCxvhZ5eFXG/MYxGCLQvjhr1juAm05C+/SlFhAgYXgZp
UqvqIHSeRwzdS7OexE25+qb4pcrt4FPSqwE/6+x8S2myP9Xg/DIr7hWdouU3N3dB2+62I83PiV8d
jYsBQYTC+LyiccR13iJ93UMugny+BHIf4Jx7EH1pnbBXk0YC0TC45z8VI0usYDuo6Qis0exSkLR+
iDZx7OcUt1U25aLDi09u3uVn8j4kuGVMStt72pH1prQqFUuZT2P/FUcLh9i3KKVFwTSEoPEY7Jt3
FTPkPuJC8lcZoJcve0jecmw1DY936wfMXPHuFGYHezq/3sI8ftijn+/bUTzumr/iE2kXiKSQdFHT
OdchFWkfLi9e7um00LNRK/WQzVU+G59Zxah8ugXFbew0jPyRFrKL7oYsR7cyDHodk7rcwgLthy0j
9LPB+YwbZNfefTqaQadDtJXwmpG2l2+KMn0rm9msvj7JacTzkrJ5whzmmfgSNAGUjlZWrVcksfmt
VXyDQMKrbc3WHJr0SCsWaIKHmJmMsKMJvdNDwa+Y7vWFj1UzisSbYKmGWA5LJVWc8MJfPCJkv4zt
Tkg/x47myt4FUxqpk7zQtWMPpN4beZkqLnFj5i0V+koKORHbav6ck8dpXIy0WYysYFA8ZaANLMnT
WoKRRMnFLT5kywBDrESIIDz4YRftbHIwymVT0sRpoOqUmXAiRDAdJ3D9moTls+iiwwDKpbSStHlC
R2yM/ACEoEzHxOoR93DQRiNxNjGwjIKz2wCAysonZVsEozBvaXFl+Uf9P+aDe0KLGVk5PptehlON
u/R7PiBb9poD80emBNPAvIsTT5frjOkSE9u5A8QlDUqMaBcaJRNHid5jUtQpDZ3hR+FllJLstOc6
UuuO6ea9n29GzxzJqCEUsNeqNi/8LqmSEB2JpPgVWw8m/S1cQoNJ0uYbU2P1QU1ulyVH6FZ4xpnK
3rRD16y6l7y3MwHRTOqqQjfTx9WTNJNVrA6B+ajlhs7OfoW/cE74GG4THhzAzmPdzTb7lw/kns8X
bU5S07fsSJTt4aRUzWnaw77srCjBmsc5PLBRaQZUpBC7ZeET/sNHdvLTDsX34p/gEKTqPFINJQz+
fvERbKHC/zDn3biOKFWu4GpHbnCYCTfTiDjDhBPet5crXazAiEjAhBUVUAHC9WBJx7Pbp84OlQpM
/YEgVqpzZ38Sw/JQNAdUf2XjO4n8iQ0N5uwuY4R7Pgz4eSr5PGhjV+QVVi9BCU7Kb/vPfYfYKm4K
8Cwz6DN4sGkoPNRSl/Csm6TgTTrfvAE0y1kLbqZWaUbH521vJIZqCe2O77PBUtzUlspoNLiOvmAV
vQ/6kbXOCqyjOc7AdCVWvjYWL4YyrPphblSzIb/ILvH9zK13vlWqjZAfQozBJ1LjXSJc/HeaHkWU
eKfuWlOvhePZUUcv3Giz/1mM+JZCEStAsWfGTqgqjzX3Xlq0xW4kDXeXX2iaaU8JHXXXIhFJef5C
IGiX4Psee/teYOz/nFv5G0rZesAD5sfepHWtCwAqoP6MdbplZv57mKlfQGXwSAqj1ipTRjpXeUnL
a8mxJAQpwFaEFwxm4hYVlqvT3bGW+VQ/HhLTqtJLsN9/GkYMSjOz1FUGtrs4SCwzfWFJL6gZGHMN
2si8uWMjW4nt+yLgvQ8e1yBkKhAeLi2UPUns/OB6w0izlOfZer8CPU8JBIOgttjBW5Cy6MNFQOtk
h4QlOUKTKST8SpQcF5RzG5OIbJ5JP37xT0nPdsmkHZCp06Coz/tfaHVmJq2s9+cwoXAnWVMGiUG1
2bus7mc/5DJ6oyfk44UkoTW6UtVO6Zvs9qBxZFoDjTfhTzMzWGN6AIOILmeEWHCYhLfgbawONAip
TEkpP1cTKGHe4pOn6gBfAn+0mYCsw+cKWvzdjgqNnAyh/zdo6Ka139NCuszkoY+BYggVF9uT104H
zaDI9sBo0Sy3Z4g/iwlDFqDNWMUzY1urfzYRcMk5VnM0Blgg1Mf5fXwmrch0BItdy4H+lXK5nezU
qIfOH2Yr+WOUFqEuUke6eTMSrzJEJkplmPk06IU6U+tbOchBN2M0eyCEnZfzJaCtoYjrC+TbT3nj
LL3CqcgEb5CG9Swi52ks6HLDY+H5kmr7ani3goGGUUmMxHZdQe0liBqn5uu9YQ4f1pGklQ3lBdrd
ZqO50CBSeujm8V6URLV4EfEXYoyAz7mQ/2Av1aIBC/hVzWn59o+05ZWB2f7LsrZSDDmLk3/rxYXl
vZd79rZCRj7cecyQtZsXeIFI1UVMSZuT/b35USN9EkCafRhJKHf5LgsW/M4fuLAQ9rNZW4XlGUWK
RQsu+QUbJxfQDvmUBbY/g8H1dacVo3IVuzvI7JX3GP/6MkIBovcD3+WEpnevJR9pI0eYnHHIIRLy
yBLdnddMmCj3Mb2xA46ovPYIFK2oK/TxkhcF93aMh4Z+xOal4J76GcPjw6hRA6pSWVo58Ekgu4yh
/FLM/rseKFMfZbM6ztLmT24Ok6K/N2pb2l1A+nNVengjn7PLwnZ2S42f/3npf04/7iUGi1tLfhAN
eVfwUIycPMVQ64aePpc6BVL340t7n8CBJx/avt3rzo4QhTgwZPqkcE9G84kTpu6hsDWethrP6n9h
kj7Ji8/S47Tl21FnIon+14X9ZOdCaxsNXm6ZnnuMv0nwkjEEOmyuGu9drqT5BFllPNvb3GOx5eUI
JQ9msV23Pt4GFLy1wy111JkIgqvRtnfvWrHpMlYBP5Kx5/2ZP2BUUFMUpl67LvGd8K9tqKpj/fKc
oosaxJHfC3pxXoblfMOKT3cWQHuUiJH5WEGGpBgXt8jdMkiaekgUvTwSUwYX9+00/in9V/WXKJqY
aGUugWqen5cbcNeOWMXYAhsbkIbZi5Fl8goCSrzDfTpYBiytofYdCPQc3v/quFof8prAZlvV6C4l
SC2axCp1UqJP7Se7FYkXUQl/06WQTk6gZ92suAUVaiXFglWG77CenCZp77KIV4FbN+rq0Yerggjv
1ZBwQMN4kk1LDhtV0yzkT9M1ccHbMjptWvEG/NFJSsZgiKrEbcYCaPKBhBnZYgA2S3vofBuvsv/x
MF4tWxC3Hl9WJdaIyJvoMYN6rjxju+c/cBuIkAH99ggFKU4gZa+TZp4D7KXNxHlUqF8WMoG8BAOW
pdvUGIRULsacNFyD3/WBgUt6hpQbYfhY+j3YIIWgCsF75azY/dnnN/PFdJJTqITleo5sylsL5J+3
1bHMHaKT8ooReZJfkL3Ee/+msaxPJhujufN3R6GM9Q4ZUApJGbWAy/Go5peBxad5R38Sqpom53Sv
0RVDaRjOgka9vsv/cF2eNm3d/h9dpoDwKBxU/1kERcqBHQsuLuZQK3ur1qwK1rQjlWj4qouKAhSJ
6q/ZqCVNjhV5tfZjM34K1n9AtnE+9bUiVui/erpDom2ISqSvv5NZWz8Uq5HdjONLpHSZv6JyUGGw
xSLw3w+sRtbx4Oqs9AUjFMrITuZoleVEO1BJoF0MyuAvy8sHE6uffFZfKZdT56fljcO2fMU2A8U7
YDzcBQLdL2+v0tY2SIPH3tekOZ5EjCc0V9hzDZYrnySYfOgaTZUFB0oHZcfOQRUNIgx8fao4JWD1
DOpA39l3qwMty+gr+F2xoJ1ECyayJEWIp3Viu+MxSCQ6VbX1BlmQJeKdzcFrUOqYcT3D5u/Ya0Xz
9lxRsEGwmj9DknZL0X+DlpRk/G3X1af925KLvKmlty7/K/p8GH4Pc6M7Lk/efvhf1JJwlhVNe/kc
J9bCyca9hQZLV7M2MjcbpkRyo4FhADRgMaupeomdGHEjng8E0g8ZEGImFM7KUDn2DVFKxPyaZmvj
fSkJ1ePcdqXwQzTc5vLjqvDcvKZ73zpIfGW7H08W1hAGTI057x7EWOliZLhzrTbvrn0oV6j0Kt5U
IBCSGkL6H/V5ukXSkR04bJLyiOEBT7J4n8xbp96TbVUXoKpuc7EC1Ph2nC7u+T9AluHsQvORqaSk
a6MAjHOa0h43ruag2FmLsVLCoWNUcKocbSmaU/whsr8vLort6OAK5MStHy1/y6g5bzwPUN4J9L28
Fun5k6zHpquzN10/NUp4cT/0soYkn5lAiemtKfgi7xNHgmJoIiRf/azD59wxNJv9+y6nfYimXMKh
Zw5bdncA7qu/tuaqxq4Xx7hd78sJbznaLb4OPXEE/S7k7Ac9pkSbq/0c/lvtU2IenD/EBELu9L3m
a8r43ff3sH2d2/P620bLjldUBD2Rz3lJb/rIacEMIdARls5f4wC+v53xz6c1jylsL/H4V7y7XlBi
pUPwB/WuGERvCXU9/fKMTi3+3lR3m100hTFwJa4iqBaUVUdKOEJe5gaJlqiegVB7fgPE8FTDfCzr
l5udhALs30dlxpDV8gYR7a4gUB2OmJvj8Escm6x0KkieR8fErCgCO6Q2nPqfErdGh04jgeCeOUnY
1DcLKk1+q8BEZs3UBM6oMmQR2JcRyzECj+xkSgQUIRJxOu4fKHfPJpJBiVg5GkUJZf2U1z2Ys6gQ
mC8DqNKYY1lIcUeKhemFy4vq3+2/EyMuYLYiqeJLWqOOa+SAK0F9t9xBPFLalIRtYkZcIDtC1XF9
/dSButuFn+iYAtUJtirq08h+4u4CHLY1q7XWAhl8sJI1gTN6FKHkwkaS1gAx2caSw7DUwemM5hhj
kIhih6J9G6NhnIdjx6Ot/C8U1T0NuWxQyanMGDWXRAaVXfHeu4Uft59yaeTcEoyXNUKE4H6M8UZX
uQQU2cNVNfWRijdB+i65cwOwUuFjQS2dkkxprdh+obH6lgkinujFJc+M227eQjxc8ZojPLcOdrX3
/Hlq7HtR40q6J2BhdWXh0hDxY709LXpd7mKU7FHysZL2N3/lP5/HmeF+JLc4QunoRJup/bLWavbZ
C2MH8vvI/RIcGjktONCJ/I3rqeC43FAoTNR/BpQlCWrbtM/vas4V928zxWvcr7ujn+/vBJ1DCdhd
SE6MawekxWd1VAku+KpftkJv7YtweVGLrQVq5uDBygVLIE0G7/2m73OWoMPU00JZbCG/0Zik99nO
o8RIhlykTskxc6avSBbPOs3k2gUCRvFEVEhoDdWU811J6wC/I4GZ06ZWIwGGQvMtg4jTuIpbY1m7
ia+7bjZtbPVBcKUpxWlzRL6FjSGy3PLmB73ThGOhZMolSH09ldtiUsrKtQnc8SiJ2kipxKG6iHjE
O1290FIcaGIIjRfOBmmEoqaQHMFLvDox5nugGgX4tpox6z2g28c0Upq/Hby3CYfktDuAobXUrca+
YHmY8EnIbbNAUOYOO/bk6v7UD5GGVU7QeQEo19SSsoiFoB7YjnSMCLdJEsRpgTQQGAzSAJAw1c0E
mbniFt66Aj0rbCen2YHpruC2dnn42K6aPG4OBFL+3+UJv9j5O4a/TplYBOnT2gVBFj42TYcbrvHj
s8vGPuvjDqGNG//laXWxfzobmXNrVYt4dlNbLMb52jIj0YjLK6S97gbTvNFYv51GwABL1vHsHQFA
2+FylpV6alOtbmdnemXuTgStIB0VSFswbH+tpkHoiV37p+82/sF6N6/bZt23dkLJkL8bhPhw1MK9
O6db76zzLK6OQiMURVcqUc3U7B1VQo6WY/RbotSB7zhAqME3+AW6HsaCcj9WsDvMUPFk6HPqaR/Z
MNpO3RlwwopEsQywKxCsbP45FoV8bYBwBwOFK2AgQKNGRGvlEroYLyNfMNVbvJxnDMOn+v/jamNu
YOieBNGblGAChoIGvU1X1SBVmWukP+OTt5YU//lRJaq94Ae1MutJeRqmLnhIbYQBWR08FtipKUDr
nU7fMs/BCrB8rkTASUaPlH94KD9D/EM3UwS5J1xceZo2z6hJJqM5X/mqiuK/7DXThU3LgJ/2G3SM
m4F+Sk4yl6Dh8mQPe7UVPtLWKygf8/NBsLwziWStuX6yYAslwk+OjQy1E/kAiKCrnnMQbP5lBPks
hNZMJIZt3jOf0sK3iy5sMwNip6DB2P0J4FNUTq/8jBU+10sUyh7c4uSGC7wvv7k1w74o9rbIvTQ7
h49nmZ79DvdHhGxxmVLfGV5P/TtrX9hvfPSIwhuZRNlyck3oGvD1+l1PpP+uGc6y289hpypft+4S
LUbRfNuNG0kGEHeW4NLfN+bmhu/qtjrKI+Lx/ycjVypm4oLR49/bLwm1OucrYKNAuQP3jIcAK6HA
w1ygPnmUnTrys+XPlr4PMYnzzGm2vf8QBIVUGIPj9GmJ9Z2Psg//HbQGGaIuxH04Fi3T70FA/o+D
5quMUfGWUW+HHa2Dg9n+kNkfRnZuoeMt7USen5wCGFFed7f1T0X5XmE7d7CF1mGLXPZ8n+YVgd8e
Qg5JxOqpMuuPaNhQ+GAVEQvYc7jTBZNXGM7kJEV5hOS+eDbnernP6akrP4dahHeuYLRRWWEYm6S6
LbDLDHegx4Ki1kWtnZJAXOHkZSa19kspyl2LV00USeZ9HJ0RMMLi8jlb0c0E7OHd4uHEDk53RVjc
XqLGiT5hKC4sv0sqdgy7c+l/rc+V1NSLhMyp5vT3zdu8q1vPsTvdm/Oj74/lM8JNE+HYSUDBRrbT
cu5HpkoGFwihExxEnTlGS98rbkzfBopBouiFyIMSUMWkxHwGGqdZB8gQZKFSZgLrH4isZMpKB74G
+XMPrIPC3qTwkF2tI9S6N/iWDugQFItNZUllptqFedE9NmlGvsSe2PJBKVGARWQpzFXyURy2vbbx
W5X5ekWbjG4GBvuFafFV3eZnxguwqWYMaCSqI9xcBrndzGhco1A17w+h5+MPidmFRcYzyK85X+6s
2RL5HThbDtHk9hEECvRhpVzyKPv1XBEPLo9ntgjohDjxJozPtLb9sZ0+cNRFROLHGVPOi/2jc2cx
UCsShC+tUTERc13J7llU/TNpoR29CeJAKdCfuZwdfPiUt+SyrRdYKyLhEPC1ZB6ImmImULjaUVZV
f4rH8sNABwD5aiOzHkRFyyl66H6GYHXpp2qX+Q3TIug/rdmo5wQdTTiKrUsWsWztRFYPcnEyNLQ2
1YkLNV+6o2Y0Gsq+SflBjdmnYE1xWXxW6oA6cBWFD3Ta0bMf4pEjOxFNUZnCbsaurpHc4uzZ918f
0GtNgCFCThdSxQZHDHNvHB0aGuflNNbz5kF2kCFafzCbjNuz7FEoMdJbxJg2SFfRXlGhDZosjhzK
Zj3B5+poPiWaIy49W3s3/p6VQrsNcQrAvW43ZHjxLD5WEH+hz300ldkzC5zsXZT2e+aqCeuFrQs8
he8Rf+5BJXa0SqwQM+L6Z87siXT4ZqVW4hQ5o128dma3tt4K2OQtrSL4/Ua1qs3mM9hxFRv6nX3w
W97OR5o6p7/p903jA1ArJ7VWjAAPtCMYKd4XOr2aG6pXkOLmOR+I2T1v4bPEjsk+jfaTvalEuyOR
U9DBmzxHSh9jgk1y1RAxP7RwejFuQRRDhjblAjkyKaOG2r6mBfIX48ukva0iMKw4YalsQUDUJjvs
UtB+EjSzYQnxnFJCzipVyMdEiz99pPiO/gb5R8gHztzInRZBddx3ruD6Wx1XzryBtogpE0c9pFYG
TwnSum2CB586hj59tNsjxX8wNFpeJe5kK+vpPqp+tEVZX/WY428TMm5vEjiv3411Cy5HXLvUeTDj
IlBIfKp3GuHMRpnCYfP1po1P2rwgQLcq708jfdCLDqYjOc/+Q9yVlywhsrF1aIBRfNz/I8VF32gN
CO3HensJML7R22+3LvXnZFH+wJBfkDzhmOGKB5oCAXZ9xUyGZk6IRMrhTvBJO2vHoONFzsTKwfs5
r0i2UbXtQ9YHX5Y3XXwu1y4K5omtHLM4luWVSCkRATnVfihNtsRwjPoZ0Cod1tIn5k3NDc3PANZK
8CEPuP6Kj3/ytfZGGSA/S7y7LpmXrSXeINHfWO5G2oaeixzAk6i5LFXliGHuUV6nC3wcOjyC1Vnz
lNWgib4AagvQrhB9d7bFUNu3cQGSVbtM6kXaji+dCDQXz4D7+CZNJN+/uOLepERoFi91XRbqX6rg
6WZKORk/LzpKRBFfvdJoQcuthOus+efb5K0BFUmBpkSfYtIiKpMD0bZ/Rd0o1ckhOrRoY1PaYeDR
LJxxR5cGJlWaKX95wPS+oPas/4DyG0vYyViEB8oGf9UkszIexwEzomaM1oFxQP3zKpR4a7Wlu6FB
deC7R5Djoe5ZGjEy65Swhgg72YQ5CzDRy6FC9li8vTzj6D+YnBRrIcvjoOcH/5Cl1TmXOYojlN5M
0KsLSw7Rt1ngtck+LDNyWlkd9W7EZAmNI8FF/T1UhNfYGpq1k4UEIfEG4gPWodHtA6lL8UZCHyiL
wDRht4QcjjBLZ0rHLQluls2yBVpmKUd6Zeq4ceg340UbiZUF1SpaoXY5EzmdoSRKPjTqU3Yw6iXP
f6LCeTv+SujkeqQuZpCYJ/d4Auv4r2kgqdthiYkN8GbPHXkyQe1eJUjgYvGN/5GZOHrYlc6085w/
ECY+umeuvFrJZmIqdd70dYNs6RmUlrDH77a5ojYwvNLROJzQVMwcLoo8ZxGt6KYaQqt6mup/dxD2
PR5O7WSvpu0n14mvOKVAiERdWj+SoY+JcHKpUfO4BlpEtuY/HAhj/BUJEUcbiaGq5vBwVmydkzlw
4w01CFwAm0qE62OU8cZaE9c91ThiRUw68HecWUaa2IoLY+5SibnQfhBkcBF0aeUWXeiYQadC0WMa
u0MFUbXnfzTssIjHH1TwQ36ylmC503qP/V4J3iCJQIopfywfOm5Uz1/nMHUfNgPvclqUtgkUfoRl
XrsPVSOVHB7ihmgNA+GU+MPRG7kKOYxA56o3R9BLqWAdl8KOMtV1aVOkAO/Y+1B/5y4YRejGu/aj
MU2nYUD9dvRmcsS6WS7+xLGoPx5+Lc4GocHgsiT4tpIQtyZ5qUAyfmZohEs5xnNTjwg8cw7v/lUM
U4gBsuGvNTtUBF95vcMuUcfVGW7wDRjDp+j3vLs+7y5jAu+dLE+l9E230wt8RxVB1ncuc5e4xIOm
7KWLPiGP4LAK0S8JBkFS45EOa6Cpmel8z6z4zf9OPoqjpeDktH+f8wRRgGi5IpToQLl5CjgqKS72
zAQjpVOItOZPPrfH8S6RirScj10ltoZVBCOJoNHM/Hw0XK4c3trXvmJrog+vekESLeXxt5uR1an+
szD6aAjMOUlzRy3UOSOtk5b1GGLi/tnIDgOT4fP+Bj6rgb8UHPL165w5VAJw807O4alBMTGZtA0V
HmhdDy2MpvJQdHSIDwzG7mr5Z/Z/mGakkdGZJmKKYQvfMZ8whXAuHh3qmm1QEn9AaP958b5+D1d6
s40VOtbqImcf3bPzu6J1Yj3LaeBRcxiQ1TV5+c2C+yQAZp193oVADlSiutQN1tXYMVFIvELUR8tc
cjVMiyPVJm9f7UI3A+5Njl5s1XHaOW9QOklEmEUiIX+pI3KIOqtbfbYSukLmLxQLgqbMVcv3Z5gq
4xSJvW8Wmf6DfAZ9Bb8GiovMtKDf1bAgdzQFYcAosR0W/S4cISenXLuYWc5vmec9usRQENwsdRGD
FeXoAxlVQ5aWfYOsHcAL6ZQ81Dfh5Wesl/NWfaoWJw4hnfWn5dgDJHnuF8o1xAUuH7wcZrw/IZw2
RGbSMRJ3EkD4tLRBsUUvZFof4wrWzbFgYsHVgDxVQUNeRSNuDux5AjiQ7UbEH38kBKKGtqfo3T9N
MtYKApUixFTxYBHYGrTs0otsCCmS/eat5Iuxk5EkXliT1bFBU03An6Wc2C5RJtQQf4VVUPGpfnEv
47jZnOkJssKWfEDLdR8MLPypjFyQBM1xlx0DFarmhdaR8EWoaOuqrAWT+L0I6m9eTRDs8utdguSd
5n9pb8QgZdaQKR+BMkFqBQsfZPdIpi/rWfSEt4b3IwBdb5zsOO1fqwxiU1Qvkc2GNtaWm6yhQbTZ
jhYWkLnLblshBvJvmYo4xp9BPIKm4V2pUdj0G6S0zK4E4LhhDSQNDchPmYLcezoXwFbjRRuo9NyU
oTl2nd+pkE43dNOkrY+bENARZZ4IHHamzhYBiAzSKnIAQysBRs2VqMDUyQAMcEKvccHEr4vGz250
D4JO6OgtS47bnsHSvtqKjSYfjxqzzeMtQ2CIqITLYAKogEFLKBFr00uARYPHtWp/CUbhPvrkSr/5
8dwdK/V+MtvgGhhMjxplrLaGO4NwA2bavQn8EYiJDgSd/oYZ62/MJPD8ReSBr1izpPpE5DiJLTYe
73Chq6Z0VRo1W5MvMnnrTMo9IPvc51nK2O6gVQ0D2xfYtiJpaYbqk2/9F3thFPh15eqg6ofNxu5q
ucZJMUP82KWkIny3Y6e5pZ0y0X2oos18EhR2lGRurXWT5jofYpbEM2jwPuO18h5Kr+2nwmr7CIuB
O8rd8XLGdFKvPTHwDZRH0mUedU2WblxmgVZxHQrdo9bTR5nS29XEXOCQWQ3mCvurjtij25BrndC2
wRZgQ9BoaZK5ACJmL66hf86sz6N4gg0wBCGZNwA63WSi0fRb9AubooVTMTM0Y3eG5ZuypZ2+br+o
VsQMdyABjQZb34ZMvZ9+gzXzFr4Hx34IkpA771glDAc8HuxIvunLsVIJRgJ1fVodl8oSfTyJe89X
DExb5PN6uabyFLsvMxocaJtluMs89Rqdm0atdVZhp5m3/uOhPDnUt3sTyI6VUuHKtGTbQ+I81iHo
iGFEVXS7ARHPCjx8erJmHWdRnuhNEsa6dvpMUDmWH/YgAG/hiUc5LHyUPeIQgxRXHIfMst/2m7YG
XhRCyXnADWlG9+ZhJZWrzyVsMhB/6EK8Keodwk1hbDlSybm48gEqH99Wgl0KYAhkABJcCnwywUoq
b9yNB03h6X9wFr3m1sALnOqFFlwyoN+I6FSTomgAoWLoO7vvPWXx2Ilxrmsiwho34lHHSdtpJrod
MazLM6QQi9T/c2zuGj1Jz5cQvX8wg0j9mzPWiP8sj7dXTMG7AD0Btm9bFKgFRVMDF6rT3TMFE1/r
gsWb3jFHi59xWjrJZwXfAGUnPbTMtW9L4oCDDM1p5yUwXdsf0apluV31nqhvJgAvVARkg5QzU8g0
yVmb/V06opT1klGik+lct8uwzZI48L9uRKXoN5J3OQu3TIOl5INxL8BwF39WjPzCtBZAynJFuzYl
FxxYZC/CoCaBrmigy79ohIa1y/hlUfp+2eglf9ZxHHyIkGroKG4gycoMp/HhWylk57pu+hTDwB5I
523c2vfkur5PbhV/xfwQL5O8Jvm9MivIUSGZPjjmBVRArd2J3NiulRBpJpI6CrmlifU4eo07dBtv
VYGbzpxwOzgBoDEe1Py+Yrnylp6s5ktJc7x6xdWBQMRbjK6tDUaB7H1my70OyaKv3LogR5PzQ7ag
wu4XNTAbkxR5JkmuFl4gVAtreAbw0ga5so7N+ks1tYRR4FW3iqbIiFNF2RSQNESHvw9VWPCfvL7d
6q8mTUJJcVxfmBsY9/07OSKMurIBkm1kJeTqmhnxgSt06To5c54h7FdBvQcL5e9uEFuluoBmMhiJ
ZrqiY92CfjykORbTxQu5UaLp2letcntNPvGHuhQ/vUvKoW6CBvhE13VLXOvL426nkTOU3uWikYrg
SlO5ytFCqz/G/q8azGl7iWdvW2xQ9/fCsaTKa0Lvjx54lcz3n8BS1QxU0vqWRCS4Rl0kMBDDR1Rt
miUSyDvDjeMa1fJ+4WvEJSpuqL1SCYe1HtZ/pbeOKjUGh6pYPpOsTaonhV9U0sNNDtuya/JGShfu
7kgww8ummKyOwLhBAXRnRf/FCKNvapodHQIWZdUAon9tGaTIIIqXM0G9OUqWzhHrzlaSIylsDC/s
1RBSTEWmwycW9N6tapXmL30vw+pF6hgqBP0swnEIEHlRbsmy1oHM04vTxe3aglIcKhGWrtfQ/3m8
+EpSzevdTtEvBXwpCcBoG3amg238DUHaFBmZrmWIm5SNuxvIT7hizYfSNEOTutq8BcOpl5sdT4+c
6pewnmEIGgG4hm4ZiZBNR+Zjf0a5ZYuLtIS3wCU0OYrpg+WMLNPwhLqKMuitw+0bYBWkszyBrvga
QZgH6vH6x0h/U/58IH0W7a7+HJ4kyDtSptawHvzdJM1HXrlRXXorvansT04/GC7UouKZmaYW8XJT
tsJxx+IU4fI12JYKnKAnRgNbak6owv3tunpZ3dHHsfj4bCFbyodGmSUXBaS1/16kwUxdYwsGXqDg
6esH8Z4zVkwTdD1HCswwwCuRV7vROD/av4A70TvV+8jmX2Q3F+AVLagYwEJVh0i3Ch16+Dq5DU1v
yIK3SUZVWNfdXt/0sVpzplHoKW1XOHmUiMzKPVla/7e6DZEpBShv4UQiPUdNUNd+9J60aUHpcIuL
fxg2Ey/9FFQ/HPxpoTGDqu57u6S9duXwRcEUG36iXDu916d2XaSsuI3VuwGCujS1SivxWe4td/DX
rLrRkhRtpKl5fatOO1Cz+uut/JYlcch94jPOsjgz8s4r5Ol52AW3ysJd2Omv+XCE6JziShqvtvtO
rCXaep8rkdS7sg1U3F5tddGP1e2dEH5ZWXvOmrReG2orQk1co65h2cMzCUeAvXbdY7/Ux3bye4TN
BfYpT19v3kigwEinz7KtqWGt1+6F+t5+XquygAefeiMY+OzVg+2IkdEILFcCpO8fBVHZeFgr71T9
xqnbSnKJ1fXBPGmNXVtkMdxYYx7oD2EwTm7s7HTw1Xb1oHbHpNQWBsaUIdHpR4VbeXEwMwNHWxGo
ogSVC9cjI71pt44S1DWqrZ+FfJl7sNChMhbPtT8d09yNYmtIXWd6FT2FOrvcdvW9kU9w0A8F4ZRD
vESFDwO6mvoWsO4miQ/NZune7J8D/4o3UHGz+ZjcYrevfAV4STvo95SEfUyuHey9qFiQxrg666XJ
3WTAUlh+Rx/bkyzWT9nZyUpQS0B1X82r2FePCHekar+3qhqYK/HyzGJXKm0O87AFInLmrfojX3kZ
rwwgXYFMXivlv05mFmIsN4HiFd5yC4lUlJflu1TD5c5gXc5Y98p1unltJHYZsuVVvk5QjS1d4pN5
oYFzxxreKCJTl4ABUaMfIIJ9ViI4s7AoQsDq3SFyH4bPhvtqgW+xPY+mJOs9loCC3diYCmxThnuZ
U6SKRyGLzly5eQAONgACaGsV49fqF2vEFuQGFnywlKRlxJns/SIwvhWJnmi9yRldvWCWF/CGiHzH
AMdOjFX+yjUE/2KbeLVNnxoVR/xm9Y+Cd+8n1uVUM0idqR71GbD1GmoB9PYBevc1hm5USyCIYSiA
ZGqA3ZsOuPcYDHt9GAfBOSR4JSLKco+jzW1QYlTwiYgUe7px/A4vvEAQDteCqv5orlLEtBvbkWOL
io4677g29NgfAhKN1sLz8vayISWm5d92hCj6HFdCQkuvIO+1NL8gvNGzsUWTeX7S4vCr7mUaYLaI
of0P0xfR7y9qi9e/ITkzdpeeHPXfKUSp5bmK+lFo4y7x8yRRuj7Y49CLTAjzRWTO0pe/Uieku5x8
dWmF5v3Y32YEkoch7VPxVAfgLt0kdX8GW6u01DBtb4VBQ7NZGOfTthjdfetccC8vn6urEq4g3Pxb
umI84VZxq0C+o/IUndZOrPnoF1tTmHoGFx7wV/cUPhEGtydnmlu/KXx8lkEJ/hYsbkSyNzV4f+Qp
NBy6pC0KuOnsLI9gqNI+vRJ7lVjLHKHyhfT7ikFWshG0PwfmUEE951cKHdklSM+wy2JcS5f7fEVE
BJ1PZ0y8kuJf9GT1qYbY9jP/JXyLQt1KDUsJ5ceu8+UubphfJEEXMdedy1vz2HjrWE5r5vpDXbDC
rFuYAEHdbo+JD/xg8W0F20ORACNLd5gRd74nx4sxa0XnFd7yeSElAD/7zieD4bYWIMLXpbdZvn2g
lJjucBlCxKPwdhCePm2YBNXrpUedBY/gYVYGL5rOc7lQR4Q/kqzOjj32HCBI0q/9CLsk5qw7eqjB
vz7+uuKUPw7gX42N9726qG9wvoosYY3aRCJow5o06K0ryB5oAt7PGbXaCls4WFgTlYWykwMRLVJl
JP0vrEDtJFh5YA+HN2e98uPv/J/SdwcROebic4qTxdlL+w3Zg5HOlTW2mQW5vTvh+Rsa5W0+cN1P
xwlG8dMqBdFqDC7IoRr5gZ6XWH0gwXux8CjgGn9BLKFw8yrE5+6NxVCpjKpDeWvWnav1CUflk/Ka
cxxGv6VeHv2iAyETr9wKMAinwTrAyDAbS9UQK21NTjAVFWGbOIlHlijh4S30G5SkEqvRU87tn11M
Zjua8hnkH+m0r1UHGfvrE5nvu76nKegmGABxrtfq8Lz0R9H5AouFPCfZ3EayUWOc0Vj0Gzo9Ifxm
KlSRc50P1+EdtbvfxVbFBLJGVl3O7dvfR6YMPR4snVN+RwglcWlpY94vK7dvOhMlBhSm3euGz2dL
DPEYhErSBviVFRXzj9cwfCvdY2HnKRMDaoUmr1IwnNf4Riy2t1WpVtiwftYpUIp1GpmesR22Ucaz
FyydP+1SOC4PSW51uoiqgxcyCvrfiWoIZCqemS0q0XfU+HJyqVyruSiUuPG8VfaAH6YphksUuO1r
li3AD+eo/enVPtZHwh0zidhUbcPwbyA4BzUaNS63rUYk3MCytQ6PFOkv/VsjBzBqkD/MeV/YEVhl
+kePG2JWuEn8qAcXssYu6uIr9WHDawqUtqn8z3/VJXtEZ2HVk3bwf+HBPoCvvL58FHSsVMqUfmrS
p4i2NYQLB1W2TKPvTIP/Peot0LXtDELq48IlHhZPDG3/volAxdJ6yx65Fxg2xqJC6BDXlKJZSAIt
j7614jtWxvbsuHlaA3YjThuGBsmaCoeFWnDNuBnoshSXn0JDNGkNluT5kXHwu6uTu0mXwlbjPlPi
WaiNsd4QdAjV8O0WIg4GgjTNUXZ8UIglT4dNiWJLHxS3Us6pEHBtEWmBcQlz8KsZwRNmxhYeEZXA
e70xtmxnNe2jOw7RyRdk2jGqZN9HHfo3eA06tKsYc80tRZJNVQ698kx+Ov/fmODX19DiDjE8qJ17
rVWCXJij8YGJJBWqmkDTWnWCM4gRQjd1bqL+cFTzH9BQeVNsbpyccxWakH5QC2HsOXqwpS/9zWea
xexCAPWImfEcHdbvh2PKlruAnVZkx1kzepSIIXRcPShJOIUeI8m+UJvbrMlH2vLilpsIZqGuRtje
j70L1klH6KR+vhKpWPrYfnE6u4xSjTYjPPUIdkUjZcBictyxGSfQB7Y+Yk2pm5yaBnU66rB0UV3u
BnjcKLFhP0RYGj8HPirXy9wHoN1ifJrV/TLwTXLBMtciI+O3Ob3cPqnDMMkg7kaG2Q4pD51e1HyG
UcgCrF8rqOgNkKzAGd3+rPHuOOW5cNG+T0qyj5xoEsgZgEu4MgzEt9FvZh+btZHrZS99Yebe5qCp
3+vJPwc2L8df9Gl6NDhD0txD1jhA0A2vAUfhvoKRRftATbGwD/XWPujWqfKbZc+UfPCtNBt3IoIL
GXschT6EptyWCtF0/UIK4cSffTwYLny5YJFCZLXL6ozJfluuuG0EcF0wEG+epDHvEaYY600sUIUJ
oOfdMg7SrtEpMFjaOR0nwzULJ6lRWFTTM7vfhACGep+BF8SKvjjdgIzUylozdi4XCTSe9pK08/dj
sODi12meeqIklFlSQvZHSVeZZnTcNkVc2oK4UQBieYv0ZDK/+nFlsSAxwjfoUjfZEJ362JNiz8Ki
ffqVQ2PDq81bVD/t5lXgxZNSIfsi9P/LmA1Cd3ZLcTeA9or34vPJzmHXi0w8W4oAH2K3jwp6IsJ0
uQmUEUjFy56pk0HQfSVPd5IplhzHFEgd7eAxYgQ4tjzpCwwnHLpMwhfB3dRxebyevDoKUUGqQgAb
oqH5Ph18WjQaUg7GZ6gBf7Oa7IxQbdVxqwS7maOkuX9B9lQySKPjnHdlqVs0sp7uwUDJe703J2wB
tdAHER9GHPMsky5UKqy4/xodPUPqEPo7mSQC6fgDLW0rs6IcEF4tJ6HofqB0GMkiLt5AntQgvWgQ
qqNQXKHB+2Un6Rdr2nDRBfpfW3qusYUZKcCwhkGJg534F/LnAGWoUDhwZ6Rq0OzrhPYGzw7jmD04
bqCJNEeqXB1y0ODAwztOa/mZccl6BAv3cHFYOkmGlyQ0BwMPg8fTlYxzKnGS6L9x2bSO3SNhDRen
dcdyHtkEW50DiUw4aEmSmz/+lPH1vq5wNpMuAiWZb4UKD7InpNNa+RsI8i+JafwhmzI0huZhHoUm
9YSDuyHpZx4A32TgZI1nkla2TbhRdn0zSE9MTtlXOa9hXCa5bulgz7KzNGxC0WlyOX1YoMEGLTpk
Mad3OI1oWocl3C6BvT5JIZw31GoIje5a7oztdkm3hbiFz2yareeM4KzF+yGv052RgxrOmx+S+CP6
9o4xBJrM6v1qW70dlUrg9yaf8exlMMmrBETWiX0acgUARvX3Q32BvExuMfHW5Ua8rJmqAG3h98xl
B1iQCzQIAG4G0D/gBfzKsBY8YRE+X6RKghfzIPNp2DxSCzBPSCddoeEpEjRB0kcHYepa6+BdOHxL
b8LQurnAOpChKjX1h3LER3UUiMgOz2FgtbAb19biSOzK8I9OSK9xUcj8AALmPWv0js1KdIUJC2r4
TcoKxUzK9EyGUlZrFeiNmyTQVmovKps+g44OVzR/LgBdA9UV40ytlFJSaOVQA4BSDuLWqDj+lLJg
1y1oS2kLjr6tQsnjo3TbOv5HcIK8dCJAm4GWJ8B1yiu+JfSWJj1LTS0pMnxGNthY+ATuYKU5LmxX
yk/N6susatIgBtyqMX29xThs7gX3e2Gqic36wSaTSEiLN28PlQbVvPJ6/A9LD1z8lW8gkko+9UH+
0kvofgkhxV2m+Mkbg0YxDDXk2ga+2Q/zn/BxTPvWltc8eXwViSsnld6/kQIDcR4M4QjfFva4lUhg
BGq5I6y0Nn+3cTIE9CugKeVQrmbYHkWSTjI6QuS8w8v5sNoHsGkSoXVm0humYFMI/28geWo5xvwK
4H5s672yGYqMYvB1byTnkoctzhuTnBqbIPliZrHoWCBT3Jx51paZ09qaICuHw5/tzAarPHI6yU3B
VNfgaXCuZYrjioqTshoTwlAhdrHwwb6Ph9K1I+15sKzRo1AkrI/ykJAKVnkqS4m9O+StcpK6p5/s
3o5KAwq9AXgNyUMN2/0F5lMhLBzj3+LEfUVUUTr9spOyYcyNruoSuh5L3N7VazZUmGQw0BhjI0yg
O/wmkJU966nrCebMOrKKBEGzauc+u6mk4erSgeXQk0D7RrONagzOkrImAh2SETG7nbweieGqoj7a
Iiu8A2uINEptg/U1ZNWThF6lWzTZM2AKUcuTunmZ3pt7P6TuW3J6nXkZQPDgKKr4d6/WV6gcORQc
wrRtzn1zKncmOPb+MAeJKni8qcIUVnL051jqsq1c5ENqtzZ5rqaJG7lc5gXgoQVsEcHEu3NfZsa9
u6tguXai6vubDbkXy4K3uyExBZtJRBBjd7qYAspLWPKs4amNVHAxqTrHNQgK60lpt9iZCh0YOefZ
RFLOmx7V4dAYnYFgxxN1dbsCoTab8/iT2q+THxrLs8Mmcmu37wBSF8nf5AcS3yAFU7S2KDvBZnp2
PF1HmY/jWJKDBfaS7GTnesuNptm5ca/L30yJppYF7IKxwm3o27YRaQHTxRVTlnND77/WNnDOfn0r
Y2KzlPVipotxTu3qX3mUlsR4DH7yHn9SvJgWKHNCKI1KB2YpJzObWxkTwrD1CZqEhLeTZVSa9Hlx
igigYtr2fz0221vCpYGut3ZepntFT3uexBzGQO3WwSQXb5f9fyTylvUqfo22bvRmknDxYsukYuLT
YOrRO9hqiqxXeO2P85WC/m8rFX8i2GvDxLcs/ENGQpT9usCUlXIBsJrxOffKywBPfgdrwox1BwAQ
wX0P2ioVqfid5IM2DsCKN8jheZUtF+YKpMNge3XOhf+4MnUrjzcf7rpktn057tZp+EKNyfNdHtYM
63h7tv77Arh9Pw5Mx7FqmyYCCWp+f/5XRHLr+QH8MLQhcYv5yaY+kZLcfs3ynJyTxCYK9kU7yb0h
nzyWWYgwFwaJeXl/yej3xiv8kvMLBk1Yindkvs1gMm9vF6P2c+mwLkj/3ms/Lw8JjI1AGlTeSCXU
zhF4Y2F8cjxXEtbP62i1vflY1tXjKorIihQ9fAzUeHLlKOkQRaO9w2J2TuPw3bnqZGyT2bVQ6MeO
QrO6iFchS7A1VwJ7YgGYBw/MOlJbaCAuc+xfJoqgSgopwfeXsePjpK+ncic3CGAOMdZEh5/BN2kk
rHUnCgTQiT00uJhIhwQTnwn29aQNNn7RhmF/g8OE3Y5XuQ4gFQ24zBMw9kiyvXp+GqtP9ibBfqBh
8fgL+ESV2Cev/4eTJSBpYAmbe0SYWXFD99jDp/tz1LBU9jD0dSX6M8q0+f+ZsSk7vzm6xWMrOFHw
JFmkXk31k6ymrNF+135GjOgNvNiwlYxGSRZuevpt8twzryQNOvkB1zAjpJZ/dyRSJkJMyWth13u8
N9tQsFTPuwpRdFCbILcOcuWhK+5W5ok1jW3G4Ru3+ZU2cNsc594mY/1A8HY+294GkOu5OuqAcH49
Qyopa8K/AZOh6FeALOkaRJ4pmLvLQnEQgDwutFhIFv3hs+Oe5iCNxdsBjmWFtFcCeNH5pWsz4c/z
6JRcGkDVDm4zCiAhkXQgeHTdEH89yjOm4xs8Zxmo6qnbG2BLiFWan0AwBZy4uAV/Gs3l9qN92EYQ
UKQOsAfbzaHGnEYCVe2VKr3KBFVW1iAYXm4Uw9wDOoF9hveGqCglmFKyT/3+8mnSZnsoyP2BVokz
6Qco7RRJLMM66r9LYDvxh1RizBkutyv7oDTskWsPb8UAU7klmTz+3Mb7g1iitKc4E4+Ne16iSnLQ
/D+eDk5jplbzvnLqLeS7Rxf2xMgd3tR1z79MbaCzX8LxWPj/Tj/p98TLBzxZB4uIy7Lq4Xqc/qWy
Pl13V4Gaz2O7aWetjrvMjXln1oklUsshzN2QA1rMHTVsu2t0grpUMB/p4/rhFb73syXLZ2TKRdTq
yJeTC2dfApPd8EISWEIpMabcMUA3r49b3ToD3t7XbwQPktnaChRe17/Xr3ZAByIVaHbqUxNnC7My
LElgpwXg/NOLJkE7gQgUy+CwJb2VLAm86YuGT1W7RND/OV/QL91JEs/R/LlSdbNNSXFL4SQUJKim
1oaU015tUoH6D/EETT/l11blI4TEqwZqm23ZpEFeAUUT4NM5gMpPKQ4yIAaOoLu668Ek+Cpc+E75
9A7NMNgjbVLo2qP96Shd9pMHlux3PYuYNwnbiyCnDFNXxZbvBCa9KOJONahF8aff+PPxBNcfQCUz
a8aShCgfS9nyBp4DAFz20jE+gOWWKd/u9D7khqgcl2XMjIxbGSkhjA/wWsDCeIlJItTt64SSBpnA
VL0y+19zCLCB/zQvQkG/WIfQK0fuwJq2rDv1FnIeTkXb13fYNYF3Q3zzADH1vGo/OyOl3FqAK7E7
S8qDgJojv47VCMW5kJxN3BOlM85FO39uN4Ru/EBMFCHu4ycSKNu7sz/9fmIJuiTqq0o/JiEoSM5r
K+h636LeAyW8Bh5Xgr4bir32pT1q2XsY+3oUpjQn5zZyQEd73lG9cqNsbDeC4UATudxpB8RoUSOI
qYbT9tsS8yisVCSQbEt/Qrd4QG6eUFEMWG6tz/3yq5DzqbUbUS98hu0nOw9d4+B38p/yfKpSOIBV
BrvVTTQ2oOAwitMA2GoL822dRNJ0zdqqFAjMkPn9/CQ38xLPqg+XIFTmy28J2zIgjaFcp0uo4bs1
U4SShmWtgwDKzr+xBCNGzypLyx8sAqcErGket9QNoLnaKAzciAg1cpj7vWEC+6VuAmjO0faWx5sn
/0U8fUnRUH7mTQLVMSSrL1OBZaGUOk26/whzSZMgUJb94spostP2Fz39w/XHfqo0EjGynRwySxjL
GS+nebtthAwBUfDeiLxw96BK04RkJBFYkNegN5G+4yMCuhxAL7rMKl4bGG8o61tn3x3iMBKjxZJc
RA1b6Di3kuX4enlK/kmzkKLE4Kvmj4tJt8ZBHAH4W9XB1RIJ/JWFM8IhHSeAxJA5ts/Ra1dDUG6Q
WNhwIPfQxtHCkKQz39lIdmQr4v0KGXj+EY/EXJsdRurXCnFljbFq1Cxr6M29/9AhbXvNARfgECuf
qv/6iPZcfXUaEmpSEU+nAI3FPrRy5MToUnIWSh94n7sEaKEgtbnBDETNm/7vmyUaSH7KFCBgRL7v
mTsucObTGbybOdyYRZMoaJQI+C8FmHHe6IrAXu6ZT+8D0fJaVSQkbVt6lXbfosJpD+NhnO0h7lvm
8OT2fFOnkPfqhxFzgF/afJ/no95V7rGCmhwyZzSFA+YKOpOhyjz5awEKRwWDQA9H5jt4O/q8ShoQ
21Ue2U4zNx9NUw1UtHC9kOvdNR3z9SlJviWb/0+iszvTOr6+rb6BFcrm27zMTwhm/X9GxI3ZBqOv
9a6LYcjkAAHWDmEHN/DNeCUdOlmuNQEOK4zMcy45ccQ05NOmh8uhKX7moHrc7Vaw3EbRActcJvlm
V141vYqa6avObQCIDJ5zq93OWbphC4PpXStJGPlypJHdtQoJZRvjV00XrYX80PAWqmEwAPBqWIYF
5rfA3qsAsRUc+GPfxzb46vm+aFc3S8l0k9aepSgv3XjEnppSYyxtpG2Qr2MQWV/nV6q5MMB1dgBX
DbJj71Qjt4puT6eQeLwNkdh68mlpYt3ZgCDO2o4RtXdgbcXVxk5kj2sfJc150jHq1zYI2BZ2JCqT
yxCTsg8SND5hzmAt2POziS8Yqj5uyhpCGuO2qpDu/O+3hHisgYxfKJN1c0rYCg/rYg4jsQMfdhLw
S1gQo+r1o/U/3znatXG0pkr1QIW4Cn0KSowAGDgpP/YR0biN+YtCGeIcEqSQkX6KboOwfaNh8fPD
/WF5OQN9lc8QIDbkNFZQkV08YG1SI6ijvOlOpkM2UGwdXrMpbLmza2fNuHtE0mkU8BnR9DN1zSw5
YsuACRM1T+8oHxv800ILzvNDxs0mWn1m473lpP5dyauHspHtRz+LflhSUduEUSHIaACtKhb1y0aX
3Odxc8DWTIbdZKRs1c7HP+fuvmaboh/bqgqSJtH3o+lQmZRiwMR8UT7qOVkmJhbVksumHNFZnibA
Pw16FI0iTN3fPdJBfa8U+DD6suNlH5bEwuozaDfJ98+Ka1yN4reE3WCk0Qmv+5R3UWfZAgP8otOc
k89Wn/u7usQlU9TzNeuTvjgVPDvAxjFUyvqPJ6VTI60VAMH2dPnegsAYJecrHmA0f86T7RWUQgfo
ekzoJ3pxG557lydfjeK7iNxDL0doIbf4Awq2BJoahS1XE4cgGqlN5+IPb5vRoSv6vWBi/lw89HaU
NbW1z+cGX9Ij2ZrHXiOEfx0F+gU8UDOHFH2t9DbX2rHy2ayAklloMAtiWmkhE3mftgaOVl+B5pXp
vHUs/+U7j25X/Dbw1ruwbyWqEfLtQRSM5MLd5bJPdQvCJXB6uGJMBbgakqMdP31MSAGB3XvE0pHC
7LdWk12n0/bDa3fQG7VtiGUgvnG56YEJ26/OwbFm+0olzrZhV3WPHZ7RbOcFdhO8jQtVkhaxiIEY
/vUNrDMz62gA1XNic/LMHhbbiehJz4W6omwjI9C7BPRQxE5bLR/9YifaLdIWwL3fORW+oGJYgJ7p
hzvaLWHI9hOsjXDhLFWgo2F6jAt+tuW4DZbkDdfVIcaDhQcX5QTzubJzMY6L8W8FJRLXJtjOwWpZ
x80JFu//AjWw1yuILxINt7GYQ5m+mRCwvBpCXniUXwQgBDDH6DrKvHq8l2jWfryMEefHzP92vCXK
Lnm73W8hmzMXSsN1IbITWFlTBWkDUJBskXseVKAkhc/E7Vdx+SqppGortfL3R47bhj8cspHKKNO+
w5A4TLA+kO0dlvmJWIP3WS1Lzc6mq5+sYJCoGoijBd/AXu+iHjKbduJRl7PPvl08qsxwoluU7uHN
i7z5fK+N9Dr/w4Nalp0FRXUGEuydrkZu8SwS061mqZ0ggwNhbobVX+Qwp9crbnRIp03oeIDZoZ0K
Ki8FjKsiAiS3Jp4GFsqR+6IExwmmsnsXu9arSjFzqhhOxYAZNJBfY7C7ivKYtEgU01WasvBDHckK
WKKjccDLGPiW2xbRoiUxMgZKC4F2/8VcX0uKVbqA7WssYmZvozwuz+gjtH7POf6qDptH7Y5vTDeJ
axgZzVcpkz2ppEze0vE3+LEzeq0nj2xxUZEfoG72uTaRR1Me3/pCwTsw5L0cHxYn7HyjNW5DQqjy
+lxwlLMvKXJfJNndMeFcUfttUC81RYO3OTag8Mx3vMlG5aT+zZT/VvCPl6U0wFNEE+J/a5JhkBF+
yh20EmpdFL1P1f0BTOa5pTyD90H5yOczqU/P+qJQau3j/h7ArtH9aU8CtFR+/1KnwFISXpEF5HNG
4VeqJKxMtuYQCL3vPPJPN7ZSETjL94XX6Fv84+hwmYxQKjINl/fhIG7sv3cFj6KJJt9GlEZDNugs
mgnhsMIX/3LP9kv3BCeIy+Dg3xg5frKDEmiOGXuw8HP0/QpgK1uZ4E4kHnm3/0pf9V7/tEaGFmlQ
2IEWn2WXiUSs3Gtxb0rUYzSjx8rfvc/Bp8IWhb/5AjL6H1CV4sHdz/LgtzrGD5OrCajX74SHS14x
EIJ/MaDyk3vJfcT3gTQEFtlzxIk0zv7wPVYAtCmdfNAO0YPT4MJunl5QgtWRfV/0qZ5ACp11SN78
E3NBe4WeddobPnqGv6pAmn83L/qMtHXWLqCohkYFtdHhziMGzTi0vr79/KpL+mYQ4ZQ8VqhKpW8G
Lo6pBdsjOLBdKUN+5RklH8h1UxmLnpkkd+MPi1U497D2o7qybCdkx/GgAuapZV48uGm6+whyc2fB
9DQt+9gTSfjyNG+ASukJA4Xws/yAIYfIXUPG64Va1C+cnJzZLIo+quxyroZnekszyDchWMnEz2p9
H85SNGvPtILckpk11zGwwwcHzC6/oWOyeGek0yxDmXfpDxBOj22KNEUWN7ryyNRH+ZQfOO8/MYeC
8zDh/q4ogytVHg1AdJBLm8uXa+yEGJh/5JfOEYZTOAMgsmUtCXBnWoTNUs5k38Gx+SQlW4ZLrwQX
0KuxRl6WW/jOmu3YnUsO1p6iMGgXC/IOdf55rvIQuvGxl9nEE12V/UtpUN/GJtbB5509JwLaCdYJ
bkfpL67O1nD7Tqz+aJL5WXIHibUNsMtLNoyaxF/G1aGxb0GPkTm3OT6e8hUAXlnLNXVxQrhVHAp2
E8Q5tCuHpZimRA1Ja4tVm23J3fKN0Gm8inn6aglTYUkNBA4qNFEZPwoY7gp/TNXYj4Xyg00w8aLT
ZKeEKyshb/ThfRZZNY713FT8AF8tp47eHUCYq0P9GbA/P4m3EaIsJ9N5H2ZCOjEPtCCc/peqaafs
eaHJpdqbfUWzXDZFFBa1qgZ4ZsJnrndRp6VIAhEiiJb1g4ZsySpS+24ICy1YkwfY5BLiW9Usg0/m
6QOtV/ETx0Pg+sVhTOYQpzOsEqPaTLNG60HBkSgGHnvQY8Yd1Ml4aTOtRxAAPDDCjC47vp+HuEsn
ZUWHesJs0DolHpu8pHtyIwoJe2crAxkfl8PWkmjwiO8L5S3/ZD+ymyKaDIQluWEj8WhLuXmNGnoB
LVjZRXB1mL444XnhZThjXJTx9FWnXhIydprca0EegySOVlOR3eKVZBJnVOVk8MxY8sr6R63MHzLY
N0duoVxVWgE8NB+F1ZId0a2Zn5mOun7hHrea6yvh/O4PET8/YiR+3vDeX7eGG3hFmgJdXEM0dmgo
L40a4yDX8flgUoc53r7j106Q3xp0eWOU0lvyPlcBAFjL/m0jBSnBnhJISOoVdf6lZjyYHO1c8y9k
oCwFLRNpq2GHtB39Fk8sGYOwxcvi78rPB0reJddW4SPs3TEFYOpn1dquB1/CsA5KbXgxVCfa82oB
8XCGhS9OtrMRSwyA+GX5qlxy18+MkPMojm0iU2qgbd5vuGE+e5+M7+w6yjd+3WZQkkCQi96dRB6k
MoI3VnutU3OUZY7iammMKXdgmZ1WxqQnzV6VlnQeLf8DJp7Gd+OpSWh0u8XwAZ6NrFnazlKQmJ5a
qx7WUwt1NWwx5RdyjTZbL8G+VHDjXBq0DQqS2v1MMyyuzTW9yBFQh6lnQwIwaGN83JYAJWgVjOsH
t1jxhYuURBhx+LkD7Kk+tUtxo7eimB2B46TY5BKmYTSpW1jmpyDko9C6ilo6CIHKfXzW6X2Egt/I
Qz0jYtlzjlltVA0UXDwkCif+4fDXLRwU5i/7QbUsZHYicvNnueefZT1GfDsVWNSyi+FDNFdXOUXB
VGVsg8LT0AVLDD3YBMJ7zqwUlbhfJkeB1vwI/Qlr2d/c9pr0PTdaGKOiaFuLjbp1WN+4hl9lD8MA
i/GFSnkX21RnJ0tMLSo1R3TDowEJb4TuPax7g0yLRjQo8cV0JTfg5njWpyc576sQp0UwGR5DsI/D
eUXWEvoXOKUVcpzBWC32/LPAzqtb5wwcfW0nAG5vtL1+Wd9451Hm6H8KraIMpJirUZo3BHCTUoNw
oSlqE/nGxN5blPX3/EeC927Y/D+47h+d+8xZdeZ2Dr/i+p19TEWE7iTfVy3wajfNdR7K97k0ZDKL
G0tFm8eHT0NjWmQ09e40By3FQDVsXMRtELRpIS306pnLK/Xe5mfUfTXqU+PWnEBLqAIChralb7dq
QRvUnXs/Z1L70JjnYDlEfKG2LgnWMq8m8GHUoxTCylM+MUDxw+El5CV4+zjootvz4omriZcSM//r
MvzWcM/2ucegWdzYNve25GJ0mJtmnnR1vRZbvemdL3WOYsayv/G33MjOZEuJxWqQYVIqUytSfCdv
VQF7Zmwp++a0TSXe+mSeIOkGRbOGghedpOt8kN0m5ZSpob5FITq+5naAB7T28x+TOUu/FPC0baXp
ucmZbRBmTJQlPuYKzgQkhpy1n8lrthDGr2s4mc8b85xVu12uW6+3DdRt+8tAQAb7OnIep9m/qgb/
zI7bMzBCzAGW17v/LHzkPpgQdWrrHh3lkMXDDIBMnPeqh33GIXFd1ir1SMeXHbLT9GWB+hBLjmhf
T7d+GVgE18xK9q/RY7JcyusxIWNDWTzAjsZGV2x6fLOfoE6chCGy5o0fo5zS032/hsGgaKB7xGB/
aaxcxruXnTp25hEZbhvm1M5hUo42riDNWfQccb2zdxfi+eDcZl+rEYaO2v6dij6xnIfe7MWZJLiy
VZpS7X1wBs6jwguggeFjPOvD0ihS5VCPUKf7kFmMt43BylW7g+ha1GzvcUF1jo201jCEF7Q82jyM
BJLHESYLQf4OQN2MH7hLNQRnaZZ2FXIX71I6FcGS6nxpSP4iCaQ0MlEJs7TeUQ8TAHnEngcquwUN
SmsQDNSniy9zxUAdTPp41pz03g7fGgh2jKPvUniiDfu7DVeEZijhnRqybf1jeD9za1Jb04sV/9IV
J9W6pz+HwfAw8nIG3pxZKxDrM7royazb0smr13cMc524OJzbSEnP7twY8Jek7O6qtALsvcvlsgdw
MeLzvQG+9tVEwXc+FefPCgUwc74DVBB1BEOyIckaeeBB7k4UBPJcK8Z/byPRtuPxDu3hVBWmnJxl
6Q9xtr3+kTfceLRp/bvxLH/tjSyF7nE2wF4omfpnnTljtEBNTW7HYgenjYKR0soZ4buK4WoGGqq4
2SPO9mf4sYGLchyscLtxb2Q4jTPBYYn1/Klza+wUtnAjFlSztys83mqfrZpi1JYkYLt4EnZ/ZTN7
RkXfPXnXpfXI5ZFm+AJ5GomCw4g9Yepcf2z45u05ozkqnv+VDtsnBXZcVXbiNzjwuZxFy4V2O4sc
E99RL7wYgDKIP+mIML4nGXjfCGjH+HtwYya7OsPvXQEq8O1wS4l4EH/i+lSqtWK3M3LbBN+vN+1T
pi1kLbSzwqS7abUiJsf91dna3GHyJMw8QyAwbls1OFTwU407lULpgHF6ot0mpFSGmeu8eSEGgjeY
qf98AfmkvqNCZxhtmfObIHYuRIO+d4bcxZ51XhDHY4es5yhY7N+n1l5UtE4l7L+ZPp8iod8w+Gi1
JkrMglzsTiBL5IheWxBrrPUutfERZNcdG3mX4xEkkj4aedYorP6zENM7/3O3hVVW4D7BsHFaWJKn
3OYpKx1Z4Yd+gwyg45/X/JzKRCqDjPvuYyWvE5WWMEx4y6uE+598ClJAXGGC3QYjp9n0KY9L0YCD
K7V4SGVqlDHCn4/XmUWlji0kOhehJz6Sw5CTk+X/5f3MYxJvhdFORSP87MZkdBaL/jVeSHVlVqXZ
g+4LF3HrNpccV8exGNrpKuglTnxQzC24ZvzAGLzah6TN58P9fuOagKNN5RzM4fvtFHcOlgL0cwQl
J+p6Izl2gTzO2TjznOJmfvRLUU7oiSD5qqtcQWwZs0y8UfptydnliW7iyVjRwc+OUiN/c2ZBd8eJ
aYyRHwM6nfGlY/or63mRFt4S05pCrS9cv2wrt4XAlw4/idEkOUqZYUCuss9wApXO4Q1gt71fEx7d
4bHx8C5mgb8wWOBxmrGlCQFPgmhDosuFw8u7asISdF+vQQ04GfQrtFB8nx33+LYUqugjdFj23aR1
vDbCJh7JBncrsqM5YBXgbUYmj6YGWmcrTnfCQMZOvXAmMP2WzdmIWAcZhcL5Nhjicba6Djg//fR3
mRWXk+c1MPyxKQofbMnllaBVMEaRbA2hybecRCJMidMNG5wl2FooB3tCoOpPqaQg5ZxHl0AiFak1
F4PdTsrg3idl+T+nf9xXYlvYpVnR15gSm3I6Ho7wBKe2fcjwemdp4qTikud2tyT+Luitcu2kvsps
xx2HpC6kuBzNkEepubuwFarDckzF41qk+I/cyP2X64sRdUC7MOZCagtSTVeJFoWrMFJC6dhvZH3n
PrFLtIIMt/IzDuPkrvdTYoM3DJtM42AMf4j7ut8XRpDc25BaTNeoNst1ctD5+hYmf1ueZB7RZ0l8
cnP6yn5Enh7QSLKRW69BLBtdU6+eLa0zC91zinmHXaFppVteiEAb9BFLEhSfP/7KS7P+L0ccXfhv
5juwuMGKhf0bKitnZTtkB3N3+nQypkpwlfjOYpav0u4ElAkAhnAuD8tk98qUeBqdLFIw1PT4NmIz
V6L2s2ZG8DSmOss97AkcHPOohwtDD/iQoz92wxHEVtWjNdNf99dUSlYV9VYeWdDnXbj4RlVKLLRg
IkDkvO14nS7OqxFb+qLBeh4UZGGYQvaik00t+N1hEWO9/hB7bJoUcwOb9Zk5vU7QbAclWzfMWH5g
VIyOvpTnCNxGrXruwCVSm/IQYqEA5sv2+lnpDm2GfozECPTDq6jAAs0aIcZ9+0uP4zeZQslSZ6MJ
F+ad2qT1vhD1kZjsRibax2ty/9R0E9LaDHx2KTtPyrqM9D+jYxi/ZOWS/119X72PuXEJ9y6TIdvU
pDRPZ4dypPFCYUE7oDm2NiYsV4PuJA0+gtO48fwXRwpVxwxTTiTejIhLqBOYSiViIAsbv+vugGCd
wl9pSvbdLKTJzYVlzHnZp88jpVslG7A+5E64fmTd/fxT6lRvUpcTjABTtf1Niy0D7aTAG8F5hlNj
8NHAbJn6pq3uAvCv0x7hzD6Vc+Y/XD5sAepB3fL1aDYcA8nd5NDNZMwb7BPHlokJSBbyNLYeKY7K
GGxwOLEXynTn3SqIHlSDoZRjUdcldmelWnL7vR7fKjqyaoX5l50tG+Gh8q4hbeC4VyYzihQPYnmI
wGpxpf5t3u8o5JWZ4j4KoQ+9Tv4OiHJHJh1OkvT9C/Hk1npX9X8W9MdN32Woxgm7TTBW7KBLHNWP
OLTlg1Rt0wmrJbW39q1Kq630t29asSl+DXB33dMCEqJ7exLvUvmPlFclL5uTkEWhhJznXMQvjnX8
GPTi/zC+NJnXOkobQfeD+EBB4ekHIvAV/wUsKcZcbsFi6aA6bubwpYxUnRmsW2/BkN7qb5YlJuT5
pSPXlvoqjDVlkznpeuw1O6m1Nct3Ls9xKQm1a0Ju0nUW4EJ+7vj2cfB5+h/blNI6HaOtvvfQfZoI
t+YN1733Z9pP2DcOqMsUoMNxkHRqzeFDiubWVQ2mgpgqDmZeC2F9n+LCUctUg+xcVFtF7RGEAxwn
bDs+kmgCJ+GgsZ79hUdeMRgLDh5VfeSWRRYniAfkHBs5Wc1UMciipo2pv+Ta2TcjGqh6tgOTdHgS
nXlLnMdmvGJeYvBZcgsHHwVeYAC4DuHHlypWAdtJKSYwVJIviNv1HoAH2TDOZn3AvP50y3OeEiyu
s5EjVtZ4mqwHyktONSbpHxBRANaZri4vmilOT1kWaJeHzaSSsYTAcopBSIDMq38ia37cvMWtm35R
oOhGAixKXkutnUrgUWgIEdxpOZ+e/Ub9Z9uBEmNxCewljRDbeAbdHB4NFFqLeROEXg0MfjkygCg0
hT0VkeY3J208ZXJ/mehxag0kMqvZe9fCDy9xWwqDz4seeugfo0G7G8bUn49d80thMYReTfgm7+WH
a9xi7gJGSXodB+SI+L9VobTejtRSAsn2r3nJCGCDjSy0y6ufIurVH8d3G/O1nERNORUW0z0OvWCz
VusCR/WS+/8d0aw9ztoBZM+lYa6yaYAxHoGNbgDzrC+xd+rfuKxxC1VKdNKB8KT/og1Y1hpqnNyw
E6FVl+BJ+MIXw3b6d8d/0AvNruWzsavAa77eRN+D3fmsQlounvXUjPnYN4WK6Q2Wet7Nh1sSaWxU
7dIMpgZvb3SkTej7fIfxWmfIezexNdDcA1qFuKhdhHAN93av1SEt8QSByxphLf3JdpjyihDuE0CM
zwKBlcIEVVqqYAYdGU5+hujgwd7NYcCfmPUtgkM/KevHafOYRxvA9ZK4agV7KIDn/yFliQDwGRAF
HK7TZKhBtR++igDmo2cipHL3/bKiA1IE7Q+mRUf7j7uagiexaVuLjkaSOG7J5sZH6GQJksyQV+VO
IHtTSc5bbHzUtyihGB9bXZhlpq+WAhfeLhMGota6mwes+SxzuvsoQsrnXBih4SJKyyip487GrFO8
H0YTPkdnbDdVtcVEv+ZiR+20Vg4vIR2PsqnBp62coCFD3KIybnA59KeQoBb9VcIn2WFEk/VqzP9Y
DYmRKDPVLVSTOTMv2GsSe/0gr4G4+wMmYByv5HPCVRHtUATa0vJbs7klocMfJC22N3obeZHYw0yD
l6nahu6zZxtpq66R/Eri/+Vz8XKsJXlM69JsWtzs1krrS02EQtceLbtY5xQ0R/jiuy4jeK7g/GUK
cE+pOsSEXZuP5t5JZ8yWhJHVA3j/ZBzgy9cYwxk/+qbJZKlc1UN1dpR4RjOsGa/1yR3tcBkUwmJp
uZpl2RT5NXN/+RbVVeIkFKbKxOIbspGjQ7+3WDuizM9lh9MG2onKABrWLLRy3fSffPNdDPTlg/gH
d5eoAQ7v4xIWdgXpi00S1dBwJ7WSXOWoRWx46hbn2Ab2LHjJoIJDEQGfdZQwzaluPWKP7M2dEJ1N
JyWjjplSkp3sNhB2abXjGZG9fCdAaDTufROS7VV8R9KkQscWLXsWBo6p296oxl5k0CsSgg8AqoTh
eXMA+XYSqMojEWT5xicZOAkUdfMxSqQZ0itDDhd434negpxrfTuHyBVwr2DZxRnWw1Vey3MJsgaA
9N+vTd6FK1jEIXe30OiYBtFoPRqgEEanHQa6L05mBkGWrBGB+A8djQFsbumJ0spVnyjraQ9iRXWH
7oc3eOcae0kWsHXF2FyckHKcosAt59tBpsUwZd+zHTahLzUI0BkIwb9QZxwapO4i9R3mDnW8zbm6
/XdwklpztZ22TvkfNCyuoUFuNFYYH5WeSalu8Iw/AAxDxjxQBhqVz843j4FF0M5K9HJQhQ2i829M
FGdL3g5SB4WjIP0CgYh3JsBiVGVGX1Kj4mecsOtR0rumqT3NU6s6mZPhlXKO8TL5PITa84B1TsFc
p8Jd8gskYwwKTWzX/q1MhUlbNzxh0Lb2u5xQlAYMpMNrggmlhEVarRXVT7USFrDHqquSBb6awEO4
TiOjVi/BjyvFEXgSsV4t5GQjCsxlhl80zOMRNmvMED1AUxM0Gc724CTuISk7bEbSaLxWTTiafqJn
tZAYQKGg00jJWooA8mphq5ZK5AM0pOWDmsFJCZ0QVdZiYJTXsAugQ9jjfTPvmR53u70NAzIIJ3Hg
zK8ieQiuePR52mCE0QNAKflz3T0/0Q+bWIvIOVGz688ZGN7esWZfwnNtUApvvgpQKuAJnqIIbgZ4
GkkTkMAJCzNK/qlXbyAXwMWK7SzhIR19BgyzWTWeO6EVWZnwwqsQ7XannDlS8FzgWS9mDnmdraQs
oZtTJbhiCdanWOKR5Pl57C3zz3CopBEjt6lWqx2++fVviJ4f35KYK9dydFfzJHMmRI1Y3miHZ5SN
jKfgNYSQca8jvo5ilJJ7FaeceeXlu1sPp53llm01QKxal2KU8gdFu7s4k5woqi0c6etzuQMxQM42
yMu09KVZ6De7VXbwpxMMMCLDBvRcZsbUXREMSgUMaJBiAhJ+3Fb/F4+Nail2Y0n0Xmfxnuf79bYj
vzWzcmO0XYhxmQkgFTm8FXLXK6MI0odEhldnOsxtw0931v3MIRXO6reh/0lStYU1XblWo06XXsop
0e3LcBUOeq5Q0d6q/WtHBZLNprYLLAsRTUjqsCVRVoH3i2PJ+L3reK5vfpOzfgM3YJYtNpg5M9s+
0TZtxLtt3pqicLjuFUtS5oh0gwgjWufcbEXDUj4I3m8pkV0RfhclKs+V3AcuoneI0ecmoG5r1gPr
n3iu96bW56Ne4GdbK/tpyVx3LeRAVIxkvmj0JDgANwPiGdr3Vp7g3VEvwhS8c58M6Ssb4uCkBDHe
Wo1lW3ciu0PzZTTmN7kYEzCFEY8u6RbrqvNsFl8Bc/j4mnftQ5fUqL/UqRTfMAu6Flq5jyZQD5w4
yFBNV+zdH8F8MjRfVV1Tzg+bRLRTxX2Uk8UeYwqA1tramcjeEZjK8Yo8JdkfiNWEvzKLRvoJc6xl
V7E4UusVInP47rBnGZyL91NAgx3MD0NIKc6Ds5LEBQyqBOyoDj6Nb8z2t8Okj7YqdefA0ZcRw5po
HuzZ11cvcgi6uxN+RNix1lKYycHBxvFNBwN6dxbwepq34onEimnl/16Bgf2dLa91CtazFeE31T4k
hqJ6CR0fbrQXtxycJ4PBsPeMNtXotiJQfhdHqhFDuUm5Ha673sFSL1Hx/TYi5biw/ViQgcmYtE/7
1R93u7GdICqre8WHVruWjRYCtAGdDSdj5c0IHuZTXW8rBJMqAwpVu9p5ec3SLD+SmY9/GAI8iQQa
w/wp5Rab6BaCJAcQWWqRPbAwR1DbcBUWjztEJN5ZxYM3SVWYcZJsdG3DaqwQxTEkp24uirxM4qyL
GZbjfRnB9RFrf/pjQJPuBfyk6nmE7vQLb8cAB+yjA5z54Uc3lrSWtkqH2Pfqt+aivOpWsLFkxX0I
vN6lybV3SGiBpW+gry5gGqYnV5JSfn9nb00/PgpXQSIfd0cjaHAoUbJqfHSPgibr/DNUOZk7I/3F
oLlcqtscsYUiVZ9P9RUO1cx1QRaZtYkqTza56PcH8WvQSga3FC5dKAQIZvIERzIzv/ndd38yDCxV
MGCGNAq+auedKw1l4R+WYSJ+Jqz6cvwih7/P4LQ4lhusvEA/v+tx632VleqnlIHIhk11YUxB7mVm
ka+DByeu3+nrpXgYWfXArEJSJOgUOEIsnxfaTbhyu0FKM49Qy9scfVRkV5d62bBbfaIngk46Z1aY
RteBifkmmTRnrkC3SvuaMuoflm/aSj5lyTr0LhbW1+HgwvxucArZFipI70uXPhFXutNOgvvOfRVq
Khlx7C6rER52WK47iwcuTcDJOoK3faBmkqPCIWQIBWaRYKGei7Gsyd2nKC9Y96HFIVIPZvki6vMz
0RaEtQSwXMbh5QsG/yWNWHkLvoBBv1U0p300Wf08otcQCSb0cVVR2gNlqPrmK0840AK1UvKCqLFH
iHsAS2gdBWe9sSxFO3sA/afA2GCPFxYd5L1+V06znQPk7n9hWzgRba1Wx0DSNSlkv6J9qAdht/pv
gZt0RnzxgZWz76Fry18Nf0ZIDWmuAj5xTJ4cEaJ3xqNVKICrY+e7n5kKa3ySzQxa/EL2pdOfhys3
lh6Uoolm3aVtIO6SWTguOafEKjZvtBGFdjKHiCovJYEMnjp9N5p1IFwDEU4B3BwZS7NrhiPwyISp
1Ruv8rZuD42x5I00EzGc/lkbyc8k1SOyH9XGKtUe8uV+31oSn/3MP1My1zFVOyLtNqcFWs7vJk74
sXamTIdMUEYYd27lYv6bfUAUgXbU/pOcuCUGxInYUvUmxsDVrbfFMqOCQwveea4kiA6p7E67zlVW
4euoowIjQg0tBM0JCSMSN0k7UnvumFhacXANOxOTFshO9MIk7lrEyVXJ6pQdBmh80JWXdnj2VFlU
AfaXuxQt6slp1Br903G7qUMIjfT5bO5HKA0ZX9l4TGs6L3mxMRwt10ZpYrQ+JgzPnQsKurMlbEDL
KCEbqbEwMHtRB69e0eLxbMm0VYbPbVcCz8fjwa/bLvQEXXqhkWrRTjyzaHnpwu2NcEEcrP//2HAH
nK7i1QZ0wOlAoRiZFQ7wxUP8wSX9fZRxWD1D4mWH5aa+8r3rDp3B8/rAL/qH2xfmbcONhCzBNWTF
GFns8YN/qhuMdxLrQ34BTpyvRqGcRRBia8BL+Tn4+vFlH3gQuuN8TWZiKeMXdooq3fLBToJYN8Id
K8o7Q4eLEEd9c494c9wS6/TF//dX55AkM9tTZkZtD5AFZarkIxAP6UVtT0QvyBVqyRbG81UieNWS
fScH2J5RDmJ2N8ZNAkpWf/kDMDLV0xM76wXkmeMW9EF7+mODfdhj4E9mkMogaJJA5tE/DJlFhfRp
ZlirVlQWWh0jqz3rkrc8fA8ngOYfuD/aZa3Rf0xp8PxEzMVYWbsZDefihKfpZrMHusQpi9ju0k0V
OXm2Ogz0li76pKsWzN/+OD4XgFFs3fQMtwdPsmTnCE3Q4yJBVU05dHfEM/xhRIqv7JqBJ43OjWwI
1Nu7EYvM/NpDja63x11jj4Kopz/8VVaamu2+cFlx9plANyiIi+DnUQdeTrrHC9kho2gMV+hosNmg
7LkeCUz/amcBBZqpRmxMtxE57fVuBEmbtigaojwrlM00K+l+JewCx8HIz+1TpJUr0IROwHU7+9MX
UjK4Sd2v0JgAhzJtudYayghe+EMC2ZYiHnsZWO6xKCRhu77DV0pVBrIzfYJCVX6D933G+45pG20b
lujgctGp5Cl6V0BG8aU6U7fIBI6/93MTj1JS6e4KnKZSsY5v6M2Xrl2JtzkYL9D7AHONi1CQBb3C
NqdAHGqgR2UJxTWxtPtzImm/1JYLbRre/y1DGTIhPMtTB5xO53cIwlYNSA4spJzgDNo0c7xvTj42
C4bCYA21Bm/nhMuARlV1T0T3UEr6UgUAzAHkprBMAGw+kisdxnsZ0KjqhuehXrkW0HqKj7b/v4NZ
dvupGro17n7B2KZwWo58CVPK3y63b6z5SMn3kfmVYwVtndIZ7ZzEhSaEvYAT2O1aCVc3uqLQLYPl
MT8+8bFue3AftkFg18xaW45GH+brsbXIQ2MVeekk6e1n4PELIjcj5MopfUN4ulH5jjsvlSAPmkMQ
IsFEP7/AjyrXMgNPKT8Lo4zv2FG+pEgLI99sR9+jAK8HiG3aaPKw1BkdQE2XbCwZAKW8bxb7dtat
sZvlGx7spzsXJtX4noRgGojb5RlqJUqQo4Ed4K5IpbOc6sOHPVtBQMs8oiQzSaq1dfrnTjm0SE0V
82BXC8oy0gfMzXugMZxe8O8ZvElRo5JJBTk97HaSOLkzDbi+IQyPXmgJ6QGiW2bpcQfRd0vqrkZ3
H0K3EU2K4LwuyoYCMtrnGlGM2AQ/HDR9P9dqR7CJmmCxmy3wXRrlYdiw9l5r3e1+9bXbAfZjJuCi
ePtZDHhxoYK9hjxVfG1TkdhiPZ+GlclqqWiiDZ/FNp+y6WHh0HZRU0bsT8wQNaZNa1pP6iqYBf76
T1kERU+iw2jpb5NC0Ib1xjeOmnjzxl62qorNuqXKeOs7TncfLdsZ2/VKOOFtfS4c4P67AJAMxief
Y/82NNquUnZez07Txbk+o4GAKqFP5wwe7nDMwdWSDV20T3WOULHFbx12V1B3svWZHTAmO5VZfbga
L3rrW+mNjzySQSUhAxbzcpde/Lv4Ix+eHfU1a/4Lic+kNwgDmK+PWZIixw6Jl+PfoY+uONymGEoj
qTu+w8itkpE/tKrH3XkJ3f82+BGTS/iRz9+v3OHuS5zf5yOX1Q29GxLVbKUjz0iGLnpTa4R9I66i
YtApIunr9kRJrXu3omASJN4A990Pes3RL8qWzuXx9nksFAvSNtqyzbl0jGa1+c46tODZlOqi7rcW
6B2SICIF6xE0tD3Jr6GihEfuVq3wJXvK88iNGmd38pDeReQISWa8zWRpY/jVj0D6854TeEGcsB0w
NRFoIQGOGfwFmYKO0ohR8WliSKJn5/VsxxQKxs1UrRZOfclfFMkbh4Cv+/PHCS/IgEvwhfyurjjB
XR1Zyj8LnHaMC8UOeUtSlMuDsyhrzNjqJcUTCmi46zJLlKkvm/wQtbc9rCou1QR5/0DBjtbZwIRq
S1qpO6w7JVqmHtHVeYTXbjWrTFxRg7IDDZVzsKLKqKxnvbBJScMfLe+eQwMrP8jdFSoA5ZqUGiko
BZFG1GGHzAQdzSCj+5CHElAv9hWVM0hm4zyvUEqcujENCoTzQhpLN7JMfdYesKrN0lM4PNSsvpJV
j0v4fxtV5eh4YBG6/ifkFtqC37/EbmYAwqSygzvj4Yg7wNMpsixH+DRedxulIaAUtCZR8OFcrUj5
d5ufH8VUx9jufJ2lQIoCwbN/TnjzVrLRQUWavFbPLu0qesZC9DEfc8CpFGqEC0jELK7fI8YRwCx1
Qus6wnvFIA604ITC/T2sy+0OC54obd1jaT1JqLgaPRM4KHkG8UJW8lTPAHEzwCGxXdF9lnlbtoXV
SVKbxYOPHKc6/l37/3FABV2/Tq0907ujlaN3NBcyrolmEOxpmZkKY86c0L703lMqpMURheGLQbDD
fj0eIdVvdVhfzkaDLC2GE69ZIp4HfwC/RcH1m8ZHXl05UlX4LGN+uj/ULZ9MujVbhjq5GksUzbGv
xt/+IZM2f9cgAtCMwua0hhGrLGR909sR90iOlaWp+7UYpPL6xYX0HCG9/q5P1L5l1VHIiHeXZbet
4SUv+GEs2/ShWPfSt2jR6QizD3gMYl0wgiMl9d7Qich9GhoWCuzL8eyH78djEOuHNjhmmIquOEKl
HLnkOXoMw6HqOpVrr1Q56c5z0WiGq5OTHrBAjDGTcsiy6LWao8/jtGzw2Sk6a2N0AEjzvwVET3EC
XT/sN1Jg7c97zdFF03Tyd0UzCtUPbss8yRG8HhUZ6AlI5Y+gGVNvR5glN6vxDEUvFA4Cg/U84RG5
3nzXhtMgEhbEhwc0wJnv+Q0VYkVhPTGHxhVHtuYBQXYz9or0fBJoxvQb4YxYajLzxV6CfxVF98ZN
e3SlhDazyUTpZtK6HelcvlZeIS1qT98OM8rasevvgat7T97LYNFi+FOoujCPl/3WJ2Rj5Pbiw7m8
C/NrWl0ta1WsLkLt97FuwhjZPwLJjZsl0KAMsLzTCFk3LEXdlWvgf/4BIUCnERZi7XXclw5MwbY9
NmSAMhn4aZHhBfPe2YVmpJ3lVsh6ijmCTQtsAXOY6XrbOH1OGnPah1XJtc6cqlwfNroz/+PTprWM
ynLkg2OiYgxABSb6hn0bIEgxS8sQ8wkoeBxuxLMQ3/nt8hnO++Ud81fzjg6F8cLuKVDU+nykbEDm
e21Sj2ssAu8xhbCd9pR/0DvyBdTngjXjD6Ob43CpNLbBjJDnUoxq6Myh+KVLoMUgEgXyGgFWtjLP
b9jhp2+A1RVhbSiwi7VOO4zPhT30wVviYwfv5isVUx2HsU0Qp0WAfxqO1WAmZ0mJRh6PQxSK7cRi
vWOIC3P2cLtMuLX0Un0CoQSXSVPetxNs/pNvZDKxApo1zGO1FuBssWwsNbykn/Ga3eUv7ZZ95OZY
NZDOQf2YC12Qr6o7Bbgoql8fxWOMn96W2hE45JhDNQZHu9R6lUKgb46yRevgtrJmUqfZjM81zGvW
OiYwiobRrMN4kfFBGbQEwA01lDzUvEWkS/esy08fewLcxOiTNfIqG72T4OJTlG1oZRDpMhVhckX0
dJMV/SorjAkAvMPRn8B2ugVdQOBQX17Mx0LJNgtxv+D0fTvmKLlSAMSyfUQn9Ixs7tzNTZk/akeS
/yZb4whpI7ZJcnYfW8sKE9T3ka1susRtIEnJf6iPjzY624UVjLCWGhagoZOP7V/sgmZRIy7lrA5k
j0CPQARGyUNMD3wn9HdGysSoHmw1o3hnBsjFWW/VglsjMUokhBKwt06KefDuRdrLCTltLFjwC8aA
22Ny5yXM5IEzbAxV4Y1AVKBizGcsnWAYTcAv120kPh5xtMtL4LvoHQv+sdepX2u4kyu3zOPTFETi
vf/+EDCwYmGlf6OnVndbE5jC3eXwfyXQf+dQyv2RPhWaJbxMOBEgOGsxsgQxsngk7h/D05/icRcI
05SFKd11FDHKT2oirOQ/ZIvEfO0Bc3kMvCbwDKZgvskFuOIdldV9vKYN3nOXHX+sAa5LNGdvUo4P
CdrIjf0DezMnPS4KIAJCKpqXP4mIps4CUzEIPbUJbXyWZQDcRb/etYio5WKJ64JfmCIvZ5oWgZzM
FCtcKOKew8tjpk5cx0G8qKnCx5ENVscQsAHEaWciYJwQ0LDAHdx157t5E52alfE+ST4EAoHa1IPp
ZRwyHR06GE4AuypzJzHqEWl6vIQ1UChtUQk0L4rSmfKWtT9fdr+uwPORXaItW1Q1yccbRwmuX7Vt
4QJieRU6NpW6VvCJFxC20w2wTN3AhCh0iICqEEo136C26DmNG14DI9pW1zuYZMxBDp9MbRU0bXrs
CXP73KDawpQzb03ELsSwD13QuvOfXLCGnb1HIvgSXUVdhIgviSZuTaaIvxMTbFbKDuEgzIalN+Yy
r48VpEP2xFjMUmZA8GJp1MWQMP4XMrZi8Y1bSzOZCA/LtpPRSqUdim+C5/VbvpyzPvdDYHLT2GdE
5SdMZdx85Qmqz/Ezj2KKHuy9HR3Noobra0Qg+7xIGKXYABIVfgPERF7aP3wAa9UBnUwXJWZv/Ys8
vqrBPA4RjKuT/h0sxVvRpwhTisfLlH1e1T6cVL25RrUVgYjY3czYgJbCwJx4FEV4FZxGFFdFfsAZ
7m7OhxqL3BCRHdBBXB59J9z+8JhC5ieEBGRRyXNdcBE9yaFa75tyAYQJm+9Z/7F3JL96DUB8U7NT
QUsNQo+sAACxfE51YOvhaa31mfxmrQXCTzB/nRSBTRdl2SlQtv+5A37bq409L3waogZ6c5lqg0XW
QH3etHZIMdEQzq+42LVEHGugHgj4La/nNUF5IaRL9AfEpTZBXhSlI6MRnYhOTuVhXQQoKvH+L5K2
bb97grs9k35EUNa35P31mzzQa02soKUBI4l4EnjN5slKUJlH8qcsOAnm6kTsSESd20dJmo+nnTsC
IUnJmoPJjgII9TsSfKs8n5dqfaA0A/OL2Jju9UncQeMoW1Kugd9jAgGfu/s7jgVsYqJrpJW3av8L
y7kLC5O5ykL/D7+ZsOjKO7IpG63yyVB32fFrywgjTfyerA53lJ+TVjLxVhDTjz0gU/w5EF9yoeNA
7YgAvDox+6jEs0kWSWj33P8GFczIPs09rpgyg5zXGeJzyu5kCCiAWFihTt9WVIAIC5D5GIZ02f3d
YLOHJm0sxsCpYQUYP2cMhj88kbLNS54Dvy3GCZRIHSw9A5RgIo7hNeRwa1f4rLW7Ela1078B0pOt
L8Ka2jII6F2dIWG8GFWYVE9WwhjNG+v98+tRswHW/yFWlzlRAPYnsriCXzu9sETPP0I6ocecE6UK
cD6kRiSGfuM+2iS3CAYOA/W8dXnfRDNOlHBMvN9LlfbxXlzrsRoQrIGCpKyNyMFnq7cfMy/e8w0c
NiW25Q/SVmBXkKStkaxMfuVHMKAu1eB6ikW4mf5eT2vWYm7P9V23xjoI7+JOa6XqYqpW5Ykaa+GQ
TxeWGOf5X0dsDxp5q4hIPMsDssFos8v9T37VRv7k3gRRDr7LuK0l314TRA/w5f187SYpRkNe+HrL
j7t0BrYqmWvDkMpZYryEiPZaJa5mdbugu+NOjr1Oy6RaOBaYltolRRx0H3znRC60dUNQ9GqG5oeX
4erWsbnjPKAP1VBiYtkpP38x3XjolQ8w/95tMUZBffUXzw141EjioYiW0ZnVVrEB698CbxH8GnH/
9rR3t6aKwyp8FZ+wM9rlFMCdlcAXT6KpGNFfyK2Yuu/HxdUVkDu9NuTkQKdYby2T4DD05SLYsA1L
PX7GvCr1SzZjw0Nz9M1tSHVAv1EqHn/3RPnpeiTfl2q0HYt/oSgBMpCPB9QfYTUFeoFihq+MNvL4
6X83GKZ1b86nskcendGoJbMvsSLy8MDr11rSlP8ZiLe5+B50ttzoWaFKTQ83gkN8Pn2rhFJXJ6V1
6gG5JBjXwHLlINm2QxXvPNASAwLNjt+G5AM5959m3QxiSG46+Oz7IASKInaxUwQx1doWYpVpYLca
oBRpSWpC5V78yzgQ9e3BR1am3mBQnDQtKsDGtlZqJirn451vIyOvvC1MP4nVZeGFTJsMZnbnPuBA
jEFURL5CIalsrHuGODyMe8pU8H1laPpUWHCfwS8Sz7TQKMLLyfwi9sPUm7xJoxbBD+JjiIHeHFoU
AjmUPdhkmnRhVR4ikOrUaKTUd2yZ0QpzltSADEqIGh1HgDie2FuN0K32HGolLsIJ2yQSlrCTGKHN
8i1Dvst/PzIPHJmzbPqKGCL2Stv6OEqL6QJ0dKe+IBQuOnFU8qnnguUTfHGHVyEMjfX4/OtHcZyL
gSO7YsFJXqZ88nvuNGrRUdABGdxYH/zl2MzGDsq8Xjcjy4B6NFRdV/Ms4/8iFVaQ5OPlXu7NORo0
72MoLgYnXFT14L1+KkmhkQDusweGUoqdtuTn/UN202FOKuxjyGMcPCkfWDyKrT3b/8ijqhSNqxmu
H+CtMrR4CbnAsuuXT+uPKBPHbhgL2/3/qwj7l/HvCJ7Q9mBpTOhb5CFooJfB5uTIKMjvm45a1kFY
xJHkty5ClSeV1kc5kTnZEIow0Fwbo8y4qwUTfyD04Sdnw3cUroaSG3LTkKvXxwom5PvUS2As7lgJ
iuIK+18zPvzZjlWyiZT4R5D3a18tvDUhOBrHxkb9qNfIjAKoiQl6L1Yr4kM0m4XFNCnVe1xTSnk5
38mRbUOzjiqEPcaFxoGM22G9rp7jQ+SQ8HBz/aOfDDWHCYlCzcJe07RDgbGPmu3s+T5GwPBeobZl
A0z/8FWVryVCJOD5vLaoY33GCNbg9FKxRKADBMXi0+0iPTLKB1XGQ5AFWabBM+PWOO82WDvau2m2
Qqxa4PByH4sLLt6S6BDLvjooaCP+ugBZPf8JRqweAXKeMeoNBM3OJUmMYKVULC9Ue1PiL8RHPQTN
o5UV2+wvocVR0fpJnx4yB6yg9IOJVEHY+kB+33F7jTPpT0U0VG6FaZEJz/UW8vbb5q8mKYCbquEA
k5NaFy49fumJfessAsEhEoUN601kHN6fA7HEEoY/jeXbVV0787N16ks/gpczrjezxTDl/R34g5Zd
R3O6dvJb6BPC1BMJZlwXLauJ1y99mngPbSyniNAnAJ56eQjlSCop5UiyVg36pgws4onV/8Q3vqX/
oD4h54ekh8LICNtQcIDQ7dEazGKUmtM6EKpGDwyABsHNLFQcPRRQ1w8YSPB0QSgADMQh2KVS9jLv
6PvCJgX/MM23i2kjATl/R6RREF4OjuPs+FCK5qiDWECrA8cMqDIKOJBrZwcSVHq41Jy41l9BcMvM
jwbWwUd5E2qf72JYBZf/206iDz9NzdFu+Us/qXalFeXJdI96911Q4GrV3hDEpZiZl2UjI9a09a6T
hjUsxMbVHBuMAbB/bbPGYyEESmD6+HvNyqg0LEiJ8DS6clBYQWwvCglRVm31VoRPX9V+FFwSBwjY
dRdsjbq/2aQ+ZR+dArbqWhjGEcB2LCVu73JQKP6SD41QXzr0cqSI2HmxjBExe23Yo20OX5gwlbgR
9uhnDx3pMP0TAeXiyCzLYkJXbc+cVXVMNQcOuK+lV72feHZW4m/LXK1klRXm+bZYBFvaiFymH0cm
/j+k62Kooy36/A0zzRrVA0cfR3x8AtDMP7njzzKXr34A1u0VxgYyB40oQHh4hHfXlEUQd7LB8cg7
oe2qBMPB64GHSpnMuO0LNnn2VfE7IA+ARxxcoHhszynVN7ZsfVf22B/8OjcUs1o1fK65ZxRrk8+q
nsRUqrvRZOKLAXeWWbat0CRxqcMlYMN4634BLLOg1Fw/TQLn56e7VOfWz6lBusAps9RpGKAeFiMJ
/4PmnMLrB71hHQKlT7WOP+9AMD6sJRTTRB7w35l9iT9vZ0Dl4XRPO06IbiZez+NldN1Ucs+aIgoa
zoNHA3YQBT43fjv/GXISOsEL9Z71BmcfytMg4sEQ5RfAhzDxOUK7IdceMZbMYpqn19stBhb6Qrax
+BrG/VaNArZATlOo9orncxU8arWSwG4sk57oWP8PTF6K1lz2VEbmUu1c6VZkyPIY/FhCbdaagemD
XWgZsPRr1qBaq8AeAwkc0zhcEpwYelbux4YPb3gFb66S6N4ArOVnI7JE0sXqghpDGT0ER9dO2Pst
QyZTPdIVdGE2Pe0pBZBWiWSoMk6zzpLleCS0QtdRe2RA07K4FiWbfjRwjmH/YnulDGAwzyDz8dlq
EWkubmmAUnfjizczEtpXxuDX/mc5OoboHTu6kR19NCHpNX+rwUxgFgjfDjTkW0xJ8UET9r2cNYPk
TliycrZxDhOyHFmRh8pNfO+c77eb0jx9Fr9ITsWu/+ak4e+/m+cAB0Tid/9I3FY6zP2UxgH0Yu6+
/Mz6qRnRaJWGLmy59JtGz1+hm94GZoLJTWMthIpg0SI9CZTSjL5oYY7cF27YrwyplS7uoFpvOD4e
CMZ5ptiejmXkyAAu01MvSX6YVwPgttSyQiParonwxY/RyRfaJzV+7RzFf63zxqdjTRI5H0zTToS/
7IQA2Z7E9xj+Tp0NHpJXaxGdWKf9hRMul9MKqPTB4LiNnBHGDXvNxAuuWMI8iIuQGnzrwNf7qgbA
kbT8ZxMYzIJp0eXk7+D8fYJFJgSZz4FYDZNsGWZpGq+0pKjQwlZo4JTo3VuK/iAQ/54zEYW+Wjv7
3uMu1+DTXlgjm04cS69P/8daGJvwoP8NCIfawflNpblAZGrt/roF83/yUva3gmqf1XLRgw6B5256
VqrLor6IqxTWUlHcm7cbkigSPesVHJi64427i4OW2bbLrmdgyROcCjmk/ayQgf4MuJ9qmY5Kmazw
Vw3Q6by0CDe4fZ0VMLacE9flvXEe2CEETDgXLsTYSIZl76iRxHNsYrbAXIBfYq6OxM5aJYER1n+Q
yXnDUuXAku1ph4vCe2dexQNvu4XJKFCghDWYR9hHaA78oWuFbsrPWvJBWDJJrrC/rLFGjRHvrfdt
3bVq0LiI5LVjUxjnGEwiBWUxoDJCHsuz/1VgeR9wrsNAjSxgJ1fbpPLjwRceBdFTa3OIoasjLrgb
QBYbBi876nO+AW02EC4TRS00QFd4f539U61+6jrMVH1Twff2U0nlYkfiAkK881fwk6iJIVE69tfo
c3jyw7E3HECX0taw1CTcoOzfKzn5+MO68+SPHQUtSIQfcAVrNRa4T2PEwKgtLH+ZHVQ/nMGXKYO2
W7r3eQQbWzCnordlJ9Z/3mftuXW10n89UfA8E3gx3JvbNVCHHqUq/ewLfeb3ktIEm+zuhpmOd4XT
17HmKr8oVs87RAGBMtgg11FO2BwSiO8UQdWk5T0mAO3vG1JXy1lD0DNXlgpDaX+R3GEeLmtbH6d1
pbbnN5qUaXmK3rsbT0H44e7h2flfFeIbehp46xMaUla6m1knh/5/C6EvDhT9s4E10qD0T/Eeratv
uPjZMfRr8kTiYCPSKRHz7g9AFY4pWBZJul0e/rNmcQDoBWSJuhIjTLY/5u6FqkiTcfXxzrL5AQn9
dPFIRxOXgim8oVvqZGAUQi+XH0nLO0XM0HoBu3h6SXgvQD24CArFHV1GumOoeyNoCVoqcSodyVfV
8Q40pWUZlkS4StSfjns94D/OCtDg7zhrD/NlQbSGAECDLVJI2tB8qvpkw/IlY2/QdJqoZnGvnnH/
B23WUmSealk7od16i9BrYqtv4JNb17cyYYdUbCxF8Gzw9nV7I0Z6iWAd1CRmatlzCMgmaS9JYqr1
IjGBiiaOayiZ7KEaxhFJBgNLNzmQkBTLgBWYDphL7fUP6r1Sp88A0BoVpvaaR+gls9Ewb+RNSv8A
jImsbYIg2XfYvC/GyNvuKeHravzBS2JuilDhJnVV4+pV81pcirzzVuM3G1gOV52xGznUaow1AsBV
rl1IvhBIr/f+4fKZDuc34Btb8hvQSgvuC9y5LaNgfkwC8q7GZA3Mmbh0ZjIbRTynWMzbhqqv4yci
U3PNRY8HW6U/NwL63Wfn1T4AHmluDHOKj9cL+sW47QwSnL7BAJzBzp+XEFgKHpqtEejWF9Unn8LX
31rSBOdU5cBjnHtNYdGAcV+3UVj84+OZVqOTrEAbBG7ia2rNmCSlMdaiWQnqqUXhXQ74MfYj6qzs
bcsn3ztWL8wPvVX5OGAXmr6PDhhnDOozwYcnoyMTFTeroDiDu2lO8j38EE56BiP/QRV761CtqIyb
81bs+bn4OYoEjxnpU1W6k3HHDqILiu2HWb9Kt+A1PhmIgPomrJiBh5bi2i4V+TRmZVHI9v7AgPvx
IdghvaBP4XkqO0zBwfDxzD0m/1Y5sRdETlXWustyOwq9qSu7x4aI+MvuJVw7292JheIezO4G7sQ7
q13ttRYQ+LNUzU20ZPs5dSq7z4SXXYr9+CdEUMVjGREWIfXODvBM4Frk5xIfb0W6683U/z3i4zBY
bmsSA0nnknKuRZPSkjQdU86y0udKG81qygr/XTkk+pTqhyL19dEBhCtgUFdR4VGAdF2wToNhFW/b
Kz6b4BB8JvYwVcaAQ7M3rDwirBWQnwbw2H9BV/7cBNQ1gHI/7N1rJwtZ3i3r17xux2KXp/04BrVc
3BTi6rhSpie1CgnTxHApCfQGniMc18e3m0sN7/x5jKp8kWV8ORxaPbTgsTvDnMCmw/WLYlXxmCnm
OnhSrG7QWQl1uexRvwjCqv6tw7ydewwYZ4WU6j889oXMQBsiQ0U24axJmklAj9nfGHB9wcUzRRgj
Iqz9zM1WebZY0E3lQnCbmkI6WUPLYWxnkYABE6repVwk6P9uONZQ6yobv4rGJtRmTHBiWnUXOYrH
B3x3HF5gCpAv5A05lDD/OysFRiq6zP4PffF2ALMqXxapqWuuxz1A9UkoudKSrnG69i6Y2NmcTMhK
AfB8lD60gVvzgr2CUZqbe6+mFUXPZbMn0UhhhgSRd8hZpDTqJKoSqx8IgY2uisXOH0TWg6F56jC7
2G/sTOuhlljhKDK4lquxOWWaoLmN6oyTUlGNcinGYwG6UWc2n/TywjAt+g5cXr0kO8qLYJkOs8Dz
6/cuWaUaLo2zjlQCnj+mrwCtFzCo+2oKgWX16ViR/214wcdPgR11kdTtMB9HKueTOQsSCS+iVkoC
PSdtGDnghL2tjoiOwNDzY5LBfJIZNh016SynQNXEPkBLJVW3RTp/Cjj6F+9vC9rR1NYVqTiUri8u
s+9xZDBh3trd+KmbdQzxWs23f6ZGpM9Jqcf6AJ7rrbggB9rCES2qtUEaL61VDX+JmzA3B9R7p5Ay
2CvKP9GO64upVMq4WDPfFunXH8XnAwHNduifwfs2sM82Bay87/7g3u68u3z1gaROTluj2iDekf6f
lGsZAGCR+M39J64ZsHCpddoaOVV1PYKins8obE02UJH0hOMh6MW+NsTKEpLc444l/9dYKdGhItRr
GRvts7+K+bmOxqRo2QRrxI2Nl6jlaolOcxdFZ8JieHi7347BLb3UbNHR9t0LKOf0WIRyl55OquBF
w9nXwicY1rrKLV0yo6Cej6SmPs8lvqIuVjK7BE6U5fzq8CJfuVqPGkfkDUy8hVF6Pae0L4zkLuJu
mYnDekHrpezWCqRfGVHobF71kNmylbVQFtjUhboxDmKePsSgYdfkc9rxyril/5bsE3VdN4ccfls+
AiMBykmYlqu1DSgPCVhpUjlBDT2Q1pDkO4y1vYfMH68Io5dHru1fBkFLrljWPyD8Dc6f5mMDOjCr
w5L0NQtcFMFmQ4u4ZeSVaV+NYDQathSyYIT5XXOL25273BWJ1PVLHeGFcEGyc/Nq+oOHDmvAbqLR
PjOT15o2SL5mrW1Z23gT97s5KzsCk9fK1I+T51HkBtZSvRhrlq9xGcu9UDpz7ldupnHcXyHvzyLC
88+q3VkXDLW+6pBhH9qpVGZkiPl8jCBvH3uI0cljxEiOE7udtpr7JXe0UlvXswCjQghmH2668pYG
V20TSGVGQKZVMf93hzROhGvkwE51FU5/IphesfLO/sEO6YJ2CM2ATZSBzJPujxYIq8WmjyvJj8/g
3DQ76KuRy6Dbz+TRXDPDkHqPO2YjXs+TKkREf9qjE/noKjsnh9XGlM+NSRccGYCbWc2MUPXnM1mN
hS1oO34z2vOyYlBUB4CgmnEfAwq0VtM9O+m6mIUXwuEXp80aVtIg5AqbConelJaH2btJsFi/ZcQA
/5Z985Z/IUPFJPAs242ugSP1aSfMG/xQcwZ2dKV4DOYtWHq7JgSjI2NfA/YWJfKk3Wm/3gCRQ8H1
6oBSrjnS3X0zg2Ab+6nlJvrMzxG+pNZFE1BUjXXipqplfLvw6qntYVvO4zjRGLTfaH8DbUiyDnkm
Cf4oBQFBUN7649U1GaDDGjpejgq1mEh0btE8fsFhF5rGGIxn1qCpOEsQ/AKs/oJ9A8q4YSeFeyYb
TL1z3CW4S5AjluP1PI9w6yzsxcZA/cvVoZ2CIWNjUKBZTDX4dRkm5FqWcrZ/3rmsoI5AUhHmP6vp
KC+X1JNrsHbrc0MgHj0U6vFExkAPdrHvmH/D3E1D0/eVDQTqH5bwp6sXfPmVusSBJ95YauZcqv1G
FN/hYnFgAYexIyRqfcohe9ErokPj8twDprrOO6J80BHpix5bAudVFJ5561zbmOCKj7AxhpwyLyqK
cmlqsR0nJZ0puSamMNCY6PJAD/QiM5BT6bEg+JWuU0HKVF+2ITwI0mTNSSRnZS4A3Mq8vpkRcqEi
+Kr8TgUEwExeNXhGW9ztUi3AhNFjei1i+N01wqtrKLFDRaa5wNkoJ8LxhOt9F47jZ5NCIRva+qMa
tgaYrhwXOe41n/RSeqPK5MCKTUMMVRGzVrWaEii14aVqJ5alMzYNLdUPPB8DDpmYo5ZpPNBTeep5
ty1nfvfAOi+cB80BkSgw32M1e6ukfD7oLAnsNGtjvabC44AQND1xi2mOkv9srM28rNg0WiCaXzMc
Wk3TzAbW37Tg71INydAP5vdpWe8L+jl7nfX9w25lb9Op1kCWm7149Uji01xgwibqJCtFXtBgYlB9
tFl43r7BNnAq6/o5eFx+TtcVkhThZutXsiBLDeCSlaZtdxqJ+buyBXO9Tf8iZezpqQYV0OyMf+dl
hIBzHUdJOJqCsAnJeUMwgB1m+nY4sR35u33xZ1TgYd3cnAxzrlS2QowAXc1uUz3YwK4ild9tHrib
GFnNVTmKUKJZLNcNN8PkJXTKs12bCuRNdRHKetYzdcWxGJsZrNoHADvIcJ+KAzI8iV16IIEqY/3H
AshwBAOUlmwlkkwf0f/pzGhOjvcGhl5eer8I1CxzsvvyBT/2Qoq9WtBMYq6ipySCuVgA/rujRZaa
aOoCXGcsYQKdTZUDoD2SnzlRxg+JTjBA3lmW8mMOjzY4vFqe16nY9bXQ310R7CVkCQ30TyGYIVaG
15nS+dsCZE8PfM7UDtH051Kw1zp+9Z5piHJrFVilFLMyF7w3xNdVd0+GeQdnbpmv7c1syRWuW6/+
0Ebx4kjN5HRBI3l9MeMUy777siC7VxFQrtav2ZYMquM6lgEMZ1VLCd82nGwPQUmRAGzEQMGwhjrK
RvmCkAWClsLy7R7Y8FOCvbAFM2opzu+y55BA/a2JcpV49wq/v3yrkvIPpGvVqrJi+Djw6h9Qn/Je
V7mN1UMS7DFfNLbEabPc3AujuWALs5pZocR3fMXlu1GaOWMMjqodvGyMm2fY1cS1pFdR28nutaI1
GyRGpWXfarrg8l0Gy8rCzDEnMlesiy6icP+L4pjo3paKz6vMwtDRco5VVqeIMKh8X9BVqDBIksMa
kK1kUjr/CMtdZfRG0sNKbAQVyM3RcS34u49ODUVqVpjOv2MijM8gimGFLn1oyQTaJVvsG5TkoL2N
7rkh3FhIAS0LL2Bi18ilybJi9RwhY3QoFLfTOzAoXEiUiYvFCDqUufV60eZ41pVz+REoozhOLUN3
gUpOSi706YxrelGcjlvJetOO6fFpUfk/ukhwQ53M8V7HrRu/yiXVf4eXuAHHQfedNuBDh9l5YZv8
K6i8fjYVj9CHot2H+sc+lXmrUmlXLhuZDkdLVeXJUXZxsEww0mcAjN6TCucG0eIe758XwEX8TxYD
x96iR5IW1lMurC7CcLBTdERxpT93iMKV8fymOljL85X0Gsoly+m+tuLMn9yEZvGwnsx/i9m8cqhS
olCu+0I4ZMjT1PXhRU8pbzPFLGLvJcOQ4pqSrSIbZtQDD6UJ7PqrLzqqKkvb8JQCIrbDWkmn04lS
Fn3A6lbQWjTTbwwQ1BRNcqvidEJOsT0KZV46m+158bRrb2V53MMSp7Qf+RLgz/wA2n2K8zMZ3dt+
e0KmR/BO8+X4QlwKUr1QCylLiufggZ8WWYsOqdQWQGACUv9ohrJ4jw6i2Ew7OTy4cIYdfTg7gMr3
I5ykQLpT/+a8rrBtkluaSEwupX46egisf2o6krgu2rD/A6Eyj7Bnbmgz8zpsqbNizfNSf/3Ab9zk
6Q2eGDepSugTzSS/zpIGCmrUL5N77gwX+WNaisJtunRdCTzhx88rsffRgxW6vUdKU45p7OqQvIGW
YKLPzsjEDjzW1mfbPV/ey9yMm+3rTi0CxSf4ZBOp356C1R1tD+RxQma8gFyi7IJTKGX8tdJJW5kb
Gt/mOuDEb6CAEhBBdO8zK/HtIgZygxNy+BcIhjqJPOyfPAMELN6Gw/JnIhl1ILjroBhZAf/ZD7n2
5T0G7cVrhxDJpfYlzAUqijFzMjh6fAwxo+UXfRzro0IJ+tpEYXn97d9VWnEiU2ZkOOaiJoOhFRNC
Gn5WXZ9QrInNOUJN2f7h2OIw2auPVusO01Bka6sK50rfgGeWG6rbpyhdbmNA/djdwmGMbnPNRDOS
hU37UBL3SMa5znIWLlTTxM54S8b5ZzUK19lL2P8Y28oR/qKaS9Ein1Y4oq+C0XKUahUW99l/gyPY
csOKoyXoCmgr/BtcoInmcu9SFLaU8qszDojtV+TCr7aQi5Z7idQV6/sWMa9A/40EHf9DpIUtfxii
+MeoJx8E9HattDdsCsLREptnmFpI3BEOxmZW0fkHURPA4NgLpQBOGs8q69HT1MQWWrm2c8LcAWFH
X7qpkvaMc8xKxe5BBAt+4Vhcfu4gBoJNbOdMvST8QupaZbRyX6a2+x3PJDcu309f0I4+r+SrMGRj
eozwXRZy68hwk+7mtcLiP5Pu72vmXVm8eHLUblJBsfROgDBXB2r2JstVPQltSJjUAqF5p+nXXKu0
2W9625+vhy4o0xqEeQq23UOJR9Xv8F+8ZJAIxrOfQz8pEQLKiyiX6B3TeQYe6s/VJuDfgRCFag/U
6wIhQ6RTDxgA2JSh9gpUZ/tRk4r5st7eLDSIJ+dPOSR/mn0gzEUWBOHWYJVbH81bx8WPiaGaIc9K
KStRAvV2G3GCCXUVdWM9is0sW7lYnGPI70d0LTP041vGGICieGeQKtw8iVgYFbY0HDMocRWAJ2h5
1KknmzFU9Uh20svpCW5U/xzRRTeeqZEGiNPxAy2LuD43XmErmLDh0pXLgMOHdhzk2cCFxhdcNXYR
V9SjR75Q9+vDJqLiJYkE22HMk/6cLzLFj+Qzcjm2OOka6VCqHPaMEPy8lgnln/ScXl50Lzzms3I+
7XGEseoIs+piydXeMLTBJon7hVjm5tdh+SpK/78NaFfUFQmr0iBMStKHQPAQ+ilXvbJlkmUC1Xf6
v5ByYBqdY0OkEK/9ER+siQwRmH8+rEmk+Mgvraf9BfTiDkIXYsAqVl0yDkrxkS2xj0pvAWUJ1TXh
V1vdHylJGe/tpyLIns1+PakZdLsKiaYL2ZOvn3Dueku6yvUZqg5CYApbmBRifmGbWwU8j6sIHMXZ
pzifjT54zHEI6mjiRPVwSTdPV5Tc0cefrRmLBABcllwvvm47pmf+7RZplmmuTBD8uLfKIVQhr9pn
o3IJX9QaOKTAFqkL909qReR8TO9/lWTXJzKS9/GQX8yG8z8WGX8S/4WM4bO2tDaBs/tpVpkr1Xs1
3Jd4WmiO90jHR+i60+cFEGkod/WVQ6iCOtFT+LjVusBQL3sr7Un8EGZdDK/tUMSgCF0vnaacgjdN
exNVkbgk1RY8pwMFdC75JG4cnIgmocTzn3we2/aRnjxOjcJjjD1lj4GF71NWR5fPbWXQzgPIj4lw
1TsnfLUw6f++4TTvhbTuKm7FXqQe6YuPDszsYYsXtTppn0ocEM6YaqIz+CtyLct1TC5Tvxq7v05c
x6FCyDy+ebbzGdMS+2tp17dvfKcJ+rpi8GKCPMgJXKOKwuVbjBTYzLV5jdKx4SE2UdNKOvhbuf33
xZCzzOsmwkacW2MU+sJ2R4mh3nCusgU0XiqhftwKj6UnPfJWVVK9f8p0fZfzvlS1Ksbve3YJpnsC
N6RD3kxKQnRYAvH1sh4YbfseefZ/+4FoIPn3cW5U9/6M7xOXA1XwTaDG+bsDCaW5aKk7H5mqre6M
FuH5CiwEwyXiExOs67+MLf+0hQZWx21HBmFxhVkDxJ6WfTous7vzGqG44rEQ6SZsedP4c6eof0q8
mpYSaLWV4EQD8AvqrFAlxW+fjtz4AnPm/ftvFTbXUFJqyLzl+W0Pr39LR0aslajvdh8KKpPaU9bA
hm0m8QjVeCuJkqn7rjNIL9xYoEQPw3rSjSOOrubBvxkyBi2PwQuOmMI8Zv8CEzyOZSQC6apLYj4/
mK+Go3/JbBQRAmVrhCwHcFRT/QAqiY4iWVpZ1H/UPge/KlyhYVZPnJ8Omt2jr7NmVI6zwusD1kxG
OBrW0rn/2U1u7xKBGiKrIBC8DTWOdfwjCA2rKGSlUNbTqJ4msyjQCevTYBAOPK/XgtrBxTbaGCDx
+CgyrSHJTT7h80E83NwpOkBGPVx3DKykoNCWpGVSo7a7c79s80M7cbdht2N0/AZN+8HKr4UBZJFi
Sg009CpbxubolbfGKC/wlbSqV2xWnbFml8ZUoWIG/iLaZK//mLlKxRVXCWmi0xIAfgzZcQGdP8lZ
rSYfcUcU4g1MrVmDUgC/PPKNEJG27vmtOd4+56iwmtctuiX+3mDfBk+5YRBTCZyBNIJATPc5WPJD
aCzjEaGKSmec5LFqpkZkN7QajLeKekNGcQHxOC4W87/IF2NQMxhXE8cFz0W3nSjaRauDZ4H69mnJ
v1DKwOcKnPBFw05zkjfu+GU5PJcy2ZTe0+/DZ7Y5EqhH10LWnUOtZ4V4iNhDk/68B/peHyvHI/0N
/FPaE8OTWSTVgYcWCCY8hbBc9uIDhW3j2HA/iGi3CuOoMKbbNlS/CHdDQdeeOdG6uBteWfNfpPOC
SEqMH/nd4SjMtErEquE6gRfog/p6fwOpGkD4P8hetGbSl7uPZbaoxVepefLQX+sgQTwaPVm4xMlv
EwyR/nijOzAXyiYZRmqW84ZesJvT91bV82uhB4XdfcMq9h3WWHATw/42DSRCAjoE89FV1Zuc2tnn
nwsRdeWOmlDZx8LIWdYIXIX232n9e/vDfIgjfp7WawAFAB8Ir++jv2S19Q0PciRUCaCP3CfeUqRy
fwO7/OlZ0kMD1neNLWDGTS4CUB4lzNII7SsTK6IJIvFNaLOpkaXsQUPO0Yjp+0UM+rYqvtK/Uu3W
XF4Qcwknz3Uuds2CJeeoWjWGZSz49SB0JP1BmLVpNwDwDKjmm1F5XXzaEdzqyB9pjog3+VwtO65U
goda5D4HfH50C40mAf1EaZCYRb1E2iUwYtdr6UnbHfj5+TtRaLgfls3HWEOz1mRl7jIIF5IKZLgU
fxR4yQ3Fvb+1mNIpKUzOeEeCF4ZtU9ZUCAL/7GXrmJ8Hh1KCi+mjZOJy0S4A7h11PTfGhSWwC1dB
8fBSljma7sH7exsjkQ5Cu218lJ6Fh9isIkXtZ+BNQQWvxnTQ2Lf41gDW/K/QPim+M1VD+B31FbsU
YsDwUxzUNXocjnX8Ik/FV0805qhy3rc3gA/tDbCBz2tuGvRSlZaQ321ff6YLKvcgmUJ/nzlmfvWf
dA+RQlgYUIFERmquNfD8raxOWP40IElC7PmmdL1nMpNPIP2Oao8mGqeylahDNevzxV0psanpKn23
9S96S6ax/fxNAJhEi/CnILQ2UWYFnDMWZF87dGGenx8kONco1otrfQZkq6r9BCPTeH8nbL0lCCxM
OeuK5fcqOK0fl+mu5rD6ecGnELYnqUcWEo7FCirM23KYfvBkiTiKOqux2kFiSLi+5yj/0c+U2gLZ
JKwnbJJx/3U6v3ElrtKU+lALVjvK6tHnLSkEyhz+Vgqnmu0EBQL7Kxe50ci+Tk1FS0jQyZejDh8k
8Y+o8JuQGX2GycluolHhRWpdqJThNo+ZT0QOMtFAslEIIMhFqpsHO1u5/iah1/jU+BB+ZZJEti9W
39jroUHLNkT2Sm8DSNkrqhyNNGcNWoTMoMA8rzKEbGoY4adoMQiNmDNhv0c8bU3MvYNZnY1lTeHT
88mGpR9rUyYjwL/LDjoME2K7T5uRdYaZ+8sS1o3XQbuBuRD6Yl4sV/Laot8uFeG37PfHHyQzh7ZY
PMf0Sx1ZwDNUgZmI97ZRa1URyKAGIDGvm3B+d7wbyZZcZzFjTKGQwJfI80uUByW0qwTlaettJy+X
iOnCvB3a3SpcwkAAPW1pGs4gJEb6hldYB/JP1/mZL+GWBTy2VLFYjy7QigkDP94HFXlp08vUEz6n
YESI2r0dvpPyUwvsvxQtoxgeTTrEsPvzTxbH3MCCyWftB8L0ImkOlPDEnihJ/LEFMRKYqwWhqq+7
CuLn8cOt06VEhUK9+iaUyH2Ry1TL9ol5VDM9/lRn3Wt9vkqnS6/RmzUDIofxgcp2ciOL+rrnkXM8
SYBUWJwjnO/yAEbvN/Fw2h2LvXP/3Km5MYr+EM3Utj80MCpJkGEp+cg2wrcrX3K/lKUwIB73g2ZW
7UgJmmjRW1Ga6QFFSKohP5MZAEL9lkDaIsNjUHMYypVKlvTO9Re7y2GNKpDD45czc6kQqDzyVeOS
/qFhgSqJKKbiki4QsHHr2BwU7xuwoyqgVkAxmOVarjzyNZYEi0nyYCSkuLd0/toU3XTaKH6hmGeO
T0M4v2fVppAQD9sibRqcudqQmqH5XVvmB4MqbWDT0H1SWe8gmajHLKuRpFvA/P0xrPVe9a5U3mmo
6FlzvuQ0crMAR4TwupPVBzdNDwDG3Jaz5OeqRvYFjTsdinI6dK1a3iuLpV+M4gRf9dPFDY0m/A65
wFjh2H/ttwwYebr8QKJroi+8I62ifyVPnjMYuGkVQaC7zYjHbCmAysnuKHyTsaD/FZMlinOH3CAN
HKsbKWgC7Nu++A0TGhkh/xHAprErWjoFiZ3f+Sfu5JR44CdCWZeQvmXv4tjFuT3BUrp4Bmbb8+F8
yebQobqWUkX19o52BW3Tbf4jeXAl866YTqxaxQLDzwruG/hNaJvXegqjU295+HBbLYsqKMz9cYc9
lIM421Rzf9I6PbbyKvJ/IQc+J+sVFGlNujCYrWK9jSzXS4Pd+falhxQK7eAodZS8f+VRS7HoDWW6
KGEpxTM1o347sCxpVffgKIuDXczLL7FbFjI+CztqMakHOEwJja9soahRcNEZyUFg+Hj2LsY2YdWq
KQhMOPwTf4AS3gIDBXZKPc2RLZIuw8z/1VZ485/yF5mbuU3khVn3tcBDBD1NqYqLW2ktIHeeSR9A
jvfE/xVX2TQXns39cTbHIsY5p5c2odyJDi0zZaft9AQ9cAaVqYVCbntyC4xUpRgbG8AU9Pspj9l5
Brv8VncXcZjdY4491/ECdmwPB1D6QG44M9kJ1ySE3EoauQQIKOd/ETfnluywta/vK6wCmZPrd/o/
8F2QUlTWR4gIeC85zWfJ7hxk6j7dyrbDEICgy9+9NL0lgSn3j0q6MDlNT7t17b+bGX1mZkHchQVw
bEPknLEFjQzvbyRywsQwwDebI2B012UgmmvMM+YV4sQslZtNgc8ivbYfuhYjXGV0S9pZvphzWD61
5KmR36ILcwc+7vyLWJ1Ya+FNWSbWVtym8lVNg2HcObJhFNnnYcXZbT80pY8uBY7siJ5E+KbmCcgY
nCUYxy8YLE0zhkz8HTOKvqshwmKkEMC+prg63RVsO/ZujEfE8CesZ9Ta9IhXxckQxzMfGNCXT3vr
YLEBiztSiNoIj2E8neZGyrDBYrFUY+J43RbNm87mlfPTmD7n76AN7K/gzbNil2WW0T0CllGlZb87
MyMGaNdjyImXIvpwYh9PN0X6hf4KYUUeoHdEhIF12di9owxOBMPClnyaTGDoILazlousgeviYua9
muaTclUSW1JtTdXOzDxuSmmZ+Mp+NYW6i96I6yvXrDjCsrJJ95nuWLxFFHxkwkQyKSwMpm0Qplhl
mUtKHD5ki5AluKbWBgqSS3zCE+CGbvzd+FF8UWv6g9hMuz6mXv49Iq6jhjgOP9rTqEVMAD+zOnMc
o7bUuCtIFMUoDNaSwUp7K5nxlTZTTipCTZIAYz9dIlUeiuoLzVpdjtBAd+rAjCv8v7eyeGkQc6Az
RPIrsAoIdzFnT1lb9bYB0XmJHUEFVF89jCruVIFLvMRcBHBP/My/fqEfeDPDfLaMCCWuBlhcAsxC
8xMKUBIxSOw0A7rHkBHXjiXr25r/nWVf8EvrjdPvXXZgWO5AkKtXSa1hHlrc3rpYjZXCZBt4cc5H
gtD7939rohWKrgHm17JalN79fPFegQZzpKohsH2E1JIMWxUBJljeAcRTSw1m+3fHwO6pfXm0IdOA
MRvHC5/WWzd1Dgq2yDASUNW2ZzatmrwbxsUH/D44sVPBwCFGly5lsT5GxPeFEwA6O1YSdNXs497z
EXUEsWQM4yJQja/+dToMCNgvbMqmc8NkOfOR2chn1g1FA36rhubYhraPfoCxZ1ak5IJJ35mGnSFx
cHiPUzaDWNwxXGKRzRR4ysDy3PeVe1EpJ+EPZcVJHBptKrCDbZnHnKPgJSQrmsbHQjdN5WqcFzhj
qvSoKWHEatnVkzp4go+GQuChF6qYIFM1h9MC9N5vI6fBhbRsKS4gnPJcye91dMe9pa/wdRgC3FHp
9i05Gn+04C+4+a85SZyXGdKss7fZ1UkuxsPo3ArRMbQY1yjH3q/wamOK+VEGUdWqsSG4tMeJwoGQ
6tmZH9m8geX/nxo//OSQ9JnLyV5Z4Tw0Rk9Y5CPyssdfqmhyyJlGKeBykeHs0vZg7BMSz/Y6KU3d
kQRWYZvE8yC8KjBQRcFu8sMaYWBi+LWXCOeM9PK8ObOZFx7+LZiqCRlvktFXfNIhQTRwvJOHD/9G
PLF35ukJ1mgjYw9K5hj2rVQodOT3/APvW2Q+KO8i/R2Q0iDUKEpvlNMdvuhWhqKLtkYXVT03QxRz
BomMvLOWUsBq3ppOQ2nAyzOor5PskngdF3XnJsLTszjv3Ykpyd0MSUpNmbuyIDI3lTNEEtYFIyCf
hEzUUQrnuTAYmsvq+UmY0pj80Byi8INWusGbJDu72Z6TQsqiN3UKnQmD0uycB1jxlgRqcYM8BNzC
PE2H+tlb+1W4seoYtON0YuNMAIUDyVzBYqO39wic8w9nuZ/h29hlVage4ZsqyYkrRXffTJXaBV9w
9XzTZbBzBj5GfHbggkxjLkRrEBJkPVhc395WJs4EJrN3BVtvXfgvmtaoL416AJztg8sd6ND2kXsm
z1E8W05V79TGrFZEidLOWsA9yTxjgVlCIRc19JenT76WT5WPClUjlV8u4GQC3QApliAmLEKl1Qpz
vYb7Y81BXahnP0LCiRG+7cC/id9XvXLszvJVdSdeGJeOim7WgteqyPUfoYNlCX47ihYUgPfki6W5
FHm+tLNMe6RM0Aj3MRhLo3bS40ggwWTPnMkUo8QvFAGjO+22hF3UkzoJp/zbcTb7KndafejzQEpM
7R/xiiR27nW4jixSNdpq8PL84jisfbHjDXpuvyeiRjmFOdQhergxidN6EE5B4tlE8u3LPuE/XN+v
XGKKXp30465dvS19izkciD/5vA5vig/gSgcyP6HAop0oSlFWXJP85Odai67GqtsE6fv4J2cbytW+
1sOh/5jAKecshuoGhuDlQ56bTacQbQ+hZh3VAYKEGbPgYUvpLRTOuaWnL3bwnRiKEBwwsj2NiuGc
G8A21jUlJ+ZCWc7jA6rQRY+9DLlDt32mwbrpSPieDuZ8mu9wrSflMyCIep19JmoeVVOfR3T7og6F
b5jpUBzXNtE2EGc7L2TOC1ZeM8g/yDVpe12Ds3CBNXdUBeHYCJIgeDMoviJ2NKcYCYq1GPUhI4el
y4m6Fq6w+7V8Swhnf7fuNwudrPnTi1Gf0pOTEp8SxQYFAKIIcFAhetm4nKij4W875CsgN4vwrf8h
aO7aRolnonwfFJuDyc9I8CNyuNgdMO/xhCXuzdoMsEgKLroDKdbtTyguT5iexIgsjLBbQidu0jCq
uyW9BWeRbww/gBpBFid5992G+cFDXMPVILId/7R1Nn4xJQtU8jBaKMm5V/zrLJy8RymDaudTxmcQ
KEPBD6RyiAWWVsH9y+B93U/OMR2tzkPTV+m3AVyVIKH0iD3Vg5jMvM1ha8iglcsVKJqapnM7LflJ
KqWzPeUNxRkhzC/tjaFMbIejeBLtZoqzxfcqKGbXdSpFHyl+wfV0FiPKMVImgyTFVmLLRnhPUcL4
AzrWOybtz/MGNDie5Mx/HGrz/lhyZSq4gYW0jdPXMjF+V49zSygpsQw9IL6m+DfH/LcJpG05egcN
V/d7ho2MTI/ZhHjHZs7LhIQd/i996m8moUJICGFjwxrlyxgmIRPPjb73R7YHyq+oPu+J61ZXy+ti
Df9O+OKP3rGacEsXfX6RlkKbAHXT2cA8nPL3E1YcGrB8ku62AReEv/JSgkNj5KWpoSeOiE7naHtU
eIZ9K9vEsQsg9GmXI0T7ylBnCqQ2tHZjxPkTRxSrwpieWa12uB9FjwjdfcmmY0eEW6vGFa3rnMUx
D54rtEK+1k/lQVsobHOLv+9OSng3DrcIOR0MayPVrH6j6Ib3BigcMTR7q6FdftXpIvO/CkHYnND1
5mGUBWu96rmYZ8DmPrfFV28ubVagKA1ocQqQeodkL1uiWzZtaSZGSCkDUpx1Tb/rdVb5ccGqdjVD
9JNYtzsusAFTZYhmzf+98SbOOaXJ/jEpIGjyJutdBTAdsBedSVhaI/NHq61vWwHHUF+s3oAYHV6M
J/UbYRU/z5tEk6dmpqkpNMmjsS8zEg3slQV5beAR75pOWLvG8+B/9L3l/cjSmN1Q1sGLbVuY7l9I
cNdzGY2zdSwdWyybDVyUOcm4t3MfUrrvtDSWjHNpm58Pej02Wz3Iex+URU8StsBVmcotmjzkyorx
rDjrRkafUeSjhQ5Cst6KHMgncpfnEev7lVPB8ZKUwW8qiaC0yYz3SR4XV1cRYzUvkL1QU5hWCUkH
ZnyO9l5bAnRy9zZcM+JaE2d7D1hsBIQn/lytGULG5/QSp4+Bb1DxGL5uCkqgoCNezCcYDh3K+96m
1U2GxuRM3sSS55N+s4/ojvoiUl8wjo06y+Pk/IvCA0oUZgv0ldlaq2RbJMnTqg6UIi/XcnGPA7IO
ai+8hJR9Odd41bY7Y9QxOLxdm1y9cA06tnOjik+Sx716UfYNTiZJCm4fMJXOBgb4PSAnKzO8Pu2S
fH/wQNIQR2UhWvLsKzCTBGMZOxe3lSPVIKDx5vt2rxZ8fjhvvmRc/sYx6RlxmFdPekM8O2XCiq1U
JTljf4/P1n+rQj/n7esza/JZfgzl2gDs1TOBOuatNOxjjJhhL4O+DeKeMonQLZLC9/Yls+L6MmoR
huW+C3IFOy31sWHGlWFeH5KMdvj5X3qYDP3GZe/fwhojoLIYow42IjkqAQ2OvislSxARlmVDCdmz
ddNk65lCc34dUeqmPKM3TabwH0oBQExEQStPM8Cb+s0/g5cAi88h0Br00oAPmjafaaoOj2kpgIw4
K49jM6dsGAoOo73cxZwMKiRhgq0bqKzs1JvxBUZF/JLu1GZnoaDjT6uWXnWpWVOJbwjr2s/7NVsA
JNjeAusAhzQS1gCSTQNYclY22BVr3cmR9ZwpaeBDzUW4goMXLYu7cHGWWQwooKbhiJcbMUhe04sX
ke/CoqUVjWHqkuD1S6Hbe3xVG5kLKsJ9ajGmStzfNJeKB/6fX0x00BxoAKDZqT9ymb5PVRI6QpJ2
RzjIWF8dyz6NTuxTO1z+bqj6oVpulCql7dymkmJLxb7oxSSzYjX8QucQkSMhbfScmNomGv0pPdg4
a01VVmvf3gHpf1borjBtP48S2Y4/JpJRV36LznqNRKOEA+YcTBjEekiffkM76ziO4f7lYq5pWZKB
umWK5L9gNulqDZyfG4eYrMBpC5RF/wLL5xy2kjnGlbAvuEOgQrKYlwPEYwjBsFaaUADBPp1p19+O
Hb8484QK+nDlUvsAHbMnAt/z/5mjpR3OICZHL6MpS6ZrBQbHLRC1rIL5THDeDoWln7cF8TsUOl+n
uQ9yTNibQPEtmYbcBfwRsB+zCcvEWqV8bpclagCpweRhTXqaannMO46lvmEtLfrEKIQPGcCppJiA
RX+Z6CnT7JvDO+EvDFz5D2GlknnjUgByZPPMZp/SiYSLgKhNXNQ4Tm+7sSCEyWVB7VUhVz/+8F6t
PeJ9+AOyAfXdFW0UXWcjvsdxXSUPkLgKnUIXT956f4muWH81DHDYg4J8kprhmSNK5+T/g5kFuIan
b6AYVRl8isBH6bo12sXeTQikgQES1F0YVmOgFZjJQcSTfW6FHz7DUt7AdhVUxcY3N+KqMCYB352J
dHsDU6hBU0YSTws1y67voATleGBRkFvSlSMpIn9I+dXXwtT/8UXhhS13mqVujmNnC/58SR4RR1st
sowDqLMvvdXUt9XUzUA19xZPTVm2XW943dFocKXULpN02V7O8fw9y4Pz1Yg/lIC+L0zTUAe9fZpJ
2U/H7/h7S1+YtklDNco49+fQhCL+G2hkjtpwo6/SU3TfC9EbRyA2+WCngkw9s29ChGEX2yQclpMP
HFZFJXLfejwiSqOxhjX6oYnW0vjjnJRJYbKbavcljPZ7o3U67o6rVWcBZcqXYBhUcKw0zuA8hOFz
/n3zlZetLyaMiGrrjv+pHKSdUrLIzKE8ZwMQU95VMn5mbOaRNEBVO1e44YjzogRuxX8KbDiMDgu+
wuXhPVA6j5RCMpmdVPpOBfFAXDp44j/gcQKYancI2qOCJfOpY6HZGdHab5RtjOnuhRmUqcLj4a0Y
/eeLReV5r6W2PZrH6Vuz5HNx4jt9qj3O+45aZ+7kgg4kFN3XUBr0mZafWlXfitPcZVM72EHs1YaN
SvmYWL5113k/4bVtEqCChLSe1tGGgFLaMxVJgbTUJeupPqi0JdAyLOqMws0VrSfqe/eWRYpzyryb
m/XLVqqjkJTjyvD44R6riKgD1aeJDMHodvBCCvhR7F8ap6vH4PXOyOhPOKEI5GqLNDgw7uYmfewA
gCwRAcjLBEP4e0iqORVGNqUTz4DEVT6QLXJoDmOcO/hIONdmLLWTfltjlagahcMzPFpAPUl68viF
zf8HMsvrgG1pBhZIdkG527JhCKztFC3+BbLQcuEvmZmmPoxgDfCItBFxAqWRrCvgHaDhCjimgGt+
2Twn6LPuu8bYWUxnK3ZDDcTXx48aaIbcGaWEMcjFaw1AtVyVirJXu97StntGYVueRpTROKTCoIc7
F8AHHAUSkajziARZHLvR2/JHLWFbC6VFYOzKaW11W6lMMgOz8sFRAiBtFZ3K09ebOat4aqIFishn
Yy2UMxoCR1XE2rTFPVh6zpK1MT9+lZDqGjjp5PgBpUA61BFMISG1ysNsLl0rM1rETwcs8BlMXQqs
MloSIjGsUJ4r1C0RjH1q0WmVVQ7X5230CEN/XSnbmOBAIJOwS1YioaCpeuGPAvflL1fdNsb5u0f6
AgKaL0M1ztb9fI8gGcyrEs0UYKLVfCReAjaDHJW8OkfsjVsR4Fws+3BXFNHLKBjASgYg3DKl/exP
LhderMYuzSrkJQwsi8NJU8dJzi3uTWlNoiox+ptdRFgwLQ2p+HFUYoM1BKHfZWJ8Kly548p1l3s+
ZkQCUmiKWogJxFIUmOYUjNvdPKYrVOilKSCr3tLjDpAZ4XqzuNzm8KpK8tHjoiCjF+Gnr8aoqrwa
eRbkZajTWA2v0soOhNpOPzegLZb3mLOtGFSa3amDENn71XeC8hYnhegTbIB6lwXFmno7iy/YPMfA
YIL4YlmFcmK5ujgUFnsUlcKpaIYTwr3BUJSy1rMpiIyTyIbKpIXzkT4G9E7NI7uRne/bpKKtOe6c
XG13jFivU5bAoFJqJVfGVzOJO9rx5off8OxCWtCln6hzMMh/EykCU7Fcl1k3WdQWHoxcml8yx/2M
BNUc8r50ZOPIE+oOkjVHcpztT3hWfvig7auZd9gOQ6BWWjnEgNOyrDUbnkLjbwgIlo2JtWKYLckk
1PEeK48P9em+2wCA6Eoa0NfJAYSFl1ockJzQImmfA8A0zFmKGwcw06FbhOTVkjdOWdo/CQoQfv0w
ajN75vnTUjMB5e3Y+I4CodoTIZg8Y2V4Y6pLKNsap8kPj0+5eijUJNfjwICeBgfqnoi8Tu4V/nej
iaEM/YpeMrbkD+cLcJ1HM2a7XNRIkb45uFaQsNKEZ8GiSnQoj61BgwpJ4UTTCQCJxoU1nfK8cgM2
7I6MrELYLSkd/VOBdCAl14TWVn1ZsuC7/otx6yxirXlGzk9EbSevzOQw+YUfXaQQrY8OkmWJa6P8
ZwZmcJH5/75PlgTs8Wsqz5FmVvr4/vXjyXctNUJgXYc0E+cbtB83Wo6tOGFhDsdcqhm1/yGGdr2O
7kNlW/ybBEChfwx2JtEJUC0ygSkuaT6N3A+gAO5xNeu7UDnOigRJh4Jtyb+ztnRrVs914YbuQys8
esBO5pmSpzj/y3t9e6ogfhCAikDv977dimrdV5awZBa55p8GDY0i+2LKDoO3vLPiMg6HIEik8HQx
tIJCta6tTRqPzvBnTm6FAzRKEtWmhMK+fFo5dElT/Q/SqegSGh3E77XPBxRvduYS1MBtNk1OsA+r
DsEzXkAaj06HJ7zEZ1c/sqA8/5Q8rysHZGjbTkzQo/c1kxkggHtqajFKQEDj9DGQhY380UEzpX6i
6jTkpFiUcNTlLavgjuuGktd4uaRU4WZOxoh+svrN15nVSGEslH+ayQqAgp81h6mLDSVwUotcXjIP
SQDMyTyNRfV8FzGcXkIyMOs1UA2M6aiDgmu9zdc4BubJ09w8pnInCp8flqoNPYrdnSo6gsS9E7jW
/eepIwTXYAYckm0XzoAaXJD+fRISmhj0qewZ0itDd4rbNUdJ8S/j5ViZTUW8FY5tdJ2nCsM2KmJp
NGHeunfj8a8htUnCwY3VRsiX+4rKSuwT5kP/Evp2fwj9HBWFJdtu5LvJwe1gqdI8/BVCMGrjkagv
paaPHbuj9xBI5NemXdCZi7LPMMiD0b0gN/zSU+nMOd5KyNTLyPkj4c8VCvpbLfrn2C+X+LsJBzcq
XcIGy+bn673TerSySQ/NopN70OWeIzIy5qki81Ij0oE84hx048j4/P5kNUKis5BbO7018wJDm9T2
s0+dnXO0bpGO+Qwu1ZaEjyzlYeiEDfysR/I/f1qV2RHOOcQVl7R5U69JFW3EZTbect6WLfc7Qg7L
NHjmLZA7EiJayEIiOarTOFkqBq9fW6dFR69+7Req55ZRGKivYSh1+Gb6rX7BRpL7ZbvbyjzDXkWN
f3wGAhHSXUXDLQljxM/7G5bNNydC8CknV1dRD/hg3NoJjds75J3DJVbZNM4xNJTmpCzWPaN0xuZW
Jo6UI3/0B6XIBrCi3G1n/fGbVbY0vSRA19LDx1PAWPn9TbFn6MmG8OyhWIWHB6SRDNNPBJueDzMo
69PV59Nz6j0vm1C32/Yh0r3n+qAMFfOPg/keyX0CNa9C4kXaCpqRLbhwGyAohoARtG8b5gX/IBKx
ZyO/KQRFfXz1FiNZNvRQU0xXfM/bAgOLn/8lKHupvhbvzsJaaAY3Ow0JjJ4fjCuYEw5bhllHrBl0
HhMGzkn+xHe2W6eLQ7O08PK+T6W6JQtr+JVnpnXA9fFFoScoKPFRdKQ7E2Mhl1qeICsKwZ1f6RkG
yFmMnrf66PikY6YO7ogXhsOhGDS6DN9ZxoBjlZYleb1m3EmrKHWy+crFGuU4GwgQNavErm7HXcPp
Uf5sJ0+urB5n9uEyz+inB5Sy8ZKvndhy5sX/JabGdBuQUPOIiuzMr0tth11S/5BSW+xaNLfonKq0
0KdcPo+vKIlUHUBGq+wCu5j80lFPk3+49EajpDJgGpcsvvC/hHJQywg1y1erj/HGFaBprxnzy5Cq
aGh/IXb5Dx8MivHcJB7fiH9/wpDb1bk6jsNH3Y503FESJe4LWwUPC2hyOP7xwXvbvjF+8/Nu3axm
71A511f7nPSLxyPlwq/KD/VrfD8esbyCDRnlgphlWAQc4xDrHOkmwmhH5DTQm1SG+FcA8QxnXEj9
yDnSvU8slpRzSOZ35MKG05uStQ73y7m02ttg4m60GWfpZGIMVS1mwFYCybV+G7dCdEKe1iQJUj1+
Z1hjp7LbfiVgF1VRqhY4DYaBmWZ2keuLFQYA6j3HUVpPhIHhDK1aFvnu+tz0CZ7HYTfc/mN320Gi
p+obZMNT2abJ1Y1wtusTSJULn0G5/p5KteVkZzOlhg4M6uegbT3ph2QAJhJU0GwgsPS2upXFiw96
v7/63XN4q7i/XOqo+K9TQsoVzMvFZsRHGXy3XxRKrxJlXFv1g0qbZ8/DQPdvaG2OsHj4WujOAm5W
+wLpfUuQTmUxzx9uxQHYigLFI7giJY77K2KhbNVyr3/wnVY7a7de9xT03Jk0z/UkGXoGfntNbluR
ojgT3OS+9hUeftOS4jh7gtsk+YpXyXud34iHI5qzdgkZwX4Uo+OX0q7q7BAH4OIsxYzpGZS4ssWY
wsExyjqsPc+ZCgIOopaavwQkhzof7eb+k4a7MhrYQ1+Whn5u1PXJbLxplxktEIMXhhSTeyORTFVT
hqAep2HojT0woBLve1j4dbeVYbrHO+mS3fjwywiq1W4zYELBTwGt3WtFQVSvOl/3F/V75QKxgXY3
DMoWKCCX3hFD5J0DUxoegAfVD5NQ8sPGPsL/ei2WrOp+AO4EirKHBTT6lPf2K50W0mzjYpLLz8KN
/O0J6okk5GM2HRMi5sho26ofT2fRpgX2Xe/qgbWHCao8tZUKhq3BQryq9h5rtAd4SOAzoThH9yI5
VEr1g22uV9RRMBzsep/DCnjDQaa/7e5RDg/xfHWOMOYXP41Hv0fK0hfRrI8vxxk4ua0LgKMKa4u5
hJq2ZTy13bCgIN9Wy1al3uBvgVIw3F/9FShzQMn1nLCTSTrieh2rG6MeygBKa8gcxGy6yDjFHPkF
oWjn7lrBZoUo+wvfDFg60cXrmRKzMgs1h/SZo2hIm2ICYGmSwxrVJVtgTp0uuwbJWcnr+dpyhGW0
Tktn8x4DFySyEv/3fidqgbTgvsou2jBdlaaBTslAXg+cVK2gwQntI3wM08unY7jVpsUqitW7DR/H
eNYjipcAH/XVGkx8RWhV2mwnVLfLBEJ4bWlEpceCJdXn2JN/cbWXS3E7/4Z2oqJj7NbRG7OrOELa
ORIBDSIexAr8oGDqH1MU27KE2lDqodZqDoXS9gKaWekyamXQyzcKYPlW+1Kzan5hQo72El8GX8z+
rRPfHp0XxBlJdI6QMciwhtIUWnf80csxdJF+XzO4gdpYoNF9zjM4f+HrW8ywPJA/yoG1Tob6BleO
7x9bclNSJg8V3EkCma+MQkNwggvI/7ipv4PFj9ljmVxblETgsAhfyQoajF7vcxtMkGO6Iv6hI8W9
eX2NYWHpwPO0iA3P7KuJS+jAlMAYkNiQ0/NRYH/qhGbTHQx6rsXRBitrIzAeNgx3fX/WUMAdLyNu
c9sLElU8JT34CE2gMRKcyKTCJHdC3J1fyPemMZCVruEISWJY4DCjqcn5FJkFSvX3NLeC6WlKN4VM
c8jgujsh3x8rXqT3pIoMeLcBTZDR/svc4EH/lWGafKjBMij8s3evV4gCqBQkVobEFcvbL6DlLjo5
vKmRX3/IxsNcnBb7ZcO8jaZ9uxaYJQJjSMFidxqjnq6/Pf7KDfs6ej3EqVeyUfzHUFOjjpPxT+PG
pLaTS+hWg0Q6hv4iRkFwMIhQt7vtlCSZvY9ETryDx9v1Blr39XNn9+gfyqe3sO3QoXYoMRj9ZhqY
kM4evpolpDY1jyRlr1apsQ78En6B/VT2In4T7nVl/vCsB91j6cYPbsrPsrj6exF8TCv4/XtUy6tG
x3M0XRclTcdiiOYeZbHM6s6C1sSjNbkLix/lJvHzZWw90CkS1GDzThGIKK7utUi4pkoi1GqvugqI
UeXoU5I1y5o9hGxeDuyJiv1cEXgLlVHRn+SfQb+476BHR6z+T9sPv9vfvDnJLURats7kfILOBJ50
7zF6WTBEvM7cSIPDbB74fxYr91oiL8L6TmTnPqXGUZ1XjPHE/IGEbuyMs1KopArF1iy/h54uXBfJ
Mh6owehhv/LJdT3W2QbV6cQMd1gnjXCejfIWYwP614dRlr5KNqIho+T55pV4JBuToNSuXJSLwH0V
tkFLmGg2lTeonOv1dkuiBN6/iL/TsSDRL2wgpzIC4i5wdKf/H5oEb4sz9wy/uwcGR6NoVBoa1xCf
24nXQsycSq1yC6kMOrLq3ReXN46STp/ep2hGhbyH+bUkOMzSQHkm12zr0zkAmNlmL8MUVeVyaWxo
3CYHPXAycD/h/q78V3ZuN058PLbXVav1zTLcrvuP+98lCcAM9cPthA76ANCsgSIOEtExeHTW0YP8
2VmUuW1WP0gVoj8OA70xe5z5eoBf7GGKv2ozh2mZ7d4zDbDbRDIeV6L1mzBEB+aWWM9bQUSZFWUn
WXIQHqEtDm2INPnlmaxcm7viyb3rysNPBY/DDGQSLQqzpJAxdRdOrOID7JixUAmB7PYa2JkdB3T1
hDhpDOjuAqGE5DkzN+Vx6VhOaQLXMLHB2cXns0a+AQ8E8HPdiFZKF1p17mVNZFPtJ/CY48iVa5TS
nskSRRfjiKhTjPGYmc1I8X1hvAMRUH9BS/1I41lGfpstpR2NqRJdaCoLHfDds6tfW0bmHfyijOwM
6Dxh8fNLsYSscO2sMtquS5Zf1lHGXUP5DAlaaaSZBDo+DG+kyjBc4j9KoojvajA6cmwGVgJoACUP
79bLBSkNk8dbWp/YcKo1YhjDMJbE/WPAmDV/sCPS8lpyymwRxjRjkxDrLy7p0qj8pIFeHWKBABQU
FDNTyhzhx+7vXQlgEPEqmT5KHOz/3yXbM/q5s/PKjPg3IGVCMnwIWX82dR6bBE2RqQ3w6sGviWRU
erOllSpPBX0Hfs/Zdatlr9qAGwZbWvw27eNYqEI5dRXMmWW+rXx9KKQ2VDEchwkbO4VwRe6ZyP1q
Hk2fiMFQWy73PWUkXb3nuUkv9wLn/sc81imbXbiuZeCUpgO/kVnrxzRXCb8njJV0DzWkzJAHG9eH
KOyVQ8w2YRwWVQZ7J7ipUAVSdMNTCtnBE4r+nUORjWVdrp2ZPD/jStrbVh73r4VdCuVZ4lWP9491
k3gSbOVV+C5VU5o9QvUZvLI4upL8m8HgHTE8EreBfs5UEX1TSqYCTZ0UCk4VIyHkbhinMCuHyC04
1NKCu/rSdrDxuPD3XH+ES7OJp1XvQ+XtT+8v5LiaSTQI7XlcbT2IrJ8AO32A748hatxhwM/U5X1y
6YLAAebnulj3Yg0+wATSsLZhGeTucUc7FsZqNKIxs2YdPUcjraa1BawJIpaevRegID6vyZ2+2i0Q
J5+1/J3Pnb4JGtqlUag8Vkp2TZRYI/8VGSljGYLdunonsr21QtfS8zIJoszUueNRQdZSOAluXlj4
fMTMijT2yo5Vvo2bChNkQDau1sLt2cVL9VsogC3riFYfYpAhcYBUZnYrOY4A49+/2l7EQPQkXtiX
t/v4R9+9afieNhm4X95raLSTUELm5iWFghX4KWz3H2Iw8y2U2zuZOItvQOeiLVtVGGM4amy4uM67
f+Bg+FavEhXp/Y/JZMAYhy0a5nY84cZQp4S0QmZzM1U1KxaZxWmpLOBJMuzU13G6m70h1TIA8RIF
KEujY7xcm4OYW8tDl6qWv/bdXB0pYD6IqX7SBsHN2itXQheJsiT4X8k79bHHyQ4676FPmTQAEU4T
c4cDc/eyEt+F6ApqD+7U+Arc44JtJePU/rb5Rn7nQv8soTyQM/KYF9tv3MrPMTIYFYDclfVlvLFW
ASEtmLKa2tHFDZal26UA0O3bZH7pvrEr00Wz0+je5Ug/RRf6LrGo8y7jKZkgUAYYpeV8gLxoeK4l
sKJBFGesvo/N2BH5fRbYqgwJucx4EmKpO0nvwJqVb52TzNGun2EiTaAzpXIjDXQ3vsv15O9jPYcO
/ZNLBwFaYnVH057o0uodMFu4sxaWUy0RWYYms6W+X1mOr00aCGHv7csQ9ysGWHvbl9xTmAM0rHCP
WnkIcBQykrOczZlEmUZEBA+kQ68qn9WcVyjNjLnGUcU1qO6ZKI3p/IbXJCjErbFqvmS4rYf6cUJB
2SfGC/avQB/euQt8WoXijfE5iRDjHwjHOyfM9YiTymmhQ7P2JRFfziaEFd8MNLAmZ6eaULErbwHN
FfVaSirNLpA1iIbyRbkQBYUUq+gzxDxIPBieRfU7EMXAX9oGOsneZyV6Z8+YNKyVBYJ54+VYSHX3
i3lAAFWmzp+VTarRDKBXhkCBK4Mir4lBtn7ARynzoJb1qYX8VxEV/veH8c6szPqR+syJ80m42yQq
12io0uZ+NmBFlbpfFsAtHIUY24iW0utM/H8VWbQupPMn+/jEx1mtfkxSIv9Tffj10Un1g5kTWDGS
dSjIxX3wff0a8j0PWBOoKZkcltkKpeRPfFBZWtemOpJE8VHOtyaEWqJJNhyjb1igRS6V3xo1QOXe
AjM1JqmYWupd7GPfV4NKfpEuWoOWJfDjIqAKCf5ICdqxYVeXRsIku+LKEqrhxgUCwBSUwAXUt8vX
Nq1WFg9zPBSAB4d2jxjswHtNDP4Bgtakm3Ix8Fa6vU85HhbMOmKrEWkWaz6kC05/Mgo7BS2mcaAU
ctbkPyiS/Lv98wyH/xRTorFPlphMd8BIHXZYLGxp4wrGvQ7QxHuBAshC564Kqlj1dhF/8AHDper7
FjhjAHwEUtML9QVvgmXxzvayitVuIHNou1EAV4Xam0tl6TrIxQ2KSSxr2VNZ5GMC8jgg21jtH1DL
mCKsTvCrSNOF9UHeOwKSMSStVjTflJ6Bks7iMK+Lr8fpabx3S574d/x+uHTbT72zGUk3b/hWyBZU
q9Y/iomks71wpIJ4irjsVFepNeXBmvwX+QiPWAAzsLMoljqs3ZgEJpv2/l7nDY9VCsEgWqi+ovYs
o530Un5BAqYeRMZ+b9wPaS+zzo1O/VTsktyvasLtvGomRj+byWZNZvQtJm8U8OFjq+rAyp0RyQu0
zL5SUpjJ5ezKPTewUQt89BkU6kmcH29SBILHCFgLREj/MafQkX2ER0Ecbq8q1gjSWitLyfDscMdW
yMdtQ8MKUYNmgDjs/kQM+yPq4xa82uUfwhJseLqBE+YhvQlVgG45PngiEVRWHG6iatxce1cX3WvY
I1HDPANmJYY+EDGkJFLdVfcOOzhL1N6Hn7/PimmDcONiGa3a9zM+biKZHkiUNXUU0Csn17opPzde
+roTPzwBl4YSloZFEA4u7PsqoOrRCgUa+MY+Zp/LBWJ6S2NbdSKA8LbG0H9PQpwJfcqOupIO1Nw5
aEG19VYLHa/SHGSUAKak+wla+NvwcqpHSkmX4Api200eSzjy7hVvn52QknDPVfkc3SPd6hb3bu1V
b2/8TN1TdrKmKPv7cr/WQK0HSR9DiyJWKjNTGieuJGQGqfAHOuTQMsKVPGKNDVdJSA/FE6KvnEPg
KMx5Z1LtCE3329XjMlp417Y3BNmTljm3vulsp+e4ToprTmxN87ksNHFE+I6s0da1kXdtx9ggbusk
t1y1RAtM0RBEa54DY3tZ2vO4PM4hN9OrJ7na8EU5y5Wh6bZn90ncHjV4pWD1B+zfFHfikqmhBVAD
LXiGMPCnZX+rJnoQ57tGAneUw+ackdC20Z/qXs44gqqQ8/V3/CyFS55JnYMAlI1NcNk0BeWisy8E
xIDbPUpZHIwogxdPJwj/HWurJSiL96ymVjCHg/wvm1nepTqJNyfTFZ7J3LKe7Rxau88VtPdWYJ35
bvbL7Ao5OP1rPkpUZh/Pj07IsnK+Im/8vk6lysDRxkUXaieC7XAjFNOpPkxgRqFvaw2hHyBcv6QE
SfsGRaIlx/KdsE37q94Oj5NsSO8MHLTc4ziLIDIusV6+BUpdMfs8v5+ri9iKmpGbJrQUOxIh5BLK
iuDW//tW7ljmI1rZv/364co5MkCgNiQHUkKFQwCMcX/fs0xldwFldmpdGCya9pNYnoAJy/R8LD1j
THsBZugZM7Bxm7hFIe/WHqKvjPKDu87p3G+pXlqZM26dxHKrSHGq0SZBqHsIrdxx/3qBSJyUXOKg
tdr3cj/XLGUs+VJnfI8ykorY6zungco4LsFSAMfF1jmbfRAWzQT5tkpMS32XdyEM3TDPYzubnizG
X9t5NaiZ1dKci8sjTgN9TJRwlRbkzIXK0ahVO1Vp4A1OY/n/Niyhnbh4aEgBINqXpM5E54vWzzI7
SuRXGnnyqXw37tQFWT5D2FLdB8DeRCWHdSHpFRT/LofI2/MHOe54D/r+4+FPED/7TmRVU5wxxXuC
IJVNeIJw3Br31MGfrJ5YRqrb8nvevytynfLyyQtApT3OW4rOGpPbwi8YHGBsTZF8JokD6VV/JxOF
4JVVYE83SlpQBqxmzq8oyWm16LzH0thGmrtGQM0TOGWhb3NKAmjC/IEuS4NxfUsLydeomW1D+TLO
6kE8Al20Dl7vd9dNoJ07L8cXlewm76ARm08xfGc39VNCVCIYVY5Qa5+VwwP74kkF7B1mPm/NuiW3
QYq3yo//7wUPQJCPq5Gu8/g+4h/P9HRYSEDtJrQ8IYDkSmRXYveXsxix0jlfMQYEMf7XITOWTr9Y
YeKYP7xXrY6sm2KwUJZATGiAI3HuMslffJlcoRsA52s6205EE9jME7OqIL6HuQeg+kPl7luu0c7J
PBzS0X4YlLtpdbPG6JnC+cQ34MEVaaIVQqIUSKszhDr2sSP4HKo+NoWmKtuv3HTHSfdfd0B92lqT
yrExpivUUVeWDEvbEjKRIyXoGr9PwaKEV8QqCTGbVMvIR5x4/moCX9n3d0B8VFan0gWb/AdZBp9R
edqJDJIOPb9a5b4SQVSDnwqoo4i+KomUK487jKXdUiXWXZuQce/Y2UmCt6evqHcB2CNyAK4sGU4Q
1YtdNuiAKmZIqgrhMN3TfSfmQZRUqX5UU0ZTMi4vPN9p5wwa3LIXA7cQ8sEDBrkw+Gu4Fx8l7gFg
Hs6yzesydSfLbkiD7dtETPeYuIhLvvkf6e0IM7ETINWSybBI5ZoZyqG+sLfEu2/zeBuI9Adni4A3
+Wrau19D4pXPcymZhKclYB+Yw2mCsUHMnSbZFjPLHi7PT1Q56KusUDf7xKa8FnohMVGU5sJxzr8U
Zbmy7GFHKD1NgKHv111kXJXPkLjT5i45Mjj/0MGhTXInB/wzD4M1CWQNsCZ/8FCmSsdQTdlsm5ZU
1oSSAG/gpiqTPSaaq23jUFy0RWq8PfwYmkOpNzLsTOt6UmEoNwlXKlVhXlBW7+GekJBPpbQeNdKN
ZnyJXbeyFaLdMyb+iOUonVo7bScuafW1enL3ohbLXOnPCVtTsLwQcaLQhpXfmKfu5jGQ0fXvzRBw
jiG85vhj69DgqWqYpcZVI9IRXjRml6eYtDcbm1+5sTRzkxsZgUnlBRWJdmCzVvcM9r1nuY6IBxC9
rDBhzDGjIR7/FbaSCJdDtwkl0EVi+5d+u7X0LVwix6eT47Ms2b4V6RUp3NN/glMbkGqAEOQI491f
XvU/ljeynVeeN6yMHLBlp3pZuL9qC4ECMUrSWagNTVRV5lJdJixIi93fqtNW2cBUotQw4WcdbrTS
+8Om7ZkbSSIgwEgXXEkw1hqvX6tDlUOKSq1RUCE3MkP0mUGZZI9qWjuUyUTvtGfcc0N2W/xxenfk
IrLPvRTIZVllu7rlTfqt/jSZxzO8FT5+YeSFk9vdv1UFXrfZGs+MbpLJRA1fiyfD9Q8NUGx4x/Fr
AJrFtclyMACkCnFh4MnAyAZbUDNxp33po45jCLY1+qh7lXNCzOzVBZEAkNaTf0hr2ltkBLySYrBW
ysCvzdzOslT2gAJdR2Jck72Uysq1dRNNILLlR2V0MDjv542uSrNmUJGKgWr1dkHh4k/IXeSwF1U+
xquXjz3l3LqvYyJ/4/MGmma+8X9fOWtlfJxmNIqkbKuJGyu5gUdMdQ5mC20ghhDg4W9tNeBogmIk
B1wPO0iLrO1SV6LDiVxZfblMSpf+jCeFCUgeckltF+/naXFSpLQF0ymvsGaYekNpnBbpvs65IyiC
btzU+ViTuo8GhC47D0tlXFv8mZtfewS2wqZKIr5SIi/J1Nwe98oi/0LfjE79diBs3dOg1AfNSTLB
4Hi44r8slZBcS9vB5Tws0ReDC6ITxiPpffG//NBkGB+d2EWLUR7X80YlgZEM+0vJk4rUX/nV+5Y6
DYPUHBetE/nUH83ksytT2DWibrhKnMSaEJV4ly2z0TVluW3PZpxdHcDml706NqxU1zfbnz7S1PR+
1R2QhuramYDeV5ajcl00myCfZ6XP8bhMLMj80hIAQ4ISQAtF4XHTKfrxRiTeYHFM6BTDeKqF0As9
lHhF+JallUbMlfBcEjBuflBeekNyp5GfezyBiVjZOp14Z961NFf9TiRGhlECbosORQF1Rxg6p5Vl
4Wi9Jy9OTAvP2x4TFTfBRf9xoeaSfe7kpQRw6mYjrhBkfIcufLhrneAYuBdZrRqCYuVD37bcRKE3
h+6UUjJnvQPhEnPjnBOxTwZK9yJv7rsnjRBkzsVzta+rGsJPK22Puz0/jM1QMaGuH47DtONIKrSV
+aMEX3NhOi9SOmILRijadp/s6vfG6fTGV7oJT3HZTb29Ew2S8Pq4sV5esIvJ7OwTNMDQ1kHsry3Y
3hemLoz9YrrSoI8uBCCMyh96CHOEyFhVUpxaL/PWzA7Hb7WQhL5IM5o7hP4vrPfVPdZoiADuYyJ/
MobkjV92CEbuB4yVkz+VPUECvz8jG4k5F2f0/Q1u5H2ojwP0PuP2Bf7CthT2RMs++jwW62+RNmmz
mt6nmqON/vZ9gHlichyyvZ9xPAwqZBCQfMS2dNDWnLcCnrA7CIoWhiG7Q5qxNnt7yecD9R7PhXEI
qIfCTpCYPVUqdwlEdDzkrxJ4DwnJVv8dxomyWTVw/zXO9J8JHtPpIj1xaZLXKbs1m53nZxwgzWrm
8DL/PYlX2vxVstJctbceCfYBO+EI2jpH/I98LTThdwhs7bc1l3uDWqbz2E0oVMnoanIZNRvd7j4a
qtsTJta2l4pkbc40ISpMpByFUm9iOXWKxu7gIARBvvNvubqBorYkWvfzyBD/W77cT/dcYlA1V/p3
95s1gJXoSL+3ZhQsXJDIeb13wG6zKnCdlNcydFdKooJw59Ltxzacen6hjWPlPsIiCR/l5JU7BA2l
Kib+u00ZDLZdfi4TJWR+qkblGVbvd+tt2gNl+1aPvHUv7K2sfkVrJOIykpGClZsR/l1yPQ9T8HJi
+FeqhqpVlKFDA3yf6L6UbUCgjINlajPnoYX7VSmH1hRK4ExHc2lVLjeR6xP30axs1AFwp3PtjCuJ
N45LWA/j1BCLJTEVBtx2yNKapAiOhJU5eiZgc3ge4J7ZKBNtBqpjBZ1Idhzwq+FPZsOwXuNbEdKc
d7GvEVd+0M0Ap5HwwmTvkTm9BX5fLcn1tqDNiY3ANetM+N8JuhjHU/xFp2pdRzrybYrKewTXvZ9G
i2ou3tmfkCUTtfIflnDWF+UlZ6I1A497bUsHxjcWJz6fIwzE6k0+5W3+ZISD3UhsX6jgrun+fxBi
nvFrKNA2ZNRiCDl0+c7blnlX72aGyC8sqmlQQTRhXx2eMeEXKo9tbLAHWwOmCb5C5dLUWhqbjLuj
AzdgsK5EWPIiVK1SDI6SCBSRzzMqrSTlsGEYr331jhadpvwWr3Tpb828rX86M/1C5kHLlXBZnWXj
LnWPqXEipLcUjQM7LPs4Yq2HNFaQDj5R3W2YmT4r4qiVegEP3LR2yizPaQFeZ3FxVs6dYFbhaeE1
ZrJ4OoYwFGtQxf5jU9D1zN4HNsBhH0Qns1LmxUhV2Afg/AHzsCU3P+G5u/tx1t8fl/xRiHYJTlz0
oOQfXMohL2YEsEVyDJFGY4G/VIm5k4nOsjwfwwWzojF5IuNZJ8TxsH77v09WJJVaV50rqbVvU1cP
8+ASNVqsfi/DuFhT9Pkh67d/Rt4UOv53dpBnI4PgThlMzT/UoeO5w6wvTWkcVoId5AMvk39LfH1d
Rj5qEIWl9d6qMkMnFQDUOiXbv92AWtt593QBQyjwn9/sDQdRHE+oC+5vU1dMy5L9n95vaSEyL1IY
HCV6x4Fv/Cc6S1F0gvTfQoanjMWdPFXlX52KZ2KAkILUo9/GrTr0dpAPpHSUuTc5ZNjlXR5iwho+
HYUiGW4M3dotVu0R/x3Zwom9IwQLzGuEmJEjg/QkRCoET+IpW1sB8zwWlshkg6kgG8O3OLANc2NG
Uu1KcBAMpgXq0yWLP0KgSEfQJehtQzekAc0eb0eD2BbT7Qpcb0+Y7Fza6idreXMxoL3cn43XdagR
WASXXuDutvzrgFCC96pwnMaMQxcE2LHGgcR0nb3WsjcCDUYsPsTsn6q02akKloLk29/CpT/UJIKu
pFcMXvqQh9HlYQ9gJXCbqliFIEBhal/z96PbH5qBf6dUOOKOPrZmk/4xQ05pbYTlKkFLPCoagXu9
ktwxS61D+hIZikBKY7PlHZjK2olEtIOn4AFYv2oAu6J6dJ+7+V8Pg7FvQiGoUs616pN+8rHsyIaB
S/7UIQtt6AZQ4J76u/jbmeVFqADTobQfRyVQ2y/0S0IbEPe0bAOCAkP06P/Dv5LbYYka9KMiUNLs
kNsbdzqsucAohRS+ZsFu897Cayv5Vf8TZJrCiDYsdrT6LYIISgo9UpSYSPwgetKUKWpfGoZX4Hgn
iumtbJNJKNiHFaMRtnI4Ska8J3Vv1orC8iI4YniDXQVy3QEDSoJBydfPzeDra4PAJ0SRs8JbLecd
m61FtLcnv2YycOG8Y3Uny+X7yrLSn8W3U3WCTmBz0o1Zz7vfdIMGH/98uJQhtNlPvUsxqKn4iTyB
dEeSO2XczVcHt25MhcnQrCTXsPNIUWazual+p4T5Uh6a36vEEr6MC01FeOC5YAPaVM/WXjEM9VTo
UX1tLek7t5cP7wFuUFooM0rLdS1CLRLp/IMb2W7WileN8JoE8tibVgQv20s5o2pO/YWhyc9LJnIR
lU0DGfFj6+Ad9KPB165GzB8K76RZQWCx+8PAY9W8Qr3pOOSft4X7HLbjumO1YskG9B3cyH1wKh02
AuAIeEfOxH2jloBe7DnP2s9XUjNppG5FG1501rNzw7c5QiXARn/YDfhHOIRpgn5YQIObhWUkDc4V
qF25JcOgqVQM3UPoGtwOLuOWlfBxqRZ+Kb70bJ71HMn0hIkmgL+Y2lzhYeX43Fzgih2tgimYi4km
IJOvjL6EBD+t2q6TpLDj3tnKu9pzFjApexVs/Wxvd9BrCNsXksc6N5E7e6xFRw2Vo5+rq8tCe9La
ajrxPFMNFfxbw5fOhnuqiLdnFj88+oXb+7BwGND4ZKE7XoJLO/yO6paQ7uTVA+eaZjH4Fvu4kAfF
K8eM143g5V67tA/ecKApVMGZhFujs9I8VS6cstDAsO8Tiz93ucWFYaJyf3t/82Aoc7TALG/offOA
W+Kf/DfLxQjqSpXBGqPcRqTSABOurotZ2UNVsNbT1WSwk/5pz6ZSEGyQAlD/Tts+NrLR9SADRrX1
ojDtQvKydiXNkCeewSNKx1etB6YlOAxXC+Nawxd+9L1uzBwN83LLBkxRCYSdgUgiCTBzv4bkeZEt
VEk77vVsqoZvIZi0pRsUgpEZXo0QlGwsZHxa5ammqerZuW7ESE1F3dHglctz3BdsHYoegW58phn9
q4JVNsrJ1TfDSQ1L53lVp8nqom0XVZ58g7/MHM1YMmhlEES2h+hUYHh5uO0UAC5tzn8uXBnHQYX3
EGpHKmoJd8NB4ubXRm9Y/lNXbI6SiGpKZwT7k4E50XStNw9P3WaYoJy/osMtJj/VOqsDc97VlESz
vIDwm+cBnx7HKmVpRYWLrlToq8jmFqXdFOLI6dZSe0r64xl6LxjtCLTQH7639Q38bu7FC0DIxxs8
FUL1jOczTXaN1i/WuHqiIJDdLa1cdrHsHIiL62u/5EYzmrJiWMycjmCAE4J851IM5Fd9nvDfstww
kHYT2LLQkbHdxsCZql9GRLsudIZpeGr5X6ZQtcCA7E74GeHCbGM1mE/HSo7UrZAuYUXQVkj2Sab1
GXYtMuW20FlEh8E0jRAe7tA2bdY6MO10DKUs/jVOUjyjW6IsRQC8js7DPr0RnPapIOCi58FiPks1
I3DtuuQqiR15txs4mlXnPXlfgul+Ul6UDOOVzZ1BLVhXtk0NLn5Wz4bFKRhhPz3CxseARAF/bK6M
GWQMSkzrk17+0Rl0IXTYhiKoXihOBDzORcfD8efUoSTvEigsh8ITsxH6M7RvD+lOo0I6yTN3tqvf
QbDZP3QMBIKaHWyMrk3akuBYKqiDkogfZYLafjzCAhXgfCs0zmV9tvaTOM1zwPff8BO/11d9qANP
CetH4sbiTO+6KhRQOolSI/5XuuzUGkpcPZmcLDga17nPOnZFWcvQXsujD8hNuUxnrNWgH+E0etq7
0ZgNsGcJ5yu2l7AVCI2Z36/TECKIzurHaRW5C/2kn2Y5d0p9Z21+QZ47nacTqBK7jucVhuZJ1Qk1
N955PBj/BoYQ6nkoJZC8Ps1PFNRMsNWSis4eA8i1CfNZDPJY2GIKmFri6YA3WDRJzSNUykfZ2AzH
OtXc1ml0jjShDYN4BCFrDcatGyfoNeakNcDFnI3Byfb3bETwBhJrI5YHMw3YX8NKdqllN7x5PRUC
8ZJVSKBZrAPZ87pkev7sRo8kl0Xi+iRYaVa/sRddK9Of8O+WO4fSCh09trHMDLoVuGOkBKVArh2E
DkUwZrf9WGIrySejrgLBqdZQpLFP/V7d1QKi4i41i0E1h6OE5zIpRQ9tmvpxhGQksuEUn9k4B85G
P3sPJ64mP6P5DNdr3iOM0QpY3xlDoiJ8mgyXdcUZ+xHwrgTP6tQI9a97MTw4jjvwLplmtfs7v6pb
kJXTDK/ruEeU96MPdoGX8pTryzGjKDVq25r4883OL+z0QdbEFlqa+D5beOg8GuD7eV7aq4vjwAD3
4jrktTeR8OzbYNFdruBdFen3WdtD0VmPfFA+O2YOFbqfBLbjl6rVcVN20s8paifdG2kWudX/LC4O
RYzMWHMS3cdf9nOcw8jzJ1qAwXmsViuQKz1Kqa1pqTrgef12n8vJQmB0EWLfwQahzmJ45wtE2VXy
pi6HFPbwQObAVRrTOQ7nb1sC47JbHrJ44FbomyxkptXsFYYU3LbJE3MULQboka5TmdRoSN9a9B3U
SbBOzKMagqaKAqh/G70KQnuTaD1CYgBBl9Wk7j83K8slOiruQE6+mvRwn3gDxF9dZkPAorWNhqxt
Aao37sK06cLCJ1L7/5Y3D1oDF1r5E+5qGy5xUEQSD7opNiG9QopczMdC9dZzBkevp/qIhD15sT2L
/xUFNf5EOkWslkKm+75HLF4e8hO6UEAfseBDQAGzONi/sqFkdF+mJqhcG8UIh8A3KsK9NnBkkETQ
2Zy1yET6gKJqTe8DoD+zShGc73qRNXV2JuZi7c0MQ/jK9itkNl4a6qdU5p7+gdZqLpmJe6RIXzya
PyQ9rTLKJYMm26x2FCm4YY7QnS0cJsgb6wiP03fDh0ZWKctsy06lhDQX4tZb6aEKFm6f+k4zCfRT
oh2QZE+yolNnXJoHF2ipDNKEA46Dp037iq3UanWCUVCbdJjqhfd8KyBwifjqm9FMIRul+oB3dKBV
fSvkpyJQt1iSHJVYXbfyMUad7L+D7kezMH0YFj77HlL3zzMIr64pJAggb0Euurja3ytCcdZffOkM
kPjsWdxLNAvYEoteTb4DTCqK9TgwrV+A6NOvC5WQtV2iutUolYTVGo/t92pbMbgqq64szSIea+zm
9VnbhYb8qF4nsksLtbOBHfPfGTH97l5qbLu6BqT4ZLgUkpWkByYCFDTjB2owGVrE4UEPhqrAr/uB
WNVP/U2MfNBg+uBm+wm2CC2o+f+rfoQ8v4RlH4Glax+mwqlLH7xxBxJpiZad+Wsb40V2ZxGwp5m2
hNi3ta20GBKXoxS1P7qa0bWIybkuQ/e04hUsO/4EqQ0dur+fqktfYy88tuO3mT3JIig0uE9hoNeI
wj/L0L7p9FWJmpnBWDmdSMO+sYQOUs94bdJe7zup5TiWRDgUBQqX9/7X0FQBrqhoav02gOvizp1Q
VRzXQHHwuuotMj47HjAJ+RrR6i5xBj/OdbP/cqJ2r8Zr8MIFvaXIeFTxuynCblY1/MDyuFpRGgcv
NNEl41hh/QyKOWwQhbpCs+IpCA9IFnz2lAgXXVn80j2rpQHiOW0wS7uHG4pqN9Jr6lblkc0HML2S
MGjQR3VJoDRy5sgQgN0D2w0rDTJgYqKWsaHy5Zf4KFH8D5gAFuw3/FwKzVj8pWkB365BpcVqADx/
4x/Tt7VD1kDNmHvSSihupZEaryP+O+RRLnsMdZYQOapfPWiaiezMqnLDBJHZb5TFY5hoZhoaNtQq
H0MzXXIPPSpw+HCdj0qvpXU8P3ucQwXxL+Ezsggd7sjQV3dSjcLOudpX7gXaagoGfgtf1WOSIIPH
iyQGzqlnB+RWVyu74IsfWWSSuqoZUtWDq2Mu+0EwZG/OCKTkI8mm5hi0W37LY/1WO/Q3Y+MqKPgM
7E/+19DYpO3paCDw1+4LIHXg/EsBVD191vyMWYuTN2HbBFWyYZ/8jVIzfk8dk8LLglmITvHSDQb5
j8x4OJOkvOyqEO0o/lWWmE2H8MK0DIUFolEQ9loBeVAgU7fV15olgamppnz0hg8fl93AA6gtr5Hq
bxSBkwb3xl1e0zSj3uXlwt1/ICq8siBU2mwPNllloitl7wuxV2CUWJRDtODdHGuckvNHq5hXuC5G
BA0bE4KzGbN4SOcuKYmoE12JBBdhVG+XUq6ePsfkMmQ/8uqq+MV7aFUkpo3PPB6f+Y3ARVBMy0aV
BnQthkayD5PApXgCQbu8bWgilhfDbdRwjA01BI69ILEfyhY+rR+XKi7OvahEcNdTeAWEBXMQHmPL
CxvI7TOWSKzfLWfL0luw7HUqZsTFJ5iqjFdor4jxJz+fEHna4wn55jGhr3f5/goiLaUMA3vThhu5
xMwKx6nu0RGANqVuZoMAWAT9jM08YKoYUKs4HOtW2ri9obzESWA1jcmP9uQe6CrRiQH/FbNXNM9X
CHM+oTRN7xuHPaJiCXoiQDqYCSW7KGOocGMm8jy7yNeaO0rpOnGQpx3LqRr94oJVx7GOE4TimeDQ
UThPFUxvJ2zlSZhv4p9tnkcD/K4n3demV2AH0OyIM44uG1I6LlfMBeDdAJerBlYEOzNQHlb7kWRf
6ypBhhnGUJhIBbpyD3tWVp10OYGgYH22VSIBnrZb9+hw8tDw7yCJums0hk8VG6rr2Oan8b6eRBYB
yzRaM22vy1KNNX+1oj48CgC+JOtHNpH7YI6tPST582zMffobmcG5+xiAipH60thC/8KrpMfNRcwD
G5vh+f1koQ2wp3sQ/xdA7UHgaTAoyJnuN4QtuRFdqF9k3HRMAugvS5Or5v0jhmm6rIChh3BTTlVF
+VBM2OVxrR11t4da56eLAvwoewOX99j7PxfGSbHfNpHer4K6uLHojkSCaWCatM9GFGXUKE4xd2dB
NZxCSHaS0Pg4cc/f5C8u+6EMVoKstpZcrKIOQjhZYP+3aSOPfxCI/OElxAI/eXR0eRjUX/CzWOjI
/ZhYw9qERHc6MaOKadwO2GiYL6NY4Xr1dK1Bv7MarGZoJOFh0/yCFTJXGXEfZ1IE9Pooet7umjy7
NZo0shH9zGzl+IMBrUGA5mKcpD92Qq3nU+GRPWO1MlS11oqHiUxDXtir5YHX4KiWXR83pjgs5F5h
f2PufEsBFcl0pLgHdqjgZvtjArELRM026O7BHhlimVGYdNdT6pfGmA4byRa7dGy/rdANuVbqONth
FUlEhUWRe8Q1mWmsbLwRvRTjTwuyu3MhreAC3YxXgqLBo5J3+52FvqBk/txDOmheDPHfAcZR4JdG
2HxF3CNiOyPQKlAfYwVroApdnhe/Ecs6PZLcGs25jax40kgM5RN8uN+Kko87Rk5cSysbiGi3Ud5q
jrxzswmJv5HK0Erc7fZR/L6G5Kns5W9ykhBdOrGc22IXDrYnM3urMsWY8Mi/Te62Frq8GIi75459
blwC/9fUUBNq1JFeTnvysepDgWf2HDiuQ1FAaOFEmDa5jkEeeU1I73hyapoa9kaGCpTH+ywGN0V2
0nR829STv1qhkCjDCeG7gmOGn65xllsPTcodDM0+mYmBGtl7z8NBc4QZn0FDegrSlEvrCd7jkniG
gWKiJLcBRp59Rfx6RV0of/B8Xqtty/fQf3SvRM45exEgDgJtPAU3OiXCnqnyufzN4UsoPmRBJxKJ
Ry/m3NiNxisgq8IhY3Ny6GldwIil/9xJtcHCiYFZ3FL3/sbe4Z7F5IBKTcW1p3UGQcHqVwfaZx/Z
RwlPhQBtk0+fUBf7m0TbREsbH8txAPk2AW61hsTTajks37Z3nJT8CF4HrK/WIjoXOU5ZMqQ96KQj
vXa2yaKv2XlWaNPL4APCkZKOJt4fTK2hrSKYOVxQ210j1t42HQqr5LfbN0EyWexSsBuotCucVNHR
2HXqm9XDwHPlEs9N3UAKVvOjoRGk0CyYzz/T3S06+jFCeXnEOGNeGHZYsWj3FtOk5Fa2UGGZYTA5
QxjdjtBvRz1kFvf/UY803NuZIug8lSE3v++AwgpcVZS/H/P5IzrRSGCkmUcHFKrQ/acTlHyYGMHa
sn8wULqZ+0jLzkgQkA2Gubv0nS2WEOiiz9DIFPpoicGc7YZIDaknyaN8dMZS7inelcmsP8JJgbG9
UCu7WuPSd0lwS8K6kI1VJqSwYl+He7mQyw2cBw+mFt56fdpMaZ4LiUZzocKno0lCugLeirDt2mfM
0WCC7d0n/pzT2yyRaq3LvgehIAsE1lhAfBG4WlLVfNiPKrau85mKLekGYxV7VwhO6iyDWlgeRBxR
og0DPVgQ135nSPX1znJgBEzvxZzXQINTdDB6IBBUyLVH6S17yb12GgXAdvsnWpufxTGp+k/818Q8
GCaAck7D5Z7N1EA9Tr/qqJw0BZ0qx1opnSF7+2J+fSY4kOGb6aOT9IsaBi0Rvw/X6RZr5r7mT4/S
hYuYhWc6u8/vfPvvS79one+X5GRnZJZm2vCuQoQSdblgfli7qHmWMHIzrjBGhiitoPZHip/pWxUD
XxZCIZAg43dSE3adP9Nm38djvaPDCL7jTqUjBdI07hilozFNe6AEAqSkbiSq1TdOHrEtU4I4ObsH
tu2fkt/OKdqfjo6Ei+dk8/PgVVkk8NtHAFxY1UwHzyk/gAAGsJg3+IJ/yF/7YM4ZcopU4iFbUd7E
4SDI1v2yJnGTl17H9u0XSuy0ue5oo/wOm1bi8ZOtBbXxuQQ9sblI0p8nKIaFRFXi/z66Knp6kHrF
UZsEm5Focr9CQkJptirqMlgAARzZ9shmPV7aGiD7lpyNuS/MJ7F3xauuJ4jCyz6XZsLVqtVGsYJ+
L+BvRFbOgx5Hh3zv0NUrllo1B/eTbO5xnUsL+bLldfZoHl0uho5y4ucSrAcMy+er2MpudToAB9wR
fTSD7FPwfN4Bo5iNCG84/LEmcyt56+G3FHaE5wVDvPVByLNMu/xONb3TsVJa6FOC233h4dszDR4e
6J7DUfRGYSbximo0eSO7cQ/JaiV8gQPyZEkKcItdHokT2DMBLrwty9hl65t93LGWoXYg9aziPo0b
vQpAZIYsurbtaHQNHokwI1B6zrL00dWqTEYcmW78ngDOqe9RL7JL+6STsifgV+WQxHGFEkQ6ofg9
g0JFvHDmbavrCoSRQdKl3BFySNznRdDHdJk2KzhS4AlyfRwCVAUvxLvsU30rrrFdsdeJBSMHDBhZ
herNGpR218/REd30mwMWOKYWi6m7jjcfU4zCk8vQ6n1YXbkDVTEDDSufGp68tLskx0ao5Que3Yrg
18p+PNlnd8eC7fjzzTFWur34IR6ObGRwRCMp/p+zfn5ebKQTo5PH+Q9aiOgkC/Wty6lJ8UHV9a3O
U1pwhwks+UvtXk4nX2uVV9RlfqETUyeskTK9OycnjwInIM81HV59CMwWoeeZ3GHo0QMAArbemOBW
1vdjSVRggKQpQHRep6gU9KFq6LWNQ29c11ogCHGY5hnw2aW3bdhg+IYK7Kq3JSyzFfE+iSPG+5Op
Wcm8wGjcva0HbI6JTC5LI6lQ8pOOPxlcqOAZd7befQKW7muvIdnBs8F1OvudrwWfyifSXw/foJci
pzIrx5lqd3GlLtIkvnvPKlixSne4XW8CzA3ZAXUcIlaQUgwWJ4Fv9j9kUKwsqoCMgEvB+mQTSnKW
4FpOHcjvjpQXjYIZdkLTKym3PRUZByfxFsZ0DB/+i8IwOTqBRC5Y7ojD5NxD7+6/GZPt7crp2+xb
Bs3okoqOnXpoO2lkzBHySYk1DizuorQVtMDFvZsFEku0eK0qf/MWO5iKor/+TacmWJoT1RTkWliB
a6I8v+MiBhatrqOX6ssJSv03aXcL2ELB704SMkaJky+T1ZAzQUlnEMh0ec6x1r8s0HGChtIlTKSQ
qlLfI8VxaGGvg7ln/3mmwNXwS187BAXLi5Q8FxzxRUyyVM1JTFdaRFPnND3/JbOPtYOIMuDFH5Kf
F/ExRWMwRk8tzh5BIFxYl/lClgasDw3biRDluAcS8rUQH6n48r/lFo/erAYuOQX1Qu7J1+qfggb0
b8tbNgPkd5Lnm4gvE02Moeui2PWWTER4HE9QiCjHTPbzzHyM0cexJf1PkEjtLn8CMSWVW5o8Dg6C
+JeBeZKS7Wu//l+9tgrgeB8pTm9IASui1nwVythJ3RuWh4FcBjOowcffYoIw1dcn40SqrVTqnqBh
h63hIIFBXo3PQ9AKFS90BQsvGlv6uW3zqmxt35F8d1QFC28Ssc8GUJffKx9fH/Nn4v8M4aQjm3GK
5o8nvo6Oekue0n83WTJwBWJVDA/GHyOOQDJZ29SJ56v0c0WMT1IkIScZTlx9xVfuFlLXD6swzf6K
saiWlCNgz/Lu7j9OhDOHRESp+4AoxwodbpLESsoMjA0MpyQ7iThOfk2AvLK13CdvONu6YVYY60iv
T1urobuV2TPRXW8cWCURmkYDt46CXGq5Ro8USXIpdvDoDKtb1LAeWDsqxPERz+UGiri1MeJKzOAT
32Ed/DlUBi/yi9Lb6ENM4xkvmT4foexMUTYYEfITVTmzlsmaACgNbYkBUTFEGVVEBamEORcg6Osb
eBV/Mh31oel3/fMWtpSyI/B+Ha6pSPKar4y18LdtjDlVmrRul6GsulE6ytVxhTmLJaYDGvscJx7j
wABc3f8Q8U2fnbfQ7kR1R5WESHDL2B+c8CCrclwgrAQpW087BS9G2AWrDuSXeJMXxE2U3C9E6ghs
XyeaCliwmaK8CBdgx4A2eQ5DEuNal/jAlkB3vzA4hoPfd0VQkTrMhAV9sNY6ZPgqy1HsHn9jrRxd
Qn+xHYq0VY/FGgHEQuP8tXs5BFcbjqFg+Y6x9b09QhRdd5bR7m8hQZOSf5gf1qC9OBIZc+r8kERK
biEmby9iDig2Lro4bdjIvaGK8Oi1JzTNVqhbkR5pvRWl1YCEiSZQ6+jooU0vRxlKsvZD1ApMBsGb
M3pwGRhvGUAjS/iDjMg4cxNW/a5FfgRG62H3SaZ/7Hgi7AqySpIwlCqtNUAoOpcgbsT+JXHgcCQH
gTDmwIA9ONIPyd2DLH1ucyfiW5TqVub0uKlQmFevlCTgvd/aiYW3J23IYYyGGB0O/6MRX8eDtK0y
mot/yDPnbVtpQCSzsjKC8nWBgr6utO5ft/oMJtwz/K4ZwKXaiNouJFH33u2PI8GfLlHYoLJtF37q
q68dnmBRbn8RPA4vIy4iEhWW1ienl/uUJwIbtl9uM+t8iyd6qwdTnSUVY/rstwlIz/IgbPUSoi0m
/x9gVXB0laMbtDekXJFPphLvQXV/VeZxB4CQaUPmgSxIymezeDjynglYOco2RGjFHCnQnMsX1vpu
9GJo76UBPcfCAu+4jZecbTvm8SgsDTToPIsE4Mmfh7k/XzFpfgh5QtCi1w7uqeM3RTRWPXXd0QGu
kFsDnWZcR9FlVzUoNCPNUlGJabA11Aks05C1V1g80kr6HIuyXoPlNxUyEXU6VRk826pjahebUDWq
kDXs5U2gF1qUjiWU/5x/H1bws/BvX3kMCTrewlzt5ibAGuIxd4ZOjMMDFF5YvfPrj1wE/znSSZQk
O0qkgAT2nkokG+DApmWCUc3KnmAK5reGH7ckaQKN19VldfS7g2agj4Oz7H6NMqLUa4JIdmoyF35T
+r+3NKVYJ6ffcAr4Yw1kpqu77mwgrcJthMyi6Wf0g3RHWGpVA6n5sI7/T+lBgqytZIxr+9Wm0U04
kzk2VvDgduhpdPaANePHNppaJd9lXjES3hyDXkcYiiWxEw/CXesJTHFMw2cIjmvVbfbwYTHQrTKq
Jxw1ANXFcuRZY99eOhksfvYqn5O7cJCRncEaj4372zyCmwjxRNrseZc62DBi2oxIQ5KORjiEVjWe
sId5hQDOOsbWwF6LpDblJDEG5Amjfg9hWqNSGPpRXSyCdJWNxQ7h/vtQdYYpoKLJDB8wJfG1ezSt
c2Y1/HzlkfZGVLcRDv005q0r9pgdvFq8pV1ZHH/+3wkMRJJTDFLwvf+nDrU/Yrgerv45uCa8AgIM
NiaHfhLjaUr87Av9z+QHmruuwbhX3+BSR9yrStTNgKDKD42rqJZ749POawKK6+Hs+Uh+h8sC0/JY
vWo0MbT3BkYJ8vZQEgjXbUsvHcLUvGmObmkb5Jdlnm6kTON4NVHciyasLAZoW5p1KqpAQLFM/Y8Y
8NA876J4NIrCoAFCOl6Z0w848h4/jvNLR+49UrMpuMxIwap5YQUiolhm1JcUOdTk9mCItrzN2jbR
mCHeZg0Mx3kw+grnk6U1uy+jkTMr6snPk7QkZXqzFhb+7QLgUFuhh787H/74MRGrTuZGodqqOQwl
mcrGbXV7TEun9SfinxOBEQ7IOqXSOUFWr8YDtq4wOQNvDV7dt8MdLDxe+/2hdbhyzau2Uhf512II
q87kMQwTBPplnDv4GYYTvnw91L+2mxk5TfuCBJsS9CGrLwcjg9MjoR9D7N0FfFMQfiobYN/xALCz
WtedFAk6j4jUg0tSL1pj2WqIxCJYxWPFK36mdybLnxIrn3DHfOX899TmiMcalnvK1QZTFLUHhyF5
7t0jl3tHBnDgVRd4Y4BXYYF8yyOCAEfOHr4zay7HK17jGl8/EnftqLa4qQvbqUPP78qAkIWRcePC
2q7R6ohhrgqi/ur9d4O+2ulRkSkZB+FXhlLXH1J5QoFkISOt/aHlyRAn5u1KAYqbMwQOuBLjwxru
zxnYAzgsohxXX5TV71nuCsaqCms8V04oln74bWE7NAaxI9kvOw5Hc6N48IpgYHzuPJWXEW7zDI9z
Ffw1CrqCb3lfwmmNp2WAOQ8v5W7Zx0b+2hrkF+YzhOF3c5c/LhsMldhMeJfkiiVncNthqqAlY6Rv
XVNY7HnEOzpP8LXbQpSQzi5mTjiKBR3GdfCKrH71AwkorjJmzIMoElrdlHPYUuTBeBw5wxYMgUKx
l9ypoIfCksE/2Xw2TrHxZg7U+qtKssdg4a+DxviS6ahrLjbB6xgigh2KDAC86QxaPJp0R2yfqQsy
hjXEoMfv09MzIkVV+sHtN4xLcz2shdAqwpWqG957TXYlA3eOyjlDDcas/GahRJCNXQaD5wpVSP6L
ajMa1C22Dkcrmt2T+EDkvbGT5DghjZ1wXS7BJdubK/nrPrJkvXbulk8l8+FP+x0xZEMIgltAoimJ
zVh6i/NkAax5khw6JRD4TD1DgOQNoM6PgkIwkEkGGz2Y7BtstD09YjQZ/dyOXcoCCbag4c5kcQs/
DoybUYOqf4l4DpQhcRinJil703HgZRTUmu4GuNBn65jf9+Kg7JAsBbE1MYGMXB+b5kWzVxzOvm2u
MlydykqNNuPMEl0I6VXYhcLQ4fS1kEdJPKtD3CSTXbKGTHJro9sFPzJasrnuq+W1DHTiqYYbnbSs
lTLNp/I/YYOJ6MWkNwZCBNs4L536HGTLCatsBextvytdDSecbl6+Q0dwkVwoE8eEiPxaY9jloWov
x+qPFpFNB5lbSxcNCVza5TSmNoinu0tvvj4tbpvAWq2UH3XXf1HgBjkD7AQwV+ZZGNZ30VxxyeW/
gzO5D0FYCsDzOdky4mwMFcTpmaCu2eAyaA0t/ajok5NIOqY12HE8of+u9+sOlB+hYPoUhLEoJDsR
MQYkGoP1YRNzjuon9XjNOw4EAYendmUZ8EhL4FuKkp54y/YVOlSqlN4cG7dchQhpKjzwAygiveeU
gTItFaKqPTzXEPwr6g2Y7RnmliOXZld0X1e7Jf7hrjpqq0+lk/mPUXgyhlhU4pAIP05pmJ1C4gec
Lc7i6OsHLCGNXuPLq6iq0PFzjRyLEALlYLfOtdiarK5WBitJ5qhgmSSCWkSZ3aDJUzeZRU4ouu6G
Yl0utMwOOuh6AVDfmOebYQKecyUlMgjlQkFBcxTGdEFfAHJKh2Cb1k0pqHgkNsRUeZQQFyyThT+f
UciF4aWXmEgI7tYsJnbKTF4x/42DO+n3Cko+o6i4wrbN8bRBv4/bGFlYRt6Gw4wT22BIHeVUDPlD
u58mw7yc/SeoPiij0mnEQ367gzT29a4MqpQkLczfUIYhpmnQRv3qEAcjqvZvsr7pglL6GiUXRn6n
tGA4TqBzNWUMzmTEwS5+tuUESg02eV8XKLA+mU7xWhmExBGLIualp3PNIzTZWxwkILHhY83DafM2
9RHp1JSPF6tKMEXRqU2UC6dPSzI8MG1z8nMOZoUiI2DCmirqlmZDMeZ8qx4VaW2CThkfkXhcp9UY
M4zAOiYlXWdKErMLsurm0JKm/US8IIaSXBlda769YFccjHQKT8q+Ac5NdwU3pZO3dthAj9AifFzu
L+ZDEYPlOElT5l6vy5Yun/v6EMQGBA7W2uMhyUT2f7gMTfKW7dm0wm4/wdax6R/5FFX9FiI4xVtK
SaCi10jasz5zJ3NeFpQM3oTphrd7fNpgAVaLwIOEgg+1fYNvHW5srLWsq5NS5nC9VvyO2cGtJyzh
5wXtNJGoitKDLWwdsJMDJG8nNIRzykQFUtP27S21VpUEkCcBLQssIjglxNz7/P37epH37hGncSPU
CR7Q2NhwiDB0Wu+ptQ3i2Eb9xJS9oYh1aT/1U+3EkHSWzUhlvZdzbNs7YakOGPn+ynp6EzB1NQYj
ksyZd1LQQ7PJwp35NlbWtdW0pBYS6d4swARn6Bg1YMPGu9sZ7B12/UuOiMb/C2UkWurQyU4ziZ4b
EhxoJ4HiGkPhLycOGzLj2boEhLZQYDZls/j4R5GK1zNExOfTORr9wRYwI6ItALtHcWdtPFMT1nFN
tZPkp7MiCqDxX5D3oCSuMausQYQlAMmFSHbGKk7CbshTyu5HnF2M4l0go91JRFNHYHpLHEsbd2ke
lQbp4P3xU9jITDyzXWicfic7U52K+EDQJZzJgPO92K9PX83dz4ogsntC7mS5LeUAjC7VUI8kgnMX
eb/viL6JRqIqYhXWxM9GxXAEGD96sjYUmTRPfiUA7eiyolx14hOl+XmOvIo029YLmuPsCGNUHh4r
F+rzoeDHsrQhu/v3AyXY/ElZQM9LqlvsQOH0f/5JQDZ9bKgMt6sEAECPtIt+3drqfOicyLNjNum3
K9YY/ABc6tSG9VDmE4W35SM7PSPp7B52HlQr9gjQ9C3rx+vYgekUBwDWUh85EKTxF0qPyiOYNyof
RKKlPdYq/jSxx4Yjc680O6nnNFenRHhHI7j63ENF7DxXNhM6T9p/N/2Qsum/2G6K85ZQOHPOdDQW
tIczWiinEUVGUE+nYUQOvFNdyK5WMzIJYOIiNIpJzYstxAsh0fBmEi4ErwGcpo2SjQC3/jh9mqwN
A/bJuyy+Q04eHkA//1qnqgeNarpVlW8LesSS+tNzyBqZO/eK99pSxGfuvDD0v2oR3jTyr5Is4Ost
Gt0MBK/JWmHnWA8QHIP9ieoEBc2RK8d/SlEcQd+XSK3+nU5jHCCbEvVis9zasVg2okx9abKH1ODx
9FQ5Cg7lzV+SvLs/pntH7sCdZIQwpnsM53kcgOdJ0QkGqg5gktFnYLIn/RD/2pAOXobao3bI3v3g
URulPsMSbVuK7zzGaiQ3RRq0R3OQY3P10bAu+J0/4MruCfGLQQTYk5p2DeMsFAkkwn9poLWI8K8s
J6cmoBKpP4DVcTL+Xfmdk554opEuJvBRAtv1CjSZlHrB4FupO56XpDYHD1SU27TUeuWz0O0Po8d5
GTJkvlDVXje/+zNyq61MI6b7yQnX604AR/H0cPRS4NI+7BfrJ4mGmouygWyWhw8ZBFkmEs1cbY8G
t8l6jDp7/vCRhi/WqLiCB2psrPcl/tZdZOjeVAAr6ddWGZQJwE+td0rldq5aAfPxm5CNy9nlcJ6q
ZAgvVXu7RUHjIf89D0xMZ4XOuJ/mWtdrAEc+mVSXJiQCfRsCf7psENL/znCe9TbP2NFytwwFo5Jp
qni46GM+Fiu85b/JHA4rUruGT8pRQdEnrcyrChsLdJGae7v3MYPcN1myaMNq0h9+RGyccNT58TBj
+iJTRrAbcLoazKPdWMnOqsv0lddg3LnnOeHDbuWFTE7wfvos9hN4MgdWQKaHlonHloyoOF0t1SXH
eLWWVbOT0XYGPfRR2yzh+toGGLDot4835vOJgADz0MV18J0Ac++THHag21rPLXSxh4NM9cYgxTzd
IKFXko3gk+sOOVyJ03AJvEHJ5epbryZ86pkfqSpsX1nYL59YNyt7CuPKUa6ryzDFRee8YQH6BUbi
umoHZYgTUvM5wlwnKh+XWOcbJ+EJ71OsoWf8sJ7PEG9YmKEFS0oShs0vF7LU6jyoa3065d67AatC
KdEEKeYb76t9rW2B7qHBuo46o2EQ+PDa0JQ3qe6To3J/QRRKpUTxbwveH6R9cFSzsXe7l8zdMace
O3Qx4qUn1OJMGiOh6/H3Qp/vSpEdy9X57bZBMYMd1KTyHuRdDkpAb6E+v94anNaMcGY41rGnQE6t
eJibenPgkyWvqTbbXY1O75/UC0DL6I4CmIhaLI18svclJ5F1L4Iezyj+9WgdWXWs893t/ayVp+fY
x0tJaMBabdqwp5AJPbBVBI1tvBaxCPa2Iz1dsNBvOZj6JP2HhtTK4N/NMIN+aSfHosFstgXf1r2t
XLD69uUUmQtwaf1TC+Ua3hRbTHu+QNvpic0saFSRvE41wznc8besjpyPpZ6N/2IeDIqimYzdMu4H
wGe0x5fURZLrAh9uhgRWknAVCsWJ8J0ZVucuoecV8np43NPiypqtBqi7UoEViRWCKQ+f4L5diEDo
mkE4YiPl2tLtbYBTt6Yn+UqA1shxjOhAmKL/glDjc1IHC7zaNGD5KHmISOgnO0i4Z7Z+HxVcYjkJ
tYg+utujEkrQPndc19DaA6Lqh65C/Yiam3iSbXCy2j/lJv3+G94LqA0dWVK6Kqj1j6Y/U1mRHixR
2i8in+GW6nPe6s1uFKUEw8E3jW2wgaICPWn/HAiKO0b3K/lcgpaC425Fp/UskOKN/7dGbNDNrzjJ
R2fEvxJBE2MMbSjxJ/9A8h69FxLiFieDaV7ONhZuSlUzYKpgdzQUjJI24o3eyoOD+n5JvWh/pOkj
1tcAfqZkJ+szlwd4G6pgkpJq8bE69tKU38/tKSSHqF0MMpvqGBGyg8ONjarOgQCgsNgCDqgiUffk
uzuy6Pzg5Oc59KQsSq3NF2vrMNMMUUd10SLZD37HSO8h+RGJl1OUN2uSmr6lTxBOZOMDJy4SbbGf
z3Hs7V9Iiudr7NKg25xjWEzfXqIq/P4RZ+xrVGL2IsQxPG948obrCiMpjc6D1NFSeXpX+2F6zvJB
wsqNznaZ+yPQz7l3619hwvMWM4nBYJt8O71sBFeqZAunXcfbEYXbuXtWHmClwLPspXNftbtQ3C78
WSuIJgQj/lUB3E4UQBxHVXn/DPoBIlBS15XGJA/pNeiGJxjh29FdJH+nnHxJifS0eYqSKEo8f3VK
Ewm+/tquG4QtWTJw2DLzG3s7T5PXxKED9OlK3PsIL4t7vz0z9Cws2Ux8xYpepmLzi249QmsQakpB
XZqboopSctnes3LAS6hS9BZprD2ybQQ3PMCPyuGnDJUKKZcRz52SbHod3EV3XhkqjqjoDDdUtSNj
KeLozc+AZK9cpn/pt1zEaDyVVjh9BxhsLOUWqQQ9zSURtphP1smB/XAduwwaetFNG+WZI99NWhOz
Erx0HfAxBzl5rE7WwoB3yGdH+FAkEVwK7gtkFgbBLQSqLeknYDDtavJUi5GlhU0PRv60JD3XcS8N
QR1IJ7m9wfuIrkbBMZjzTUstW0xjS2O6zohCGl3ADfYfc6eVXa+LZ22l5s4GDpox4ERKHjMfm+bv
sHfHjzS8jPusBEA8kWu+2PFAeW6yHD6rpVSPpoPtJzfzp54+ZwmNDQ50VKxcgOwEPVVfxwLHf22C
wSoUyRUDGmJMd0ylWHcw8vhUEMy6WjdY46t3zm7h6oVBW39Ih5apWDcjYO8hcPqjLJVVqmKVPoud
PWEH84GI7WDov8G5yvnNNxUFttnf2Wp0SkNz5S39gpz9qQrmS1RgdcaixmvQK1S5tCCVk6LYJKdy
giivNe1FqAkL1AmaW8IMcQzs/hWX78FKzbo8LuQG6EXsyXZuDeqwk3rvl5s7KqGrRkvo+Tf/+tJ5
IHTNQgjXqv8Qe/WwCGyWfia1+4nzNP7vEJVHHSHIK5o3/hyjlKiKGREy3NTKc+7Xr/8M8rHRpGWE
zrsLOeT7/BVmtArWFh27NJcL4nc1X9MO8NP7jU3uLMUQHOzy6ttcPuFRfw2QA4TNda2zq9mAdi2C
4duLrbsa3wASrUqmL2WqfCd4+tAXCoNhhWL03dZEPSRkaqxi500IhVvMarIDSsc8R9MK3IdLbbju
X7+kUq6k5AKTBSmjSh25gu7DTwASVEf/JpRIy/6eyM4XDaWvo04uTWPGxXftF+FMVxaZntEXL94B
9te0u9NPGYSRIfJAwc99vGaBg9OzsYbrQKR1iGYZs1orN3watpNpDVgsZhvNM9j3ZTtjj6Ox9UIh
DyZUkPfv+UNtoad15Od0stslGfxlWl/MW/KgzFHNKK5icnLfD3gJE856g/2W0GuiJO8OGQfIcXKi
/5eJcXfGQpCOqhKokqL4DGyOgCHnBqhNUIG3JeWxKD06S41VAE0YZ1HZ1Ojcs/Pw0LKp1NWcgTv4
7o0F0WsY/j4sg90m4xBVsjrFJIoWbcCswizZsA9jngh9cxljguY/snw+HI/2+mN2SCeFR66htmHz
+rCalpfqpZY/Rg5wUxFrQBbgEUzRv5/nIN4eMfb/w+b7SbWK9pmxCk1GpNl4GfJW0VvvV05EZaIL
fpNj56t10dzqOrnJZ0JR2WMZ6tOfTTQCAAnpzu9GYAhaPejrCYohpYnUwt5UTwm5H9OXO9lqe4r1
fXG0FM1pgQg9+E9s35h6cXXhO0rZJniUQb0jEz8KX8v/dAhdvjG/ZTZgbFUiGmXeK3HAXwSDp50r
XG0j6ltsAnzU78AJa2ghM8pMNZBo5c0xXK9tvfXC19HrgaRnYGgccGr12jKxHcKyg4Yzn1c+Ywtr
RiQsvTpPGZ5sY28KQsd6sBDgmzcHWp2yGM6qNgumJzQNYJsJYIQTXZYnKJxyWq4AlVL8AGlxH9Mg
95a1f197SqeEBkncZiSUytoaBhYNCPjfxjWBx2ygc9qkY+rmEwKiUnQJFGg4DsS7fTX2QYqDz8Qf
kQ5rZW+SnpoPTqp7NTkd1NkrbBjn85yuSlcJRRkakMKn1mJsZxuxZmGmE0UlMnwY+tWZYwttQCK+
pU1sK3/XBhZjk9ThmV1kUvNMF/yP6Rw1p/BNRPKCLr85TjIZEastxe3q4GaaczGC6zAUHaFxb5S0
6EfPg74sY+sndS3QVe07gAa9ocoQ8g7XzgVBDIKsfezfreDVdtPtQs0kkzGNpcTKz+R2kFYXxRF0
Iqj3eoVAkQxudmzajFZn+XwuORiWbychXGpQbR2wIqCYCBipTVbSX9eb63gw829EJZf+U7pShfwP
Is5n2odz26TnpZ3pR1AdHj1oroRCRtbJNXmoxZqHRrO8ZbXU8dPb9bd8EdfWG/8VWho1mUvyDs7P
pQSBEC7GmPrI0D440W+vkQBE+mzFgX3G/9TBY4ukl3eoLJPWJrzvq2WLT6Ixe69/FzwoI5x3C25d
aZrKPpi9aKSVZH5Z1sE1cFGvILLpAnee3XFcBi0KLz6y3Cuh7EPyjK/JxCddity6r83U0Zj4kqs+
yMkrEGYKTn1ZuyEcjICyG4JBi/2kIS/eMj9u3jfOUT2aDxxgow59HdmkQxbgWNX1/x9fNI5nB1CL
K0GcymakNyaL8DlmUJsTUhERA3Iiog/XdPIZcd+DK1c5E7exi5TtLdPjB9kKdjan3pMKkKpp1dpd
29pGsHkCKPh33qsMnnvrU2Ob67QiSQBoHShwJ/wlp7y11t+tOOVPsLZ8XcsqUDR4qsPGVyh5IZDX
QRi31qVNtKirVb4yVVD+qAifePJFwZBknoC4TYho1USURv+sC3norZWun1nZ/w1kzDR1abTFvIUC
wyfvMzpc+aHJTSDLyYX9axaXw3GEkNp+YDsNPayWTlLMTq/JMajHj0wCB42ebOX9t98LCBCvMU8o
hbiwFe/VPyhAQiL75H6aRCjwOvyROVitx0/r8bxATRzfmX+IGkMp9SntTdipHsLjNDACGmZnePO/
p3k7kNGV6FQgUXZpc14LQJNx1d4Tb+T7GH4lOG0s62Y3S06awAlV2vbYOwsPRenzknYcgSJr87E+
QblOlM7Ly8J77Ap51hpmqePjISslvupYOli/zzO7l2+nHJlwi0y4jTXQdTKxI44LmSKSIPiodCZd
HE7vd8Jzup4Cq0m/hypqZN0IwjQ3nHWBiU5n16zhb24lDDAy1wjcs0pYqyvyL9LamLNyTcmWocwD
Ez4A8g928fnrhbtsJyeIwKytGp4cC6UQ+0/QAzIRZfkkiHr7VcW4dcz+kjuw3bSx6OP5Y+u0BUjg
Gs6Ot9YbIBDg7HOgI3rFP1039PASorbnDBOKrNg7iYAIKmdYDvTkXPBNB4lEoK6O7PKVlPHG5UWz
srZqrfqAOpCntegnvVsacYW3YG0VvHeaZfmuWWu1F1WEgEcFvqfs0XaT8eFENr+f5Qvp71wax+wJ
bNG6ZpJ12to+5bsaGxm2V/nMzTniGG2uqEjeVUvmgr0HpGYchEhqQYddWcenyJ1TMhjKlAGbkw2m
WRHOqw3mZbUXk+qf7k94ceDSZ3t+j59DNWRngi2Zezh3Fy3TAyf4gWBmiZ0jX9ZiwY6CyQbX2i7v
rd+vghUo3aIUmhuqL+Z5znutaklAfzT0YnUfZmXll+zgXDOZUYRR7LOsZtpPDLss3vZhybT6VE4E
2rmq9vCp631G2S3v1u+oNkXXMOTmZQBIV1PBgvx/fXKNcDYaSWjzU5VT6q2ZpZgGPm00B+OSTO7C
RPxBrIUPTVSWqSyPOxWord9gm0XuOv6JT53pD7r/CslZ8Xmz4t6eonswU4wfcuHSH5kv/qEjn3n0
I7S232Ui+GhjpNbrJluMNouJLRODsqBE1WIpYoJyzvfjNcv71trcsuS4BOzq6lTYVhT+Demuunep
9zUPJm+hkFlc9ptqMGL2GEO415hSSntB2Bu9PsJ7BmN1Ra/UUiGf3J00ZetJM5Qs+Oh+CEYQsHCa
55obh2MaJw38Iawo4eQCE6fxW2iqhG4i++XG/lRo8Ap3ctUF2r5aPEC0/ANuflSOlM+7BNnU8qrG
21yBRiDkkqvOl7O5TwxAekOamawDrXXVudFh+RqFBMkZPgY5R458RLpDr6FQIKl0sloCiLJJ7pEB
ascJzuBgHXSWFfCo6SbMOb7qG0nOPY/rCaVSk6TQwvN40o6QJlzAM98cWPioKlnHQuCDtwrxxMnl
RyzO+So20kd2cfbNH+GOkGxG/bwZeSj2U2EWKQap8eQNsTf3c0D0nAwUlqq/ZpJBEtg9NfCCYgnu
lW31Iq8W1cMoGMSTO6enpkLXEfPsA8vuMcy4txtbloetkYreyyyxTRbjCBO+1ZPC++wnJC9/DKh0
K486B01t2Nokp7Jkzqt4hd39VdMOjQg4bhahiOEG7VZanNUE4DiaJgeXszDLWeQLmJexvZTP22b6
WSqBs8WwRFeHwwwYFIbjVvg6NjMrlLql0jJ3JZ0qnRZzBSsmpwjSJ11ZR2ifKo8xDvu4FruFkub7
5dMbLHKg+BE/UGNGWKd0AY2k3IySbzA3WrC3Bmlf2YrLMsgqVFBUCw0hB4vG0tEVQm1BDg1MzWqi
dIHoOByxuY/qVOdBoUwathc1WpoHoe2/NGlVkxV916fMQBWoUijuH04OfcVpst8KSsseOu9McIeJ
nw6qvUjknwjQmSDA3HUx9mbgcM5dUFgQE54cQwSvosbAgyf/8E4LyHGXfadutRo88xKTxbeOs8/x
/tTNqwzVSylP/xX3h3Ye84DBEeoHpH174NunQE9+KueQRgB9vPQ1TuxS5AD2ZGjukdDbx5nBuePJ
9VZnH0BvNTHmpJzY3EK01yhXQh3O7AgBPfnTBl1u+TFxSiU01ntosRFWEJIuzO6zXaLXYR2IyCEB
wWZKH+Y+KVmFqN3mPSkhIpwHjcxAKGo5b4pUC/DYubBpHfe+PmJrQBsq4Q2dO4E/IoH3IzOu5m72
fpBnErZNGxidAuc/kevSFGLoDNUz1XFIuzvG+qIyJvOGHo4nH1ijtYpRRIbA7hGBjZdXXSkv6A/c
W2eK+/vycMznj1rwUGJAFRzeRG+2rhugnjdINyfUakZaM19p4uwW7gf7noAwhhmDOI02MfL/SSsH
jKwHmPMi6LTWKYypdYK3nhom4ecq9hseeO9L+YsE1bNQYvemMXgRJ28uoOcY11Uv9CLmm/Nh3kwz
uVz5Ls/sOm6+rgAkwagX9NdjCfNFy/DyhbByQ5B3ZzyS25q2TPnuZbhPBAUlNKs+CSbv/1lGKwq0
fZTbngD+1gz8rJum2fQi+xV9oy0Fxgpv/Q876iSTXrSERMAJMLG4qr7OZ5dbLgbmi1+KlvzUTXdi
ksPMkIKA10oRRt7Ans3v50ffiBoDCxrCsoSzuyWV08SvrBK3f7xrTePr8/anXKjAGgkkJuC28gJ3
LJeO0hLLsu6aqaGGj+zvuZYiNTEZTp/xL4ASXDvnkbtKOib8/OSo6hHJ+oGAg82jQlcFQ1UR8RQ1
o0YLKxNtFmQc5jn1WPEXl/8p3s52mO14YCSAtihlJR7kCZp7Fv5UoXtgAtaRVpVSaZTiRDTSTDMc
TNCeGybMTc28/z1Q6TaKwvcW5oSTNI9+65TYSnkI/0x52pv+bid4CzAUTiYZ05rrWfS37zU4K4ej
myKQmwPrpdahZazr5WpYbVEofc0glmD+J4xTc/RDRF50TVobDpl6gg1Cdw3QYOrraGnvyWKC1+4k
l0LcnSwm4NBtleUdKfu1zCYA7LVW4kIR2YxoYHFVdQFuKiZ9npigInR17buvNBZJBzDPZWc9+cRt
FP39qwDefnpRlwblfKph0c2fejbuhCgt5ZLVd7u2Etume7uORf0K3Z9ng5Ch52W3PdsZjEfCUhFx
mVx22unmMdkEGCc2nsqhHL1UFYy1FuD602NDrKHIN8IasDBQWglDnzLTFZzVPSJl3q993cmYZi4I
XXIm89eZSbJP7ZfLijUfoLAeG5ejY8KZrP+T7E7st0UaBtmFb1SGLGMj4BbgU4MZxIF+iTYrnbnJ
UDZGp+Uca4upmdWoWCZwGnfy2jXOWuAe0X5aSUy8iBKk9ZjDCvmTke/DwwKtEJ65OpQsRhbjf7IW
tl5aEjb0kKpIhvtrmz3qEZWrvJdXxcUIRlx7sr0tnGOK0Z9sNsxWEi/TJmx5bJrelhv4KQLPk+WE
8Jfkgnit8zwCSoo2/2w8FaTzAfpE/jYXemc4Sk8Lm9oJW0/BWmYAi+PmfQqDpxc1E57Us04Rs8A/
ATALRi0FBuc48en/pLrkrUfYaK7QcVLlr+9zvEmLA/dL1A4wrpMxZ/1FGX9g9uD1hm4Z7MMbwjI1
oUV0Gns/Z00fog+HHlTBOWk5nsnDZ+iMfdIc0QEIkrz713OXHEBsOY3BuEiArYTytMKWmx2/gpAM
oYnIGtRDzoVOlcVYV5QB/2LS+Aj6qVcr+fwm3wucBrIo0rUE7ccSWZ5xtGEx51Jd5oxbZtU3JVcN
VmOi5fb1LFbhuJyYLM+uTZk1OLxiZ/JRmTgRdjiXsXSqmRr/DZ98RSvoa2vVsbXOMAdg8FNOY/ZL
2vFkGG0I51Y7kD7IxoeWTgiAQZYOrJmeXyFnx6hpXA0/jEQIFJWJqnx6ViIFXbEJ2Ghru5o1b6pL
N2a6kPftA/dhOkm9lV5Xl8ZWxHxBlVMIAxs+wkUeDxsCsFjFdpQIM87nRxWmNanX7hF81Q8CnP1H
zYYpHZ2meTo7JYqum5mjL13+b4XAvYQ0KyWJzQN60HiyCuNBEYIVbssVSTdw/D6mfWnKxJ4lhery
qG9+QnwHxf3F907scIPdNPuInxw4mIzho9Kkl+LJMi2vzwXEJblDhVzktNnUQj1mITO+RX4V6Bff
q3H/mV0kolTv8NWOCb4U/DuXVRvrUX+L+YlGsQQDh3/zX9kpen0iENd0ghIYNhyLRvy9SZRa2B2s
YtKfm6dePSU3LnlzHyHGhGMthMnb3TmaPY+p1vERe2b+AkHIYSyO2/XTRuVQDTWfjkoqeg+hWV5T
wIeSJsIXfsPKEITBpLGLnEPkj++FLiz7HFSMpI1I3hNkRxqstqQ+RmResaxvRImZx2nvUtHDnMxg
v27Z4yLh9TYSPmOojlmNm1lOClMRAP7q9zf9pBhgJDZV1g9v0dS5K58xm818cdDIsT4RzWnVWL73
hqfzClmBHS9jiVCqJ+zuqLCtUI3RC4+f5A/bSF+MRlFbhn2N4cIvt5Ta4cn8UJ2X0kSDBgsJjA+G
KZXBdXpslt0TvaQ6/NLFguY3ww2qym3XMzIatEQCEqfOBt8BuGN2R733VeSeEzNBVaR/NOh6Me7l
5WBEdj/h4aJ+HZ2K1Vz8SejJUp6tdB6aFP0x37m6sQzuFsAFNCXoP/PohwhGlwqPaVrt50wgxWIE
w/UKOzcCR6AW0CKoVjjufkRhit+vf83ED7YNV0QUnHObdDaD4Z3sBsm4gihRYNTu/nvkuWbXG/0m
Hx3sfv8rv196aEKsMHrH860GhsFEWEKSUKd/UdBWiWxjjC4RsDzA9q5etmDRrRxlURgVBVuzn1kb
2riEbAwWkbQsravFfba/TalRF0GOQDMDF0citlQBRKuR1y1MJR4d3e9X9jLVmnavlub6cLjGGwEG
b/91XpGq0dq8HktIVSfVGsOAvjJVE3Nk4flirAz2MiFTd++n9v8FBcyL6MLb+nOn4gxHOBMREsVw
O7yw617ZsK6caCQO+LRSvm8zOSfS/DyhrLKUr5j1GGwLuJqcJSoZ435B/hFwlf71FBTXh4snU1bD
ni9joBxdqmJnnQ3Pbn4pYwK2f9NLUgfRsXBYkbZHy2KuhtO2lhw97cMrki5P59jXCY80h97gxNEM
bZ5ppPTagp2/io1/EpMWDJ9FDHxEntpfbOjJk+5CsWwhRgTG6cpAo1KciN7LwNfZx/aHCmcgfVjT
eWKSVIOY54MXz3NTrigOtoLO0Z0q2nomqdWuEWMT9upsJ+9lhzSa8UMsUCRs/RCq5H8FQCsyDFYS
Jr6wPwN/rsItxixqgIyfBjt1pMrI5+mztShlSgLrJEnNq4HNZackCHDP5+o6WlScnYmbjgemHPfz
8bQ1CBW0UiGBM5920yUn4fcWNsrkkMpa7FV0wlMmMPV5I4ehcQ1jgHW8cFmOsWe6v0qG/FwhmaCm
Xt6Nzw816HDWvKQ0ZWl1TQuwzdsVQBRYxV9n+NWn+Fd0sUBrWPjX0ZOdtPUV1gxuCqd6Bd688mYR
eDugL3iTQ2uz3PmpJqjOCx+N5zN4RxTDCLQqpJSLvBIqmTiIuVFjgDqbaplLaYGNvaCuiqvSlBNO
EmX0KlqMCqBzjCl8lRC0IbyCWaI+Qbqaam8WECrogXcLGs9Nvdg87HnUSxtLBts18/hT6xoXxFA6
mx3hc7qC+gSKtuJokjAp6wNamaO2woivLpaU26Wl/1SjNSwVUe2rhF27s9svLCr1iCvj3sgDgbGN
k+nTKBFcHtM2Y9qfU4BXvrwzCtKnE1zJJeiva/FMIwt6M5jl9f+h+K9vK5j6fJhsg78p3jfZY2po
ab9aYEgtdSHKD+ncXsMtMYpcU8KZfUHuglRxfT5zZ+a84E02iSbpDUDLX7KH4IvoFJYiIV+ydUHU
j/mZem0gZFAtwwQHDqASdHip2NR9Dya/0uCCbzOzT2c4VlfhMDUkAXjcyyMu+E9qzbEggj1KaBxi
eTxrLsBJH7C5CaYwnNwmMxXw/ZLFrtFW7wZYLSj7/bfGGpF7aK7hiz71m3J19cER96eQIf0JRXQ0
qcQdLF9Ij/BbQ81UziU/6EIVOTYSy0EFVj7gHvaRIxmfcMn30BXZMyb0Dmyn47/rWpR0PWIQ4+Bh
08wZoRaWpBiQeJKr+ogQAlN9/3wNAbzNNTnNp7PjTdYZS0aAVjwKH5ptc8OBqb/c6C3t673BRjps
UKFqRGnunSkZ0uKweEPVIVJ+YRPaqleRawGJA5hsyP25o3tbhHXRO7ddwmp1s3mrEfdMcjDiPB9c
tqOUV5NbdqY2yx4x4Y+2yQ31kVqAmF/4qr6imIQ52q2toxzy/7AbDEccB4HgpeqDJtyaFFkvvkt6
JnnQmymN8Eb1fHNuCDeXcF3wHeinI55wAZBmS5Qj0EpBMEhPbbpdAlHJFq1LQO6XeUo+hH7NVzTH
hCqeNvNWbHlUZwqQE2UQDa7lJmsH/LStphBq+SU5fKu98Fk6qj/YZUStr8FPUk2uGsx7syMDmxVf
n9Z3vs7csSVgA8sq0GIXlO1ywuO8/I/pYgZbYZxpjNEJvrSsM6BaVqSej8uMXvByfZG3y2pIGBBX
l9ZrGC7u5A9eXrHD2IFZZYTOcFXE1VVAlaYEmsyw5k76z9gZkH2V03AdUFBcYKf5B1t14mLOyPQi
vBKzxJgWdrkz+dLL1h7bkJhUePohTSETNWzHZsdeAQSGbD4Y84kMlx80WshwknWpZ40UdJGFcF5h
D1VKMo6M6GhoWRnDnYX+0yw84xBfNhfuV2OSiZYHn0WQfO2qm6zP59vb5K0bkyaN7u9Nv5T9m/7T
eiQpua60D8uR3wBuXKp0Qn/OPT6Nh0yGf73P3r+mEf5oHfy/6iextlq5PDSqcBjYLvosU2iQREbP
NNGa7kv87OoiLT9dtVWrRAVhrljUVgfpBtFglnMN16Zd8h+hNk3b6vULg5sARaeQ7EWIsgslIzrv
rafYIStTovkIGX48sZXym58s7nlLa76nQkBJOYBsC3YbJW6LL60sCXxoFFYIABzk/C8x6JyIVXtn
Icde+Ad36g6S8dt5lGagc4lvv7me9pHvFLWO2T/BNOu2H+Y4wWg9lUaCKlHvETolSJKKXXRWR9qk
42fliGR8p4gzwjPh3QZdDDTQVsriIA4t50i+mo4PaQ+M2DL9YmZ9+1IIicD4k3LpIgIGmFn52/ge
hKfqNhHX0HeHyz0wJUtKkNIwM7flcNTwaljaVe2m/5L4eN+v2rbZwy6MqwF6SK92Oyq+e8kMKoXF
BiP7WVwK1w9MnxDAOeSrsHtfTFWFSXAM7gtL/6JWYqox+mWXSp6rCqjmaS8Slm+sM1MCNrrtmFge
sdQcAbRPgIgEhWE3syiSxRhQ3bfGWA0fRH+YQ2X6NaX+ogojWQD9NmCkZaiq6F61WHc+Zd2uuLte
761dMyLq7CfNMi5UrESKFTC2OLiA8I3jTPw0NIQDpn9rNOsmgUSwkYWV6Gzek8TwViDElBKBd7g1
pf1Ejw8VqCxcQkqAf2U5I1SZfNuwQLGOVK724B5oAVNww4Yf1aOzYV6T8NaM7nFUxmvcp3tLpLIl
LanWirIUelwwj8yf/K7uu3dgVyihcwcJajsvFl7oMb9/pvltvoxtfcMJ98KvGSvxyZ7+7QCtzRWt
PHWH9HA2FUGq/GTd1S1fkGUoR1eYr85AcbeFS79Jm4wvJz2dsI6ieEMT3HhYIFzsq+Pjw7YMCskG
PkVbqYLqIxKumXbgHCxK8tDE79cvt/rWjUmaNFdz9Q7t2vFev7R+Chi6OTk+OhQAjI70B7/P7ysJ
m2B1WF9WddSmlV2c1FHqqzdVyfq71gV8+9tIFn5bZEjF8a6q8NvDk1R8PP5xXFGjzpBN1bVaKXNo
/hX75TLJ9Y6J4fiJ+Hld+O7z95TFltnubuxB5HkS3L7HCAmBVGve9+A1QMtkfDIFft0FLb6/0HgZ
du7z0MfvM7tly58YEO7zDdM7MBTPMLXvMcAqmczts6+F1nr8kAjdfe+4h1lZVHFlhJezM2XkqFYt
ipzIYMq/jWx0ZphKv7ZWyRGv0G+Q8vwkSldodKLIOHtmYQC5+awtKDZVWlYt2uxeNz4AyxGv7exz
A6alaN8ZOY/XzDIJvUkBnXzIBuUKXM5KCt+Qt7wLtvkrRczvtayHLu4v76mfRwhAhq3q2wcfYEYz
fXaq6flbUr7rjKyfCNT/Vtcr2pfYCryeasT7WHDn97xg3C0mZH4TVHDer+IYOuQntMPeDEudCWWg
yNmD24/Kn6NQPXCF7nYWqoTfvTdzhAQgtThQAisyd4Hk7W9wt+qP59LjdM8j2Gzpa+HSW9ZR31Jj
kmk5/V4+XjjYrSyPjP4fZZ2nVPG2rNv7acwa8Pm99B8pn9T9kbDpZdHsbMme3kl3U+87KAfBLPaL
JNPWKpdXfwnaXUzmgthObIcu52Vd0+GM74DpVOH4SqsK6IVyzn9KDpc+m1fHiRyfrNbdkMlBPrPP
r/GDic+qyE/yGPqhYy1P9E0p1Lm/B9mwMZ6H1Y+KtcbHLfWHWmp0pTOebLMHi+kpse3OTus87w+z
EO95qzo8SJR58bg/nZm9UxLBFXqUqXagfHuAUdxFwfbC9JeOjJkDOhOQpLj4t+hACTJtUNWMvx37
/6Tolx0KPyDazLxYwthX6w32Unc5QkkMDEPU/F4HIChEI12oRetXVJuOr1J6mrSNw5jncblJ8yq/
WLQqwYa6xp9PW1b5FmOE0psQtHM61qDOGHkRH33TO9cC+HyAiByQfRid/Z83FnB9uiQPhd4pKezU
Ek+1oYA7VQnaCF2dI/17wGB8wkHepAFwvUDqGokmLdn3zGrhGdYhKAZsQiwBfO+vmz2YQ8CyU0LJ
74rQ/cy4Yx7e1HRSO4MSsj6dbUR9j6zgmiNo597zhp6WclUId4BlAeMiitSEtLdi5ViFMNVsZ4ZS
uxGgYWJoM65BK4sG3F3zka9VebEqDY346jD7F+M/jKQoKKJhkFF1kDEwBcohuaue8KHhXpB56yBy
YlZmiilvqdDCKQVq3hiaTjN32kw4lLuCWEZVoOdIKR8hz4yTWqNFcr5murr6iTy9hJNE7B9VIcse
QCZb9dRQvqSoBK6ohfj6sb1rXLKr4A9oi5F03bWHvj3D3KSQJorO8GDHgDUvYst46fmdX3Kc5ozT
AIfpNxrDpB00VVy0a0vVhn3beTn6v2+d+LdASKhDPXT0yY01ELQDVP+zJhk9j2+GW56YNf9faoNO
dfug5OiQ3X5Qg+4WpE8KYzJKnLwCj2dMzBHYmduqGkRMyWbpPjNwqx3juW4jk9pDUJJXLQ/4AcZL
kRxVgtk/4ofP2Dr532ZqZXcVDqsO07Mr3ORAr1nMsYvN42Nt3PJvZjLX16Q7afwndtlSJuB7ozv8
6kh6NjzMQ7/hF1h9/cy4sTCL+TGWRzijaCbYOOoyfaOvkKDYKuB9BE8Ot1Ai2Lh2RH9N+unKrFuZ
ne8wP55k7ge1WyQ+9WSpGX1kIVWNpn9qHbXkmH5jKDcUqDebwLSTTbS06H3UNiahB1kA/3SPG8Ri
/e2C/2CtjGo5zDVAZUbbFujbeeaA7Euj8Vx7WMSOreqHotQUbztns7qL02etRUOIGLTeVd8o7gcg
XkGALEP3MrOpMsIc5LdQg4l8snsM2c3uPGZkqvR2mMPuu6DPPZ8f23K65IYIT/ye9cWh11GfaJdm
Y7ytj5Mlwk59j+VomYI+l5HTCy2sFx/d9M4Mu4evl2PNhM/x13KoC1fNyY7txr5yhpoVKwBubtqV
hpvlWW6zXjBtotJXANw3elLv1Ku7062gHeIABOIVkXFQ7qlVNZtQMpIQ164e0YrpLArRAXV1Lfxi
JYvwxRvbna4de8XaO/OvX4QR0PK1NQs3mN1LLQRKIiCM4LpSB11OOVP0eFlWwQ10qui3ugaTaUgr
zSvtF6hjsvaEsuUT3gd55botkL6j/KMyHvNfdYSMC49XK0ln3Y9YY/AmtayzjcVFfYaH0Upt0c9C
iejGPSS8ialR5inXSVUVX9Yra2N/imHUi3vy9TFIcSGBTZePBuQNN/G6DEgek2dYjanv21EAr9c9
PU5xkv+HpIY375jf7419Ls1HESg9B3IXyR6K/NriRSFKuY0Us3B/tffGKDDo3DL6fM2aae6LLAZW
Ncp6yCws992yqR/8ABKtz41XLvVjUTf7N3r39BxP5kIRQimGhRmBW6/2xmcXczHnlmyA8Ly4iU0g
ALiQ+wAwpNQ47s9GorDoEZtWOHkzxo6VxmVwfCr8Tz0KHwkoqPum6mLrzBAXTmEBJtibQoksRNjG
eVsV6pDI4vmRKBPbfQqAsM0QcFPhSsk1d3H/XgPoDcECPYTGmjpseutrEHmpd1is5IXTp6la2G8Q
AFhdCRjw0TEoqBlUO1C7vgFXb8cuPsSeSoNJ8GF41z2IgCOuIazciicG9foRpvcOFED5rPQOGzuq
sniBaTLdacx9BIoHo4h9Tscas02J6iWnGagpcOlRoYVIdkwe12JnFz6rRpD+fgSocvqD6T5soIrL
SM7+cbkyuE7o0H375IrpvA5fycGnwqYHYxxbM6eXIfsdULyMTv/AOu3odFAUNJiMg7jXxGgvFM3Z
XIpMBUcGMFPPCvtKO/4pmq41L2ZqHtfvMiP3o3HzV8NG4Z2rHoNxI/GI0Iy4RnQigBMgtoK89dzl
hsEJQ/R3h7CGwsZRjKy+LjbMW6vYQPmA0+iL7Uj/LdYNjeVLeda85cMVVsre0xUxy9IWkg/MQOwt
0+u4e/x6+Eexh6PZcRXAXCau1TDDqo/5nxIkk0ghK1BPndgdlNGMWcV1Azi2RAj/GYR0pNGlJINg
z+wxgxOCjmoKnOlxYOPyroryufLpuxr6Sc+XmDDYF77C236yZ/JJrI9yVUKDLpBiAGw6jl6gCS56
zRdBbKI6nuFT6STcx6DmexRNslru2ThPbIeSpopVjO9zqCVsrcSuxBkwQW2/289lAHKatZHyzZol
XS9h1xnW5KUJfSEN3eL4EjugeFvijy4/N+QBXYFZRIfpxZocGCjo1Skqm86eLLc8c9cf0nteQwZQ
akWXw7V28S2A92IPBYSx1Tj9rSe+f1bk24kWh7QKEH7xkn/Yd1GiFlLC9OEO8zxh03s9tkDEvj5s
VZdjtv8ZgCKyKGV5/30IM0l9YHfgEP+WGgIxypsJqRNHpb5PmutmYMyiBU4X6Ll1ApwDvKrbWPlC
kDs0A5lcShGtHhKMNDf3sd5k5HsnjMrficXsF7mtQ5Uio9XaBK/evLQnt5Ohn3mEqMSOTPi2zwxq
WfxvYHjIxshIr/w07c5oDDND5n6OLk13I7Wf+m92dvTcJbYYbUtll+ExemPN6D/gaopa/V2UDpTp
JVP9YYQOHL8/wgrxEP4P1Edds5iOQx2fAziDLvF7sbxaPpGHIY8eIX4Fq4XAZwxK1UuyU99VOwTi
pm98fPvp0PQJIdlnGclTGKGdTV0oio8Em0bbZYJ6tTf+tSq4OtdsMHBDyQAp3oIYgRm9KTonGlsX
tZfnXIPiJTbbwu74gZqYPbpon+ADOKJvgGeTiEXRfQZ5sAbPKtpKbWXsWFUgSWo1kyKZNGRPCGYy
TBuoeCMFG/v3pwF14Po89ymuzgoJkIUC0Fll1f7IRYEFgX0rR0LCfp4r+WMhtGBGXPbKCtXEnncK
TBBw+cHch7bUZzq/qanUHsnGqXGAw7wcZiukJWG5fJ0qq6EPUhcol5adqEYeBtazGgPeJFjcq0NQ
2AvTOKT15ZcBUPCmX/lBC17E+89apka48HDuuQmYZ96LjDUd0HpsTDWPtFs1cR0j3l3RxUT4cZzl
w7TA6opaIRQvkFZ3NMbKJL4theEKVSkFic/PLJZz7AABEgfhtN2mVU38cuugqu9AIy+cEqORBv21
GPcKXV7oWCVEyKzCx5I0Ga3OsRw5MaImYjrzdF0Ynl+PPPihBUcG22/lqIqopb3I/ejTuej+8GE5
scvMFBPzxENq3UNrDmlz7dz4wBwRmEtipH3Uj3T/FzQFDHNlZbkMTStD8Cgx7lvGVi8QUhRjsSXk
0Ru/xNPWJGoWN3slzQpHQvouJNHpouyvIP4Tc1sx82jFuY3oDyLcEXFZ7Gy6TO4kWbUwzr9iSCJ5
buoFaZRJwMNWD0HbshGrFN+O74jTMKjmUfSXregs/ZCLybX9je6hMwwaId0lMzCSyT/O3qCdg+qa
Ud+WmPUE7GPzHqDVl5O5MPXy9UmISPoM7hA48ltp2SLK6Ri1zbkFjS88/WGR9O3eRVhjzGRsr5bh
iTSM2VQxuzhU9Z4kKaRBPANql1V6IiuWkY4h0CPCfpA4T1T0syg9yH/ktO40yHaczNNUZ7Ay+xdv
+iVIBphT/wgxxOLmqBpI20B0E+sLGWRonjIqwenLB5PibMQMjIRS/JJ4+URQjnGiVF6AKoO3c8O1
/mG8l3w8A4ZcG5eqxlvULdJLEXr0H0cIfoHFFtpnvf1VT3scQ3H5xAedvrJtru6ktAZLKnPd7sQw
MpXXh6HrWr7LLNBHmwGdFonF0qhJvF0jWH2hRtaAVPywsLHuPN38fWYxWaFc9aBdsmoW4gV4RNC/
JByemIL3W4V7Qds9G+B6egC09lA9dhUwNJ0qkNHrKQqSyoP1bEfbTjWBaspsH5Vt18V9Ix9321Jh
SdgeTkvX+eHqNCqqF9vuBSFQKOVXqZTPSd3ZTqFwLMQDmfNZ8ynwpIaorxvErWCwNWohjZySyxxn
n5LSesMOol/IiViYXnPduuQVF0CiG7C8uv1DmKou4Jrxfg9aItvcmwI8BEN8SkilfilDX23Fj7NI
kEhMLdcw/NZvxNMeOC6V4vvuFbD+xZZrDN0bdbTEQRi7PKSd42kCN/76jmHpZHZ4ynerlc9c0EmE
PUHcA1TKu/nlUPKxDbPXFZytYjFeS+8PSwMM55oc7gOwbwESlhJ3ImCoQ7hderYQmey+6fdZW2mG
7c2VR29Sq4hTOZfK89vUlLI3u76IGVqfNLs1XOLFAacG0V7e1RWgTgwx1zc+Rnz3YY78we1i4ADZ
hMH8dRFZh8prWQEn/BaTmFC1E5jAdL6VkQ04QxgKwxSI694ODUpibfO6eIx7fM90NUBZlcoSLKlg
4H3nYhCjddKA8c+zHRvw+l/0op0yMmcp/WH3p1W94QhMuxuBOE1tsIE3dx7Xqcy6IYnLO9KgTx9Z
SPeTq4wGPyoGt9nP9yw0UTsZczYJBWcaINZNk8RIc26XRvRz5AkBrPpEH8Q/fRgs2BKFqP78Fjic
UQZq5odOCouVEEcsc1DUEVhmaf+Tl8wyMU9gVpopCx4tBDz+TLYYT4afZdunh/UwktSAm6mRJ2PF
JXhXoNkoziHe1HtOFk6A11J8pFhSFJdpyIPMJyJB1AxH8vJVHIT9VQj+CgkQqIHpXu49ELkaxv7H
9rfCtE2yF8OVyozUhSjJh4w3ADTdZZ/VtWEbEZmAhZqdKhJj5VWyo2jDyxGhKPouAJ06abpPat0A
NauI7Va5SNu1NBCq+z1V6WemJ1Wilg3H8FUYkD48h58nCHUkolqzJurbzlVa7oUWOD0uXLKZ6ke7
cEWY+Zww7bUd+hGE7gw03+6dkOMHU5RUzun8H9XOCgzGm73BJCLUhsbTxKrzFfJfc0RxjMeA3zmU
q5rgUuRGwW87SB/7p6LptbCkbhORhuClVxVHmTkuLEtbqn7mjbmfen65qs/oPtJgxuLKjzycS6/i
sO0gjVj0ecVTiM2/wdGWkHH9+0UMpJe+EU9kSDWol+U56wCmhYXe3dBsL3B1qi2um7BtsP/cTFdP
8EBV3NMsF3hBWln1N8vG7ITPfxj3B1J8kTMYJE9sJPN4HcfpSH+VwDEbb3AC72H+Lr6DIbca3ceB
wifQKybvoO7A8iEwUvwflSmHuu86U0wsaktFLlVeGQWD/sWqi5qqJA/cY5ZAnS8DTyP7+UXQu4RA
H8CAgkqa7s+03TfebipCRPwUXQPJv2mj4y4CEDJ0DyHzKDyh7IkFFqwEQ1pm9TKR5UC7dtWmS3xh
sUwoDTEGJ10Dtd8aYmIBbcnjEdQ7OFFUaSQWztd4VXqx/XXY0rkmGZWGXg97w4ScFb7C8H59Ws0Y
T4OUVldSW1ncWx7mjrAVkXhRORk2jvjHq70tAZWSAazidqEmXdWmrdeGdf9uXwy8Xiz5j/fYjajB
j88GuMrKii13dQOC8dhijdQh9lVYwI8rOYA53fy17y4KAFQ64nfGTbWSqNqjQHw5fHz0SVq6QX41
/co0l1x/QfIZhtpXxiBXzcfDZurwOXAT++A6NUdehh5W5IQ5lE5kC6BJuEDihJMbZqjMHhSdHz8w
hj6GJ0487oBBgJDQtvVR1owURKJyLFztpFnvPARZdM2x6iJoYCZxF+tSburI3njjmZrv3kY8t2sS
q2sUIgXe1188ojG+ubh1lf/9V5+lsB3tjcQG/qdoytjh8FQKEYvcWKWFW2eHWhDSzJDJkueqXPW0
aRlfYQIuWdqXFBFZ7/s1tYjlGpaj+9NYiH2NoJJdXfNSEAIPcvirAtT/SPGoG0L6gdL8CYlTF0Lk
pp5zY9x3gAIuKPN4Ovip49nUbdetbr+4cHXCUkOEsmMXVuwIF+4pkvO09xw/cHSSxaSdAqIxoymn
j4WW50ocz4JiWH5NCZVTsyKYzknre6VAtgcYFS21tRkJA2+qA4HFFJeUNWYG/sxfsXsYAOfnbAfC
LV8J6o4Il5qDuBoH2Ptv3nP2yYrxweG4iNttZoFV+JY6nubDW9Alg+l7BLBbfZjo6kbV/ZccmYMj
VrJzOr5L4ycvGIQjCI4IHVGS4uqax9THy2rEQDVtt6JFhC0+JwSOMW4vH3liDw7XvKiVMgNuG0XH
eomqmlGMLiu0qxfFUyP0HKyQMhFeuuC8tRRK0x3Q6NGNvPXDyZqU0VR8W+Qrc3rXfW5+S/E8nyvn
gLMLzaB5p9cDaySd9s0aOvmRqOxOkv1zIKYabEXXccpnU7QGr27Hp/G5v2T0YD9eiwpski9jBZ5e
l7dLy/Paes/6vAbgw4+V1mPGz77qvinnEbYpuP686NpiUrzUT/Cw8ZL9Oexh1YOznMTq5Cx217hV
ABYFbLmAPyDuWLUkOKBPnv4Dmm/GTtTCpQX7NxNriUi1xlDhcO0efYxaaBDXdYKtJteF1O1T02II
q+f+bOB3yGrPij8bs36tRoYb/m7oXsmZZnfMit7Zy+zYt+L80ltqIawufqwWHk5IaZ25zJmVNOmO
1eDRsIxlZ9WIoDBXOWJHIsr8mHVt/rrzXllVQOzl7DlP2aww0P9M1EDpdq5/aEA8ju3pOdtgZ/fI
0GIFCNVDPuYDeCBqTJmwv5PSMBjBfc6UXlNVpNpcQIrV6RrcGq/MD0FiDbJZS+x3xb2cdRjT45RW
X1OqwBnZJEeHIZRIhkASLX8dcXeX+hqbUvtwB0SisyI1MhZ8ZlJ8Yy2Ef17i7FmCkyuo/GgPmjFI
CZurfUa9OHldm7nbLTCDLJGSv8YhfGCfui+O+lqOImfG2v1e+gVEd7Ngu+HRW7gCSvjEvTI91uG3
uxfiw1+24r7Zp5k3+6L9R7DeSsdxU73dfk91KI+39N/Pva0hJuOAiYHvN6B/GtAlgWxXWdTKcEto
CO8u+DdlUYV+7JSrQEdNlvh7qRjoAw7NMhQA8Ntf8WTvz09iO5lJkJpu27at8MAPqKaf0b9OUJSS
vZo+6Ov3yJZZkdPu9OVBGTEPODUoSCSWjEZjb7s8ucwnf8LF1b85W0+i/SOumcSBRUvI5Gee2vPH
0KXaW/PWFsVw7NMcBqrXGBZqEJ1iMuGtfxJwpf7J3bEksqvN5l/ZS58WoGMKx33MesudKw5j+GtB
+KGli4xfZxUYDjoEdcTw1IEQk1vOiJxUIN9Yny4Wm38tuPA2hzDRi/enb7/L86UkOFhH1RJUp9ji
kA+WJCl8HixF0xrRCWrJjtLwmRPFv1etcJ/siOYExXS/ZQHZzeI2cZpHaaXHTPFONVdtj4xbyGIE
bjjbSdBv0i7GUuUwumflHJJRpq+EhIILm1DrfQVlBFJMXghoeDPOXdAo6sMtYXY5iJUybV8VuyWf
RUls2mN71s7GcwPcRTPrSRCR6i63bvdxN2vFfy0R9a30z2mib4B4/meRaTTT2vemCB5h2N3boSa0
z6HlWg9d6bf0UBAPf0YHOc0MKTBJMiQeUTT66DhdSuYcX3sImMhK2Tb0K/rd65EsxhYrM2KgjTtz
F3aNOPa49TuxBo0cEcl0acwbvOqmn9pZswr34fNpoF3DfBxfMaglvf0Rip3R/mzjZsv9E6eHOF9X
G+BEocvlFhaXs2Jafe/0WOEvWt6WXOIasS5KZqsrzczXCnxKlUNu0fSUu6GtwRb5wTHLGRwup7lp
ac0LMp/LS8eTxcXJ5B1uahwCYBrOhNfcd6iAUMXEVav27Zz1avd/On0etINMdLfRX8rVLUkzaJ5O
nsdU7DoAd5V569xxvsyz5fOkLNgcjK+E9IninEmSdZZCfXvPjcQ0zwDPc9VewXmYe4UqySuhW2DB
vOkrXBKwYPDtdDtuooEWDZ1lCzPqYV98OSwYkdeSWQaBkAcnK/ueuxGq5jW5YIm2LEUHs3iqz2Fo
Mj6JClgZX8JhVJIBtXEAAsUigFUtoJ1ENKiGS9VAVff1tP3Uee6EJihALQ0iAZiJr/xxy1rPd/zj
LoV35HeiiFK9PvuyvD+Cxb9kadHYuj6IW8q1oGbexAqZAJJfv5eMGjs2gDa5f1oV3sV74wquW0CU
WNjWCQELOjMzHvzbs0SXspVv43Vel9zhZmZvZzhoSkjutWxzuyKeCGccXTHGEj2XlwurNB3SfOZE
K+xlLz/7gqx6N2aM4PqghSM/CzYfjDt8io/TNBDriH6WntqYi6C2O5GFQx6qY5yakbsZcx4zg5tF
WeD5d9eDnccyGRG9GO6l7Xq/sSTU69pJ5d0QgmjXBnbvj99DiOE8W7T7T7TkSX6bXNFA4NTc68IR
dO3qjzanPa4ckpOLKHk1QjjHm7ISCb+CY9bV0Mol1rwlYi8774w35VrANrnB/CpCxHwM9BzbjU2t
OhlM4HIGkBV7MNMETSnnafO7SyVn5+H604gaoxO9oDjimOzx1G7Py57VRX9mz1y8fkiHNRgJ4pyA
/3SQFdvVYF+Jp4y/nWlogSDHgi0ZxdZLhGFNr2COTEDu9wXnHjirHfI9/mcvdGh8A3QnaYCgBxuZ
scMNuh1MOoT8nRz38mOeDpSbyut7ZrjvjiV6AGvlh2LanKWaRAzUigG3QJruAPhH5wn5wXjlZBNw
YNxPysrFRKumcmUCUBHcZUQaGmKv+0af2q/t+L1BLVHrdiuxxkhg61bSTzgQKbcslFmRTunOABJD
NiD9sZF5vwkkhrDQz/6Y1XCq9nW9xMeVBC26rLNvt5S/gLAeJCEQDm+Yoar01BAxnQ/SANNKPiu3
jliKYTHv7CJTEzCo7ufvPKgoOmCFxf0qOyqUmK+EJrbws/rN6c4qorwiL9JTCtXdWt4WQOUZUDVp
WYsWV6VnZkuOtHRXRviBZhOtIFstJIyF8KljHnYykGrxjnig2gppipQwShX5p4mR3NK6YDueZEit
Mx6y7tCyans/IZmb7EMSqI9m1ljwSZzpFsg1b6xlx5a2crz4zMsGn9q0hRNrmL+93RBrd7a4Dvsk
wjLf/+G/uNWeeAnJSdwtfKYwyBFVj+7qBWppTkJA3X4gOgdhBcOekxO5U25+wHTyFR1zowZMYm6m
qxlVqHyCDldRZAGYlR4Byuo/zV9wi0R2T7FYJ528gu6LO3KcSJpOlO1BRMczK8Zf2Lx4rTVtCdeD
u6SisDQuZXCeHptsHuuMzU4Yk63dpGNUgGKUz/h1DoOZqO2v2VwfSArrihVvSg9dq+S9oKDq8SvH
al9s0icCdnvskgO0/YLlrHVklR9BL7CjcsGpVcPZCE5fucA+uRlURaCWUKS8guLPqcKytTDumOP3
fhjV0xtxVk8hDqP+auG9qqp/JAo0DHWMKT7qzNfdH1sRu6N00na8zU14ZEXk4AbDbP410dJhmjNe
bmpicyxCId2y0uTgmANKnj4u99J747SFUT/yotZjic1IsyO3S6ff0ozRTyUC6fP9jZlYaOjcob36
r1wPtJACcpef39JA1XKc8yHEFVIkIfvCCPd4ulWy9RwmVzyjPvgkYdi93pPT+Im/EzRjdOSNYEOh
yb6QBa0zsYe/1m8BBAnlE5JptjX0xmWXEmmCViTCVGpS4ocPz6ydYA1IDTxWrC8i8N9z/Vvx7N5o
yIzDOYkV7kTqdfMv/h6qTuC2WNkRbb3Gs2poGQMZCDTdrrShwc3CK1KZckFg9NtB3PQTrWVgoEaG
cNVgYPwBmSrbp1iJRx8nsNdYvTnWTlnmVQgQZWyUdfSfyRfsRoKkdKgz+5pGIx9XfwzOUhKyKWkR
wJ2m3V5a/Lj7vVkO716PIrmT7veq3R5yRdE+h9Gwlm6m+cdh2hM/rcelmP7hCau26sv4vXuAfFVK
maRK80bq3JhqN6WANB+zpmHAXaijvnu/61xmit6ZnVcGiY5B9MAAR/0+R2OAEXs4L8oUXH8oibJW
gZTyDOIGmTziTK0zHvT08xDx4vvNpaMIn2BCPnCYQ96szrAKE68TrxV5FaJsClVmnL2rCeyeC8fy
hoevHYpyeeNAHj0Jx5MEmu7NKrzk85uzNQLpRM6C75ng9jAX4MK5FdgcVUYeZJxlvxnch0I1SU6d
yqlqprA3FO7QDGtzVp18AY93hBDecbFh3NI2ysgbpUVeKdja4IXQoGGdT7WAzyhYJ/6aQKG/8jZK
96B6ERU1UBm+zEkfafMwk8mrPHcfHebZAJsVlpEb4M9x5sQeUTJJzjAYyZOVR6QxzTyMlJT9erRY
oY4k7lTXii5YJ9JM5RG9Pgdohx9rS1KrTg+kCkakppBBayMtJis5DY70wPpfr2F28WbqbOUzqdlM
VjcGDHZ0bP1QhCxteOQ86g2iIoY08AT1gTV/8UnpPudOqFSuo9QXa1/AneNUUVhZUY2B/SG2V2Zq
UkIGFoaZk0F6uBd9X3ldzLtWbrjec/K72KndNvkJd/WNm2oz43BsWHfzguksKdjhxB95BUkCjZyH
XmrF/358D164aCzncjTRYlx+94Yc4VKEz9Y9XT4NRs7WWOvpMnP+qZKyH1XZgShnc6vieJ02p+ZV
dZ+5VOPbCuwcL0dJ4U26m5lX1cvJb3A13EpYimNlMWSwJRciGbhaqw25EL4fp6cFp3y1p1Kxt95e
TM3tZGJMdQdG4offAQyKlhAzkAuPXxO/ZdqHUZjEswgINmisYTFekqRWp6Ac8yFC8NlqDLTJNKwr
MMcqGMa3hdhcPQsWPVHtX+02MsDS1XdEgGJtejC/Q+tAODk8CD81z3wf30Em6RIlhWEi3mQqxRso
XcFDtU7GboALJPTgqKmO3kccGNtgoGmWDpie0RrJbkoi++316cDuwLOt17xHvZ1LMM1Lhx0zs7bp
Y7TvikpjVkDkkTu/Qa1pt4wmTGrd4LB2ByRJpuCfEmdI0CSHUyR9YzUwsNFQidd4u3Q+lxYsv9fP
RnCAENI2MmzPHN1Zuf5SKTREdP0d+nddyVWVKmgxA57hcA8pdg5GVsUjBokYdl0VBVEbSD2hZVI2
3hyFoMp/rbgaKMFUkfaWTnEcQxTIztTff6hLgEoxSAH7DPfYi0UkD9TKVwafIgC2vtEOD5CKAC5n
v6RmqIEZPpeQy3+YG0QPj5oPdiuXwfDJStbHBVzVo4cM9nSkoWedLOJY6pLJvGbXzu+JTJoXuye7
6jWGxv6iVDMtFT5pBz6LiGWCqeR0yM/KpXp89j4VLaYmzU3sqLiSXbSr8QUo1c2OmgnDf55M0dHo
36+QJu+qJgiXdR30dmKCN1tmv4qWjcneCLlXG7TFu5YDIp+bNnCDJQCWZ653A9GZqtVBPleK2NsQ
GlVvgZPnwSvgtjriWzgsg/R2VwGGQxrjQsihjkgHOfTYmtTA4bPFdrN2XPIUkmpsjxLOl+phVGBM
OGqpTqQ2RquAGb5PmF2P70maf0jGTG9U0kw5yI7kP+141Lamq5zc72mjAiQVb9BQhMsKYuH0PiPR
z5MneMSm/PYkm8hoF2CnF9LsAqFMzMBWc0hAs9zTfSzoByDfJ3hVSZiaTJiF3/otcncf7YSv/Kic
Q1nmb1RX4RrYJ5BcWkuBmOctln/Ij4KHnLldjPBXXzqpc//l3eN9nUHAsewisVsWbQ656lm1Qd0j
cfnLsHB02NKVBgoPmUXjV0uMloWxfcfm1axZWiaiszs6fhpY+gVNkFY0lnczXvWmnGRLCiazt6Y+
Q+90C5fCJjIfocZwIrqd8IrE9rC/vCuTbHmjeG7qDPqu+EzjNk2oTX42m2g1MPUo0E2yq968nMnV
3KLET5xtVNV2Y6mPmbNnv+Gf7sUcMpW9otvlBT3k3PufVkbchy7Vy+J+++tAFno23ooX0DD5jUfq
NgnISYM7DkXpDPWKyOuOUIV/X4SsaSVWsM6RJ5jTt5D5ZKf+BUoTHqDNMRu7FatrhAxs0dKEHiKZ
uIrdF9m46ulCVogwEb9Ai3QYHAfP35D+Ym8PufH472sprMmQbR6THl5tnjxlIQHeIXHeu+xLarhn
JQeKu/UxEmXIp7LYCn95szmRmKBpjSUWbUr7Mc/cbqGmS8lQQNO2uLyy7ptgjm1JUdRLDBXeIWJt
S3HFH1tSUm5ERhe4/aQUQkg30smnP2Sibf5k8cut9Ycri6ttesr33FCCx4XWrFCIDodYeqVbkf80
RSN83Aw2/SmAVwMqgHB/ZSIx/aeDGXYmprd2n9LLgRImh6LV1d+4naBGz7WiAMMWTTwFaP3NBPpV
W89mpBwc8QLm+LI2ka6x1c13FxZw1JD2vHOPFv5+3xeIcY6j+1LvqJ9lgjh1S7eU3W5Vk/F3PZfy
3e2s5anDF1o+F3wdcSOwlIdzgcDm5NN5sH3B8Ur+LnHmA8exE9RRTW4c4/kma5VqO0JPitO5tpLI
GSzXeC2l+d6K+g/CQtcHq/1mOL/3RWjwbPIxOkMPGgJfjtfYiBIfAVe+DSii2EfgKLMq2Q5+Aa/z
tO4wTl23nlL1QZccPeymVCCHQq0f38g7qoUSZBc50WFKvqqos6tGvzuLfMXQwjrz7kxAYKkkGOHY
MPHHmn1mF9RXoI8IQDUalbhbrqJeqSkQRm+jrKktrudgY+o7Vv6vtGm8E677jp0V20OCIUNR7ct1
Paae5Hq6T6eUqXGx2/Hv+v2Xv3qmQdUCWzN2v9et2TFvaEwFjZ7a173gjz4AzeWKsoKhG5rt6aBC
FtbBUaovBK+Pl3kaEhkWkz5imUpnduY0/LP0/HRVk4pVHYYveC5oseOP+0vVqkSRCO7zK6U1viT/
Bj3kOrlqaoaKwpOykwiP47OJS+VE3xC5tz6usv1hWmnM/QqbpMRS8aTOB5827yoIIWWoAOH6rf6S
0Jhzqd4lD/opvgvl0VL2aDNrYGsB2uNVcARFmATYCCNOm3/jg63EJdiXSVTFtob0SdGx/Nr0yPmp
6Dkp7+4L8/hhbrOW326z/TlyCRVOPNuFNzZFtOVxywyraxkEBV205Yzqutd7bdCQUC69BjydlkAm
qJfRYQYQ7oGiO3nMCVyO+vfpkYsb4oq0FZlD6tkZxDe75O7g2CZtJAymtmnUawG1CCQFzcGE9Dry
P4qrZolXPGGVZqX3XzqS5QOta/zmGiTkj0tgfsDGjskFEz6Ouk+i5uClgFlte7HHp+DzMTNx7W5X
egX/r9awDPcPo/g5p85QE8zx36przndHpHPVW9sGxg6Udt0Rz+CDWXmZ79OLG2ReJ+uAyADzGNZQ
3W2vsTZFNxfSL0PO+HOuUdJlDwMEySrk/pV0VVbjVi09RkPIe2ODDEJEw6f/EOJ7WfmdBlS9gfnL
kOH2S3d2KTGCAf0V4hC3qrXs16cnVmPY5+hsunRfw1RGEp8J44eLXsXE8RdzTmteTOqlAtOtTf85
YJPexsZ14k5dgFW84zXgW621dIJ2F5Q/EzVEbVyFFWciECtce9XAgW5xXe4F3VOY4uPLyLKT+QPX
R7OP4rxrLnGmcQeun9yDeg1qVbomEGpPRnLPAOCtGwy9McFVIeoWbdck/RusG9+oMkhJdzKHmSd5
hrqGjHFvpJozZJAL07YylS+Or7zXLXsi7+XoMuvgkgwGWapb/G+3izXwlEeRMZ+VHFOOO/Ku/9Dk
l68ya5z952mHmTzBbJlvauEFodHhgEMlSZJ7FH+0MWNvOx3DIOmwcnSSenNIHOTZ/td1W/RiP0ZD
e/KxQG8CujqQXnI2z+iCuQ4DcNBeuPcxRS/mRWW0YSlUAAEQ1DAUUsCNkWX136XXPFl2TQz78EMx
PWv22pQ+6xj3TPI6GaUkRA+XH8MWmvta74WB5JDZV3ooKU3r63SsTF/YtpEPgyYpDJuQ1dpgXp0l
iCXv7wlbzwL1DHrFraGNOFZ7r0W7zQcXdHM8GVpJd4T10Ngp1suQDNbmQI3z8MH+ciH72ohc5B2V
c9WyyMsBLu0LteZccmt59IYLplgUDexeGrh87b/G/ssAMj8d85R4YvwcSjBV2AxNnuInzdA4MANc
JWcEp20r+ouNUyrvXqdHv7pOz1NHMBLT6v3y9RQj2/rweC+NLoX69B45tzXvFKlwETu7st8wtGbh
h7EX5Zh4UygU2FL7dNb6jdOIZ/ajvWCYwkvN4UJPMjrRLaAciK+0QFjE5Dup621vp/RPQhd7sKl4
EvEZLhuHvlDhhiecz6rxOIcMF4U3pjUYEU6V9YVe5+3ghHjApADOj86cu8yDDs3/4iwusBDuWkrO
stMA2bwsx02mJu4bYCJrhWoAtGMDO700EWrjiifO96lyZOlPxzwYfjkah+Vr1T2Z7P9Ub1h2nxQp
pCW8heJ5RkE4Di+L8AhGpbLxCUzCSiPUp1q2z2ZX4XKRocesCa+N7JoVBDpZDKiImQEoIfosY57D
A90i0yprRpePdEEsgpDDPxJEH/sFYn1VVgdYouyc0KKosh1LB3kSMPdaZ/WebAwkQfxhsFqTYpQj
Z3L6jKGin3I7MtOd8CfMyXlUCL0gGWblN7J9x5hsc09u9AGKM5dgTV0Xi3hoUoq/9Ir453kgfpjx
w4OJDHKJS6UiZR4iwxl6UmVpEN1o8s1iEVy4/++o7kIDf3qen06GrtqyaQVXaC+Xma6DPvR81Usk
W9ytMROpX9UmEkLxlxUYc6t8+TFiRAhsJHPSuwZem71m//t8BkhYb+qDPvwX3mkn5f9W2REXjwMU
fNs7mmnnC/S4htwsI2Nf0ka+lBM53pQkoYdPKHBtvguL5YPNcoJ2lMW3oWQE2EYbxBfvS4DYRd0V
lL6I2uuujIZYysm6hy+HUCxDK5Pu/VtxVB0dLj0/l8gVszBQjbDgbhfGgAlLcbEMZwvrohFg8YMG
6/WTEbKBw2bmxnCH/qUOPqfSM9er9Rb/Xa5IEpXJa7JQTA7XInIhrqOR3YKkyyRwAFE2+aLo1Gek
OcQpdOc0jS1N7Z5bA+DZltBKltBMmrsLDKxiEA/9tJBr57MAMOHA3VWWeOii5g/4W2decmcNvjay
3fy/KWnpMeMeY22RPl/JvEEwHA4q8ZwtLy7p7EtkAA928XqC7z//6Q6oZ55eak2gu2oh/wZ/N/Y9
HI+KbrPmHfIoFUqrthog0CVLt4jRhguW9mVNhEs9kHSmB4uj1ncaMw8Yecy38C6BxQlwZvcGJVtv
IerpbmTiNR7ATtflFXs0Y+Ix2zybp6ZOixzb4HsZ2s1pEVQ6nbSXNID+mRd10kUcK+zH9vDXwEzc
bDcFbM5/J+0q5cQGvlgZP/cUKymGWor1Zr8h44OnkrEPbh+enUgw8ghFzJRnObbrs3ZMMv+kaPne
7V7tkVAXLmxx6Nyqc8pA/bklbC8kGbfM7uoPFtYNpHZu5GEIADXxBhD4KBM8Ggox9q7oH3EVCLZl
UbqDPFXToAmMs2GCVHphN5MeDHgtgRiKeIQPLHqGFZ3ClQ5M8hwNTYJqTx80htNmQCIJcZHTqiMs
XXYugDuPweknObE/eLz1EHPs7ZIWRJQ9tS7jRJ9euGox2PNQNiw53lCCf8GwHdyc99qDmIZbm+mc
fIKSTcZgC0SRbjTlW+V5Slgx2yoOfIjnDKtIRBJIiviCqXwLYtdQRhKLh6M4wAWGquGHMt55xwoc
23uXYYc/uSQ/VDxluYavkbeozdCl5vw6qM+8fUwlNquyEPlsFD4l+M7TXWnT3MkDQ5xWjkBupYzL
svvRbq6+9mlFcJ4XMMLZjCKzh/SnvNJKhOp+9ffm+W4rxEEKK5Q22dpScM9aB5LJlUf34HcwY5NZ
sEtKv2FF85qXz13NdnJHAU0P/lz27H3BGGF2+4hRJfH2i+XnzTgbg1rXN9xxkLwDgV6SWQgNWtKo
jq5MDoIvVL5RHrM+GAbj2odIiR1w4+VS0kohmzHSE9GP/HHRk9SbEYfuSUSYcs7hlv/uncLVTeV7
3M0u7Q4LvM7C84gLStZ4nLcq4B5gqsy8eI6FFB8bIOWFXAw3a91zweNygjW6YqmnQdICIkJMFLuB
YSTMGbSLKY2ohJB+BIedgnWS/9Gu2PPU9TDsAEyJYafpwzFNdSrtVh06wqE4/VbVFSXUC1Sb2F4Q
Nq2hbbuBmgIRZJRBY4yu/jP/DW85hReBw17AzhmWdLqkb6QIYdIpZvmNoGoeHUi1eiDqJe8lVNNs
Jhf6y7v1IDX3FeZGdgjDNQdvDOaRQsOcEScz+uNy0HykWvKy/ROD4W8zwrYDAMg9ymiLgPaVPvXy
fIukn9cfri+zemJyGeYh4IztpRvdMJkYKfs0/8AF4yqTkWN/TCw2OgpgS7gfLgqGQLsiBLbXjmFG
BXswr4lKVMXV++tZmRmRuxT/e0/FKl+E2gkS/lT/GAIo7X8nY4vKegyOgLadJtdIV/QTsBbYRVG+
o+yO/cR5nrXPGP0ei9mg6QodGX3OCP7wK+/MZChd80JOyN88zO3GG8b8R4U7g36XTf2G3+XorGzD
A1dCEDHyogiI0iAc9e+zh5Mfg5Mjupt4cZ7eWAG69CNyN5KxRsemrvV5Eu/IZYZI+u/4w1PX//B1
C8AW3abJKTdnAgmSBsY6eF0UGej+1oRLy1PyoXn4xTP3z+c+c5tAbJYL73jtpn+gGfek/Gtc92Gn
9joYLrVgGMmRIa7FiRonBqzKEgLP5QslNjWUBgiEDHmUR6TMl5d+8GRNQyET0IFgqU5SckehiPmq
XXw5D4Ir38Py5JRjIeoq7nfsknkArcfQdVia1rvG6PEJ8Gwb8r1uy0B5/EODgpGeecAAAWTMgxU+
zpRYNKeTDGSY616YODij5S3X+2GeSaAKdT5kQSLw6fXGMZ2CNNcEPzRJzjb+IiBPognVnMGWL8UV
Fb9/nzjbvMAN73SjCso5dbR6DrLc0Kh0s1OCHYXtusAd34k/8HeCW+ejPueQUiHNr7trQQlFcqTt
/ogzMn4abT9n0hddnyUkJeKr3BoLmkZFcGgXYFKPmtPXXIErzVgm76ljMPJaGw2RjPYZMF+wt2s1
bPQ/BN4GWnq0inoh9CBngq4mf40CnNbeuHjaLcHa0iWF1pBcawo5UhV+96dqIHmhEIXHswAr6+hZ
AwTTNi9b0oJbSsoJ1EjAx/8Cj/aeS0biULtiogYDqz5V7SYsa8EsFUBoXjGL6yALbGQK3HirT89V
LIe3JYw3KTicbzvATWiBmYkYoj28b1NdgzjEy4EgeFwNjMjemyq4RWcECZ5M9TN3eYuNq1Wp9PDL
Lbv1jxyJEOpUmZwiBCSoXiboDTryZ7nRxEn73HhXGY0yATSaE5VjKIjmHiqoPXeIjt/WEI2EBsms
0HIhvZlcnIC7ijR9NjxzJ2WD+b6O2mB3vxA2DY1mzk967cXLE6lTCuUIbGooVfEqiehweRitdvpA
eL1+KPxppHkeE5o9MVf0rVbhUvZlw5+mYFyXzSZHeor2mR2Rhl0zKmXiUVRWQM+Ch/iXvzFes/Xo
8wc6k3yCbAb3F1wMN07e2DZHa+sf5bhdV/O5JH1NmG4rfSk6c6RY9t4hrzv8VrGifI7YLfSLJBQf
ev6I7k6INJfeIjCzPuzRyertkRQ09+EtqsCw45ru6lLgLlmeuNdyTXOxQMmIr9+gW6r6pFN+S9jM
+hKI5hw7sHzk5VW580RWw7yQQtEigfhiSxApvxuOjRbm5qDwc5m+fS/xDe+zblFRZcTCQ/j9Vikt
GKkS65jYd/BecylyiYAKuTon51dQbxQ40HoLrWjvCowzZO4awUmHIix1NOMSGjbvFcjOmyz6AJZZ
ck0sv0H4UJg8GweH/41FjT7eV4As6r9DrEWRB9moR++q9i0T5cuBPJ2+aPwBzqdswNf3ObnOoGN8
d+N+b9CQtlRmE9Tv1lC3yu4NMuqKyWMw04l1bwPJdd3YYjte3mTcu2sr0aEPKxUN/4mI1E7ZRKYj
s+ul+/SQag9WtGS2O2yOBGCmQKHD/Ez2zggmZEx69wxCt0t7JMFNFrPPz2RCstYn81easbNyj8pG
H7EyWatTuU5uc/Zzpu3iQt/By7cZZ99e8wf+zV/kFJHJi5AI1r0iyKDL0+foLtCmhBU5dbqFnlE+
7l6wGcTWaBpnNc3GMf+WxUh+WINdmx0+k4DefjB4yPvV9/qxdVLmKWBGJ99X9Qes6JtPmEse0vzU
+bc5UO3vOgChR1BGIQXQhtwO/J4NGJK4we6Dh6jQHIoAlxxF/6CQkI9w/bJDf5WRa85D8fvQt56B
Tj/wZFTXb4CoibnR6Ns/kvi6UUnaur8M79N5PUslhqqnkd+yJuW3zMeT56/IMH1P/B2Qi+G6zv8r
CXVjTTkYv9k9HeFyadbv7y0wWfcC28MGMAIsul0haL6EL3I7CT4Fjq7s/W/fZYpZj031AQT/DoIw
EUMBYCcaSPGU2AG63oQnMhPikirVrqIXqxLREQydJVzvdQY0GcFfjH2vOD5/WfOA9RcDbImZ9tYe
1pt7Ogj5+KMynYEaadkZSs2O1RQhBbstLmOkYePd9sMoIxSgTyu/SoNuQGDHaBRo28qGP1YxOWAY
zmEk3YnvMT8pRGBJO7pVs/7Tl8NwVju/dtp+SL5jsTQQjGCAIntGfx/CeQL71aTk0fxlJPGfALnq
taxbrGkugwmqnkEU0AebzmcBQ4hz8gDCW8DknsV8drCqSPA/c8ZaEApWOkus1ab3vuf4wqUme2+y
Q0kOt/WysQez39csSW7AJNm+BtfgF7BWFt026UvOVTkoYcisKQT+ysBSNrdbJTUovlUpTtX7cK0s
yPuuAgT9IKV5s+iUEc8eYOyLNR5NiQe1m4vy9Wn7kPsS3j4xHFwI8DX8kXDuwX911rEuvJW0wb7e
NtN4bKYpvbRXIdxulTEr4t+F0HLPVZ+WjfLSE1MCh492nnyd6MxETGymoKvpb5Agahds6Bk4ZWQw
YwyEs2TvanGnELgj9nF0eYG+ftw20pfczkK7ggjCEh39Erwnsy4De8DLDka1q+TaKCQeNt7uSIzq
9MGW4NhtRRnA1zrqdcQ42gi+c/YXhhVad90EDlW2OxCv311ZR8+zF5+wrl1nDiG1Qjyzicv+eUax
WCP2koI85Ij1guwCeHCeT6D48Q3KCyID7MNPTtUgMNt2a8TL3IKX0QnOPko8hc8Otqvql1Oz6l2I
16A41qDG9CuVzFM5RLCHx/6ffoLq9PTijeRsKF9Zev9UTtiKBaLcfmpH/xkyOYtXeDZFMq2qJ4OA
ckAIz0SY81FtQ8MDtJ2NW2dlujqrPVJ4l7hwjGFG4hnuEPyp5GbjkPKLUeG7BEz8cr3BQVSU40SA
5Jjl7aogjxDB1XFNOLQkwMN1E7TCGwdZi7jp68ZpJTBovQiMYSPvA3bZqu55H8fX0qq+k4XVlVGo
idUYOAB4o0coCtDxEFr6LfbTkup/jzpLry4T4EmGVwavMnCQ8tmPw55iVL8BZtuI6x/zO6c8BsyU
gXq3E0V1K5YsJtzQK8cUhkd2Ze553kgkMeALvhOr2YmrcWBszjM2ouCn6jZRSmU5RZv8VMqItOmt
K6JVGfJOqqWapRgqdAI8QYmpt0O0vAJlp58Tgx+QDj3TYp39h9x2jDbvsZmsqTCaBeExfFTjgNKZ
fCO8lZ5jjNlSghiPko7HpRoaJ/Lh8/jA4Rk6aqhmhUyP4y1nJ7BqEGIwlQqNAWa7P2gFgOZkkHxB
9wm3afCYZk6qxJ2Jf3ZYcmvvBpGKKJGoWbQGGZFq89z5bgtnt8zdZ1geHw2VMEd5xLiz6BK7SQpn
6IkRKYcn441vIzLcik8od5tRRwUxn713YiEY90mUbKGp+eoSOshUMcy7i3UQqST8q/UKFRGFzqQy
0HXR56073fuz6vIEkCnH6iPhV2lpJUQyUTuxjtpX/YJutV19saaC3kuMJzWOC0VjXmKy2KvqVmS8
3K2jTqkghdA4Jc7v7LBATqUTaaKC9ucccuRDg4wsJssIbMyFHmVo/GJRy6g5Ntzcslvxxdld9RcF
2dkYi4CF4Af54aSe+KvXAB6MGdABfAv4ENd3y+W2XfnW+LVJUIdUYFj9ZLZy9YFfIO0df1H8TQK1
LQje9HEPJc6CrS781/5ktZz14s25VE5Lb05cwrz5p2kchUp7bV+0ABPlKuksz9lfQ5Vi5DHb9Gq7
uhoNctGfrh81PPBdVeRoua4jIsqSs/N+1fOFNHeLP49oTBMcEVjox7dHRmLHXUaQm7oTPZ0/ycq2
HcEqhKf40QwDdq5Q/gdndB+7IW1CwXzvPYALkBeh+2I7kIbl5wr8l+miyNvsgU6GDKZvwc46Ry8T
9z8qVTWQRwudlCHzx3gXv8vAMovViODOqflf/gJrwkk8pdV1DDoa+Dhk4O+UA9bccj5pxuR/pW3D
yIsjpRFNXAyqVolVUqaqTLL6k2lXQuQnTGFMmQEszXxz79TBlxHvcZM+WGbx38pmChez7PabZltu
X2W6C9yVioEcBRTSJBuBn1FxXM8y5Z9lkN01cZc2yZH261R1nT8/uV8M9ZP5V/6UOIgwAqSa10eS
ZO6Lq4rzlC+f+ozj/oFC/a5jmQXZ2X5YZ+HoOREnjt+J/pRmXK/Kb0zXWGeM3bgQht1RZs/jF7Ar
XD5eb0pa1qIRig3fIMKc6IDdhSQE6+GH2SyHMDdjzyI65+YnV2clvavzllW9b36+80gA8GhHFeVf
BTyX0efTl/USJRnUwYRzqHaNIn/Jw0GJvBTjc/yuORhE32LL/mgpyhsU+2FFzQarnbR9uuuuK65/
sY/kSQQYVAoLGzLXIjHc7FFkOAP38+lWRAPIFfcA6ZgWz//enNoOnMAGlk4nq3kf4jwMBD4SmJY8
Fu20GrJNko0VR1IvminwJx/2g8gBb6cPp6Up3HNgoy7/XpE9hnVb7hYGOfSE2a8VJWmgv8cnwUDc
clyRvS89VZGW4J+GiRbOsmabM4C9W2Dlj2/yWYEvQGzOiRjDpGBpKV8stzkmDO1mlTY5KSbSDQ0X
0tNT9onOAwVU/PQAnNYGLfifV1xzVIHmLYArbxqMpWSNtZimrGco1YDEPFghUvzHRwxoC5+PFk5k
M72lRHUy3sxJNh8qoPLDMwmimkk4HyxQC1mXTGf/v5fWDiYWPEJqbazixQg8jjl/fPSdytyg9rHC
bx16MFA/taJh5m6aXv+x6qkiO1uGSUFO4y9vVE3+UFhN2nLSEthL4JLDhZFgohaYiKWUmt63LiiE
/P01MeVRdVuUx8jJ+CVGKKgP6Meme+1DqBh/h87UHX1IG3kUulWQiqSL0MZARZG4iPkwF9Jr2Qa8
WXgfrwGK+BiByIlo3HBtNAdJpV4dPvMNBi+nL75q6l6Jmswk7uBhueHLpOkZQpxvUbst3q3d9Wjt
IqyPUN8XCxAENupUVAwETWAMRVCuD+/jrHzLtZ+2pL2UWgUj+LcMQ4vQwxRm/ykC9YCnQOMwXsd8
bArbv6uKV/KmY6C+aTbVDSoYX+lCHG5FkIG4p2fCitT2tfOJaiMfKasbkm4REccQUCDnNrxTFvRZ
FvF7Eqm9jNH4rICIdVThXNxIx30g4RR6gUwN+K1Fbo/LEkJFILrVj3mjL7lwt3RQZIr0APEAxBoh
0VS/r1h9DHovlMukYsP2ByNaZga+v910X7GN/mA1sSfco9i6kvO4aP7AEB0FevXj75Bg3aq2xC9T
Y9bRqvvNtHQzyNzuJeAaYVufLn5lhEXNwQ2cNqLArt//US4rkmXjwRHxrCvw7JTV20lLpzKR91tS
oaX8ED/J1qXiXY0iLBKevbr3hJ8w9TeSmg4GoeMn63lAWYSFZexlvdrlMvXm1rvPBCDxwIcmuPm0
Euw20eO63C/mxNxEQS/rJpBRQ7oW5/KKd0KXJYISikGSGrU3Dnm/2ZjKBnnCX7NZSBcfDTYsUbGN
mLsn7ezFXUAqP3R2Jr9ML/39S4Z3E3PIztUja7RsCvfbwa6HkA//9EqYgkyFlyfsCUvB6SMHCRAZ
egiqXY0ikFScuL3QRqnkI/7xQjOgbAybOpJf9SmAEYRKty4EeIXAAahcprNglgCUwnJ2LlXEV6a1
4QH6vA5kK9qZISOv0agxVg+h4MRNI/Rkz4PAb4na8OftQbUCdXIKc/2PPr6Q34lksILRzbyZlyzN
bJoRFa9KU20HiU3UfHy7180QFCNr27SAgdkHWUW+budM1cGS+nZ/krJe95X5nZgOewOb/A71gwVx
vggFJgnkhl+w8YmobKe9spE1LBbQWR+Y7B25VbGUqjHf28T8Fzqjlp5ZXcvNC292eGBV1hPhSZtX
N2ZcGy8qFD1l8VSJC+IbJYPa5ofloMvkzllQldHUnG4dO+A5Pq9wIzQa9ZaeZGrXNNGnK62asjPi
b21v3EaPRAxOt1Jz8yRJveKTkDMcCJlqzB6xw7JuCD3yrsQNIgLprj7WtvZuW8MXVo6CUJEkSW6o
8zPaScCsECR9tZMAyQ8ic8Uh5uoqS5sgdJymRRf7epksRZ2PLmP7tT+C6W0bKLp2qshoA8fe8v7p
OyTYZ6naWmis33zvGElOWakpXQbE0oJx/xXIHaVX+RTxi+3+AWvCqpQS4alkc8fZghmGM9KQ+Yl2
RroC9r3wqUvJ30LBVHFqk1mRN53Vp336AYXA4KfRWJW9NPWlU1NWRC15K88Q9JOxTYelUVBI3Sgk
Z6CIXVv3KKxs15IDJLANBNOwuXWenw64sERMILyX7BbNBbnpdsCCBDV5js37EIyQqIKUcZsmee1j
tYWvHUuscK+YFgkImQ6fw6gG51zuIraN0e4nPR9zzmpuXM3YI0c7qPorZAXAF1HP8HV9K19N8WZi
q/iwFmDmWvU5mgt1Bqpqy4pAsK4k3kjFtNXFscnETwVpqvC9imoqnoXxHlu4goHCdttWRK2Lcnj2
zRVBl4BijvElbYmAYDhlHAOrfM1bTka2G+N9c9G6w+MTRUBqw5Nr5mkCO58hiPA6PXliwkK0iwQD
TMrHBcRRS/ZcTNkVjrjLRwhLpl4HmuHtuBzn/D/13iKuDSXEQkNRBnh2GGWE6RafN8oMIw8GSmHH
XD7wL+hkcyWwPdHvPbOTF2QixvjjssE4oy1yzrM8Rl+L9qDXDmha/wJwE6kq1mMJwDdN6gUDf7kk
0IF+Liqx2ShBh+FFUHCm5nGyC7sBWl/+aWyozIqTcbttqA9Ho6YOF38wIGa54pipXRaw8WM26j9D
rV5dqOoMCNCmOikBLLS6n+o2Y+6eBk38tqPLVHEi9s3rmGarXmI50b8ks1h38KYVLExFO7xdjK7y
j0ILObQFRElt4TedXJZP2gIARd4xRKNwezdJjelxh3hBcX2v1FRcns3B6Sd7xvkn9n2CGKmyzH1N
FiIj/DLbO6pHhN/NZxL6vOvBt0xbbmyA+PZSdhvReEGNjhb8qkPmbrBfFsFuUXujSDGU+b8lvCfN
kse6OsREJdQj3XY+1JlUk9FCYy/t9VlGdrC6Xd6Q54yA1kR9Dm6WRrMBGGXwHVc0GEYhO5fcvZ0X
CR6Sb+yAuixNSgtm0YJ/+PsT88G9WtnJB5OFnlJ1i+RqTUoF6Bih3j51bhhlZWdWs0kJ7k0AHUAF
j1e3FD/iQcb7qzhiQOT5vGUfZJhuFAtt1j6gD+P0tFieACZePvBg8m9BFoujm0XPO/PxiPsoP4+/
XK09EjvkRh9e9m4rcdlEdGpG+BC+68qAjh1DkxSkJ2J5MX1d6IgvE+ldZogfWKCsG+glOwaEtAT0
PD8MueVXZhRtW1OuqCOkG6eFB5cWA8SUYredVrbWTg8KbcUGK00IJYtun7pQkmo3rKctZd8yKTgZ
Dn4sWiMNqsTBP2uDvh1F72EyyrYEQgHSTu9Izjgn/b98WAEYOpav0fox6yLeCcdCReJ1jONW58Qa
4kwpNlH4jam1QCkXYpyCuJOD9JAdvz+NYgOdJdcO+JYFdjosaDIh4xgeomHAnapbE3Gvk78Adppv
78RTC8m90doaFdNFslCYU43N35xsLquZUCaemkooH7XPXD+ePH6nUgxakYuWeUiMNuowLFCD+9vt
haORqoQbWsYZvg2apuNJN8mxXIT3GCOsNws32OwDB22r/Xs4x70FhWCAjKIUzDkrkL3yZ/JaYrrr
su/btRJAJKdnUr7lyWkLgvSqC3y68J/tY4xllo1cNzhKgndkWwk8PO8fkFLuc/H4e5IEwznEanAQ
qw1lNt3DaiqUQpHGWmj/ZP/l5Iy3gX89W58C1qBDA/Ozom5KzE/wz85ijJ7FCWW98BNFmVeHtuTl
AEV6txnEQRMhnDLAwodOdpVzmbmjGniTjA3eWvHOBvGiEu8vu8FbJkTYe2f2rG18+z2LMqNm6Jz6
VggOyZEv5e7bAouRH/ho1mDLNSgNDUkRPyJUTFUr3Ca/gUnqcLB7NsJ0RQ5OLPvCwhnU+73I7voC
p5/XBVJ+WyiKYnNdxgQbgp7n5qrx+zbICiLCPi96X7mIll4WFdULRJa+vhSL6l79BVKszXPXPJYX
EYpv0QogOnZT3STMd12PTFrGODRs54P2vLnqkh3+ysFpKVsig9eiv8TEfGbBzGBxPkXgXXUTYbWs
gs2C+4XwSQGakKAKVZr2JMlRWEJezGFkPI7sRixnGh60VHGRSMeg4v1aJgb49XZ2WGemYP8rDOrk
NYPh3sgbV2NoAZfpRt5E3mKZUsOPN9RVZRRq0skkJcJw4Znay1PVaDWg3TPhzOdhw08C8EHGNZ0F
PKuk7H4QwKQb52t+J2eUAmVoLM3fI3/fkFZFfUgPzs0PwkcytW9NWLuXvbqRz/2hS49FT+UaFbQy
J+GFQsB86kffWniXu6gDVHAhc1WWnTCDywN73IF4Fs/x3mZ/YeBODlaDaKahN5RhpoMX/rCIW6Tz
rV08tLijEIAwPm3JmFZF1HPGKKxqpzZ52CwifCG2VtEIIRlxLqywYYwbwzVaECctW7q68u31FZLZ
An3BTXXiMtn82iIqgP0vhb/mo8niwYlzbJGS8Fizpo+s60krfDe/YntHnharsF5q2tyucd4xhMZi
8NGQ02SZP1vgqnhrjUF4Px1tRAagx7dBrm1G+zCC4jJMyhaZsi1JHx8d6SmCVc2fXNXtwjXk/MmT
3dodkb2vuqAnfWzHjxtaidNtDpRr/AU+y3IaPvMe8pwCyUDObXTOmU+dTpMat6XFcv41Oh+ayQ5S
+IlAbbMu7KCCTLBD1Ej+W2TMbxuplMbJo18gphCHC52tinvbi1iEhUpqbiXgP8A/RnlGCtjm4h1P
NDzAO7dW2JpkLOzbELjWD9P2JsjV3CvpgKoxRHhE5S+r38IAHNpFdfV3Rc3V5F9OUlxpeIhFQaPX
KE8OOl3wOYYom/pKsmsbaeyH+U5/LepE+kTRLw3A0OGg6uaMtx0nXSxojDzzXDRNh/WmHfx373W5
7o/iMb6Snfwy9foJGaklJ+sx4jm4PajV8rf7I1CGQRR2ytV7seP6gDgDIm6gbOaeMLkFUfG429/5
56GT/tm1ilL3n2albttG/F1gMatBy2Z7tk4vj+bb3LwJf+VrxokGJDF2cUaCupWAc6KBcHDA6MVV
ROpOwXdt4kFiOv08UQIKYbcR+uZmGloBJXXuQiH4kcCxeFXGqfmFNYwIS1V9th/WKW/Vun6L2SXH
oDI6nLWVXh1AYWzxXDjBsJ3b/NxirDQNeKbAQjfH0CheLJq3Xoiov02xBxyKwkEC9KZ6KQ6Mt5Uy
YhLVUGZrs4+41kYoNeEshLGOX9IkYDWkxq7VQEklEXmTE7nIOforO6MWYitp9gvxCcsaXMWWnIVv
eOGiD+tR3M8SAWsC8wQ4nH7Pc0ky7N1ogkQwHO/4WD5/OA40GIRRfj+txberilvH0AKcDPKXXIMo
fPL4CQgQKGQbAzNoRc7x4liIlWyFQnNHfEh3m3rJjwqbLvOiAHvKXJy1ttyF2dtY4BOSjSdMj93N
QbzYMfkG5m+iU+mvmpLt3WxLeKq2radoemDqbR3P5BvAbwSu8jBzLPkUuHSKK+Kbt26yjxA+idH4
78bD94uDkjlZpwnfriWzirKaKdr6AOycSPWEvcELrZsRuaLmG1TkyUvQvOakDfyuhzFCl3yypt8y
kTPbVymQsM7wZyNgNC6wyBOGrY5jWbNYZRYOROD2almDA7oCg1Xvxn6xcbuFgnYAc8C1OyF/rdrs
dWUIjRZnmBqujH+PBu102erOW5CCEAp5GGLAW3gtqtZtOFpRo+SRW6xCQlWEtkKc6RlA+k5w/a5Q
8Zqfgs4PcTkxfEsZ7M3r5/beSS/C/85NWmwVQHngHRqzcDH3d22+PEOkGDt7LMiy/YHpY1fbQZGo
U2w9IT/AQmvA3HtP24wKjm9w/04sNsAiSatZZbtcdIudm5IT0TEQbwz4rQnzMAjHUj/tKRFiIGYu
dK6G+X/QyfaFYGPMnSdC0y7R+HTQKueVVUEWuQIGZJtHgSlAgk6zyrVxxx5luRBbdC6RA9Ag+vh4
vda4ToTDXVyLEdcOZ2PeIBia9FQYFiBFBAHxJCWRP7TqyqvmwoXq2e7vaAygsi4xVSOv5ZdbJjUe
kU1bej95oqwevm2PG69OL/MMsfu/se3u1jj84g+oWl2dh0u7WsviKQdivO4VZLRbfjVxlrth7e7r
wTAkq1fiEsPoxBB/mypMhofh/R0Eusli+jJ6MDkzyI9DCE5CZjIgN9EPZvbcIP1nI+Z8tB+ku/ox
o7IftvJqIfWjtQl1Ieg6YEK59JLbg0i+YzZTTyIDwoBoOs96Y75d3kVSXEger2F+mRnWN/FILEzv
Gbn0mvW45WaGAFgsFjpdi35cal5fHt3Ic1mXKQfqz0lIGIFK/WrkyR7jynYovUQSkch/Pyms5A72
A7RN4Nx1q+vynPSKAjwz+bMkWaB1TNcU7R7tgtwulZ2xlLYelaHHPMwfVD2pcdStHyfWLlr5zuWt
ZMfZ0UMkun/T+rO7WeYg7iuPDKEwcj8/kbjoMe3R0zLduP44QEvnifu6HD8/5fKpcjMO6P1KtGqM
ZdWgauCTyxDqrdkldhM9Sk9lSAjaBdfKQEcXvy/Mdf3I8VK8L1to5zYSUfbWC16H9Qi3MbvbfCzd
0XQul6Q29mlkjotL8HZilpc+sO447XzvD7audl6LQ08+66BrFTUX3qff/9PMvrMFMoAorZSWzG9v
ZShYOmWsFEHuS5391hkkt3wTDmmLKo1FwyO+rs5yHs4Gk0FtKgtF+3z0o2n+CM1Nm0P+/dhFCX+g
NKIgDFLiqxJQV0l2ypkAe58qM7S2EHNdelEgH0985wPeuGhcpMaFS/6/m8KQP1MtW98IDs8flDYl
zpFk5fViyylB3W/uQjC4rtr/8T3BmZtH2fvnxMnz8/YoRhiM1yOQx4mk6p7F4QAClEIzfIKtefym
guC1cUNZsRS22Awbmigez1D+h0nEXM6mJjmH+Wwh9+annQLIDG/ApmnKLj33ze+rZfYm4ZCiCIE1
beyedsarFeHXWWq/zJTTVuOsB9sT2qfz7voAWhuC9FaT41fGNP+877Sg0BXVIKgzHr3zeYAKJzBJ
dewUprBFMORMVPO2NC75Vdel6n5lPdHkZlg2ymBTr09y8Dt7x496cHTKzX6VTV8NmmbYodVl+xq9
KkbzzQCXKWh/8EnWIqDieILa6h3AI1wBjs07WB13pEfS8xFnPXMMg63m0Bf7Lejn974Uh9kHSlwB
qFf0TU0sa+ePWGU/KzbERleq9+FeFsuKIjJp9zBrR/P4D34z4H9cQJje+JVkQPktvMFKcsUXoMef
LPkS3BwZ7L3hg+s1LHjfctfoXn1piNArpwwNjibU/Pt3SIZTl6DiB5R/sXVfNO29kzV2TJy6VUpu
R7Hut7gGeMf3Hy+9fZyJgjtnhSJpyj2j75oZ5gDdkhKI+aV5iA1THjDDNwvK8pjoVEYzhyq5U1F8
Sr+TNXfHz+saSGxXrB5Ykm8C+bsevCg+SIxEYENMd0JAgi4mKsRgLA02xHCLChhS5kwtolCoCjOS
2da/C9ggOAOJZ8XVzfX5HFbrSEMFoEA9yQzKam2EtKIHxSWz/JdKa8DypeXxa86kxeDlOYuRbsF/
JkycNP1zuIgMZby4tRpcuNTOH3LC3Wdl7XOPn4LfF3FMlC1dB9CB2nPata2fDkPQ3lpokhCHl9a8
dkvyw1jDfMXksyvxusrHRrJPBmajb7ITnvrvBhR3oslMbSBrZ9Y/jWg/DWqz9rTQIAcV0rkcgZQd
l2+8WbhTAhHxFIE3g8nztpELSN2/yZrtVvaGqhsd8z5yhEYNSBVfizR10ziGmZhRBlCrDy1nGPp5
+fOFWMZlldKV35afn2g2Dh0Q2SOerT9gPKXefbFIekQVS7jOZlQss3rFPFLjmFYI1/N7SKGpA0jL
VXjEUYTCcfvy4GwKmnr9tkqtNAZFpdcB0MhrZ+2gsR9yqmY5A2izu1qEhJlXhQKIEi/m5IZ79FRu
6GSVefaSnXuk84dlc+rRYOjtq09/60UzcFAlrsadnC5zkzRD6RhEcLkAPIKj4C7woFRaz+Jvw4FT
4wqjgFsAimWxmpQdVCbUGiHekHg0l8s31llNuWgAYiMb4sljbYZ+yiIcKurKln3fgqtDtomjgRnH
6MA8ZxpqSKTm9F09qyt5VUxD+AQ5himY3elUE2yY5eTNybxcpSZeQLKenGKPvltZ7RCT6Nqxjxkh
bznrLCJpwzdkragX7aLxlWcE/P5XkldPaFEqSFhht3rpntuirwMz0BfHKKaTWTt2eAHo0h3mRL/x
ZhJ+L+Hl+EJeVRa29BoWVgP5KqfiU/lS+J7bk0wA6V/Bl15dMiND3oEMtcJZT/CQOosPs0J/Vs+D
nah0TazTZmC+DzoW1dy6Zpiwm5gw8uFJ2ll/G8Vw1d5fgK/6Kz0R4mfDwub4es4CpnYj3Ao1LMZk
p3VGASBY7Io+ghgJ0mgAYPUIUAQALx9tzgiFscPn+dB+47fUMOvYv1nsRcRT5Km2ItIlqF/vCVC1
cIpIif9aEvGHH/6BNi2m8Q6lYTdVCeyJfOv38RpfZot2UAJGHe4NzzJFuG5HzHC6c1keTO3ddD3k
B1ADzRPvf54xaE8pHSTrBTRwDWyD3ct7tR2xsHlVx1s0eBt9/QAb0fZmeBUqOwXSvBKLMQGbu895
2fK1SKaM2XFryQL2qqvwEaIffTQaOElqQrjJ6Uwa5A8W/JR586xDCLfjMZgyIT9SZb2szioZ7Vcf
x889VhXEN/RZHfIkDWGnqMl3QAiN+GMXPhGBtRoaz9Yvs+EBMg2i/3M7VxAuZZCQn+CbZmoIEsaj
/XFUt9eti+b77Pxb7mlmbzTFLkj6R85qEu/Ornm5Q10fBExJ93atqo+HfpmBJH/dDmGQpDiI8dGK
/7JUzuY3rDslmPk1NwLUTzVghAStQxItBSj5QEojr+FgnOmkYIzlVLu5s8ktumRrql06tNxqTLUT
VZ4Pqx66eZu9KhanZLBqi0ln4qpEux2bcPV5fDsBg6n6XgJPAc/Zgd5fnYw7qfDKAg9OocwQPBtE
kqavc0EJ/TdUuUkaLi6evjKP7ObZ41yH9d4PNJC/WvJbpsGhW+sUn4xqyq77x89+uqMzfVDINGlB
+DtF3zh4WXMX0elKfUNiGA+BfPQxrhBuC1WQsIrmFxD64uFLzM7zOc42a4iUjHyDz1Q8uw4fXySp
P+VyMdhoeBczZHP3q2XvzfKx3hQ5AUs7kVEeHHqN+YU7S3GzDhXfIT3tcZJxTgOCern8aNJPowX6
yJQzAeo1xr9HJXBD/tcLALzQLQF9x81hzVDdfkTz7Nl8wGNOhGNrM91lnL4Vo23w7Yi2FD3iLRxI
R12uuqoKMt1V3GWo+Gg7XwNTn82UmQ6F8xwTwK+nmTHiCHiNiJxN43OH0c6FoBeG8GUnmvvj20Rw
T0k60ApsnoX2GIQZDh1QUafE00evGUDsO97trOBGpJgp3f0MENSh2oiSRA2NQ41Yg4LVfRGm+yQk
RIJnStjS1925Oz6xID89+8DW4Ilizy8B4vGwPRk46dCgISTjoXztgdoaXPolvGOch2lYSSegTZ8P
HO5OTCfW1YOO80kkYRg6rX7yJNcXWIUVcuJqolkSCp1S/IXVxhtbBayOwznbnDzh4n77IzhyH3ix
NvLEs7rNXT5xMErtXi5OmYqYfBJb+ShYmqJBm4royWrsNP4ST9FhDuQ5dtOrHJ9lXYsZYazHP+KN
XA1xz+YX23TGcwZkcgjQdZrwtnCKV7hE2dv3uTbMc1OaUQY2iUyQRHTXrYWzUnnNyInxIDJ3ojEx
Z7FuinvYoeQtoX7xi9h/Prs38GP36D1OIxPA1Nf25nnrZbZrr92WcQhoPFesJs/h1dyU/mkJZPXb
njFhcu+CAqYrSUObr5AqwvQx+Xt2Gk46QOlXN2GsJ6ZDomEGWo0QZ2FfryaoOWwUWAb1upHVcicw
UbtVfqlgm/4ILUy9tImgMI0CC6pSl9b9nkgEtTl7qiSWQLGnDRJ62U0ulyGXShj5HMaEBRz8Rq6n
rrDDm48Bu1qKhmmRt3asg3jDAnz7scsLvdbzWoEJ+X2HnHBdt0X7h9SDiCW2XMQmtm7ZPryyAIVy
0visUMd3W72IHTHtw7mg7OJZ6sC/bkaxcToz5pnjY98Gxnug9S2NyAy3MhoCFUMLT28xHghi8bYt
ihUQzEZsBiuTmYiHX7vRhVPL8uaz5RdUTAL1shB0iEOWg13h/k2dT0Kvx89/OKOiACiSWohZ34UR
hNH/EUjhWuDaY546nDhTsi+jX6Tzurggz6uJIkHU3vhQyNESmWbNi7Fo5GnlVCANNeatq6kBoxiN
F6N53V2bnva+44LjyK7QeoXqeMS7jafXl/QBHaeU8pEdb0cCE5Z7WJ9ocswtmXfx1fOMSYosx/Q6
oqbYdiklFFgG4yn88xMhRIj9z8ZhO1BqaQ1rxBVjLeyydDywEZe+CCXZpPpmJzj876fpYfXBl0O9
WxudOngX/hmD0ecYy/NQNSrdv0YWCH1tEQFSugh+R92V5+RGsZWFumrPIwwir+jUa/DwNd/HbOch
9fcARO9qPK0mlobZWMakQmyo+rgduhhZhMX6YRWIizqSDjCbWK9FA8H6cKf0IneLLEl+RZIvxNm9
bl6Zu1mN0/Q9w/e1NhhZ2Mlus2d2AAvzmfzAAh0fYl+llvRCFTGSiA9m5gY6JTGzc7GbO5pSzOTo
rz3oEcH7O6mFrAEMdkKx0iDJYM5m0JhJVJ2ffXE9yM4ri4hvOVrvtW18htvg1gl7oXrHiR3UCSy7
81FpdQ/xi2qshS0Y1FBXA2MTHDgGlRVa5Q+jIV1JzFjzspB7o9adqeZCLUKgD0ly6PquR/yjJbwl
HJeCzsips8zcCF/5oeW4M4u3kDi3qA8/bYbg3tCBhTcetNQqJb0L02zwxz8YHSaPoKtx/+i8In2R
loHTTxm734X5d02e4hK4ftRemXaz4ysEo8YYxHYtqYdpXgE8L3K7hkJcoTgQiK5Lt1RgSz0wL0aS
Fn0ZC7UKQppmhV8Q6SCVAUjNQvcKs49nFBU3W2IOkLH3OyvqMdrRGhSsWZxA1BkjyQw9nCx+WZik
CTEVrWq6r+IOelxv1481c+OhU68azyIUokQXMFfnjHbWpGH2Sv4y8XDhXrV8QMQToGOGrQqDk5ax
NJp9txjgtM5Y560ARJUu2j1MoB20g/DQa91ou/HvCJHiIEcLULaUQojBKccvqbJfYMYxm55dkI/d
2ll6Jz2QQLx4pv69mCRbQ//3+kEt1qVVodhCAx72qbq0OyapeDUfpv1WKzYbNgvsQmUbk+GF6pUz
MKXKpG8PWSPNBdL4yFUUMJe8M7d7kNTYMJbMYhj3PcAIL2oBdIj+72bUJ1iyR2wmvwjLNRElr6eu
4HAJ/xdXkWfJgBrGiPIHVqCZ1GbPW7q8DzWOgTIhQiNbzMQTklNLoPJHrdejlXvnR5jwlp6nSeDU
CFHzpKsMeK+DW8z0EAMNBTn/Kv0M2569wS87/Ql15oAFjc+bzyYp56z05qniPvHGWwb8EtyJbQhR
LRAele5TkD6VL6oWYO3AAL6jqmpGWZcHATouTqu7ZjuanWMbXyfkDTsqnpIdG7tXJOtulAHHD06v
7JQPKp6SQsL8WErJGsm98xsvIGp5+MO/O26jp8hCHibei6Uo3/MOlkHHaDvW4jIHADMT9KUXW39Z
mXEA3cyuhHyQeOaHDGZ83G89fR2EB9xCMAVFUOWDV6YuY2XWqkQ1b0vKfb+j0qTY8YHNQan6zHTM
lrh+oc7mCVHj+BCWPIjcCtK+gwIbSpSWc+r41h0JVTHHiDzVM7VDPZvNzMrtJIRdapBx9BMQAzOv
2ckS67+yML4SR7m6fkS5YaNFdmbGPGdcpc1WI33M8dRvRDlJEce5cIrQ50e1Adv6Y27TnFtSfFWA
xZfQWX0Sd5F+81tif8U3Rs/8JnQDV6xRdHVWMKRmTeUePDKb6ZMqMgDXh/4V8VNQdIsNDfeAFmRK
Fwg0G1tdVpqbGeGH8uv2XNVi1EVBK8g7XTeSN2BPBpyh6xvpQmiMRg19y+9RONxySBOof+Dg09Jl
/G41UcFpGkIGnah0IsIKjkQJeJic89QFn/Dxn/Uns3ZninBd/eppi13dserlnsWwmI/34qhSNHT3
Q9tstynwiTt9mbK80W/UqM/Z+F9V/n4NWNRP4LvANxxL9GisOZHYAozuJDN1aZVa2/ovXtfuVoLE
otm0FjPKIU9egEBY9Y3fNM1detYhc8hydomp2+5gttv5nH4+ad/rm6vtlMCU/L/ys/yeCDauFNDr
8LkcQI9RFe//W9hpxfEAuZiahYWhBaPzjUqe7+hkHbsFNb8tdPtatHavj+ZcgQD1zLpi/xSD2VDi
IZxXZv3M0+mcDLBT3FcAfRrUU89fZGz0srOJp6IXo8KMtfxKjC/az3R21BDvm62Xi3yEZcO0VHJ5
0cvz0SuYJQVtoHviCpPPfuF4JKXRMpHsoxXR43NnPff4esz3ZYuF1zvIV4U7yOyDPTavuSWxmY2X
tAhnMmKg0cWgGwtfHqMcBKxL4GmgXgor3wl+svFzgrYq+QmYyEIYsOv9OM9DSsEfY6nrlCvSFlvr
BD0V9I8d2cE0paaknbnYW0JL68bSPqRqy0M2E+ewQfwHGtC9EZD5+D7D47WPzAQG65YOE8pAI/oF
c2UulRVTewxNyDh8ckz8mJeL/NUQX6uXE1eZa1z3UKYPsi+r5HmshuTIsphsQ2OtOV5WQl1nDLr9
I5+OIzMiWg805MVTHrH18mmtE1UUcfB2Lk5jCrRpSO3ph04S6noM77PPztvI5kRJ8upv6M/ab2lh
RhcZJKYKCCC3IC+ihvsSt8KUKBrjsaxhnuBP0Un230R2vou4MtUPBNeOf9Zw2CJ2UIFo+vbNdION
QWTbMjt0otUqf6eXxYLCntYdJgDtlmA8i/GjfNqN//WIDSvByt+RXZXvBQempjr0p1YIAeOaeHRQ
Jds534kJvwzcliT5kjkjkuNfqGExclmK8W3nW/QrKiKyxVSxLfIKyJOUOsBA8bLf4/5QrKjTYaS2
GtZ04y71oO3GZlnMQHd+IE8xVMfHJR1zV2C0FM4KOC33ST7V0ZTeT1bdVDc3rc8S7/4skIalzjO3
qnqXqt6SIzWMlZeBJhHe3OiqtfWuD7zimyys64G4quuHpOcdBYohu6Ss/BeZSlxMjPO433Qs/Vek
/OGpMmAT6NZBXVQPV9HoXySaHXESMngH/xPBaf3ezxiMYaAaVem9ytL6kQJO43TPCn4B/C3GWlaf
k44Bbn/quughxY4B+BNWIgqmR7DP0+UMJWAbLjLxdUR7yO/M1vzEsHDL5/twrDuGHkvh+WvFxeGW
W/GAH0dWRd0e4QmQ31flCh0R/stR+58kJO/J+m0WiYloNcgaBNPoD+uFS+cOPRIL5HrBpJr1d+wf
icxZHtxquY6AFeI25iV6FG0hdr9muiVJBeMdylSx/VPPobO8GJ5xJ8qNsoInWFx6aCsbWfHot+dw
Q5eBU/sjRSkvuaMIyrrWFQweOIs0LwooH2fBv5igiLGh1YLsA438xJ596KfvpjqRK3s6pkpFMHC6
4iJRtfTzo+/CZieLh2/ond54sPDUdEMYZkbHSaEbe28b4BWzqWWDzoHuUxTOQ8b9/sNwJqMiMu66
QalB8cCkSqqYZtyRRfLl4UtcC3a0lYPaLbRZMflkVBZ78ndzkVGhNoWGT/f2eQfpO2xPEAgY9BN4
JVIQ7GirsX0e59t8k3dpQSCTQwKdAb/sjdj6TLp5hEiicPUjEBGhL9K0fTPdkcM18XNV0crLI6iS
J0hVJzcBY9cT/tZy4pQOK9wFWxhxfpmOQ0URZAhxdx1fMsdCfpYGX6g72zgYIpRf8oDvbEZXJSkr
NZ6qE6dZVKvA9fcu6I9vyWA49gxemCPN+6DUHvaemPsPwVzUruA/rXoCdNqoYQhmbCt2OWAym/vT
jqtj00YBvSjWoPPyMriSkLzARt0rMPgtemkwAKzYXXZgrdVNz9na32kT/fiaxbxKyYPB3qGQzX45
wNeaPf53vMSMToWpgW+gM1UQeTDuFOV8l015MQ5NX+9RzENUxU+V1wgymjmNKigB3whAfw9C+fcI
xVQvuYtn0eE62Qk0dUu+E51l8Fle0uUm5Q87GzayYfyKdwD4jfafRPwXwhhxNWHEIN2pmxtA98ie
Ic+atxN2ecEFFTZ9Ofx5CCA6cgqRQmWJlVQ93GAxsCSerqj9Nibtjp4Fy1mFxGo4DMUyx8RR5KkQ
UioYtsnB8pI3rcZW+6uEd3Jf31qAg27cUXyMKxFgINV6jW9E9rx/ObXVqPEmLdnC+llTlBog+I+a
iFvMDkvVwis3ctivHVQCWmgiYs0iiwKZLas3hsJgvwt7gCssI4EzWntmENHS4FsIFP4rzqDa2CpN
prr4CYjo08lGZEADd2gQp41Pqz2QfZCNiZiq3YcTxYtz37wjiCGAqhD3rfyDor/dZckEmzyp6MvU
iI5OLTetNlr8dKCBFhk9l8xp4QCezcccuYRcyJRQB2dcAPcFbXVIZHgGHghgd8RPjR34MjJhDp6u
lz5TpP1R6a/fxiLK/qJg3LicyRCpFDn3KXaMTY8Nh2RJEbs+p6cdwdg4kiEUn6PyaCo6+vcBGghi
xFNfM7h+XrJ+bGgrO8TmI/KaMYIY9wKqm9HVTLa11OJyfyw0Z6iRmv/cjxlI+hUErMKPbD8y2SSr
jkWdvl1G+bPbZuU4E7O4lQ/nj6QjDWGc5eIy8HwxAF1OG8dLaMtKCiMxsDZxV8OiUfDZNBxjBO4d
VFhHHB0rdnMbZQDkTlS3L6pe0e2xxHkFmH/TRj82/yakjirczotJ3upjZHyx6ANfdO3K0NfUiNX8
9wGbUj7pRbJICF1/QeLFYAggBGZJf9rXCqZmqtaClv1fT3uXeN6FUrb4+P8B3Cym71IQBq5DN1t0
szb57xiXDkxVSkkLrf3TpuOYjGHbCaT0r23FKKaTFVQxeZ3qDo8hrVkn7msIvNhWd2Z5OlE0HVmB
+3AwewMjIpcA1g88VWi12UCwhnrlijsMJIVOrtYT5zJvjl3Fr3SMzKnMia/01QY2I73ugTA3YxHc
EEugtrIGFeJ/FqpTVpjF+rMdmr7oLXRfqQMKxIvb4+q6vK9fW2sVKg903EeItM0Gbyl6CZq97t32
Vc4nJvZ+ksh2yAziM0dGamtDX/dqChGfDIjcVJg2DzRTSSMJNNpngBAa4dkBmGPDtcj/qcDdQgf5
28XQwCURDGoR/QqpX26JdFGk2OYX+D6QOLFX0i/MwK0gWNoRLN6vddY99+eKfUeUedacQc17gXzD
NALC8ny1+fqm/GKN/5d6UY8HGhFlJipZ10ow8BZTdV3rvh7klIpkndPvOdovnwHEUjYdZ66Ffuqg
8VizytYEe35KaBRPyP9lOUQtBWJojPYUFQ/Gx6pPID5eddqpwQ6ctyhagwvD7SLT1Z6kmt98/io5
r99652kabPM+tK6IYN4kxdDO/GDK5E0RFUfQUTbb23e/aWTQyix7ivGb87tu6+RkSy9yZveaxa5j
kyWCbQu541EgQR3lZGiq6wlTxKwslG0Zhe8aVIDAfkRKQrUJpPgXhf5u2jSP/HtFz55MirmGo1lP
3edEL6Y8AIiS6rauWBxQH5KLGKOMjyARZDVIT7bSuBj7VROO44tR0J4N4bdEABMVAkkXKw/HdcVr
DjMBeQEnWumJ5TpTmHonH5hv2DqCp1k83BKJM8RG73SEaL15KFPRD6cVj2U0YeddenMnGz+fJ6yu
VxD22IxSDvvMYd2P1RGB/exsC1kg33d2ikVRztJYofY8k9812gJXQlDStncwIbTLSh0vMRPPUoYA
E+0jPnd+dydMo55qMzsXswpyv+0/K9MdoPnWeAhNzDHDLGJdv/WtfSqQMgM7PYeQy9kZ/hUn+bmb
8fOKCe3r2o+3NBghEtMDR6g51zmdzB5D9W+P8T9hsGEdA4akQQxsbJCIA4NkuqNHZKN/23rRCVnt
nrhM5b11Rc5ESmZT1YkAGI5whAQcGnGHLL7lQsytv6JKfVnMtYV/SPezpm6+/6zbtwcN/vjIn4he
qBYfQPihwF6T/Vm9CLMd+MNo5Rd1wMkCgbBXQcKKop+v6olHdlFWKjUMbUPzzBAXM8STfOnFxHQ/
LjAw22aq9XAOZRA4t2hnqnsSRP9UqLa6iuRb5/RoKZ7R0Xbvn9X7Tp/Ytclsa7PwQe5iiBDcyVhd
z7iYq3skyFPQF8Eiu8jzRyHWsnjbqjFqX1iunUC4bx8EBCud1YRyoYc1jNyYDxx6SYxDcwAgA9Qi
qlhZPqYDjotf09D2yQau6dTr5Rf+SpngxIryIe3eYP4oKevnTZl1kt0g4O3ITccLrluqpBIrzJz6
1xSeuSmRyxDZHb9j97GWPRzrci0FxK1v38n8oQfY5QgqFlQZ3ef4PqUZlp70/7C//aMniSdDmFBp
uxmm7ODtnNRZZA51apW1bSzppowGxAItKQ2AttuizU5XXmI+ELPUV463pqJLWITe3FmheQp1Q7wI
w2k1QJ+ZBEIoiRxTcnyONlzYMZ6kLeGaUEFHmT9XwrZvUNMWNe3BIP30WEi8LFcVoWBOWdBsKJsd
Rp5BGk8r+o0z/2s2fBcGiP93KVM6+jGpu9V9vptM6XVLD+uSJLtfj7Ut+Kpw26obfk3G9mvQqy4E
GRQtaF41XvYg9xmcF5+id6lfpHndPp6JHlCiMvH5e3TRSpDXHmvEp1sMyIGDV49SZBXkgVavcnrD
oyp/JXVFplflZ2iNkq2bfyj1AhmopBsXEo3TSpt61TmhDlgQ/tBdGVmiVbervucIQqHvU5l4Gj5g
XDFSv9qdFWmCcSZrbyF0wg1QaTYtfotw//nw60ZYU1x1cHzdUzX4eXJUfSwWplcLJhGX/9qux6sF
UlFzyfSMS/5cHit6SpeLuZ9Sq2ifzVdyEOXoCsXyrSokSo9C1OJraoI14XxQfwZjXnfyj0/Qpeph
pRkkziPAtzRcl0m3EfFXfQfEYJOF6KkTANdqNRC4EaUwK4AolerWRWCaNmgsWciH/UHF81WFdYHp
S+yZ+V896OkwRH2jaNQKG0AX1ANNk5qZjqi9ASks0ZHspOme/Cl3iFGaXw1S1eUX/NTD90RLpgJh
CCmvrRHwbcLXPjdrmHVFhWCWNlkCyG9I3NjxUK5/WzayjQtiMuGffQBsMKHqDyqrsNeZofY5iKLq
qSg+jvKugKPPwDo4hToHhJClqf4rsQGBqC3ME/wLEtvpbnrWR8r6N5W0LaYJ6/VvY6LJbhSvzG20
LwFEgOHn0O35CUpnhL6wFGbZ46XkyaqMttPH1gRosqX2nd+Bk+S6bY2qtpWbIaIuloX1KRxYwlXD
vx91z29z+/9QhtjVNiTmmqvRNkfrNzJfWB367YPAKK1bTbQ6JJ6ioQ7mf7ZyauSF+kDtXZIpq/lo
rslj5a+N/7qlM3bQrKBZaewF4KeLq/PFCq2VQ2hgyIFVVR8jVwEAhtFu2F6nr8G7JbXTv9X41PAW
cl9M/wVaRKz+cOhBWfp6HxT6Nlw8fE/dbJH37D7rJzUveAn46fqj2qqxmOEUTn6xSAjZuBFcvFYs
at+HvqgmTlF51UItdbaFEwfIE8Va5wjMAS+6DkSWHXt/QQ0BS47MuKccUidt9unt78WOhskOg9Vz
oa8pAzcHSpWGDPTMwwheYze5w97GwQf/neKHtDSuwoFEMzv/XVZwEPeusZl3bNw2ggekjpS/HEjd
sLUKYz35mGD40MtJ2w2QNnVK990oQ9KQOi8j9gNX8e0y/0YqFOdmIXRi7HcZb7lc5BAN7dvp5kb7
47ikPCp2YVWIWn8AwvpI42J8UtnJ9RQaABPdjafnOe4nnMItlq38rLC+1ff7UKJHTR5yZB+C0kLT
t//Xv2g0wE0xBK3JXg02CFpnlP1L2LpZ/PS/9QSfQIrgqG+rnP9k1Oqtw26H4o5eZATC/XIYKRlo
gPA6DSdEJPTlmjVja0qTnxuyWQh6gCpTTfNkNdxVx2Y/NJJCWiE4RBn/UPjNR65uKC9fhvzUK4tk
2cHRUai5l6oI+PsuUHIndo/qurDxZgvaOcJIuIcurmqSnl5+vH2zUuMbInWL7kPGK8QRWIbk5zHZ
V+ZNjtQOOJyfj0inmaeP8XzRvZtBX84YmPFPpS9nU2qNiHYvnNFqtCD0BpEAv0tmlbm0X97/oHT3
vOIVAxF1QrG3V2nNZqJ3cXvdHc0iJO/QiGYmnYMSCs4cv69/j1WBO2xNXeHLzABuqUjW9DdrkXNm
kv7dkZ2DuyKujOVCfUSYq9KI13HK9UjCAuLppflwaTEsakPwdFDtVa9UkHgPzpQQl7CRlW+fA0yO
VX+9Y/FpcYoqoMS2vbTRNHP8vWJmyNAqJBzjHQytHdPkeLm1hWCVuE2/jyYJ4Mv32vRPXV6tdG0A
4Jd9N/Iuhv8aIghdAfs8mk5+pgWyLoPjIcGQH1p1dWRT5hOqbH0Rv5sBdKjQUSi633Ke7dkIwVhd
jsfgx8JGlXF+zC+PCkGMPG70c3VEP15FurrzBeuYoyxibqYvJMjc3ny/SBhWkqXh6gr2u701TGG7
5nW9bFLrXj+KDTqvbORTS4o913ES1LTBBBjFo2xu7eZApPX9JDidx/KsHFl38toxtODsziXSrRNC
ceMfnz2nDFF2ECMIB5QupeKFh4D4lMnbTdO/R/+pOBhZACPpN4qbQnE/I65OX7Gz97nNpbPQ/ki2
Yhnmj657V8zAKCoc02JHSUG2P/u5xBIGPpRdRXyZSARu24BS5LI36vMyMmW7VFrL+pbvOEII29zS
LK3qhdH9+CMNmZWL9TjAQN42XxDsNjph3jZ8SseAQqaXWiQ82HyDlFbau+BaBfGHyPSMT4Cco39s
x5LqgDK+QY/RAfe4oDgI1RSVhg4/vzm08FGhZIrorhfF5oWfqm/0w4jqpBl5I0Oc8waGbFf2+TX6
v69m0IYhaoESJi8yc4M28/NDP/vgurIcg0FaECPyE9jTEN0zWuJSAtEIVK4VTpfBtVDpxdabmBoa
fRlcYB0/G/DqyxMrZpBzDofKyXxZDNkHISsXNrjJBl7ZsM7OhBTLYWgu4SZmsQv8ey8lxFrD+l/S
w7EnJJV6MMzq6TBgJPWfFkkGKN8hq1CffQR7rctpK5e5bN2Ko79TaF9t5yzwg1WXjGqx+MwHsAJC
pzmGN5BX3VbL4liHa5HtA7/G3PRd4X8B3cdtlUHwlfdWunZhTtcxkDjmRjDELpDTeE8bje/Yv3dI
fcq5najSXY/UOjf5lApEmMvc2l4IaeXTgUDboyX5A2W9XFSNJNH89v0EF5Vcb4Uj4G6jOIfhO7Hq
pJhzIBpdqgDiLtNkGUeOHnyFXzeOYRESTBMbv6nvh/AUUTmmZbMvVAwGkaQxgmW9zitNP7wENMu9
HLjDg36mg9OBhWn4WGQ2bESPZeF/M3bDGjZQd5uRYj58cmn4+QPgbW+lWnhpqAGDEdMB22937GQr
n4l6UaX0k2cGRZ6QPjB4ptQn7N04SqO98ht0iPW0lWzfFl3aXVbEqkuOUzhDLYqnwChqNizXgQT9
YbHfPHc0PxUo7bNIWk2BIbBtgKm5hdypuR/2gaHDSIyf1MWsLpJLpLTYX4n7m/sENWuuUBHmvpZw
8glP46Vu8Z7ZwCUYz9vj0FpnOU7OUctxb9q80PuG8x07J7PGpyeASvlQNd8x+H4tgBlMulzCdLOj
ehy9+33L98At+65kU5wnI+DNqtXUwGm9znH6pMK0tnDVwfpVcyWGSGTNARqpjR3pXpj3HklSAyuY
LsMlhm4hHAXXj0wzKaZz7JUK4iHj52HSXvdy8YmOCmUjfx71wdUvfwngX/PsXgmMJsmXsv6wlnTL
hdM6JZc24euzB8uBGi9RU5cd123zA4UbV6Am2f6hcdpmynGhPDgRvGcp78hqUwc+VSPTdp1ah+R9
cgz7o34wjdpkotSmXVWxXLJxUc33cFpxIX1WfAmuVYeX6xSZZKb6mH7nLDn+w6oyloSKe/uMRHIH
n7B73sXG5+yjTH8BAaa81YczxbGFwfdP2eENidJYdIBud3WI9JWtZOYDpMCtksbl3WgcvZt9iPMR
PlocCSqZ1k/ta8JB/OhSs6w2Vx/1W/7aVtbNdxq+hPPOc+gJLuNGPMWGHAsvmLblc3AIiMVE6VzC
GzP1S08hb/gO2lM1+wxVBKUbQUNUyZpIoij4eZ1K9pfbBzY2rRL54yEZqF9BQeOpSPnKEg0XUC0U
IMoJ8Oxh4wUFz1/Z6n7l5/NmlYuaA8MrAOl4NDzDNlfNoMX57t8axUuQbVzFXM3qX/x9RYv0jmNI
XfOtXiZJrWxBtnO7iIm+kBvHN4REyv9QihuJ6sooKSkGbkXd+EQ4dwryFJwXR6sGrun+PQEAajYB
rvE0eNNiNJXb9mgowOITl0uIFn3BIV79CEwGDmUPvZdcSm3mnmsmiciP1IgjMePpdq/2V3RZZxuA
RnfwOIIKAtoE9CY+Zrw211m+zHSAKhdaeGRVatTkFdH8eyBnbXyj8c2pdTQqlUsDTW1Od1TDqCmh
acI21zIP6yhc12pl+ach45a9HQ4ph3LH26HN8jLJ9f3661rOv98yRtQyV4B1nCHL8nafBGx+bqip
jmc5e+kcMJz23LligXxq216Lqc+vHS3XXHDrTgREHhiRoW3MtWKHJvPCvf9u1lPMi3mpf5mhk0xe
atxS+5Ibyt+n0tNxI0yVZxXx9vYCC+MU0h3yleA30PjqP+FW9bhxyCs4JaQWCy5JOjZLrqnRDZSk
OHcpTmBxGp6RuHtWbdhJRTra8LF6kQ62h7EgrNa0aGpVpafwev9J0lt2ii6WXVU6+heS9UEZTdE/
dx387ARJ6is0XdUgTGjnvxCLvrMEdkEFb44DwXu33e1WhnGjIOBAM0KSQez9JdtE3JwobBFh790L
bxQBjM3aHB7Rgx77OSmqbqs6+GQDnP/u+0tWZrhEY1kc28cO1RRllRxzPs8e5eRp6Qop2mAHbA1j
BrxBKi0QOi12SId7qGriV45/Axux0xfYIIkzsRatmCCQLbCxGby3z1YyJtEQzQHYdoFoxkj84r2h
jCIOU+VlUsdQUHqvBTJkyU1jFzk4S39STk+8uoxcnEKeCcMIwMTMm6IZ/RA7FP1gdE4J5fD5yBkY
S0rWIJIjCN/P7onUTWClom9bs7G+s8VcqeadojwmQyiAP88R0dQ7DUW2q7sptiSolQUre7+KMof0
HS0/eOL7mjoCPfsD978jaHeXq1844SYpZ3RQzHJnZz9uQheUHpd/52vqPKr+qgIENUYDprYX1331
zjbK8niF1s+c+rPcPIS36b+D1BrTxlxnF6p0gKB1NuO/2g0LLngeRBNn4Rjj4IcCJbEvnscExRgd
KQRQzHWgLoPP8cR7y7dL9bhku03NKIlPKdIeJ1lhJETHY8f8QWHFeXX7MMLQAR4kvwRAxzM9FClp
CBW+sRUILSrl8H8HQPaxrpsOnVCbsLsd8lXJSS7EN1h1+PoWEKm/FSukMythn9ElqWiFox7haRTy
amrix/W/EV02TnfLYBZ7X60NKsrrKvnh9XaUf3NXTNEIdkm7+c+7EIHWW6L8haaaAIt5zCaSoVBZ
3zJyMZE0mjBVVayv9F7nH1Kr9xSt6y4XbO8YoRh62jtZTULwMuQUsNgoJRP8GwA4MFENWVrxvSHB
rwYQJ3Fg4OqbYF+rEiRfY3lNdc9ZkQTNgwhBA3JL+Sk89MIrEbnG65pMQP498YKV3moo25WVO1Ka
MfZwT/8sST5sliUOaQOXs8cabS7bIHeQgzc1V2+go7Kj4kuZ6kgKGGHRHT5wVFQZozlQyVHtL1XP
U6EbgJy8Xg3qnOrDiwaH/Rc+rckInbGN+DRJ9eGQCVHdo42ISr1pwHN5fHGOkl6QbYAsbYOaC7Ru
gvntJOfD/O/QTm9sEvFsSl4ftMpHkSmBJhB6aXXNZjKgj1SswJLyS+Ha26o/daGcvndBsQaQkI+s
cEnKXvTWgNxrPzIF43Eky1PseSRzw1k5UlRlXheXK3y4NK5S4dO6xBgp1DsRuEdM3jdZVTm+P7/0
2m6lbfu0Psx6XZGld7DsAWni6rJwqw17YAI48wEkIelc8tET++kTg78O2VChiGcCboe8J8XZeUP5
FvqxYKBrN8Syp4Wgzz+nFuq1LdEw5n+iuActs9mxYiWWapGVtLmbaRNYPfDj4JqGeRnY218Dil6q
UyB/xa5p+eh5OskU0rPJmSy8/3EUcKLs+F11Rw0HqSC+H0JqnSrX+n/yqS9CNEroiSztj3BeC0fN
sendyW3dwhEi/Hn9xpqLqrh2QRLKJ3s7yxdnXPflmdc5BdhfORyCiBzyCEVg2uP+Yc6HsRDAKzvR
MC4prHBPRlOAphh8fCYg5/TCRIKBcHB5GltaJZt6zLkU5gMkYTdag//SBsS1jMJLz/bb4BaXyudC
F7reS0ACC3rwweI9K5muNOtpY+KDhKFs8a/GWICCw8B7xb5BkutPmia9jnx0ittjoJKsD+8au4DJ
y+mEehJ5yJZ+65yhqN4ZcKBLU8SMcnrcxcd0/W/V+wFVg/UMceoLBVaFugQY9n4XTL/QGwd1Btzn
Mk3xLsK6qabu6DiMqhKfDPhYjBRlTcpKLWuikoGgL71oCaLKHTOpv6W+IADmOnV6fqQhnZgbrc1e
2zgez1HZMLPVJYjB2e30zW9PwxCL4QQ1IfOZyeNSNOqU4izoNRqQTBwp5ejrvy1jYnloRQLW8uZk
SX+ezImxkZxARFxHk/t1refu9bQim9Zcu3ew1rFrtxbhFcqoK5bbslHTnsr654sZOa24LJv2Xs4q
Qj4SUv5EKwkqZWxiUaop1kOeHtfMi9yVsqICGTsueiRvlTCDed+wTIYcDUHWR1l4QH0F4gsgv1ZN
/A2RvTH8ULetTLyrDJJ1FTy+wVkuxD9eJMsRqaRcLpRR1g3by2e+mZa7u+IdAP2vEggXqkX7Rwxh
m08sxKs0Rb0cz+1mTFVAKOfPFitdHQ9ny7FbD+71yvY4Ctuiz/WYEnmSgA7QQGkwx8mb4xIH/h7h
9WNq9Tvuau1gXHhkdqbsC8sh/6vqD04yvp4M0nFL7xOHAxhRGpkFotRlY+J96rjRUD4X5ezPrJ9K
fxKHpezEGuHJhMZi3yTCS1dRWHOILXSFcc3XKHmxARZo1xs8NFnG4fTBfHr5Ml+pcwfHGo+34lC5
8V4DMs45L1DT8sIG3AXRG/w+pmE8d2rdI26yxNsVk3+0tetk5WYOxFKC8JbEc07+W1ncnBMI+z+s
DoiwZRnwSHJSyimlbXcMKFY1qRzhEEv4cOVe4aZtb322avKxyeWIiaJDIZ3jBvGWXMg62/eSM7Fe
69tmhujruiTmpOoWEQT4hu3qw6zHjCgo62Y62HBf79iS5U/Z4UWgjIQK4PFiC8w99ZXtKbc1FneW
/Xni9rqZmXOD2E9EaSBNbLmwC035lGetvLXd1MKurunv8C+XTDHyZ+3AGuUJdUXnpu/OyUAAGx8r
20luLSO5BO0peVa0yhBVo2KpKMRXNjn3TVQGDkTDrAW3C2IHJKrABFxY9Ogk4zz3cVkyQL4XAfLB
GRYd7/UxONZopFOPDMPSHb4FNyx93mn7tuFDVT5+6SFibPAabY3iXxL4EgkZXYlOPxdZSCMhA2GZ
2jQyexgvgoyaNT8S3LpSpqRraDD0kK84dYf/Re6UKVrkGCyX/t/VJsqiybnZ4yW4DXOSQQbKuqKo
ZDsqV+igV3UVTX5kFwejjCE5OHl1l9eroRGRFRXTQq5XrKS+BFzB5fmFhnyM+mn2XX+Yqu+L+tZk
CI1y7Ih+9EigT/3oNZLOy5SYbhyN9fsxOEppvC4tNDNws7bc1+tJ5E4JbIfxwo+NevYdIojArwRa
aCfG8GmYxJ7h974Cwfrud3W+LoLX8my3v0MLZBTNq9MP8bNaqoq+F0bHfsjdExsN14YAZHWY+ZqE
SbMOkGj0QY+zmOFO21bRz8kcpLNWdNkkfjthRPdt2Wgah/1DhEC+zB55QeTlSdNQZCE4jggcUQcR
5bIzIEFcNG4prf2iCKULhyUz6dFkTWQyJWelQ2s0C6frOMupMjG7Y6vmSstyODf4oeO1AMMCkrb4
Ghcdi+/UTLERY/Sk2DpQkyQhTVon0inAWUlT8sDl6WQs0bKs3mbg+EunE8LwwMyJtnr6ZSwubyf7
PDkeP4VOJWUXFBd5jbZLWBd8LT5rbnVySlpWkHoApCwB2aDkAE15YDO7W5Akvj56G7cJwOvm2VXm
VXHStL566MVFPfwDoFUE36bIW4Z9MVsRYwU/SuyGDoDEvnkHvO92C+QBe241rUg0fKYdhTpUslTu
fhmfO9N4t6tjkTAUYffkhjcK+in8hZ01j0aBzYalSrCpJY1Oh8POtsnOWYNDZ2ukVDgFmsmwAqeN
aNLxM/RzM9IDkT8WHo5flGL0LyKOreL5eXTfI8UCakss6D1dpvXxE6Ius01d6P0xW2zyqfiqDsFm
BNsbKTDIx5V34K0qiG1iDcmpfBAwI/wOwYFKXUAxua1vOmH+jpdhfrKGXuXE6k9QIRkscLP0naIt
xE14XhWmlaC27rtyzwK9kcLZwLRDP6KB8agZSRKHGzRjM4gZIn7qIEqO4bY6qP1oXd/0F/CpPFsE
qj4hofDLQYUMGk7KUwPtXi59EVhDltnrbW0qy1WJzosud6ptm6+5Jd7ejCFQo5DZYvq1Gz9N5a7D
U0UdauHNP2+Iwf01ZyzjfEI+zidGhXIJDS7GT4U6xFPZPwDdGvTlMdGL2qVSZber9f9sm9G5E63F
J1pESXcKComX65ctKsPaLXA6B6ZlOYF7bNJn5C4nv0Q/Q/yVdvSjAIFXhchoxUnko+aS2AgXIP2u
5RE6HUvnN5k8O39iadpvq8SaaGfjZH2U1ro3Ca1eSo1L65hRFanwUlusblO1ulZ/qbj1dcAjhoTZ
QmeHeWvjFnR5aBFacATz8YkoFavEcmBsfdrScuU5iDUTWlsZnoJZraze27Vn62rCrAWDutgSCzDz
Kn4qQlzpqJQw4TM2oS3Cv3Fe91ibqgx0LTpkp/R9dgI/BRh7VXDdSjFcrUHNuFoXPIJZuGAxNBlG
M+BFy+4fjfe8BPFNr/jRHPNf3kArnMUovc2tHN9XbMiUb7zFcwFQXoEwU44DxD7eKdEFTGn9StgC
gl4bxfyHloAVU3Yol34yfjKhUIB860VJPRcMYlh88cSuj6H2J/PEFQ10KohlI88nbLID81Hu4P2l
C6UymCAhQOiNKFIERmz/E6jRuukrPTy/zksYtk4ymquMQHK2Qwx05G10HTf5h0dNGzmknS9Vvb7w
jX0fpzxv5+eI16qlZ91GTw0+DePlfRBpR6kXKV3apiGpGDDGDtAGVEAYQl9F8SXqUU41Vcl1vZST
8IWTXfdDRZTSKHaF9CgkD+Pqos5zHuNhvr/1KGHEdAbED8s8skSHPkxevdrWN0+RscQf3jr2y+rR
8Kgqv0U2/Kl0yDO7qW/Fw54GNa/zv2GNFDVowtKrkJ968LqCSvxF1CPeeXr2LBso5aOlEbF/sJSf
a330tLAKpjB86DTBPDc95nblhmWlg1mCrsklkfDx9++LusPV4fRUkN5bKJy+gbLtUzv6i2Wlmirx
aActPvtExEiLCeOrAnhMJ1PiOwH9Qtl22wfNr+TE9wEDlBvLfLEQ6WOFRieJf2nTgrXLAh1LI4u1
m4IBfJWgw2bDuiD5t4FUAV+DgrzjWsvPH0h4QRf9Ka/VjuNBGEHo/AVaLH22INX4E/g6KE2LllZZ
fZ59043WQTaVxxrLu+8QvuLUDlKWZFY4T7khJk3umgHb5Cg8GUh7ukPO18RYKJaiu03sxgwrXNwY
+cUKISuJ7LptVhTtii8xKKaAw5xemIwdkslm3l+x4u9RhG+pOG7OJuzNMa+kt7yDYwEUAr36d2RZ
TYFLAOr1uhR5dXFJdVl+HG6pU47cfrqMlC1G2wu/l3KaC+U8xbWAVrAKm9JwHbOUKl4e3+++2ruR
3SVLEHYSzmkFrOEothhcSYOfkgEkOUy3P6/xBP20nHxCrXR7Lfq0wk2fOGTNqZnLoeC8zZEo+UhF
HeWDDrtrKqZHc7+6DOV9QRdwv4lT4F/QEhamVOER+LXr8ZfXbWR1GeFRwQZdwYUMdftylSRxnoO7
xKBb3vjx05e1ecq8Ui5zxieZiX3rxhKfJWLWBeNOZtJO7cQ7amS0BDIfa/R/bQbatrYbhgbzmU5M
3JFQI0WawNDlFr30eFvPFpDsn0gH082eNe5oaTtTHUffBy9nXzQJl03ujWvGTWeNTJoZ1jkln9Q8
+lfUnw6B+pWFZq1dsO1PkRVpUFKHObfiVYJJiDcKxMeXHPByIgJA1BZL57GIndG3azFZX95a1+Px
3hqdQ1NmyNT3kLVMqmLL245KlzMbSurbD9lU1ToAWYU/uqljSK8g5Xx3t8qZ4KyfNo5hczWZskj7
nK/GQ79jE90ZNPBRDfbEz1b7/jhyK+Sy4p3VJlvaEl7Y4ZPeiJ+q8b/AVikSgUqiQ9dD0uQuLT+5
/Shq3ymqrGHToIO18gI2DJX7ywOMFK64juM8swvk82pN56VMi+9wxbWfs6p+4JDF1ViJRj4lr/zt
oo0nsK85fK8D15HsOLTEsMwJOXGz2MHj4B5oyHQkvnmtCg4d4e7tl3wo03ZIjHJWB3FH6iL4mfkX
Rdwj/8SOv7fQf7aezR8OJ9BU1+iKskLHehXIu/gag4GWSceIySHCIPbz0dQJJy6cTeJRAj7EaHX2
ojOyhdLF3rNti/C1jGT5CxkBDAzFCuEoqG+PcRbJNjEfPhLvhJ38OXjVg7Kw7oywZ1OH9b/D05h1
Wr7iWhtjucG9UhkwC5QORg7bJRKCNEzyaeALwAwLDNakrfLtYe5m7MiszSZ1Y2drEKfqsjLeVUEB
dKZsunsgS/TwyTsCIwnsqZ9iFht6Y5WC6KFqo8bmAtLJogNqHEujbSUapoN115lH0zoHgZFNxLdG
S7XGEFCHm/HZRr8bRwpOWnm1uM30AY+85wV14vnDdN88XMPuUSRYlhHNbuZy95vmP6vS8nsq4yF+
vW4obYHB1aXrEvSPl52ktfYDqBZfigTiDLsp6hlVhhgN6PqG/wmI69ACaPPoykTUrCB63cblc0Fw
Qi+tlKEfTy7Au0brcvp23mcYSOiBSQ02z7QsQqx7nfUMgNobut85KsMuOjna6V6r088Etv+OMXNl
vkB+Ald4doeAQxCW0Dv8ngiD0hWuSlAiuMQEKqJE00YG0r0klqjFWQyu3ZX9A9OFWLSqlx+nPoNo
OporF2HLt8NqbdEd/74Q4bfqcW7XDbDyBdnOm0SzknD9ME58f17UVEpycugxptXeH6es3hBkIXlc
JfCLrqtFCp/0uuCr2nBlAb2E1En76XzfWYiYCyPtH6YPi0LtEUF55IaMhFEJAc2cdwB/HhLdeml4
FvpCkBErdW06KGPHKnk0sZXyli96RxPFLopkyxXv0IwcTSPi6FRj0N7abqJCkHdK0bEbjCkpxm31
7kMeX/TEUHINJjHI40/8TXIG1/C4LVV1CsXOGYb5yUheAEtY2kjXizb7s5FHSwRgpzc2MDEP2YHD
JXH8JzB1PU0oPIp0tXv9uMlSDXOfqeqGN9yDWWXG7zEbqkgAJYBuNZO4XmfXsLul3aeSAlyrb2bc
HihhsdLcsB1D1haywWFx0298outNuCTS5mMm+phdowLp8kWZeDWmNhctCK/Ne9mncAEqJIyiCpv4
4F7oPK546FDTMWtJwtlS2JKEexdgjH6TyV3WN/YRSWT2UZxfYssUwtsq/kf2pVrMXfWy/nR3Qdns
hyragFBXnITmUPVuz5VcXGKJgTCeU1PKOJGkktxX3KDxedhZw4u3LHSoswO9c7e1uvdYXUfV5eA9
5Umzbnj0CZomFwx0JM1qYohsgVsJgapYzMhPgbvednRuvF9FKtlSYf1KugORiGbK719GIEqR+CVK
w+YJKJUglJUSsxHsBl1uVdDVQzOJYujqcWw6G2B25JCDrS/aGOXxqRCSSxd7bKPCj6ceqhh6wCKu
Gp04zHSs6UQ0t15RGyw2qloZseYvrz5YF+fVb0ZaTaFPeROTcJPvIDYX82FghTzrdoAx2egmlNYX
lEvBOSg2gmcFKW2h4mxaqE0OACBB9jgdIMDTQ6l6EJZTJ/R10HE3IRjSBCWlViGi48mjHS7OElni
fM+QTY8gMMKDhbIDGveLEjXPUgUcE7Z3rE727w4g3eRy34nWcrzW2M/NmGVFOHhud0XnlhOVWYG9
OcEkP59fwfFN0rIZk8lrVENpi3CaBS0UYRdckYv++O4b0yB4OvhbEsbu16T1ld6OhcvGasWEBWal
BKx2K2KKT1megHUkla+X+sZ5NTJfm46sKAlqk8c4WsrW1M5mXhLLRGuLmc3gW7kPG4r1muAllQDt
u2JJqQFo30cCVuCq2OeZ8rjIg7VcZnX4sqWJzsAeXf97RjuJro6iv5A2Cp6UxcPXep8mGOmWmdiy
RtcsksHSIAU7jYvE7t3Xt7JFw0T+ulp8O59FOY3JXhGyuSL1w0rca0kQUH4hIVCCiEDXRDrGuKKu
42ktNshqUIuF2PTlJvjhixn8ZsTG3wp9b1w/Hg2c8TLvS168SNRcNzy8XZWwbG2gq5m6FvvCceLS
m3DzqT3gkJU5lqgl9mE36C4NKWxN1pcb4GLwAkRUrwcJyvt6YtsJoFYsNAjDDLptSMRsz1fBkoLx
m6kdC451sFrRoQjf5vI6o2U+5nik3puYf8EgcmeZdn+4q13V6TTdAmDK8XtiOAPQm9tfj484mumI
52aPlkgI7rRe1NEgWnLcW1kowxyQx17EI09XW92Iz0yPRt0OvN/OEo/zFMsU+qezGrfN4jRDyV6y
t1KbMcn/0zfuQTgbcrMJBCj5IwDrrwEGi6W69Y9BEsu6B4QdlfxpZII1fBJ344QiDt3t0rpZeK4X
4RnDoBaKOfGYgzYMb/WwIJpkbGkTBAAPy7Xr/TRo3NASLnmNdB9erUWpiNrmb0b8oEkgPhxrxyqp
YcAXYaFBoXF1UMR2w1nllAxuJBj1g6MQkdJHD+ddYQkvNsf9wJXtJxTwAwRp576WgXm3Gos3iTi5
50nkgfZVKPoUW2ekm41dgJmEPUHxGclPMLECUqAhfwfMNMfWMGmwLENCcdkz3M2h2H6eU5tlO/HX
eLC0A8wusOou23i3eI4asEUL5VHARYMvIiEjvjx5k1lR4dFl+BrGLuJw5SzYe7vsmJrYmbwl/na6
epIo9QB/QNOsj7Zf2KiOtHGKAc4vRFDsO8VrGnis2GNPIns/e5VvUlS0U2dszkcGTg16NdshujyZ
m9ZXJ729MsBQBpa61CeTp5k7TOf+RvceAgRPUo8oAXDOtGzWUWkcr7m4biYRMO0jxxTWHEcCSK1G
RTyWejI1e7o5UJhQECO5qB4hmJE58rpDIMsijDM9q2KPbz/C8FTYB23dfPkq6wPAjHzEjWvDe6br
YCGA7p8oAWkEeYneLVCcBtcgUUNz316pkeH8Vvg6i1hLHsFw0MPv0/szhaMVeRBfrT4l0l3dHeps
4m6fPISsfrQECkrWP5NylXHJ0Ml1dn47rZyw1au2EFSbkzSawlsgNqFMdgIZYZu/3p9jN8bJZ30F
TkpSq2D5J1typ02il/Payrp1pCW2O7CZu/EB3veW6w58LH/BJeSiaL7EUsJuAAVLfGgtKDiCCUsr
gDmBZfrsLRlnaNRhHA6na6mgCH56pasj6YVc5Rh6YBODlGeR9KfEJW2vpX1jNi17F7I/23QInIq7
jXEQv4t5CPTYHbgFZlg0NeXsVw9lI6DkCaw9zmX//9/CMRum2JpGonz1m19dL313sPOOHdDziteI
T8WMohCwehc9EfBhOMMlQZeKemBPDN9bUqsjBOcIS5wE+kmEr+Z6dvCjuPSOt/tloXlJj+qVvj3r
GFIk0AZwbhKSYAYps+kI1Ucn2fHKkz4bcJzNvbM2+aZ9Ziph9iZb2tHhlx69lc/cnrMdQAMoUS93
VTCTppcl3jij/jj0HPWC8MbPJl+inUgiB5VNU80C2ZAdls5rEGzxI5GpClfQ2U+dC+h2I2eBpCiY
54Ll+o72tJ9VTBvzsEraaZt2A+pWszKevOk84M0a16R/zDXdwx5equ9tzvv1FhWh2UwYEoxCyCoX
Zs/kmh56Gyh5jkym8I2mjJ3hEwNtae8k9H2YO4KAb4GPJ1NOdVevIaic2vf6R5XhrKgjxwuCtkfo
0gR8KYAWP2fc8Zktj7Ectx7p1FM5/g/yD05ncUu6AXOUGURDp1QOgbfoB+qSrRbaxCP1GxfzC9W2
mk/4N6vlKkCVIFiRoKDjSm2QyNRSEF8i8vx/skESOojV1eC8CbX3gyZWu5Hj2kulhBOA/VWkj3+u
sSW+PUbqbI8UjDJmWRcD/iAMIMrg0IWxo1H15tdxNIY19NpWHcqh8CFS92ji6XMA0RWWbL5wOjqc
+SYKvzHUrtNAAmO30KNPvsUlwHr0JI+TpBDCUsP1wCHYP5ij/1cQ7Is2UDZhmdWOW2OPxkuEde2V
1FqvC/Zl6l1+5qujNE1NQrGy0SkkNankb9LJ7R9PPuKZVBaYHMPiXXbT5DULIzWOw/kzOu9oYj9k
lB3Y/PCwNnofZQJccgcjK6hhIGu039ody8MgF2AAWl47J5qkPyFNBhlhemO/08TC58nFPzM/LmT2
/Ty4MfGr1gG8Xu8j4/iGMqhChoGPzuTwR4F4FTXLsUgfz8pte/r/tZxokejYuEqnjOsL3g2ZTsri
mVRtacslJbPawVbIzU2GpNhnk1te/rnLUN56M1jEG8PWfz+gwlUbklasvWJGarEuV3Sdrq2Glnhc
jFWHRFE9HuaVxsBFocR3rFxNY6QHDvfbrxrcLeItjnXruhoiRStHcy6pUSnUVyxtwOPdMFjmXz9k
EKaaHcs+zNGohsu1MRB21ijbtR427/q7PlmlX03dD4EcLbciibwqVYnlKPppTtIqq76YMEFuwhrA
1fq9Tys7c4w1e5cqN8DbX84NgrWVnQGIY+ATt2l9o4bnupvuJR/UeIl1B10mtdyiVjR4jja3GiGH
ctL3pV56BdvPDv4LnMh+OssrU4IJDEWwmmq/I+QugXmpWWZRYMeaUMziwZb9FMswxmsY2KR9IysZ
UCqnp/VVJioCQ3ar443r7NdomC/jT+I7qZh3h6AnqiaCd6+FO+5AkIizgoZRcqEsvbR+JZzaBolI
h0C8XdRgKzCfIJNrMK5KB3TdgVeTjxr/7zSpZAokVSRzlNqSG70ltoSmZfyaePtgPwZVXkM2T91H
omyzS1bR6Sg8p7ilZiXVjjq8Cp2wUJQhUtHOsvJqItmYX5V7bbmWY0X+GrSwVUZPK3DqhvBed5rZ
wiy3pdkCiCCHzGLibyCt2f9xjbVxJcphyqIVwjpL9/eBUe18ssppxe4O4oSNMU9upn4UCUiEsKgw
469rllrWPtamLa3gfiI1KjmNk0EVgoNIq5P5wQ+9+RH0wR51loJcy6bxUCG6Y9nc5adr+vzSn+Lu
q+Y53A8fobsxp8y0XoBBPulN6nW8V4b7YdwwiL5VLA4TBjMpTf0ItcUwUEap9wArmdQF0kUhJG/Z
BLjJJHwaGO0tOuR6tNhIeCqqpSuM96cRtRgkuMUgf1tmbkzGdN5y0+aK0yZ1MkOumPMK379viQEQ
f2nTJyrnV2VOZNNEitrm1A7NCty6jbXWe+GBpzv2Kdp4Is1gbpXhyGKis74FVGsRw88cDY53cJcq
YzZU8B75UtcJuwv6Taq2kovMPQ+p+W3wCkc8skKlpJkey5JMpfuP6cRfh0a51q9bWsmrbsJPrFXf
XMhzFDpNqojZE/zCdmjezncs/sT5xS0fSiAzWdKBBWCZJs2zSeN0yfmxoVP5jZ8AaS2ISUs32cY1
XcIoQDdWTb5RwnCk9BLbfn9uWMsdhWUycUfws9rYdPINaPgoZZLwXnSblcH+cIAKi5xUtV8Kxusy
Ny84jtKL1ZrDGvwodOwSR4Huw9M6Pf198rK7Tr/90SCDXS1p3Vn+OeeY+RlhAs3Df3FdHR5I3xQ0
uU4Hc06v+5sZG2zVaTfBDgFe84/1tkN09lOHnlV0XGZGrUnDUTEN+etqysTUo2T7DU3ZCbB3W16Y
xBVsjarNxUmKgWsZMuQnVni46tDGwxmlIOz7XbGEYlcUzVPN49YdcdLLLwQag7EDuDTfhYt/uD65
Wt4Oo2QmxUxaoxYIU4HI5/DTrzufNxNbk/LShFfRLBa84Pm46q14lnCid6EOjxKqa0hoM6deKio1
KZUdn8/Kbav/e0gXd0DRcVhJqJQcB8aB4wD7fmN343ZPOq18DXPBSf3Tcbl5D2iffjfwjrO92hjl
2X6r1RK9u5xF0g6YGLAT5U48w8u/1YNn9RUTQE9OJw/e+6TGPyBNNNZjCyWob3v/SGBi/0KkfBXX
EgB9CvE7Cs5AAH8t5Eg4gWAsuX4Uwds91VMWW2L9aY2mYYonTGYalR4jI6NZ/8dkuwmL5gFH5NCV
b3Mgq3C2mCbpYbh309rNpB7NSrbZZxchIOTpXnV7j6hW4W+3rO062wbancz2kptz1eTfp71i+odl
8wejzw16VmW6BvKTGeHGsk8H5zk5yhT1YrpkBhWl0yCxHRFXx6QnXiKzrDcWe+VkKc0m/LA4T5uz
2TK/fygXwkRWzkt9crALV0am1n/Q8lIwcx/0SsglJ+h5oQ43xH0a0Q8puDOkRK1lRN5VRcJEeiWr
W2MlO21CkvtrkDGqStedVfKYZzYG1nqYPbyd0Bzh8I2iHM0BrMKBEDHoQmuz0u3bySJpG5Z+2IAB
QgEtCB+rkuc6Zen9VOfe6oXG0kZ8mIqMsTWmpfb7awPgFsjszr7tZ83Zp4iaMmDZlRriDRNx/a5L
9uRpkFO/3hJiAXYygtcURFeh/DDmlK5CCJnfRM953QDW/U+VRILLXCSEhd7OElb4nXhorlvyE8R+
ttUndSexomDTWRPY2kn4mkWMQu0xgizEGXBV61VO06wr02S6V7Yp2+KTMw2VM3EZHBoIfQEhbqYR
sPUDZ8cQPmEBsapYZo/IWdSSP2KutKt0UI5MckoCnMO8fpxvfXpZmhqsp94HoyczJbkllJy6LKEq
izqsR8z4m9Y2kP3XdNquHBW4JxWKMTDXmGgZsgweM+VA9lz2sg9858uB9hjRKhjE0dXq8pisFYGQ
gXav1gpQY+1u2l9OP0urmWoh0sYJNxNCqjFKNexsxO9+WYEB0st/6VqpyBSrp8s97fehYo5mNb5T
I+nZ9pikoGI2fFoqaeRDzz8LZ0YGCKm+zgOBVQoeUPI7/t2knz64CYBBk4S9m1BXNPnU3W7Fc1OC
rRbcyWXnifS3KwvpmPkt8I74JyOMSYkTiarolJN8w3JxZYTArBMqkwMD78qtdTxw2wahOxyLxBJ7
0WceBv/AFAh8jfxG5f1EEzkdD5H72ZniDLANOfIcptTKseLCXpFEwenqo2TFJsxW48FtodEboNH7
s5yDSTpHY2q+DWBfJvQP4CFDjEpl3iAcT9ZuGCPoYLlRa/70NnX3VH3uojqt9yLFa5r0RrnQAiSM
GqWlztNce+MPRx4VQp9pI6es+hBntqNEWiQQctrjctYOb4otSiMfJYA6KFQx5+84DvAmSzmCp0xK
hFmd+9LfLmzHrQ6/n6FF3I4JlgbmwPuG1qHuwctohjQFKwNB4i/waNqCbwIILiFyVDXYcXaBt4Mx
5f0GOEpZ3OZ8YWU1SpxEFLDkGvw9f2+e0yg10rFJZjqNbI2bNsWUrZLoUXkMGv9S31esVzh1/eF3
GjB6GR/YPCTLd9Mqmb8jboZXyZBBlUe4Rguop6SeztQ2oV1gwgg2F++/jUUhC9tTtruAIXQ1zqU4
vcfpnU9vWW+MZfwJe/pa2R4y6USgc/KviZKUBnnURVHDDaxur3bujFBhloJV6w80wVa4bCeAhyu5
a4ZHX8KZbVlMYZMSUHk4jmNGri/DUwwkeA0q5bZT511nxbb1WnzuaPUqp+AtRAAsOkeOepoiZLe9
as4cFH1lxUoAyLOTl/sgy235lCTtp26kkZkAMTvujFWwj/QXntJd7U96w01rxaEaO7CAYR6EODhY
xj9rF+I4AfDQ1d0JS9IJm9OVMlj1RxluNjvTVRkUUK1tENIj89ZgEYyPo8kzIjUr4Mj/wjdr32pM
Br1l3VCh/1di3MxV20zD8vllWkSZRAKN/7ba7KSB7rWJZQ653xIMh4TXMzbOOHaqd031rqVt56BO
M1QsC1j4tWS0OVjdGlZy5EU7OZ1704PFzAVc8RIke37V4sD4hL3xhD3RaniRzHAFT9D8SLJqDdrx
PAN/94K8ljQvpippVZhDJAkIkUmGUtB8bpxsg/EBrKiACvK1rOogmHKFuuvgIiSNSi6RRYx7POfw
VNxEA6/vcHAq7Sk8eO+qhP3rUJFPWTit1JwSp4i1QgtieHaoJDXaznwNDczETT+aTZtfMM/6tlBd
8yQtptanCpnsHbdrO6dFELTwp6JuzZCsYQVKx2TsVrq+R3k0QljCegJnJvHHbOhq1gKeTEyLnUxH
RLLET4G1UnnaYyvxI9U9jg4dGEmJouSAgvJUL9FBU/Vzenre9oDsZGwmfN2rdUPV2Ml35og2N1ld
fPhuObYeeEZtNy0arwLC1u6PzuMHxC1aJioDUNOXtz82OWIWP0lNPv4QkD+gxeyLSSmFKK1TG5YH
6NhUWIbpeVULOAGKerWscMrT7tHIHoeO7YqcLgE55pbin12nMvCrth6nqvx63t3KqYFP9fjNHsoY
BogYkEpSE4qyv3PswVTLtafQJqVeblOWYu0eAbaEgooUe99/8X6yTP2OEXNxal/LU/SPhBYHnGRW
G35frEcz4gTB6nbDaaYYHYRvR/IZNWDOXeTAKRlMM8JpUpSzAXAJvqmCIwBvX7kV652bt6hkJzny
dgQ+o1aeyVxsRPyVs+0g75JrD+ZTDVONJW3SZEmNEGGvNHtBObbmKkqOdiqh62XDXlXn6CO7OfX6
DbkvzkPPoYKFu1YDCeJD8AGTn1yq+Q6H1rLvHzQuLrXFiqMzunPWuPq/5iMYmh43bUpBPH2bMbN9
GMnhhhFA/aFSDNGKm9J1waArPfkN7rOf0vfphzaGKc/R6updP9Kp+NP8Am5j+16kbQgCSUZa0OmT
QpRbqTwBwOSP+6AvR8Pr7/79XiXRWxbZKWExoxwe9IGcuzR7M27IB4+ApNYU0yfsp5FLjMZ06OEX
xBV4XBygEg2O4aBcO42OpSfkNCz/uy0+ntsevf9Sh6pTOp+1OAnwIjgS8+qmwsZkWtutSdnO7YwK
yRrz5XHlP8tWdl83hCsmewFgmnZ/pKP+VBqUc864o6tnGMw+zR/SMFysCYJeZGQLo+1+NqrBZuie
VP2gJJ3fEqLlvGy0bHTFdN1o4bsByvmeXLrPrMIQC+kW1ynzbxIqfdiuLKsst4BS0aOsaGZYCobv
pMslxXU4zErTAJeQKN9ffVJFjeHAA4YJg02l3XWNzyhixIT8d0Bhyofm1xoTyK1eLZxlI2PLCv/L
lzsa64jk39cRT6gjlemaeSwpaPUOcbEx2MpwxkDY8AvjIqg9Y2GZJ4APwKPJUfI9T8ADIex/anYE
bRHRKxzc83fomPQhVwZ+oDt/aNcMW8fOTOplo/r1RVabag9k7T8tupRQPpWkeYDuMklbXALHIeOM
PHktEq3beeiCH4qVK0X7iY+UJTwJ4AdC4DsWalp3F6e/lJ++2X2ignbBnCLrE0xhr9fdyD1CVByY
oCbpsL6lNuMke3vUBV9yD/Ic09LneiznYKhvCWoxiUPX4uMEqANYDzSCAVfnp6jmIiN0luqZHFuV
/PA7NFPPblzOMaH0rlx/LyrWzo6hE+iQJ4MsrV89p1PGAlgkq7x6nyxNuab1NAkETKhCY43dXA3d
EhU5zcLnZwblH88LZyfZRpfkKPy1g0ReMldKI5luJdyDWmpjqUTi+f5VGg3+zKY95pSx7aucW+Pp
a0zBjwUB3w6soPG9yTgJvkmIl54jdtB8qkz2p9h8siyhnYtC3jtUZL13XwTy6FqYR97vMZ8ivZ5s
mttwvhV9wcxbHx6FLe1EuQcZrDA+i0ZkFnT+lQbJ7cfgCZc1W9Uc5ydSxaXCZsSivQ9CBwKGRKsW
rsqyx2MNURSz5bPT7uLIxlNBooeIOjBk3TzbxCqlfUXB0G1soFdPeCweKvgf+hi3zqzQZkRwbrjC
OnqJkfsMEtp1LTJarXYYawRHfzg2aHtGDoCHVHYuzbUzokYI2a9vJ9vxKElv+AgLK7UgUk3hHqgI
UAkbEe5clsEmC7FOt/mThPg+X2THb2GLxqoaDokk/nNj4pZDNC+Y9xCZXSQ1lCKqfybSii2N5x9I
Eg5g5tKM5K9HSxXjoVD9vSd82zPRUNE+gySob4IX2qMx0jNa40tPIw64rG/oX6UaSB4eMHmfM4Kd
xKBkbx5Y+w4F/hUzU/BWbwQve1YsC1HJQSwNK9aBvj91MfOeXSbFr3P/l5Ecm4M6Iqmr0Y9/Bbc2
pV+rnG/6HAV7PRmYk/Qn1c+K/h5pxvuBSI1rPNfNUPBdbjPmbOgRmiZpNb2Ph5ZrGw0GoBDC5/HM
yR/OH0AjuDxSEjvAF0cGxmGH8UPiyadqMTJ9+puD6jFKfgzqOg/MRvIBTx1aXoshn3LzI3JjIdwd
Mr67gnB5tBD9uzhFWod5KT7tkqfRAbR4wyBSsq95aYG6C6xhOoYmnANgbRSIdsz+vffGptI5JUYf
Ej4m4wteH8YnqGbz+qksVSA3J6L3ADNFlaD3XpU9aNOOE03imVjv5ceByB4t7vtmp/a1ikkvo7Me
HDtnJeGd4uC/tiORGmQy5vKNQ4XP5Rd8BPmLLaZCvkUP38H/06nHcqzsFj4zcWWWRTQ+R8mRklWY
aYY+Yur3ENatXe3YP3GbLUWCUpgM33PRkGlHBCDumxziqn+DyUXxW5NEzNplBWt4jFzcdIJQv3JT
6ME1GnZzM/0CJVexpaUfw4pUBBhVLc83EULLZp3sJ9B7qDxxzAWwVS/k0TRposy7m6cwmQFZqg32
hu64gnV9R84/kLngkChjJi8kk4x25opS3ptwHUyLdovndqhDGJCYcql2neyAaJaH4LPImBNMr9Gf
t8+M1hxtjvNCciq9RUkrrzqorzPTXbLPslb0UgPKNJIpdvRaxRoDJ0OUNmI0DavJGl0gvErk6Ldz
oGM+IFxealZde1MeefN23vNMTk57mCNbRMfJejCngaSmGPEmlJNMAzur/FLT6HY+jDeNvzBf57rX
m9BSzbB1k5lCcWvZBNpilTadC4rHFS/WTd40+uq2hVQ6uH84f9/mp+uZ9PfqcjFh7u0TEYDnagIF
YFDgSOzHHKQbs77DdkSFq7UIJggM7RkIG7Op/DpRxp1zN9uRbIpPYGm7uisrW7lTZQnrojuDrGmf
HYuFtmgnJ7YwiguEviYzMjs7wb8ztJy1+QX8cKwRsk3Wcy8ppR6/HKha4icPA6xOgMDe67m3aL4b
C3MJpsfX+hs5GCMH9s2KKf2C3kZuyzgSPknrqrVw+RijMf8HvnAfaYJgjSisaCmpe5aX8RyQ8TF5
InPgK3WeK/0LGyhPbUMDNMtlyX5b9qgaYTdCjDjXRbG0zX4mrkj2wkAKzmzKVA+myqonr6+T2CzG
CZCd3QtwCvk3ALKVSsSzuJV/Xz+NZPVYAidIjEDdXHPA2+S96tEH7XuibWmxhd0Oh7gVfvBl1kIe
P6J2fQErI6eAENFK2hIbkU216VNrTxCxrCYsZNsQtrldyxwiarpiUpns7D/OIwH0bUjb6MovaJ3i
AGycyB74UwnSfiGFZsfYk4nYQVJsrzWvRhFkXc+OyhYcxWhszLZsynrxjp+KoRAxHWHOH4jnRVUh
cvfY3XlOSX/72bmwPLebVZu1O0nf32nRNYlDDCGkQB7YCxAwHIzhJCetwcv27itAz28NGmm99403
pTIodxRucFxMiCILwb/K6kIoa2120dY9b0/YLx1mmnZDfN4AkxfGhTpaSQTQ1P2yfx0vsaultdQd
pgfVCKRigG3zVBznewgj7NVzYMBRrAK97MUWqcuDp9QJirQb9AyKKATfMzQTXEnJ/EgEEgYfqkLA
XRSxju1HXlb5+YpfbU+mNCvcQSmLW5hlhcoEl/qhGeRNPyrGf1YWieWQR5GfPxWxP2WSjsU+KOsf
vBgpbBkL3sVnOFv9O76p/3bCBO6MLR9QODg7gnjkYGONHzs3/1V0CdXnqQQQJdNYf8hQJjAMQb+K
pVXvPxeu5g8Ty877uhe+qRk13ByMX1ZREXFCY1db1IL4X78PPNfgBXrxqgyq/Q2hKA8SnjZ8hSh6
gs1U8mPJ9HRZFp+0VIGFwQqswNEl3PHZN3pN6ZOVyvWh941ycd9H4z1cuExVNQ2B5+5Hx6dj5GOt
ee5aq4zI6PVMt6w8hI74QI1VxnAKMEUiBCr9DQrPHBdOLdf9IuZkOmGZtc7I190Nvxi6pwuYaUMJ
+XmXavorIRxfz4o91UnW8Z/lDd2zo2hGoXDgZx5UmiIhBpRMPQFGWZZnDbCllzd0iobDXUfXB4AP
Ev68j+Am70zkITUlsvlT189aPzK8L59gkEcKYbsNaqdT7vqD4Jcg6X+hq0L8RB7IE/co37et/aMj
CmEdiZuEco8M0vfBRN5b/A0CfnyjeRgsEcoOaVIDHwKyAbVrEgPRZTKPCgOFQHJJAhou0IuZ9XNV
dCohvxEns2ocQq8cDEoU/lnecu1Fb6m1Sl5/ESnx/le93+eaU21kPNrn3tvmwHnDP0A6KKN7nirJ
CuebkmztV4qK5dMEp7Dz8qxNz4ycY4C8DJBiRrUNYDfT8GECf8DoTqKHj4lyeL0NlZStQJjeR1WH
SZlevu4VHXy/xT4Wj+lUP1Dc+bkg7ueMRllPI8ozsdfIm6vL2u3nPZ03XnPjq5yuR8ca5ybBAeRV
CSpWiyxg+o6R1DJsF7jj5U2dXTfsaDAhiBwnPwayz9zBm94pnwCzcUfvZh4SYK+Pa7McByUhljdS
M5LYcck6sXdprc9ml3W649yJkh26OJBKs11pNP3hFnQQiG69ZnXAY0yLZZCZPLW0JxCQ4WKApc7V
faxHb1NdfDYBnlyn0PkQvg7OClR/eCRPiJYjxOB4NttuT7pmcZhVDnx+SRU8+g3vZTJJjgsjNEaP
zYK5XF+Mf2CoEDUpe8ZwNKPhPxrhemvZRYO494lwItIrCseVx0XoInMcoA4HsX79v870LOUKo7UI
3BE2M+o0wC+KLu92tz93VHJ1Hp5rwbV/PqoAWFm3PDKq6kLBlBKPR+O1RTmRv9SIYctlLDDdvTzC
y4bjNpGEhEGlOyTyBWpYo/8VoWNdoNgpYCx2JciuNERMnUj8kZqsNNtk7zxmaMNOy7ZbutiMyvNL
l5O1uCsunBqoXLKqZHoShUD9I6j6ne31wLHp0fWWSqb1M+9YnEPPYkSbclxjV2xTliSnLFGQ6ZEX
U9FaTyHj0capapQiPBoYJjXhP29zD/DRuvAK9rBwG8A+w2JBz1aG88ej7r1P9DA9T1OA+iPVQnNO
AFtQrjdgKkRWyKIvBXNqYJaoke/WSTNSmWkX/D7LTPHNIQRpZcOd345bKCQHu37mMF5qUbSxXg/i
k2VDtGDq1dI/2z4b9ykosWz+OrSeWwDRKrIL5/orhyfU0Spc605uOM9WgoZe+wvs14e262fv6x+y
u5q3t8ww92TxWNSAXC+3pTC7RoeWYkX51IzjwJg9CrKIIuKazZJ+3/7LbHgiMp4rDBmmmDhJVOPU
+5d1OTmsxldB44qcwiASWrlRRmdjoFyvMqs/3VatExdjjBXpseDZsYw5Se97B+mwBUaSS1dsHM0Z
ObzJUkN5t2wEImomJX7JEndqk8H4LBG2czT6WOnYiV1FSwZkf+HfboSElMERkXp6cPi1PmXYx6ph
FyFXoCevBCxofvW/BgdSb64500ku/ynRETln4m4O7ypH9ncp/nLURHZrUY+qgTMI9CGqI2QtKpwj
npvV0H96CSLPP1vcn7ig/Dr7AvbsVL38rwePUcj7GsH9JP8URaHuYb1LfTYj1VcMMuVrTid+DECV
ugP6sdwVt6L5J0epWF06n1dvF3aJH3JON9HS9aw33xyHuRrlZE5CTK+Byx8BEie6AyNDlsJLDQnO
XxuS1tBI+I0v8DY7M10F0VWWGgzAWWHLrzpwt/2aeeCmpYIPWcy3wg2zfL61wjp4NSqueOAcyJrE
f3ZY/UuNvbCNysm76y/PVLQ9DcNKhrACuBOyZV/Njqg6FBhvjPhxjLVS3Sx8eXFOz1GyxOg0OBsw
Je4BkF0zIdIPYnr+/XBFGLNeFfgwhEa8JCK7XxgqNNCgF4t7nvXSqB8+pw54zZooRfPj0cfC5/pC
lXYVsKBG1RaOGFCu3RTGXezTbhDIGtSCBuVPncJXrcwgWNNbr9ddFfaBDI4iAK58EA/rDPW2/YZN
UMekS6xYz8H8/pHhQxhpF/5epcIGPbcSD91O9v+bMKPfykPJWxgNReN0KAEo5WQ5Ler5v7atBggv
iGV6AH1RUKcYPSeUZX/9iExqlci5JVAcEBdee4PX14cs8frWz9hiwOCOA4ugSTLbdIPvqlK5ULfy
UdERdANIal9XuqoanWFv5uEcJVDa8C5ASWt0d9MlDarRCg4vUcEtK7TfgEYBnbpG9c5n2SDrS1Wd
92nq5UctPJmPCEL0hsjOmd84QHIcPc0tlr+lTG16lNA7ZlEQWLr1UbhdGoMD81z6oLU4rotcuz1u
kKQdsgcUqqL13DwUJUvLyhNhtGpXULzBk8BHt24RGrnnkICay+SPSPfG7C22cssM/jNwRg8BA0+Y
ppiAaQW+BKCHT/XfwNY9TmM6pCkvOcsZXBKblBIAoZbn2KV7zhzxu57u8vXgATyUBrYKClN5tW7U
JpDdoXHxGdEsl/ccydTi+3Pcl3OY3JJLW6D1y4fVkZ/GqPZeTLBHotVMSSWfFhSAF+CuzwAXA4Re
eKqQusr/OOkdy0NtQre5tmJiUMDj2TO7KuHyfhojFJHWYDaHDOWMKeM0V9ZJr/XAuRwK21uxoQaY
mG4V8Ew8Lwl9n1z86nMYbR0eNeOiE0KB4DU7zpDmqIqIEEtnC+j9en++DJO2NVf/cWcto3rUC1ef
07nCPmzLFgQAalMsDCYoyrbHuMT9wRmJ3PWUALYeMWyib7p+jhA6OGPmJDt7uWTbD7mGaNPOb+kL
RamJNlAnziJPDuCtiuQJ0X/C+Fvaf2gtaLoQoU1plwl4cYKipG1KypyDtdprmAHGaOpHH9ECCqsc
9DbPsLZaePHVDxsF5VpiWEk/hLJBXzxByf4f8fugQagOGeQEqnbNcV4rxeIpa9ejo2mkg2Ggm8cS
d6mAHVOeD96HLZEkJQveXeboL+EvB7sMKANcv9J6mDcOXAo8l4zRH9cLypAy51rO9RcKvISFsg/I
UJFeT1Uit0xAPoPNicISrwWSmymV7JwdznUQSfKYk4nE339qZKjkPdWv4YoiTh02TTI0HUpwelwy
J+nfbY67MeB0wygPWSxkfh3d9btlzG/2QgW9nCIqOfY6/XQioHfMejPRuReHWNUxnwDDgbEHhyYY
3P0gc25oyEho43hae5gA84KQowDcLw+3cdKFZuCa2SERVLC0pf5wVV2CHgaXQ0/X3/hqqBviZJ4p
in7ZWHfSCKBqJKeQfEzWmkF99REOCthmx/mtyf42OmyV+3vklzpXJlhQifBI13IGPruokt/oJCBf
5mA5NULcmGkgb2S+tn9/Gg8r3s3FEHT0pH0lVT25nIn1rBcEB4CgaQ15eqMIl6/cvvE5brYIUN21
Fe4ZQDvhnTwg1Tt0+NLKsOCdQEjyfsTOyKzDKzgs5ZML39rEwVmbEy8UGsd/T7/v0lzzMiPd4TkF
/ZuxsR2r0wqyD0afIaY3R3VhcAIX7U/ftGOn4kfAg113ybDzozhkOzDa3u+WC5J2FN9x93QGEeah
kLj64pknlTBscFnGvocXGmvxiC66GoI4GyYPHOpbeaJiSS31GgzFvuCxPjyNaRRWPR601ScyiLy5
EsURFKhnKkkCgnpBQKak8XChaZ7REQZo3vSlyHNro1NW7DxBDfk93RdEfcOWbc6EIYFcCt0sfM9K
MOSWRJgUTy+H7iwLcib1zmecoeJNcqaKdZsjB7MXc67B3jY9u9Gq6suE3zLaoaX9nFITuZxv64bm
3+1hyP+4rnv7D1t3vbZRDuTVRzR0bLze1+ZZDA+vGk0TrggSVdD+E2qXiCcbFpjQmIu6PwZ1HI2V
deY3yOF3O8+T8JlSbhjktDaD2S07xv50rR17Sxcp6rAR2ZHK03F62QIyimRU33NJT2mcBagnD11o
EZIVBJeTlV8SCVZ7qiGARkRVDtPI3S4OvZtSRK27Ovt448SpHYKfIHxk8xtnsCmobLbQBmYzGQp1
1odXQLwVMPmaMYlQdrLA9bxp8pYae301HnmcbeDwCpa0CKvnw51Y2ldc3X080l790HhcfNLILCl3
xd///zT9KRDbMKrICAZu9p1rBqhabMYIAju+EVaXV9vRM3Jk4EMfguiQi+WJTXHxI/AoIlvl7R8T
FfL2jJ1OoZZnM+OdeoI6uvVKda78OIP5AX2TAP9dQdAiYD5NvF615opofzI0lbUkgWed5s/wPCIu
KWDto5OgCMy179vPGynHLcqc8g+d31pZb0QHT49J2NG0Xr4H0rR9TGlDhPyiUQsQ16qJ1vKdXjj+
ySH3bQQtPPRwumIv263WUxAoXgwsVk0N0hZAtq44wdwM8HpuwVDMWt3VfUCrSBY+2pGpFirECsF9
jAFMvvnY27Sjem08US0m1ymb3x3laXimjUAVKmX59u+Rw+C+mKZrJBTN01MUGcUE30+0tcc+39mk
gAdTAYWGBBwsurmsNuvmhcywxcRKKdkC7vlReZv7okGuJJhopYKfvWFm2JSLuvoLpGtmziGk7Ym2
pBwXHKxFhFuIGdG5Ums2axABnuAq8/CdSmWhUE69XV9lW030FYakTxojc7p3C6N1CDm+jj5GzMV3
55DsZT2t+qhv3iJOiiCvVmokrCGCrg7aGGkHoqyHh+B6b1LlVRm8zCZavqMYN3dVZ2ld/7dRamIl
wj1wa4KIQTx/lJJXzR+Gc2GM4PU4JJIk6+mFgRpfFw9G/AlXQgegAl79uaVW6ff6HNF7d+P3MIeN
g40rHBjzX5+2jhwYVnittwP8TuuTGPhnVIqNI5Y/fOBihxKdT7ZWE33ls3Qi7LBqEhsQbtbqww1U
cjQ+ocNvhlOjSFd9lYG1Kg7aUzhAgWCgF1Vc21Qj4VO9fO93wqtr0s+n3/pPXqmnLKFIPgo4pBS5
iTllhGjJQ+ZXGtDcb+VFiURmNqmkL2EHXWrmOZ5Z+T0p96WxuFvKOLYk99qHw8XYbKslWmlXDui0
E7qHg2c3XqY0eO2hxFxTbWVQuPNbHFNgB+sT36YRDd0c4dPH0XNgchU/WUEne58mTtJQWiSSlaYH
tJP6KjkOSb/BLnUViV+L3opAbZW2B9hK4UpaxFkHbVzVhjpX6J2gs0LB0vg59qQpouCZsF2Rakka
tOMdjLNXQQuqqmjdsh2oDxi6WPT3w/oicgE1oNMRpleyat0IQ2a5LCL4FWHRryIJ2PfAr4XVugep
HmnWPpHCgzmvVv7cV/LbObRQkRiwBp496fgwcuhEJFgwpwRF4OH95rQujwyXVFjglDA5wFw+EtAK
cNQtYl1WpiNMavnLtMd6WBT+nLLwxptQnMz+K4N70nwffrHglQg5aoVwCFsr3EUQjiKngc4Z826Y
VLZN0hamavfczptNTAXg6S8lSnDWBQx/QBnujmYV5B2m9M2AmXErtakFWUzDRn439Je6rqBnX3yy
TFyqirrqEO6CRHhBTnIxk5OyOX1A6wP/cPDP/+SBl0k9COBKhu2JmxSnnDEKHyPINoke/8gknuBF
RAUuiPOK50VlF2QXumhK6/0LXH/i/E8UpF2RxACHq5F7kVsEs8cvUC1l+V3NPSrq3wzfXbVQ9PJS
Qy6ntriYV9Bok9gWNkPVLMGES7njLGWN7MKuIkaZj1HnFtXfO/jqpTRwQTgON/ZZvU+zPQnq2V8e
v0E0+kwDl1obbB2AX1NZ+l4J/1hxPY6uWfUSvgfPlpLHiMRTWb0Lnm5Llx19KG7/l8L5MydXyH1F
vNOlXh3LBkHSbVGS9ozqD3VLLMK49M+W8KCGC+PIJIFVLQL6lSFSyI94o/TOu3NpoLUTphGcuCK1
0wmuBQvaGiR5r91BKvbYIHYmc1Tlb2XoplADGaKqaJzA3OwlFPzAXbLpcg23fDOkebd1sJnvQJMC
/rD//GayBODMhbJUJJnHDO07G017TM6eLGE+d6a/pl2M0ODDVOPVDx8xUa04tE9ftngKvgMRj+3G
pTxKTI5rdl4t6g7jCPe0hIl7EfGbR26uqRHe4voVTJWLDlHN67GbS0Gaqa6IbSJNFW+EYcvqfclX
sgHU3olt1+ZE7+6u/DmGq4LCD88Ry7VY+nJflFcmoQVtkrKdOku9V0zhkIKrVSQwoMuHpMBfk+2/
VuZFwcfp/UEciGJMlGppwN15s22QLvf/zS3Uys7y/QDgssQ4WtlVw8zEHTE0OXrnlY7qNBeghN+J
nWXvQrolqRPkiYb4vCqOLBzv/ujXXcn7rBEEGBZGJF8irLVSleR0DqwBd6NvmdSwEABAuoaBiDVJ
pv1cCl7OR1rUcvcgUbvugKc2VFFIA/U0cq5ri29RIFy7lKDyaIGi+8zBtedEyo0n5n1D3zsjeDEI
1meH/D2XxOU9rdhiyFeBfA3fHxbfvmBD2pu3205rUkjuXa+o9noQy/DDZESjUrvT1tC9KnD+iZAl
464WlkZhNhcGAENfrnDIAgXVq6S3v1KwXJzx+ijLnG/chuHm6YuIlEtJIiLgUJWLouujaXZUD6WZ
DvzcDnit+3MHf30qSdhKyEiZj2dK9ONtS3J30AE66hcmYCgBuhtDgHBS4UYlZn/ClpWUKB4a/tIJ
O5F6mYlCbRv57aLqv4+7pGTkiocC3KJ3tZ1PNGNVO0bcXbg9VyOzKuGQWkWQ36N/kzWPXenC12Ep
PSX6FLVyA9+Ioo2XtPdxzAMUaBPhXH1pLTkiAg1FWDTfxDXWxSpAswKVlUzJbHxZZ/4sRe7rAshj
gImRixGdJJ5/aaEPfn3GheL8EKSRl3CgPlLsPaL1c7QeF0JLiXo/hmQvqS9MsE/VDmZ+4/82tpBu
4fOurpvHcNBE00iGgiEmPoTkBhWbp6UtPp2dCWhI6UneU5EZDYFvsq0mao0576K7QMKcdBeGXlsn
LMnG/Jtgh2PAKSqbyD16WHelCX0BnOdffke7zuhQ1y+pdex75FJJ1/f8XjamHqmk/8n1SBpXClEq
n73z0gpIa9bzq4xv4mOaydPGkREv07Ab3cZt75Kx6bSVhKJtpBDBSfMyi/HnkVAUDp9B04tuBJoV
66qN8ziNdrqQuO9MzFsVTntmiCM73Fxtk/0J3l4l+wpIOLRLRf5bzbVEMtWVGWkUWzuC9ReosxvW
6gONZ05kqBpG53B2RHEOOdW7RKrhf5wCdSTVKhBD6HS6nNCMVLSpXFb6Thoyv/AIvqRKVy9Fp77+
EzyJh2NoSLmZ9Z6aVhfRzBEcv5y31EOt3Umb/YZVBnTYM82LcEcRgNOZBOU87JL5MYfyvZQpsBPN
7rQ3dj/h1YZI81bolXcmrmYhj/ImpssfOXK1EvQ6J9Quz2AU8BUoLyEGIOSRQZHs1u8z9OCGcfJ6
6Fue00TlJ//2zotJ1bg0oe0P4RRUSOSB7owscV069Kr0itnLGqsSOwOg0UyrAmbTuEdRNObzNd4F
/bX9Ls1hChViv4HvL5ORajSB2idMovHjEnJBogWH8e1wfG2kLgX3U/YpgMeII5VZgYfXDO/yY10w
Bwv9BbgOgVwNlNrd2Xr7akI6WZyOA8zjFzkgbhLoZK/NiTw1UcV3b63D31UgaQrdj3wA25Yjy6wY
DSDwVMpiOEEJMbLyrEv5EzM7VUnEU+bApS+//RPkYOyiZ1gZNCdVYFsN3eS9YPEc5xXBQs219+J2
RanmFtKk3/caU0fv6RkUoCH+6cUmqftfVlZdzV9v3eqMEI3GVYn7fLW89ft8Qy1WeOabzr6v3QUt
a2njy9tBWwFQpjcRolSNTkvPDTsqu0RA32NRK1SObkzCL7ZHMeawifkR81J73XFT1cHBGoJWrC1Q
s6S5MLXUxXKbFVBah4gBAsR8TcWgsNZtm9HSTHWRgUuUBtk6b7QBX9Nqd1TRU4kCaaaQTS7MbQQC
PuzStCDEEh8lgHWYNp+R5OQeVE97osOu1jgcX4Fr4Ta5Ok9D0N46gi1d3NFRJJkcCt7+c3db4zZj
T2MVDI4zsmfZDoG/yA32POSnPBXpj4IeAySUOweVzlfz3lb08E40xtBgjI2hePXOVDU4vCVB82nA
9WN3FKJ7/4pEK2ZTQj27ZAY9Mb36C6ZUYtgJ0MxeT0WaB8zKYay1D57EmCSuH90wHclTW6SOuLiS
OjsVLU5pMlaNRAAKqyOct92oWRO5fgKBkM+nTGLa2REhsjSBaj10Jso72v17lmAnwCPi7m8ovFCy
Ex+NuGJTWT4BLPZDRliIKH72RkWYEIVkz6M7ky3Y+okv0OAGTmHdvIUjtOaY3SVnf0PxPeale2IU
x0EAXh5hP5dM8ISp5ZgZtZ9w8ouaBO8FqBO1xJ3z+HkKT/hWSB1DvV79Zvj2KKkFX3b0uYI+pihk
BcTezaiZlnrW8f1U1CjFpuLa7glOHBlY/zUfywFOAOde29echeGcso3xJKmNpbuGpzjODH1c9WT1
9Oc5GZNWxEzYyLGForVHAZ38NMMNbpjTwpbMpU0ooirT1zmLJrasXPcTo3s+OpfMJ8CevnCIG0HH
MkJg282MLYgkZqRlXbfriekh09BDOYA4Iw/eUrB+VMDFYV9IUwjNB2aN9ro2qSzZOlNdFOJkpK46
Zum5mZ1WhzVQs0+4Y7w5OZ3SUXumAfi3UJqzRiWM83sYg45Xv5sbx5DDSWD42rAnwXyECc1Pf6SK
/lA56vx49YqwZBo5fzJI7zUeoSGcL/2WDODj4e1BxFZXeOC2MbsNBiklU/nYLZpgIMLVUQVcMwR6
B825pG69cDggn88jUegOS+CtJ6061LB1yZ1dID9O6d2xsu+C5sFyZVqdykuoORCuaK1UVLc474tZ
0BAMVJ/T9ggExE7mp/7mHxaqyTUzJzSEpqPt02K6cNF1/6CEygPlc62/nXj5pdrZHdpw4zYwkzei
HyV5bGl0706IQnHLhiSt04UhJtNAhu0knF1BF1/i4xKY5jN9OMetTW0kBPSHl90wG5N21Ln7jdR3
73reBzzOjq0MNpzpgpNkXDf64Dta/ZqzZG77wxK4er/TXp0a5yV3ZKcnwjMjtIbzrmK2s5hZ3UwN
wYT4SgUxUnoXwbztAf4AiUCln4VCeMAfikt9S8SIjw+yjjpLwu16+rEVNFr0FgYoBRkk1z6+2ngy
JJFOCToxau9OvjaBlyBPX1//LgwKXHcuacBX0RS7tAyplhqFt2GUJHlphIO4QcF1PEieRb68VjAi
3fNsNUlspdD+F273zwvpPuZUOlaXm6Qsa1ZNYd3yjsC7jGcZ/sDgBFsWnpdKuJmwKz7cl9jnnVKm
PUXlTws0cqZCyAm1NwLKrBA4MYLW+w+9bmPoa+fhFe+CmSc7fokAl6jMx3717R2l6Og4eWityTBA
Vj3g9KTSafNj9cf+wRequDjuFyUODML5zfTbPeWkVuhDCLOGKQMt4RzIpPJ8sErd/zATZd5eqbG1
/6TswQxRgA9OZJ4hw7P5OHqHzK09ji+m6f+wLzK0bnx0PJgQpx0V9zAcR+6EkqiSP9KQ4E0u1vom
pQEvvBcz9Z3Bh+jkRHRTE7yWjSKNFEiQh8KrPGiWYqZ+VK8VlmcrgU46EZKuQChhdwszfjsk3qlV
cQR6AyTIYfTIQFf4YJ+BeJoFbOrnrSTT2AyGRhIavBb6TaH5Y/sGVbAke0JAGwNDVVDX9WOXHAJ9
DGIvGIv9uElGiprGhD8bfd4Uu90Pu4gZwL8dTYIzvAXXfFY6PCLh7Ei9Vx8Yl0veinzcvj1z3Lw4
FzA19oyfFchGQLtOCu61OmUpujmW05bq1KJ5gstG9yrNVSolWhAqtq9ydj7+dZairGuLzHEZh1W6
wOAFyPvYvf8QFIWFcF3DFeJ5CTQAi05hJgxQXOUUOL9/g1Nn7CKvmy8ECmS0i8A+28ErScKSEGpu
Lp5FYJpt1wjg54Lhavjnqrq5n1IquOAvpcY4t0AooU5G3FQACu+xGNjOHnI50rRU2htag4foun0e
MidlDtTqUI3BL+ogmUQ3Nf4P0a2Rnl9DS/Qy4+A2NUO5w3GiuhABZNtnaS99eE+PEqr0xr/RxQRL
CKa8ZcQLGO47Py5KVd1/nE0PcGOE17q1a+uXrV61NyZWn9IQHMOoAAwGVRVIkNC0TgQ3QgEOSq+o
pfiQ8zZvOa04Xua/rbsvSUHtQVcTIRC01TSf6vfZKyeRhujtU1713rtYT+bHXOB+gYUlBO/Z7MHR
shSvhkO+xq/lkZNkMcoNlxziYY8XVEZjFUr3pS3DP6JmYWFyrq/GMJX1Bj8AVU13wR+1+tujw221
YiTvtmOTqtbJY08EwFFv0On/zu48W5rkNGgtjV4+mzmIz5v7hwequm0I1ibCN3kfRpO0LDb7YCIl
49AEzdo+HXYGTp2eP83wM+aantDJkSDc+jx7nFXka6DC8TNCwmU0rPGzV8nNik1dyr97kdDsCpL6
veQgElQxv1QweLZetg33LF3HWbrjYsAZE1lObvJiP86c4T5TQd4yCEN5AFVS2H2KHbt05+xqzkOS
Zyh1rdCEIxx3P2DGudKZaepgltJjPI/cKrLKZUQVCqAOy8by+QMiWKIURtjNgrY//UdOkWetpu9l
v4+qu0eQmbnqzz6OKvVa5IpBrEicVKwmb9ix2vS+XVSiC4dehreHuf5Kc5ceNjdVMIb0HNo/yYHC
ZMZt614ilMW9PmDtVsOnk+69BIJAfX4996LVE3wLbav2VZT8IfZOaM8VyVjrAHJ2jsKzg+zlinqH
LnGtKhJ5RXbRiAvFHqO8l0OVl5P7WD8ymzZtIsyEpI2OOOtPr8jTnB1njOSxp0YpADWB4Nihsg+w
+jaqfByS/zMsfNdJK5/KtioLqaXyPOi+flZUnzRzrYNZcBaki4KbQvZo8NYZZSmZwvz1iaHoEfqj
CJsa+dnarZQlmKRQ6LZPU9xu7YjF0p46m+zrHy25ReCzDKBd3AYiLlpoRlV/XXRpVjkS+iMdqyNt
bjkUqutYl0ev2X1Y6iVrK/qgLZRgTW1WzbMtlB9LLjRMbNG/57d6dl3sX3IvmhGrFef4vYBGqqaE
x+o9dZok2QpP0nj1nYJRG0ZuVk+NoEqkAnLoLrJDZ5Oph+56oM8ZUEVz+6At7Jvao/UwgUQSS28s
aJe2TGXczuD7xKFDyRc3rnvZ+a1JenryJkIa+mXtASIq9WVi3nc2Yd/ha50VMcVfVXy8PBNDT0eZ
MEILGkLy2/aDarxHuuhZdZFSCmDqvbf095shAzN7FSgnZBjXfF1uSupT584zLINnsYhet2SJX1o4
aD3n7XkUAgb9FqzrYSB/kQIURpN1XMJa3GIWPQHq0Bt8RBpHpkyOFFYJZl1xSXFReQopXKqucsjE
1kQ1CKwerR/M+ElIiHtGERIADHtbOAL2ri7vsBepwbkxq/4bijvvCx83IqPKmfCn19h9cW/ZY/CB
PoLYWbfRHVRDH5ufEgMZoB477/oGj2OMqzFJ9IgO9PK6CYS95GzQUVGBncb169du5U5kyXrhJdo9
0kEl+KWo0B1OXAeKQ+YNCDShQx0ZK6UWKbBU+uHJw/OqR/9lT01Mg/4RFts+xhmRSdcwfCoE/Owy
zsAuTmDaHRfr80oIjMKkvljItZ+rGgh3FRjGZmZzyxyLc0HH8lMkEPn4xZWRpLdz6cdwEW3+ZVWI
hzg6gUGkMDt5RoYA02n0htsNPt7fJqOJns3QM1ZJJdnQK25363x6JeNaysnY+zl6z2aAwkpKPqkQ
KVStEGPoIvttrsnAHoNe1yq5k7UW62eZXD0Bq9HvJA4/JXknat3AmuKnaoEyuJLZMfeWzFtYKZk/
zglcq60jOHMx9BVOdBGWYDqAeqFZuLrAXs8rDaxq0olLLWC/N+6L9tX1lBcihD/eeDqG9uQ/vpjF
vqHooLNM/pdin7QUewv8HY3XQir7MphQGHY1Jm0BPh4865SmakKweY0/gFNL6ImRGsMTc9DftxS5
e/CxvEUr0hmM1n/D4B+Lo5WjdSn/82uJ8E8Cpx/7yMNisY74qHp9G/9YCKFqKcsdC/MzHJUJI3hW
A3cU+nj3Ftsc4P7fNLEkBgi14CHtJPByVON7tlE5tIHbu6gK3Y/YM5sStm3coekAcqNCH9f4Eizt
K0LkjnM0JAzgYY7zXABe317WGtcg+PIKC7EcI5vfK0pMlfma+1HR541epLK77fZj6I+urgKkY0dJ
39ddGHR9BdkRn8fpG9cJO8gAheP29t3ZhH1KveQup2HrAf7SyyIup7R4tP6stnUGwS1pYyW1SyL2
aGnRyBr6vY4Kr1LcCfffU1E2HZhwyz0aTYSAgHjFnbjlFfHBgq+I/0rkWpLtxr3523ABLSv/5nXe
OfoqS4TkvPl6pYi8uAvYIEoj+nSony+1+C4Qvlf1liGJzzgyrrEUZIOYtjK+dM/qlidHr+35r2qp
JUDT8d9GQnsfA9nRgTln1vY3KvpCkQHdzIcs2wGIpn3v/yd2L6XfpcO2BvbdYhlPNEr6vrvuhUMF
vyvptEvhkSkgJIT1csTRjPVTFFbvf+4WaVhLv97n51PBWxfRkOq8h/FBK0zberaQ0Y7PPgnxCJik
qWx2wZpXzGe/r5G0N0AzFsV/onjkiI/NCf2KSrhhCtLwEp7eWA6VtC7Jmm7QzW5oYfOH4z6ty8DP
3Te9Hcle36PGAG3lfTkHL+W4D7+RtOtWnQ3yxT66ut/R7ud2rQTHbMwczP3EsU/MuqrRdqcGLLyr
wYEt0g+MebMfaGKoJmBgJuAZGJv/c1TjQayH90oIiyXxA6KpLWSCEmTBXY8SxEHHDmN0dFZrO/eU
DuCaF/pNHI4KJx3uEVy8l3wMuUrBX+RlhN3WuV8H0SDFiiY+FUIqrKqsSK8iBkYYUuOl6s3OJ+O6
5kwG11WszRvtBBeMIA1abPY4MGLHp05T7AgqXAPK5vDmiSKL90TAwDft66TCprYTaEJ5+1QyeAAd
8tdlWdhC/7wnBsCWP8L/Oz0PaIi4koLzdYW6AsP8QzxIcfUL7NL3uPJA3/PQJ1ZneQUZK6jnvCC+
MfzlGiysPcKMQHunatL7b0DOWgQFM7tXIDVIVVsdUL67F0+zvsusK+1a31rL+JhXC20sz6nMpgc/
aBN5oBtTXoyQw++9BYIbFR5mxWoCyzggCpdm+CQEquaSGEFkt3j3k4JRvIELZzu65ujKnsitN9LR
50AkxFLwOEKYjAID0z9A8XRq7AZazXl3VQQlya2V5WvH0T3iZcvWOLcqicK9HRg1z7g8qABqM20o
uf4CQb8Gcog2Ru1vxUnJ2dHjzYHBKf7kN6aoX69ulKZBLQPO7MhTV7LShKP0WPrtn+bNSFrS4P/4
BdpFSuwWZgH8vzMIl+h+ZTvE0w2SRF2kWfr/xIosVXPykgNwpU9yh1Y3S049ijzL2tDORbk9Pl8j
6qKVwyzYCy+NikInGRuT01wih0RGQ9J+cEwTOgArdEGn/LvoRMp7so84ekoUDp82iGdOqLuxpSbL
1S8AlwJWE7Bgi06bbODj4mIN2ArJ3a40BCb95J86KYSFeCIpGVHP/zwGlisuUPG953pDbpe6fhVO
Hv6aofTe+IpTgdH3FTwC5igQurJC0eDu44S6l3e9MKRvQTnLqb4hWXHDchXLRCrmYzgajQNPqUbe
7LIxLQGSvcHN1eHBgVFOVohoNCU9Z1S+v/J36rhPr0Jvz8z04Cl7CbDU6ndDHzak3cXe9SV16CPX
8LOzkDnW4Kr7meAqGzQB3D6tkxnAy/Oa6tIpTf9N21vU732+cMek6Y8O0LIcltRZsqQtamWhGZNj
vzdEo3tvQ0F4P2LuLIzBxQgHsgnRuiBGshh0xNAcrQeHMaTvaRimSce3UeAuqV8W0BWsneD78E++
j3AeEtnGNMshFZVYhkJBxG/ZUvVe2TQaMmlMyAeU6jWeTxxo34ygwNHJgwFZtRD+Kn3CMbpGNWt7
CrNesI7K9Vg4llZLqu49qsdlU/ddxMsykHuLjm1SC5rRyb6p5JhNO1MJAxPHRooqmTNdacg1EDGB
OnV8Jc4DISwcZSashpXm8oDm5Sczcj4xqbWlu7JaNmMuc9gCMwLoj3nY2kRXtOhexUf/0au0uokm
x3IrenRuXNmkpAeNepEV4u1wfRYZvOik92+jv7CQIa/zt3kmHgLyFtTdB+a42rqNSBijACJrj4eO
hW9cAauIBr+7DjnZEJG2bn58euQQDDOYXvKxr/rdzywgzhkmNZURy1FoQCWyNWuEvLOP4wbRP33C
DIqyaBwMcfvH3wr4/YXYPZDk5gheLUgyghfPHRo6+0DxVjpCf5naQD02ImiT210LSs43EiRVvTCu
mwd7LalBBeJQaapYvdBWmhb2k7NDfkINbq45aKiadjZ3FYski38hwUUh5sUL+46509ehc/80Cq7Y
Peu/99hSJ6FaD8gAueaAyns/W6Eef0nIjRABziCtRJXKRS3Y1YP+qC/9zvl3XOfQphss9PV7cOv5
6c4K+QgtPcpPF312cmioD6/bLaXI5pga2TKoMWmQ54f6mXyC0TA43zf9X8d0snHFn3yz/riFnJmt
pkcEXVEZTKBAbkCBao36BUySSrHxgNbfZpFF6HaWhXIIaXg7OUD5+N05XfktZK5XRPhzjJxt8ugO
fIW7qIcd80VCpZd/nNqwK0Iep3YdT2d9Czx8W76h1RmAxAMh2eJihsaAYHDM50iQlsQxYP3xXIeN
qK0PtTh2Gd3JBk5JmehZ4Uu8VdhbZuGqKrH8JzluIShPdYT1AJC46g9RMGqxg/JX+OMDt+xZHkoU
yI13URB3JnSKEXGiE3o8n2y2uktiiA8FYEqsuvFDRWns2RkCq4ZEp0frBF9sPRph1oKWq0FPCMlN
UiPa/JYhJKORQFx5pStReFyqX/9AyegTMDq26l3ZgTIXrK+KytGnqv0+Z2Yn/XwVMBRndB6R/1tG
4sW4t4l9hEIdpY2VMmhmw35TUjXp9qIX5i0ieqVwOHrbTERenFbkP0QBiO75g7o2DODPnaeVXtog
kmaGu006+fV/m3Pabq+vT652UQg99nZdR2MT52hkR7SOijcVl0rO2q05uQcxn91eCs0IcoYFtBbG
kB7NJgmNVR64+CLDeuVtd6JLm5biAPGeQTlJ42wjb9J9GyE2AF2Pfe5UAT7ISFOIfVCSkUzPeE/0
qZpJJJQSNYLEQ/b7F8Kej3/CBHyPD8nWIQhmOwiOIHwVG7bBnoa2iLc4rhYL5gtmB1wMR67NPcmo
NEq7HMz/SGn7ES8R4cN5mEMI8Adr+rtCw9/HnIjJVPO3nH5KDu8RUmnCFfFo9/v4fqjGT9quQDmL
ea+LtNdY9gA0dvJtxoxgBviy5+DfdV6VAsLggP2PW02i/wXHVLIGc3rcG7LmyO0mHnUb1c7GxzMu
skt9n8vMbykFcweHvDp91PbtMafKgbZY7u7ItA2JLzbflLAiCg+a7uxvMhiasi+ud1dYAaUHbTqb
nwijPLxfq5zm7vi+xeCwuN6sCaibPcAZDiGPXllEciPDRyA7e9doNtdRCXnnVYcEJYpcVBZEBPe3
wcMg/mpxXooy2ogzhu4Y0QCkBd3Ue4hObGYxQLcltjfu3rw8K+Wr5s68CcNMRw4+gjJzK94vhyR1
9k4MwpdwN1jcnrBNqeLSBul+nk+JnpCOQeBkiyDJuVq/67unDSWcRHhsrbKIq06zI7vB8zJ/oual
YbNCgQ2yQh8lvlIzMYMZ+lCRrLORdXEH69d5m9b4ZHQz2aLPrltwIn+DlAhU3tm2dHpHHG8OAu9M
X1edNwspq3XQv9qNverXq5PhORxAWoXailkfrf+8+cOz2FCxarcSTgD0ixdl+TQJsq5EG0Z+M/fd
zl69fh14FkkSxhJrk8Luwovtm8puEppHXjbiCd/CxElVxkFhcV2NexKynGQz1vl8uq0UowY35eJu
kB6fe8qg55LZwtlDhPGRtdyPUrSOISrroIrV5zp/zdaczrc29vAA8BlWyTZEEMyzPFPVoxAuCQv0
vOoIJxxYDTlz3ZCoO81KnGKCiTZ5a0fiA5Zr8OilGQiuiA6kO7c8+Ioh1g/BmEQ+5RFSb/EDJlN5
IG1hGu25XIVzn8hAwzWwXP793QkIJeeOs9cVz+0O9gferb3S72IU5oo5Mf6C89gA2P3U+hOwu6BD
mx5eIIWTsU4Yc9tRRMxUv4U/F+GLqUglLR1TEBUxsGLrzQYAelX0EchOAER0O/H83HTC3Kc1xunr
buNH2ha9/jpllwcp3PVqs9TGJTWcCf4odonEwqmcgeORr2C4q0ZlHKugcYyxlfq2UrhxlONovRiA
cJtuxDcWLEFTZtzJ8wIUlx79HreI4vpG40AJBawtDhEEaJr61ihaW7ygDcAZCcCE8FZs9hy+yZU5
dkfp96rmHwC1HURUGjYwHMoH1shU1szmL3UsNBFaFcgdbG0+0tAnqJCBRcAO4BntxzOTjezYpcoH
bmyDxKuA40v7QTmru7AEDHWGfKc07S0uDh+F7lphgQdPVuBH7TRJt6BKQ6bgVOkIQiSPnwyOiQJg
cFa1wal0mwXvyZWDt+c1eU3Xs+h3VvKp9noR97qZzdS/AohRsmzjSQoxkaqW7HD066hSIbZcsGEV
SCyFPPoIXA7ck9U7E7vjLnhFxqwkwN0ckh+/CQnx3TlMQUNijS3d3QmktuIc2WFjJ6aSXYoWHF5J
UCib2NE+tY0IFIUYvU41jlNWHtqOigLjwnpXFw0+nGtzOcdrdzBTytwFj4NI1Wu0ZWUdcqcdPzQ8
z2f2k8zm9d/hj2QH8BT1sfDtqAKYOIF+/PvDoPDis1+RUO8Lsiewnsw1jk7mDUAFeoPVXVXseOQ+
/sA3rZ9zNhOHQob6k3uxvumPhrZdcEsr86YNl3LjW3gIcxveScUUH09YjDRvDuqKV4WLoirtNeeu
E80rZ5mtusoW6bB20/TXl0jQ1/Cs8hUWqBZ2BL0MMekKktLEig2GdUX8asp+J+1UFSx5zW72yCsv
p7LWoaS3buGgXbaakmr1BFLua5iyNtMavdQpBXLTl+B0g/gy/cYnqvyLEtH4QArvzEHxv3z8kQdN
pGU2fkzraCF//pP3uJeAxwbPAPGPzaXfa7vMgoxuz1Iokc5B4UmqpjpSy0K7Ow59Q9nHXwEVCxXD
qwQphTBPvVA3H7EHeq5v+Ucbj9/N9c5BI0IubAKtCD7ZkBYBqPM16/Z+Df+SYjtMAHp++rJstaRa
fQ2vs/kljpIaQuEQ6le0Dlscls0m3xaz4s0tAO386gFrcjbMacm+sKHGaDLHnuh9fu/asnSs0kHu
UsJkxVHdj1oO1qz9dvsO/mXffSRpgw+3OZwwyJifICkvQJnC8vZYcfY+HawZUMtq2LvjwfuVbldC
u7PKBAkOAopeNqZTmuZXo+t6tmGQXutYGXHDkCAE+9mZSNMcQpmFnjLhWQowur+nLaWKswUTToCe
mHJpnogjTq/QmrxOdhJpXBsJKDVWk+ql6g5iTjz/hthHWk8lEJFmh33KYVohB0e5ZoKqBjV3WF5W
C0KwztZfFKygzg4OklDaD/7/mP2sPm1XXTyge0JXrgKTUugeou3Wq5oi27kdo3ddpWbZaQiBFaGy
zLSPRHbuxduT5wOBB5aioFya5TsCWw3sWQ0D0GLtXBVKWtCO6qyEyGXjmUFSDgXksJJdKucf2eB2
L2lJgFsbgGHPFz06RVoMcgxWafHG7IcTY4vRoPhllCQPHhjDuqcfuilxVk6x/jNlF2RO0/o4vh7G
8g5/xWVtQyD9Ud8YNI+wyiWdUasB7/HYr6DTxgdvwTgJyNGU+Gwx6wgDyXLv6fF5Q8X+0KhKn0/C
e2rqYI10s8v00qMRppuBQsDKmhNQNFXmtyTM/CqKVNsgbEFTyC55SIzhHp0MZxaCswbQXjrEM4RO
pUvgE+Cl8MnRLh6zGUmpxVzGjN0J2wuxwL7yyKxN+BVfe4VNMAQbZxwqJWST8ViJMw69ceaT5a8P
REgdO/LACNXNPbGKkGPKfJIK+YOdbW2X7Uj+ZiHX7yus5Df1UWbMoDRzJC/6fuHDiXR6tC3kREbs
87XvixFKJ7fNv1IC0zEzc28Bgr6BWJnmXXVQCi2YhlMj+lwhp9S+H54tKwNu54mg1ImLikqT2PKT
wuIbJ2qRVehBnxsG5kvcbqYqDSTXw8nXNlbCgUIiWfH7zU3sSaykUq+uY8/zph/CBGw79fH1VEWb
j1h06ZdO4hcULZ8yNFCUsACO19VS1xCwR2FiT12HFk4kXZvuwWlbp8pUqj1C/SKkqMoYSPnMUNk0
/9CSIOmbmIhkyhQNswK+Sv7PdmWPakDfTrOkBmowjTWtOJpze1gjDiD/cmoH+U5PKn6V4EgGQuX1
EexPdP05r6n1K8s8qCoxPhw/CvH4QVHJGqvNAr2bD4nRlniOjAE8Ov5yaTt56DY0Ey5rlTdOsERM
MfKRGTmWX5wj7YSidU25DnFCyRXA8WBwm88nsdSD9qUCbTwThBa7i4os3WpvNLMghqQh8bUiIZrr
0OW9B2rbbmy1NhhXImMxX07jzr3ySXoA1pYs5fucE0zpgkuANAOetUqWLc+hYq/FEme8ScDxqMXA
SSQiddgCH7hIsXEU8zp62WlMDZj5WVIwc1p+kPU0mRUaUSJPfDr3pNjYuiXxIgnvnVnjL4o64rBM
37nt+nlWYsq3dKRFsPllksFvYPLRzVpWE5Tu0Jdtc7lEo/H1fYnK1Me5vh9kjNXE1we5k7VWmEVZ
vrsakoKvOzPnX3KYMAuU+9h/bddFrSoyJYjS6SMt3sEOjncw9N/WuhEvjPSg2n/t0lBrssBaZYYm
3+eTBAhDVCBFxYxyIp7puyjqT00ywBg4WZQ+EVfHj0YcowmcX8lcHh5LBt8MTVpU01jHas/yxaOI
RFgpbWC4vuB3aiN3/S0ZwVi37uChW2TtA3d3GwDmPDTwzNPAd4E0W2HldlKoh6GYpv3H2FHWj3O3
CLLpkWBkCvh57qGvWJQzfnmN3up9OPslPLHeMBwjjmgHNpluq89bxjcSQr+gTEa3fZmeIDgLxIex
5t3v02bkxxK1lFenEfzc1s/QrU3HjuJMrbvvpKYH6FzbmVbTivcVbZZQcYMu3PY3zLKU5E6RzeVZ
mFGFCtBhGVRlD2PIsjHmXBUnY9KpY80eRYY0W77akoSvkpcXnFHN7p1bfV8EABgv9S9Fm81PFl7x
hGW5/4qPmL+KYIKlLos0Hy+g3zzb2yXmai7YMd5OR77HNPekq4vvni/6cLG/0O2wSK259PfwBPwg
R2i9RZmMmccc7orLuT0pK2ZKEYb5+Iq0Tzlr36QEhp451qCeBqdAH5ohBp1sqNMdfHbNfM/6lkuS
dPpFLZ+4jPe9zfeXsqFpmQxZwsDJ0KzzRSCNw8GTfR3J6RSHmgux8BnHiwp9fudBtJ7/LH4b8d/Q
fhz53jwaF9lS1r5R9Pk4ZWGaUG1rUeVoiww1WGBqanR8J4MLXZMDHNzInEkxApGNtkoHCKP33BD9
oFD5c5ctiX/pHSKK5YwLvrPoSlJldFUdCMgZJxSFQmqPvPaULcj6pdAnWBFLQ5NSqG8D+XRMGd8W
dJ+U46jUSVsIBM/c+IUv/x8TL97Ndifhbc797AN8RWUPqK4JtZU5KVkPHdj2ZKz1wcoIoGt/XO13
B7MM6vrqSdjiouVh4ugBGzT+SDF3csS3RUF40B6OqtfCl7+buSqufIxBzsCw+m2FtfwPTcmP03/Z
2ehRTYcEyjMAHkIzGNpvhWHP54NPUgRKhpX8W7O8rsbWj4ZXjj2SCxh+wt/RHcy1nT9y2dehxeXG
IO0pyD/KRtR2kNQnXCSw5ObNCUF4blyOEQ8bmAQwz1lLqlTmdtKInKPPFekamRfUvmWodxZnIyit
8+tBFCwe2KnwQQcIIQzccMk2SYDIuJfbjGZ7nL5MSdUPtMWDc4HwDbeAz/MX+YA521sEngXRVAeu
pQB2Rr3SEnZ1ERYORuwHrIusNmE+CbvfGmOmBt7oJRBmAD33O1uhD8amqAHl6Vpr3IRzTjJM0DwW
OzcO0zvlcsaYxdBSHaHNoxr+olWXkaijSz66Gh7soGiILyOj0cSNLT0XMzgTbWv+2ehBRUZAx0lm
/RJF4IBWL933FPr4UjaFFEPK9HkzjJgoLIWF/n2YNQxGHHV0ou6rboPbPUKDdMATsJT3Y+K8+dJc
aGftnObWH1AtIiOufyOJF4j6gZX2bDrP8RbSfOQWQ5tvMgsmxIW7/6f1y/LFishAfLrbdhZvNbjB
ynYWKrj1VHwOevPzB8vsV2L+tYIe4kvbphf6SivklpLTjmQfF0hNCBu2YYfpjk9BJ/KMeeJq4UJ9
FSrOq4aIQP4kmJn0e9nUGebWFjecthDXUKNXZuLSjRDFLCQkzPNGBKGa9Wql8AUixKR8+7UgInUb
XCRyrRlZWrhAXhVDSpsjxfwBugXYEN84qx7T3wQa5sMo1gfNc4qC4sL3BHenJO+LwfrL0lPUIwrQ
oW7faoU+D/qKtYUjVESOF7tU+BxQONQ/EiV0l6nDDdWQoRNva0ayma7J7QC1Feq4e5RykDSKSvHd
1GbGuIBCNXUJPePpnB9l4ObskP/UwdUPXokCro2E3kNoWxIl+UkTus6oTv8i5i+Kz/2vlGCQ7Enh
iZnIfFG0Yd7JQNgoZU9gWubbmV3TDXMApVfOYd8Z+xGO9w57OppzbRV78N8qyOHNM5IaDQFVnDEr
zTBIig2+awdoJ8jrsqWjn1RKTXSRZe59nYa5yiL/HG1Ue50IyKAZR3lv8a5YSHZ/grM9Spe4qFXi
0NzMYsO0Ig/DPr4e7JtSi/PeRnubdz5MljgOLe0ToEoro/9Jrs7KS994vtms41w9MOGUK0/Ngp8J
vH2hYnuWWXJZ4rppf2+fUx/rnCOzCPnV7GWVDVT75K38oj9wzT8N3ExofGDiqigPqbGQ462DH1HL
2saksJQmE1V5YMGeSfb3Wrj+FqQmnnIsHd4LVtWfpSoYxMjm2Vpl3XEOK+NdXU5LEfOm7zRprg6G
BMD7IWusBcYfqhzao5+SFup0hZWUpya70rrXvaDZCK1YluOyoPfwqtXV58n91I2iFUwuM6s+LHV3
DqFYqkfn1pF0Cq+aHS4ULO3qtYfpiUls76gXQYNi6Q6FGerrmHIIbZ/nJxoNtl9viUxUHHKiIA8w
kN6AsHK5ULEEPCiOk/9iAZ2Xo/thVAhRyq0DzINw9bCt3VNWgfNQ6gDDP/f8+fQe528Jfxncm0Ya
2eWaMdTiwhFyS3y8yzqeYqKGvvufif4mWqnrlGtiaIYZWix7+Oga1CmLBEEnMEdnt8KU34RT2ps3
DW+JwV82vp3s8UX3d1b8YSOiJXpUih8jxpwoon08BdKidRgejF3qrCnInlCcHmHc5P4GMThSSYpt
vpwwA5qPHKDuhctvs8sWsdDHoGlziEFnv4aEBBZEj567nwnjPaO/aaPm8tIwnyas4oaDDaDodMRP
VxCXLSlPIVzBPpiaDZRSRLybfjHy64pRPJJfdqXq7IcpNea2uChAdNv3BjJFCDDHmDKMJCfW3HGM
iHtQ3g1OoVk8gDidQRyEjhVPhQQxOKq7vFqO9JYj7FCOGAmrL8JgEhUWExY62txdHadab1wYhori
DRDOA1RV5BUPBcQQjkIqYB2HMXA3Lps/zZubKzB1328keHYh61QLCA+W0iVR7zRDBDs7scrLH5/E
0i1gbPhlIL64tqZo5xl5XA59ckloTWULhy7WotTC2KiHYv7bUfqiOQy6R+EbPlQm5oO+lc7NyPVX
1SB6kmfI7ZAVfCPxLeqYK9cs6v9JGIuaXiUo3tkbylWmNvlVWf3nHDzs5DKZvDBlv3PPDO2MivM8
rkakg/uk9xfYHrB/kpURFS4fqeXdaYOZL66sNHI5RkLpfGzqs5przFKZ0nvfZMAwJh8GmSsdgCyj
cgJ3hgMkZKcL+kgaVBV7VLibnXWLgbuTEooJIZ3TCKe/h7G7nm1QvPfdG0MvlzJRUnrKMU8JMOYx
RmL8QXupL5fX96Kn86KGF4iygMKdr8f2OF1TCr4bVANqMjzqjIMdabwgaR1OEaia7jH+CECJFvHj
1TF/g36OXSBYEYY26CVY2m9SlGZswHTJr1qJkOtC2vPxQPolIGMBWZdYUUk2AUnf9+lxDR2Oa1Xz
JK/A+lAF+jillFE2pofQgzUZXQV43uIete26RA4k+ywEvuoMeQ367Dg6DGF+uvNVXqJ8dUSfZ9IT
lbx1OEYEM+vyS+nlXH5CtT9vohacTqkITuV/YJtJOOWDKB2Gmaf7ZDskQSioH8tEoyZd1tSjK/fl
450K5yh1Vv/jVq/RY/1ijRdurOsKOuYjR0BIrJ7sgOUhKIpOokkL70oB6AC8LbVlVJWqzhZMnGNz
FCoEAfcokeAQliPuZJk8QLvBIOm1g5irbihcvDNtN4WdEabG7uIbBm7WMTxFTWl5fXTAMFAzxmQh
mS3DGzJz5+7NfWtZXCt+06CNb6sZaMipQMj/OolljexG+jykDk3k2ghTM5XpPeiLhAuwZaGMiUrf
jMdjcE1ZAja1qGcxmxkbIVcKLuZEhoO9E7ItPyy0N2PvXEIt8ofED45pPq97fZsSXxsED8PTKeBo
Ctc+KEeEvhs8yNAEB0EVDpskVDQGuvQWj/i2ddERhVL6qsOw+nPYpOpUso5ax1zvAG6cL95PAhpa
y+TYPzIGtpX7bZjLsmqyFJWcBHRNWCajfzJOXl+FZ75jQgADUbtxdcdc6aYdLhK8W/oP8fD2tUQn
eyascnocwxPJP8BlvmnniAxdIWa0NT+AJ2t2XjaOVisnlvMKPeVt795fRMgK6vDjkfjAthaijqVN
5x0aSgdQ81HYuM1YOi6B4mg7eAkWjqmqCcj9rAgA4BwxIaF2dNmmfrA0NTct6jLY1DEUVkPQcQ7N
mhf7LGP2OYEeXyfU+0kg8K+Qzf++hkGssRA53UDXPf4yLCQNWOi7ahpFtnaVY85xxT6XdbsuSlII
BscG0NrqZGdbi1JAixzx9RrL9n6CvRQre7vxAVRrlLE9tUw3U9hzHA9MxdzZdYNkHOJQmjvT5feY
9T307y57I8y1cX2fuuuhEXTczN3uZLZeSWKEpxulV7unVeO6Zxf2kqr3qtBLfdRSLxVhLuU2EVAa
4+kvf8k2nXiDTKXKrinsCdC2I4hO96/F4IWO0s7Lj8bH9VcP5tzmuENfxHW6n6BYVlxBjQ1O0h45
DYzZb6uhiJyjZjTBEpnlJituQ6ZWTQAoGDnTTHo9xd0v+IrcQHOM2NzmuCtqsUyZ3n/UMBnOa+nD
tl3NGTEH/i8A7Q+nvd92B2/tVTG/3YV++2Gv+ib532oqyk4lCdbcJJTaIJixp6oLg3oTKy5BhjO8
qo+FHwpanXfhp7F2zE4hxI1mhfwoPsaLGpU3TDkxUd4GUGbdfTv0AaCb75XwvKCuhhFwaYIBcEK5
8SCZF1ebzSmvsAHg1R4g0LlK4tNW2zeY9bdJJBA1aUrneVudzi2q/eevPFHu8U11yDRl7MJhZMm6
yaMlZUqBDSw1daC0EOh9YINUvubtN1RnomCHVgBsORkdgZ1/0mjq+jE+5VZyb3Q15VRHrwN7hEu9
FTx2q4OsaUnYW/bMf4zq1gXMoYdKYuF3USfqhwrpmlHaMiT0gKcFl2WsSuY/fXzjMt82QgQ49132
ahftxLeGsniAaf9xhZyxBrhQ2j1zy3TMOYoBF+lqNSfvrlaHaGeD1MotYqhfJd/PSTGuMDD6n+mf
94AvVDyUtIF+REx1Wkm33qNUpA0yk+MsThG/6gMIaAlk6MOGAUZh91GsjOUM7NQwgYMLuHCcJdUy
OqMVdm9kx3eMTIuJAk3XaiznqiffvXfs4H+nnCkHx5fEFeO5WeubeDbj9slVk8hfEYvmh3xan5El
mXYwDCuJLCajVcBvePrsaIjLi8ldxktuRueh6i+ypKVTXWtzwvm8fyTHDYx/xGoW8wSeT9sL5Ffq
lrEiZjBavL/CCnr93H/eUqen7jrs2H8cr7IPWO98HGPc3VdpmjAVY8SDuETpsjAdHpy9AXBCdlLT
RVtM5u2lFMJBk65p8rr3KJUo+NTyl3+fShG7hdS5kWitRWZOMFVSSp8vsKXOK1NuMCe4MM7jKrqk
jmPo2yyLycorte/esTKzQkROihmGYDdMvs1qWsqE/606wYZkaH3bUD9n43+y54/EQ0Wnf7jF43oW
LMQgvcKniI8RSS/84w3qdhlHpVEAqQlKtFPBBfios+wnj6ptDUOCHhnpoZuMg6450eszGmxgRQVm
4nh6g8/f2bn9r+8okG8LPqY4Y9S3XWtcBgVTDQzXxvTtEuETcvnAH6yZWItuz2hfoNVp80liTxCJ
aWpg3N+cuhIVSIz1p152M1SwVXySyRj+L5EccNMKKm/lXM8Ti8OSelDLCMVQrBm05M1e9atWM7xY
J9yBJhCAV75cQNHqli3fhfZ1fY0sSruVth5HBiEIzBXSgGbU19mankKfY8njZlV80d81BpFj6X1q
C2uzVoEg+M9NZtAB7gg5ZscRoNKrr27G3kLbTa/j7Hu8nUhkRoPnpbftZP1LeQFMFKREeW/KKHr1
fXI3lfBg6yvTL2DzHq7OTXc9jAT9wpeT8jVg6AAcnm5uTdfwRtPxBOhtXY2RvIWVUFhR+2epUIXL
AvJuWK2xVqz1ApPYOF5qDUHdIpjS1oJ5bjeOHMDTvQ9e1KyKhCO6R4GezCJE9bpVd8QbsZ4rksPu
jVNyJypphE4XDIek+YBvPbZ1BTfAyhwOMI7O1ns4Xd2iigf0lW1ix0/F22K8ORb4pWkv2IxeZJCk
E/xLj94QIJ5TIasXgwJTQ0Ja9+WWIlKsIHG1CjODYa57XLAEqc1CdBO+FHG/zegLFqLSF+p6B9ji
nJR2RI8VY3pEKGfG2WoEJ5ArSiuQBi7ErKV8adsdMW0EMpWnxVnlSOcnJU+6QpdVHvTrUHYXASZD
rTnZ1A1Bs4YpOAevXiXK+zdwP9SQFiGX76A7PIu4sm2ntPCJs+bHU6/aqJayikMxdAU8SigZ8/L2
h/p1IcuaAo+658ob5UGol/SxC7t3kn2+ZTjHpDnd3kLfarJPjGjnppymfYUkpR6J9mSlwKdCzJS8
/MeaLXIi6bxIspd/CPQNLRkxLVSEB/4cQDp6T2jhcM+sxBLXhHz+NIwFwEjo6NBv7kJGs5XwZI5l
12z575Bh0EBGyZFn3v9z/oOTqq8xwPMnCZ8OyE+IsJHVFGT/r6k79cKR9oyC2wH3hfQ2GNKm9oke
qvALE8/Nz9PTdwXQjqkEBkDdcOFM2cLliiyOaiJ7V8WOrOxndoXU5fMXxjtH9iDx0dKhmeGqRpxJ
meUZSUOJ6uPdxJG/EKUjaAdCq4Nok5hzK5QSI0zbknTffF6KvP/WywH0dwXJVCZFj19H53SzP1/h
Hu8c+4CbNubkgZnZiH5Hg6dDuldQl+mpQlSI/YIGrlleKa9G4Thr0mtAey+MrYtt99wr/PDG3i9Z
t9UlvspTA7u9H62oMjwnfaFxlChn7R52BG6oESLrtBrW+xgAPtT1o9CMjQfl/5cI3xLx11CrG61s
dfQCGeNl9flZa7qpT7gMUcpDg88Zhs9lwvWowSxEdtiw/x2V706RZvZPzhSoUqc+P/fy6lJ3AFJJ
BcDgAGlJoyML197JBYchcF9NcwJ1hlhedteAt4UZh87c0xPjLFSZRKVI2mbQpsAROJzPranqQLjk
JwFDGqtWxP84HnSp2E3cPSr9bY5qaOSJuGzUI1ItnZABD6XA81bV+U5IWR7Oy1NWFsgpFDky3tHi
x5Tn+9+9iyU+wzMpnRoYkYn0VGOW0Re4oCfhPKZEBfVp6SqN1hDMGjR1MNk4eMRqEgj3cSsy4dG6
x/vT2af+JBU0+A5K8pNyoBiVRCbuMx4MMBkSU998SNJH1URVWinCcxN7mEIwZpDghv9zGct4IGsN
3Fv0LJWy5JCkvDTwMtj7AV5XwrBU2hDiMLWCsVa528KaOAbYk8yNdoy00WpzdSMxdwzTdgSJd8nh
BziOU6Nil6jFcDAEwNLmMXjER/kDkPwo9hesTZ7jDq97TLsWvz/JJ7Xb0KTCV+Yjc/d18zJwmr1u
OOUiOQL0+6wLgt5o+d9BDjqbL0czGqoiF1FjRH82Pl9l3isdSHCYtoyr3bclVI/5q7ln8TpF+Tup
Qtat5sE49b75FFYl7yRKhAmYa2PozDFxmbQwuZH2I8gUimKZEnTm/dDakReEFUdq6KkptKlYL4Rc
lYFcOX0EfqttE2gdIeD8UhXT0II63mDB7tmq14dEC3gY0hom03DImamcSsX0ZhrfIg5dEhxoIvYN
YcJRKn9HN4VCScyqWYUtUHCxED3W4HC7pFo/l2uTLCZW8bkzKZtaBoCYpt2Nn8PidH0XN32/yav5
wpmNXVlrAoQ0KEHLNqwi+3DbpWauZXQYPsGRsTtZ5lJne2rhuWymq8g1rGklleJqsZ/paIT8aQmF
+/If2qJIlF00UXYEU3ZFNAa4zdA2RIoQwhw5rJ+U5Mznq1InI488dcgV/QaW5sHo8S8m/HWUDeA6
o5pfk1sU0BLJCMp5v5gPlT20fPkZ8ouHGgHvDQZJfQ4uCOkHsmcCQ5HUHc4QDJ+6oEKdChlsgyoE
ADQIr/wEjnJT9X0x4XLyGfp8RxznNJiuhO6qoCP2xP5oCCpTaZhR8kl041kJwOvYiH2TXnNrCF94
T8H5Mm9reFOL1ft2Tg5R58e0QA+Hlx98pehapt+Ia3Q0HCozN9a9uuKxupqT6UGJbpT2vOgRiXVD
mkurIQTYEEpm86lDI5ES0O0US071hyRNWFJbixnS10Sao87gRaJF7HlsQQq8QHrJg7CBKhc1dRtK
8p8z1yIA9BqHxAR4u2mw3eZCyUMUj442ep0sq1JQhp1RuZtUWuxtdv2SXKD0CngaFnc5xbw/Bl3f
MRC0RlGa3oSDK0BiE5dz35QrrTOpZAi1Xj0k/JxbpN6slF3h4jOz/+Y7JNXHEkLTA4FloXamFoFo
vuplYa6vlQwyZfZZNEh6kMe71vbu5fLQNrMfuGv4jGjhpaethGteUbvqbMQg9sf+cZlAEpE+cRUD
nvQCFpaMq3kvJKDJnELY6oAP3mxLOZfO0MmpFueqSPLB0FV9bZzYokYYEgK/KSQTk10ZQb+rlSWD
DY0xyu3vaS5Q+YiqnyN4+MO2q81HNljy58vGimJV+sPdR7XASmA2Xozylv9S5GaHqqHAChwe/4QB
qFblR7hTtIbrVtc41o1+JwRkdQ3LdT3Uj12pLZUWG2imBh8bmroYtC+HtZGy2Efv6LCmmqGqitsB
Os60aiGgPXZk0DldnP31nm3CWWxSjDeye2P6IMXaWUxGIKh/7MC355Wyd1IamXZNZbdk6o/kRNe+
JEyUEYAWfo0lJeWlW2y12xaZmwwDAK6DXi98NSLBWkyTfJ/7xLzhh6BuuyBwksNYG2tYHz8U6gkr
CpUYnj5zxZwbjitwC/jdX/4Hyw+bECSQTQUSIEfUFL7JpFEsE7RmXKw1LTyoVqQXhc07jXMAGcoZ
FmgjGv3wDlY9vqe5zZBr2AhEId+eoDb/1dtNfHMNva3aoyeRyWduiqQzQfS9poz+9/JvsCveV6sj
TTTWizWU3F5nn9FYeQKpDecfedC93uemVb97SX6zj9MR8Q2sq27senRVAHe8vWsCoHPVXThXedKU
QlFyAPrEWHZNgx2z5WhHxsZLgI0OnuwsATEVOtNtWGXbiriEZFp1GA3Y7O/aNBhueFsn+n/FgHzs
qCMtap+H7CoEc/WEHHuHdNdopHTnIFa7ikppRS7/RAwgDv9tMfrZD/fQyfhwcCSBkNuxuYZeuSUK
Vf/jNh0plXOVgmVoBdkoK9Q/IBvCYVUvezVsUH8sgljKq/OJL1bmZz+RVKVvEhZXx5f8RmEVZ3FM
q7m0AfSSnlwVGbdFWkP2JjoJNhoNVOQnMqNKDw7xqL5Qnuqmj6Nt+ACS4yiqGiorIAvZS/rc7/1t
PuWhSGi9zILCteBFgf6nF7IEF3dZtsxnL6+o9LnrOFgh1E/rQgE08C/fpsGzv+jI1Taihe60lvr7
rH+UX47Q4OBfwnpnMUta0bOaro6ISNCdcXKEbFztQfJiUkLlpN7qfcAFf59BDbP5o1lPFvLoQL02
/4drJSv29Vtztj8u+AdoztO8ys/eh7ex9a+YVkLqwYxv8lypbSwgpUv/Nm59YZp0FbLBKpynwrzc
BQwjw6fUsIvdasOQPKbNYDuGzuYVIgmIzfi9R58dKOS65zlQCprISCMzhB/D00mJJ+OdHh2zt46c
oIzQZGvR19giuh3pV9qsZ2Hp7eMkyXg++Zygh+ONJd2CNTjXgmW2r8jgk8HAwGCbvhh6qGN12lPr
tLPLzoNBk52YAwI1zvP+LerALeRsGmA2OvRlgDSJdGY3HsyyX6ZLrCKFE1GOMqhosd2akqClXutk
GvpeZRxuIeGq/EEMqJmIZF+Wg9Wgz+B13WrfXHnMACJRMk8ZlHSn1MEcgZpsY4kc4O2rVvUEmQ7q
EgHvtQ1duFubZYxGT4Zmx9+psIlK9/gCuQhZy+Ghx12iYwGKlrVUWHtIRp+S8UQjOrLZxhIOFTtN
qhE6m189HYu0bzgACmpwdZqtvujYfo0CbEx5u4SKJp1uSqL/Cncw9M+ZUHb+dYV6E24rvLmAzMWU
Ea+wcqNhyvt8O7PsYc0AZj+Ktb1eAcCFw7KzkdIAPMxTwuw9eFgCK9QJ08krszZdz3peSpPwi9oT
l/oJGV40flQYuMyShqdXdBmR0nl+qzDSMZno0lGI6S2XGySIFgd1BMNK1VND+zuVx19HlC/fs3Qx
gRcTzk92Nfz2qksmhXqxtbRrFnK18X65Est4IFZkciyi7x31QQUti6e+V70RJayVWSctMnbA+Ugu
xCiggKo5X70Cp0pdopumknZe9l9vHB34r9l2HROoyJTFX0UHL58zvTueraeQvOhRTjtseSmCi1NU
drjMH9uc13HKLPyF7EqZwWB5JVv6mrf25+1yafltougAS9q7tdGufQrq/CP67s4ubocyGtgkT1rF
QdzsG/oMiDcoTKUkaaatIsejfa1lbtO2tAFzRKv9VJ51GzxTib+Zm7znaoqtmQW8tSxbPrDwb/HL
uist7Sgusvt3tpg0zP9VLYdqD5jACDD7EYFATjPA6jLxv6RfxLHSll7j0zj9Ohv4oMUds+OhuGiC
176hvO62jI9XJ6kLLJlDlc45pDQgh9n4VuGO3+qOPJj2rg2tvODslrUzmLPy5QrpWTAvvJBEuKCG
B7P/znWO0Mkoi6csVHrfLtW4yDRoWlQaQ7BTxlTpER+IkKrpHf8plQnX4dE2uefjtazb3zHuJfj1
1QiPpJCl4FHuQs9K61gFzalkoK0c5tazVLtzFwmaGJawOlfirCU90ffYX1Et8Ij5HilBLGFQsxMD
Qhdf9AzHx8wLTFlUOU0Yximc4quPSkc1fu1tEpiXJfeFj4bReiaxFZAUg90S+vxWEeHdkFPkGkZM
IGtbNt+Y9YN2FyAQu57hqQ91qEP+OmNhInL9TridcwjhaQw7831H2o2ZA57kfao+cm67NqQBwUjJ
nV2VQc7EPPIX7uMiROH43VHM5jlr0QCoNrZFSkp6ysv3jivzEGqwo9xj+jASI5/LplVwZeORjhNi
GaxD2ikDLB6tUZOlDRMuxtJxWnj0XlZi/yc15oryZWivd1yjlVd4KDZCYY3Oe2JGh/Wvtl+zrX+S
yMqcQCxrlX0vdUsUsJw6P2Mr5fZV8nvhxJH1BbLI8JEvcMzNCWfXgeOR8V+nQF82JXvupldAdnrZ
ZopQwfi+XB2OopnYcxb6sXz/MKqm9BFsne47vuGL6BKKHnIjmiycD9Dp2HMXnBs6MLraL4ruFT2u
twiwZe3kSJmWmqxMqQQ3utgBTLxUeyvK5usJRfanOWFIr9z/hxURCb1LIUxt2Z+HMuOiCeEZCugw
Mf0z+hg9py5Zxw+1FSGUHVh9tu2U/20gzQ1/hupeuVg7ErxA1TX8WvTN+F8NDmbypgaWEG/KX3c0
GBdkw4pR5k3lI56OgUsod7wuGlCARwfbHhrIOz6TbqmLYDbNvjLxVpSjYk5fvyH2OhnUX+GWyfdd
ICEIB8/wUCizIlkaPkc8WfLtC0iA9tI6FODneTGzWKXABcrKiPJdfZFd9+T9BQ8/jJORTjLfi+ty
HVdPeAkus5PP24n1nFQc50qDv46WIC4J0m6BEblSj81IjYipxD4jIn3Pq50h8nSYpwkdh5u7NAPO
PpQZHXR2RcwViiYP884+opB/8sjx4yvdvDH7u6UiBx4L435ngWIsr1ddPbt2/PdO6q1oe4/vrmCs
vwYNEyWhAWwgCuBzbAgZFcnCWTcM6rWQy/kb+MvMtfJ5yU9vvW09nWx2KpaTGUKJHKliPDT5h5v6
uFHXzOPKo3749dxXkLY0LyPhTh7yWTMS7VcrSGUmCledISG4oe+G5KDTyeAhY4z0+Esd59WPE5Ym
d13NVDfuOSQ1iSeIJRVlS8t+CcHbcn+Zv7KnbIsS4Aqzqk3LeJk+03ZnnpP8I6XCubE+UzjMbqk0
JFN2qh538TTrccJiDprd+SSz1rCcjiAGoKm6GrUZUsuWiu6i3Vl6sCdWY8QVtIT/KzjbQmcjWv6H
V1WXDUVR/HheWNt+AqLFniA5sTy7/Jg8BrJzph29s6rcoXe5AqjsCSh+OPVxP5f5NR89K8qvDg2C
a071j/EKpUKvw8pZVKoI0WxfZ6QiOJPq7o3R6O+fD2gLSNC1wvY8CImNPDYIrCzJBMKRUpI+xq/a
mJX28yffevvB6a/WG1xcYSFlcBF9XW9r2mfBebHpCt7p13EajS8LhAdBTPBFguXw5++QqScH3c4Y
GGAv+Btxo5m8YTFwHxu8sSuB/KBiI5HT1B5VNt5LBPVt+tl++61j65a863gFlI7vy7NCwo6QjqCu
15JN0XJVQZpBXncf008U9VdobCE6drVSqF6iUKVt+crmeidj+KJ2ZNSKzpFBuym7juL0qf3Hj2jQ
T4qDLXyWQt1b1kUq7DjbTPFvna8TgfjCAEm+zxFLwfNdRqja9Ao1W/6iRvcyl9qpqKc7XdgKIvsi
rQXQpu1P14Z0Y2+MY2zPlaPiMxCF7J2LOmxW3NzvvmZCXtcbobjqQypyPPiwjIYP+bwn0RwU+U4g
9ZhDW0pqKDH0WfsSTOQtbyQvo8zC2mA7cVlVTD53eYRewJ1XfK8+nolZVtXKb98wsMBsRRM7Pd1s
zKDav9VxS69NGXKx9ij+b8cTys04XahLMjfCZUJZUUiGPZKilKbFnPShT2vR7g4fBI/C7c/DeRgU
Ip424DCisDP0N/PzT2mAQz4G76nQHAaiCkFFrLPRH1Zs+1eUgNP35g+P7HmGAB3rMMseOw82vt6O
rPwawaJ2Ih+SrfiUkqgcNXRFG2XSzEskQg2KhRhjv0bkYidFI1vDSwKCQLp2FrEhgq4dAoEYf2Yq
AOsrcjHb7di5e/azt4Jns8etWola2Buff8YDZl4rQy5lp2SBqR/4ikwYZfd+DC2HXgVIl0Dz8QdB
kUkSCoyOJ/N6qCsV2dDioFSE8Mzt8xp8fzk1j8fG/Il4Yw032Ypt+RQ/N0Y8kQkNk3AB1VXpTuCY
/eFVQzOfCLop1Z52QGvsIRPwLz9U3aFp0K+ZAJWxHeWo4RHyQHk5y4vqZDcJ0jS7TnSemquUT8dL
IfflGcth41pygYJxBKiWyHIsJUbe4Sg+OvBSqG1WqBHy6NiheZyBrN6FdtkEIrqnOXsSwf0y2VWX
tZ2sjDUIfnpkE5ANl5xKxGMTImNZ+Bki66XrU3MDTdT1arezAGc5sxwCj8x95utIPN1CyO9tgr02
f5ZnKgOpJ9GcFs2v8UktupLyJopwxBTj0RvkTzbAcabFCoENJl4jyIcAr4dePtAl/WG4HNKqRH1v
AiUUkT6mgHjqjamGtpYBiUMGEhGyRyy5/7iNArPBVp5lCUEnS+BU3fPCGIEq0jJZ0QJAY5ejWhq2
IiSHWhlCtBHxC4fDfYjG/f3kRJS0Kz+C/iwVTolPHtqKJdVNwncHVDncjkcb70rwlB+cyj6AOeKh
/5YQiQMXv8ZH4QE5zBH8JKXdC13NwDl6GztceJcVEhswCVfpIK0cXc2KEC8yEhIMWMuwYxfnbscN
JlWGvoeAV3YvUrYmnRklMP5+0g8AH39psjfYkoiAivlo7fCgLFWhNVz7oohHdC9RZeBDBhCMEYHi
5kRBP3K45Zb/6FYrLfRoB1aZQ3ojx2UpxHML+8h+nDAlXRHhgeTt1MZkcQdDu9WzWZkRj7BNe7mV
3+x/pyL9RkEDikLnR8wseTBHWmQBZv8rDq+K+oVkOyv6Jf38Vz/gj8hY0GlmhUoSaAijoA5nrvHv
IQl3oIZPVInTFNnzyo9t5oxiB0qsb26nHlbu/sKrCV6neTms1xYmI5b0ZYKgcYLLhHyZ3e3xiGuP
ohxCU20IIFd08GUzvjegSbZTrgm2Cd8kPBndG1l2JZcTZ9Mk2OYvijTPox5QuRnDCdzSRVaE+INn
b4w1Uw0xPT+qE6ZFX1vJAD1m0cPDKS+FJ/bOSUTyy9nH6KjAk78oITyaZqejMNHgc/z6a0XGHO1i
4K8wC6cM+WTKxupDcq2oG27i+j4aOmVyApAttDQPg0DBrT09dfh72HSPiHDRwN6Alz7khZpY7iZF
5ynGxqmpbqGJIRo03sTEjIzkBI8XMQmPfecqIYB3+4K1vqJvJZ7QkQcaYlxw63UEhE4PqRul/vEt
QCBA8PpGXnfb9qOha0lkQz/6QTmE4nEzQWjaGiRq0MX8vMowkaPyszPtF6lW2KMCeySqgWpoWfTc
TtKQnXRTwag4QRporlsSMkmS0Wdr4B1oU+cM41AKoKGfJwicz8ToY+rCTYHbXKJX/oOfpqktsna9
sqUePMxqwcJnVF+pWwPipzz463vZPXwyGRHGxjnyfTs+C3OoTHuimn6R6RCx7SNRbKugGCSUW/p8
+xfu8tXDq+4ildsv4yv66B3N/CxfO4iUFPePqeXUeuIE7YdI4hLF07WkmVHdFU982MVxb9hX/Y8i
7tb0l+7AH+jNx/GEe5+91t24mRj0H4+LhDcHVXCZf2G+eoQk0Jzhj8ck6ukt1xNkz8ZzssOMLObV
ZYwGuXvIfnCWFU76QAJnSOg29KlmBdYoYsYKLt6aQzhTcRNYdDCvjDAHb48cPDQC2WtylSI+Myr1
doZWiH3oTmDU2Mw46DqgvHjfZZ8d/7jPCyp0xGWEtEvq2rD1cVxidG71MWTDj0rLYwYMKg93qfV5
XxNKV/g9k50pfV4nhZ0KB3fNiFaOukBVunyMKEpw03M/Z4W8l0pD+NGFUQpA0J1dUTiK+zPqUQZi
JBnS/EdgWyQ0ERvY7Ye2Gu/Wp+q8SDvNfRkZWerIN1OGSnZ8qvB9RJzVo6U7/S0VOerYtz/8hGvx
02cSkrn69tVI6ppwEEJGCSsJDi+h/pImGNI7DxY/F6qDMSFXjb1FmZS0dElFTHXRqB75QcdGdQsu
iaYNbSIvm4RWc01U1rIfqWuWk1rZk8hqzGLI63aaiP2n6F4M96+mM0tJBboJDVUYKZCO5xr0/prQ
olV2D9Hxd6joYnukxEKIHhq9IZUw7e09NlnDH2Qukuz86XrsQh0Yb/SsdoDOM93avfdsTV8Ialne
KMd+GkXzGv+ZbZEHtM/nvI20+MD9bIXNbLWPkj1NkeMB3IQwVsmdlU8IAbsxWt0r1oroHSKwTPXu
vV+WGkvxQetx2RPivxPOLU16gLUSFosBp/AtrEfFKNYKI67qgxYv/zDm2wE3Y+91ULDbcJhk65qE
wMsRk7dR4xlm379KwylUeaPneWKfUHuiUcpmnJ98oyJsgRV9uIbF0MrOgcsWFaWL4YWkguXvUg8P
k1pqh6nd8VTbPLCanhBktOLemvxgSN0yF41rOa5Gy6ktuq35IDqAPbesaVLIei4LVmZqXEyTn+bW
tNIXQX5YIrcV0XIYQnbCkJIlDL2aHAVfCK7U5lbm0Ga9TCEMWf0dau/35nqJkPIKjD2/4QEXBMua
oG5trX2cb5yY7+SQgd4M7PqNXJJsSWX41t2HeEJjECJ56adcH1w32IMZevmecIT/YEoVDCQTfNzV
Xf/xsy62BEZiRzU8tjG3R9e/aEagvwk0e3QtpWR5PRANrJZ0AkPHuYm11noloJXiRjvX1eByLmmr
N0zpvLApf+s3AYTNW3u29WdemoPGFD0+v+AFsYV3J8gLhcEiluEk04DO1Dyj4xo9kXDjoWK3/cvy
PKWLItiwqxbtPOndMUiDO3ea+wpQYhVS5BfEreZCE2uMzdjaBpH5S4nz3TdUgLQCwxBx1UUTnFDO
Lx6qs6Xq6sdGZgBtNxgOL2QJU8BzmXFWeQYpJ/EXqIntpQUQ/OFnf0PEa3nPdWqOR3K7QKCl1T9G
5hCvYoIDdt84WuG6T0vTcJE7mwj94umHGNt8/Of+ICH47pe10U2sHXBunKQz+7oqzdR0ZXSbqh4i
WrHfhKF328QNo4cE5oDJy0dK46VP90JL2YIditB2MVyGSqRWTZ6wzXUFXv09aJKpUlmNHWQjMAA6
O92F5YogbSSJUO/tdS9nU0kbxj4o6hIcH1yLR62yTt0kafGV5dujy+5gmzR1GBgK7SzPtCoaD9vy
zGInj2K/AaOWITrwdXvvDwEbH5HCmrTOFGuzXbnLao6XocQuv+9tOiG1QOu2k2KAw6seOL0us3oz
ZpGnuIhVj7Xa6M+n5XviMqxKGS6S9ML2JnvD87amSQEx3CvCZGoLlMRlcB6ckFWe5BsVM4ILCcNA
j+B+Pt0x9MLdjFMYuKJ77Tz4R64YMWWJ8URdNCwYGTBBBNGLsXBWSkXZ2hMBsAcurWpnJ09WLrCe
3xx0wF6HJXw3tBxqU4bNU2h4FwsLdF+IfRdiiyiAAuDMgQvebpZzM2nYEnVHV7Uh2nuMfXnV8NrC
JvgkTFsfM7KZStWiyPvF51KMEt9HcheyWWAQ/OCxe+cAP1Q7oIEZPZUnIYgGBG7X3kDhdb/zTk7B
KpArPFMdCp05SogKDOozHzWpPxZj9S2+l7UwuK6mcplltWQ2u71H4ZCjB5TFUKdryEqqRkI6qWNk
/6CwL6eyE3iHGUWj0QSAea+UXPgndNMKoCPVnpPGs/S37VhOJggEBAxgHwHMRdtByHJslWWXk2WY
V7Nzwe5nsLPNpXYX+gE+uDunYbeyV+mpl/5GCjHTxZ2xM4Ik7W37njn/gVTsGfV6EnaJ6Iz5QhjN
/FJYklHSyyZLYvdUL5RHpkzfov/0pHxAWJJ0EZjf+7rbHej/M5Hr8wvCFk8cIJJ1yEGG4cuwYy02
iPc2GIJ7R493/WAvWOaqRdfgfFDZoV7iZawoNHJSlvXWRv8R7aqM4Rbi2qtsrxNgy/ye0uYRo3+C
rHtKg+h6s58N7AG7SI5UyVHqa2JAW/kc/r757uH7+rjD2qXidqQkssJWdeafcLqMNjkze0VEr4pS
NExM6sWRayaTM8LG2qwmgz0vHjDHjVp7Xv/3kvFqQSKaOJOTF3p3rqMY7H+XvU9vSsHRIN0X28QK
ItmywKvUAXfE8TAaft+iVO5cTYVlhZCTFUTVNrPdWDeLXwGSYxk1kA3p18uf+2rpi/VAbMMnGOBj
mkO6POR0wyaDcP4EoViZ2CIIqJOoPyvBu8Um681tED8Q46gwhu0YphP2BpB20vycH0CwQcDxcSfC
s/ZUQX2B0MVG5MiSUem5Mc8qocw3b6oEUUjkkhTadEV195ifjzWovsiz7veMqoVML90neLqsQSHB
fjluxkzvU7P4GK9zsqiX5wpO85AHYhfix5TpO1bR00u1EWCoq0/XIZLWXsZ6Gyiq9cpwlhAimVzQ
kYdoaC0kncnK5h6Mgea+1eYFrqjqfbEBUtQ3yGH78feECFlAepdjJPbZtV8e2xgIqsDDx/dXApwc
4m5RMY9wtRRd3i3+ZLtCJEBwNwUKTX6ybmxGygubjRR2UJBIM5cTmd+TigVjpWAtGo0UgfeQ+mq1
lfK9aKsdYctsDnNz77lRGX3VX9bqiI8gIT626+edvsLPXvZ3ZMe6i1R95QSGCzXC8ebu8zRDn8DF
4tUoHnBryEQFFPqlvmNYoziTiag6BflS2U1j3MUCjePKZm4UJFFW04/2LTNk4ZuC41sNtj3dwxxj
SBjT3z005onlbOJLiudNdIS3lELID5vAtD3F++v0KoeEKr6d+74eP6bi2AvMu2OMuURqSJU/Cg8e
KajqL+QBEQw4iNi50WmYaMk5CxW6CkH9gv83Ft1dp2z5qa+iUalNVjKzYhLWiMA4VhkF2uX14RYd
2y8ckA+5/YfauuSHXvAXUMLMAKUBiHzNvBWf5NmTxMqN8Ev05BGunql7XfC69Dn3rB4altCSe30l
2HFySredEt2bGuUyiktw6/TfsbY5k0bvXz9FNLjR1twoheH6I4CS6K4htKLJOv7Hb7KaLPno5CkL
ydWgTvUm2YmcMFVK5YSYp/+cSxCr8kyWDIs1XwelUxM9+eK1pbCWWaEBgyMPbk3xffiRGwnd4FYB
mwq/kjx/RCtvJU8gbJg+yN+/INy/YgIOYpyTiSa/lL+bwJgiCtAkiriVvajMKWd6HdCWu1nhIf3I
LSCncdeErVBFrIFb8ytP4ewOFwQ4iEyNzTky4teYh22nzxg3TC6V1wgVUnN1bFa7ZfKmG+zLPAKW
P52c68OBIsu8nLzKwnN0Sohmh4rkD7aggzfIiueUrfHfy4UukyXHesBPyVxxQAMntHZtsNw6pHiI
rIvOawaEtxdmMJV7aWLXoCku896dqLYYvMlQVbDrxasNxWUjI1BGfuS3tcDAWJKKrh7gYCaBRXxP
rXZaPcct0o0uOERAMAAYX8eZIJRXOIKgYIch+OCMokG/c6gTFcILx2a4qHvmlwOo3MnQQTJg5JC/
48EOzr8pfyRZA/4jcx7Uolyq3il/ZTbWjG5EKVQLCrnPhzoe3QsB7sep1yIwMBJTm6NIYe7wvquT
gWnevBjndbgyPD3Dyi+jR+wlQ0VCXy1lECPX5VVFHA+a/IRjowvbHKV3sIHhr3rqnieIqMqDFIvu
CCN8taMa5hzenIVaBDBiWIP0Kf00w2+ngTB6NKAiV3un3F9mYovacrRlsP03woZIoe6kwrK7HEHX
y4ew5N8/L2jrGB7KG0UAv4y0isrhVlz0MnLUtKTx3q84o5LkV1WV5FwC01Gwfr5HX6d2KWjPeK/C
9bH4jRBjKPbLRu6GEQChE3qU+yVV3fJqzwluWjKB9eC5rFxGMGc+3c89qu/BAP5nwzYEpMAc1/ZA
8jNC1E7bwQaSq4N0XanjzTJTG9d3D6qCGRt/EXm7rTJ7K1kI/BfvQDjim0bDUq5VC32/5lfvp8m7
7UYIByYQAjFtWM0XWlMUiiPg+dt9ycPTQyLlmC87vx7T6FdrbiOyvDs8y2O0rYWNqLTex7KlUdHg
WMBN33uRJ0qRsB+S5zUftgYcEUzKK8D931KPpAVkKovmqIHKG3ID86m8jTX/pSqbqrHnpCwy8gOb
nKATV0sEO0Enf8u31i7fYGeBbojNlKqItSwWIxMUdJc5wjmyG5ho5Qlx/VeJRtx03OY0v7LXI+YS
Sf99am6xP/L22+urJf+6s49IvvJmw55dXEgYUgE2LKQ7QkYTlIHnB4VKB8fo6mnqxZUR5isibDX9
ldBkDXSL+MB2tVO6oeMsY/d9/S5Z6W0yEvw9FdaXUbFOtrmFSAHKgNhSRlHiNWe9nOO6Dvf0iZiP
JStBfcBGQzWjnvivDsJLqXLt3ZR0UGoux11gtnyJhUUNVyy2XLLiYACqTE8S13xL5J3L2B9/g+wK
Xm5IIvn48bOtXYpSKp/1YR/jdyymmnqlTzUTgnYRU5ZJywt+lcySe1nd6iYGlMNz4rXORcI8US/i
AV15aBFzsrWgIxS1B5A2PFkvKQIFgQeNbROOMbllxENQOVE40viy0JCTxns6jd4nxmn9ojEDtRyn
YidGsAmpzys/s6CHPPTQaWhu/ytblLs+CWg3rI8NDEroItLuKM0RPPkiIpRgyddC3+BMmPqVjuI0
eRPreVG3cVMj1VsET6/R9RBh4XtILOjVIOAXF8lu3EFW8Er+ehPwTe4PqmBHIird0vrEay9ISwcr
c7XhLBgZh8Z9BRllhyo9wurW0vkzHl0JOdlS2Hk0sCAd1nT4G/GOHXPm/NleqSYV5RN7GfbEidEq
d6ZeTXreD7v5ybZG6OwvGUSjpDFXSzxt9EoR0fMPpE5oCgV9dBBZf0bXDl+89D+3gYwNG2SdjX5C
YCWoe8J/PbeH9/DAT3GlHF9sgTztHgc+uF40dJeiZyIk1ALByyyVo/TS5Wsur8sLe1u9xBXinMXI
XcoYYOKcJzllclVUb8ew+3PCM/PhGESnPx9n9LS2M7zL+qviK8HIFEpGQOvK2Xc6S+g+B9v2hUDM
qx8xwYAOtVnwA4qVo92yotPsVU/Kyx0aWpxOSl9eMPfx6Q1kK2OPLBgLyd/Yoh44rqBcvTgHphBY
qQy2mf9aFqROE7XHvKjH9FJJtfmPwCBkamJZySJwCV55MZ/dNcb233th6jWJVNZ/gbmZBS88FioG
L/VYgftYOn7LA+y6PSU2Pphl2oD0xmc3OoIYe3LyiRr8OsYKwjZKBUW75e/9kUnOUD8s2g5EkitE
TGcpye5lHwJF2mjO7EpxM2Ns49uuWCZAXMIA8tQ2xiZSS+AUNI3OaBY4DOTRxkBjykqPPCa1ASu8
sOkbezRfGc9FMkUSXaA/qpbPBfyxA2jGbICzqQt7jq7krLAl4VY+lbwJEv82qWtKXo5FDyiEZA4/
bXjbHr7+1oZCKOj//jeOi3jwgEH9q6ukCxN6K3sp0+raTKucLSvLuajv9rrwJlX0LM/+mKQ7wftj
DzIJYrMiZ0ffZhEWLAngq9mYInUBCrA6ujvpcl5snLFElNcW4KNqpi/3zGZNtMX1tV/jkE9SrS47
x3mGvO3Ymx+imx4IMvqu3ygCi573AGCPElasxi9HEQev/HK1MtZNlzRXnWboQEXzLxhvgqQoqnkM
/IxupbHT/0gLPYV/rQBWdFBUyy6/h9YrHNaAOFR6E1zYizT6HG5/ULZFG138bICQLIDOo2RR2iZQ
gE1G0ZXM9CxutlzJTJD6vmZSn83WKiLmiEtvrbrGsZTWA2/X7C0GOR7HPXfFcmEepoZ22BAjb9Jh
QLjPzGCd1xAEh/X5yGmd4w1iFwl+bz+sCKhsbIeE/THkHexC2l/OEHOLflS8aF5Xhdyoz6YSYp85
7GEzySud9XZLfLt64UdgWYg7/XNNLjXvrwM8Str/XhNu+ax7jit/xji+d/WL7avXCtog4s8Aoo3m
s9VLLm7AReR53WyeQaAl///o3YTvtWkic0QOr/MwagG4WvM6bFcc/G0p6hIe4cyTNFvHapjUnWUi
xLQw/kZoSXwdOayO64mLAoVcfdl8ArLxYBjzIWoaN6EQ4aIMZXC/glk0RUKBo3LgtVMxd+n0dAjQ
2NiufNb14kaSpVq2NZefcCIEjyXhSjJW5PPWS4qgx3Ho+nxFMtB5cQ6m98XfGGkBsdRdLfrDmioH
V9XrDC22KuMQ7f4zPDlswPufAKKHlsgqJpeUG9ljK8mdD0HhwiVYGbzXpQcF33cfs1wQUMWT3NyZ
Wu2E/2X7PMfAoRiGRwSej9sNoHJd911Ec5VbQM8sKvNihvIb4wn5koETcVO7Z9I3TM9LAKc4OhAM
S2o1RzrRNSOzdnBzFp7va6bdMIVdx8w7A7+MMORsAuf1WejZj4UlT5Nloe6706Lw3OokdQZfr4nj
kZ8OeP2qyzruv++WFT/xlRYfY1ZAFM201doQPLtUvwNkV+24qRYs9pMjF/D9avFprOkjUV4QDDdT
Dt74OwTLpdV1oIIZ1entnLLpxbeh1CWsL7+pmpE5NIOSQfe+sdd6bYXKQfUf6IyW3g3ZdE6p7Js+
U/T1D5fFEdvVB06anKGgItIhm9y02qNI5Aq0g4unYop2KfK6wf5z36oxBFATBD6vPOpW7z9c6hem
0QMm/6BFGlmwZ57pAH3aM2J/XLZLPHwQDnkPBgZ9dFidLgNWoH5h+ob0yQkGXsS7RRp8ZemZScio
i8c8HHlUNWRe7yaIclCSsri3xUYcClsguNvLl3EIpxWHVqDDmx9wtG0AYSH+mKX0CLpYyueYHdke
CMwa8z+Egso9g9Xu2ysloz3l5TJOcMUcuF8dacOuYMRO63IB+LmMLaYM0DLRk3Gr8IPzupZE7PxC
FA963HOK1ZiUtBzrgEyJAUVJ4ajgvht5lE2JxeTIzIonK3u53nPHrX56L1SmnrBvHtNe1L5H3uas
JfqUKYq6Cf/5xplR9PyT4WS1TT6YTdjeYRb7gPm0cxvt9drIvtto6qeWJ+dcrqtuVIhHITCN6mG/
iQs1YL7zMsQiWBIqaT2gSiplVMgsFB6YSRUG7mFDwGqoEsJVYRa5CHIvtnGe28GDSZB0DIgXGay9
t2mqB0c8+YCXWOCSjyfQDo4H1QYzb8D4ygBUBEcVsCdkysjNRNpsZ29FqCxPUsT7qIBc3s8fp7sM
qFvcCD1MoBx8FA9A2D01WrRisCjxX8g9PqJ+XKfcMVgUZ09zhSBUyIschuRJ2E4xIKq01obcBbND
31eui7ToW0yQRsHShz4hEe144+ZteHJoA4AWmQlsXeazTpyMeejA39TGFXxy7gOJJ1s0C68XGkVK
1NKgO5aqG2LviZMyCWtO9+bgb36geK7PV+fdRzuXnyggNuB2tJIGpuGCnZdjIwX+5tHvnE4jfAP7
TxZj7cMsN/puP7ktrSWmxNmrlVf4XLJWo/LxpCBlE9sWFDP6CU5aS6HSk78p8ch9ROxEafMuVHPE
qShQNaSd5IZ7qUeiIpfa0JMtMpV7gjcDrFB8nYecUrBt2cuZILZgAgA6SeT+fv91rk+azblt2sW2
Bq3PCKY714qI/6lTyyaObrZAMKAP9y/oMqiVF9BN5XPIlsmzsnwrAFi/N0rPAMV0DeNY5/I+mByk
TrAm1Y9knWulO/RiYZh4cP5UMrNwFMt7YCAzTEdRx1hgG45iCAhYVu+pCbMMk8HfrE7Uv7nL8lxl
2abGFqNapaNuyX8uo4u+L3bww3yuTaNyLMlol91G259SQ9RhHGDn1Uh+XjHqAEcE99XrS/Wx0Qab
9vwrpvWgBrgN7fgMXTPip10WaMSKEfqzcZWPFYAbfl/nLvQRVA1JDfbap8/r6EShQO/C3cVQeKvs
xkL05KXUQOLa+hv82E6xvfxMZx9hgjQ4QUzc9VyLbP2qG1ChOTVDPC0X6nbc51ZShYH6H8MGga9p
gcTiLodwlxiwjUmmFMHvOsdaVOdcx1NakE5jZ3V7qpSNT1IxzKZXG3W4AqLZpMT97x/9s5JtKNW4
LYHRgGtQY+Eoyu5mn0yoiVsBynhfh3uzw/Gzwza9UmU7W14GimnQzVMGn8NwLrXj7mViqT4geXJL
jCAo8mUtwogd8G2ZoRJHvyKlkWHx+veluwSqaHtGskwVsjvMr6b27UN97Le3HgGc8xhXoeJgMN2M
+HzR/CvgT3j7kXy72F1tbVniGljrPPQT4fVDjZD16R1GVXQp2PAUUPqI7IpH1AYIfhd9wj7Otgof
HOeb475t7fH61EjiwkrtAEMbU9atckGxh8DiVyQoL5m3MeHdzfSlQWZWt4zUJeZX5oFGFhpBGxLD
p7oVHnuwebbdmjLRS9lWxbTFqkxVnVrV6eDeYV3qxm3vUJSejY94gWsEGjf/3u/K2MyMjORwzp4u
waPRvjQcwUZgQwZJcAtPAFg6g+iwn6cjnLnktk5JVJOZ7WXvHHukRe3QdEan/0Ni6a5NJndCaHRk
OLSaYh4L8PbMPbtDeNXjb/oGLwEOB68BdIIThv3bWhCWBy9ImV6wo/x8c4goKiEhqEVv1tGpHPnP
aG+dgom9OQvBrBTvebjdWbs30p3ihAVmbWtTwbpmC8Gk3qDGR3Ux47EofQBaN26ZIr4Bcm3f/fFI
z7TJa8aN2A2McZXhYDmD3JXKvudAEnxE3rs+ISu4JzN1I1TjfcyWVEoVe2So/Peb+6KSv78PXdmk
t1TVXy09UlS6oDyHl4WzVkSfAMC5DIRYbb1n/7o6WYXRfjlr/inszNNTdSOekEDrnDz82emyI0ai
EcGs33LzT1Au7R/nScyCHw8BmKi+sCEiq4Z+gtSsDxmvotb7d3N6fUWkvOuHFl1bsZFinR2ikDiM
IrF66ENZisrgV8Drce4jP1sUU/9tBDt0i0+crF3FNqTR6XHIphQ7ad64/Df6j8KcZlU+4AKYKLJ0
w5upVcWlnmJb3NsEVbST9n1IeptuW4Jwimswotaqb6244BE+gSQRSy/HqN6ff70LV4/CKx40awxf
njf4w6ZGesWKrNE7pBTkI2kTvenDDy41aIVk9K8qxorILpq84/l1yRR+B55/sjQ4dvESaMSX9j9t
UQsg/yeOwN1v8Gx1gvvE4JIXfJNykhA/2RmMUi0qmFol0g0HxmO1l/HSkq+3wKuJK1S8PJvpCIzX
K6sqMR8j3+b17mvALm+pgqQRHXuiHe06RBJhNOdAjIpIwB9WYa6NHgBs/s/EeArULzUr5FQHg4no
A7IO9U7rYJZ5D5L4WJ1eHZRWIiZkLaeARB4NdqfWDqMcR50GUjMagYJQX7s9bOHq7oYBRi+eoPS2
9YEw2ytn8L+19+oX376oXpZEAb+gtuHJ7Wch/OnNlKUwAePAVF8odjWfE4c7KfDdNI4zO8D8HcdD
hkEHMk9dGIR251ypfhKhxal9Q4fvydM+OBTwdE99i9zqc144vVwziylUtz/eXTv+YjRpSp74o82P
TAXq/O0sbJ+bFxR/Rmp9oifFm1JIx5M0SS6IGbSkX0NZlCV6tsYklTsIHe8MaOXkf2B5gDwCjg3n
CIj6FcYn2hq1dmUpNFHnM3oDocQCSlpNsszVtPKZPZb9994LJ2/U24HGpJSGWjenfvDK4Odzzsx1
TjlmWND2MUiyfNLFEdFijFq/RK+ZK2fwimkFr5FPWXDRRYv7AB/v/SBYe+n74wbwq6chbkcBRDRi
crLkErRwqo6197LY02e6s6AuRfMGiMTQZaRGKZjx2SOnqhv6DzTECT7ad3jJ7OMuog9lnxxCwDHJ
Beo2/z2lg4eTwFfsDdXbP8ylR5ILv52WfjaKy5eCg+wu4TM9YotkabxPwa5DcWRlAcgaa9oJqB59
Fhcxq8z7LnsZzvlxk6/3zaCkyC9z0+IDaURjylj4K/p/rqegCxStnKdQNAa7nWDftR1nkgAQAqEs
aKnSZx/Te2eboVgaIch9AVea9wzX5TxYr6EJ9eY0bJU7zD/7ybFnIttMlffEOSIuqaTOVB5tfnRe
B3adyyULXWMdtc9mAVMOaC7lcedbIUd7w2dMSZ06o1xnZC7Zy3XapBM/revoEyWpznvs6uKVVE9P
BL7dxk5JlrA7NB8TUK1/W71NOgez/WwcEJheqk48uF8ck5MNEiJk5QC1HtEYrPi1ARW+nPjcayXY
iXuu0ChOAsWM5Al3jLMiBuYUa00Pac8VEseSdGIfeI0B/J7WgUIve7HNgXZH2ErfiL1hrFmH0JA5
7d0rCTgcc2c9lzvMus2MBIOnZmx+5zd0QMNkDvxyREGyRjPUACbKtEodUdcXpaJsIoqTNsRKueHi
RqOAhURtmVcSdXD5urU7O0GB4os5hq+2AiztYSQJ/Fzul4fB42YWMY6p/kUCRINCs4kJbTE1pgjO
Efvl7gnEuVLglhlaQUWV51Sz7IoYpQJgDYVQFvkmYwkiEm2YNqJRIuTW4isb1eEhMwEYo6g8Hzk8
INUOes/xc2lA78r5mlSO7744ZGowufY8R62FisP+sK9PhDNd54Xp7f8vDS8HAwXNFkC129/duVTL
DY/x0xcxq/JaSH7+8Egt5qeoCpx4AXRxD9U55TO88sWQM1l7a+rLx1hDNmnbtOqooxFEfoTFlCLv
ixx6nHSGVaAEV+6mhYNEdmEWZgwMvFuJsVnZ0C2SkBBATqVtpjTV5I2HPrK/6iQTenRkcWw9+1QL
ihOhdbsQB550vOdhcuzDZjH97DpG9lgwJcBAEzuNfcBrOqneNquHXCHZ2/mdQDso5deLHK7XZVE0
ZgmP6GQT3XniTYTuBkxf4c7P8C01WAHZVVwyE7c92HvX7Upx1Yzuqx6nW9OoDbAU+5UcSDDL+qNt
6rCi65nDuwUyfkUFOA3p/6stc0l3VTVmu/2orOa+C989g0zW0OUDV+a10DrKhnxBM9hebvxfHX57
Evehg8elbMtodvCLgcT9TlHRQGjC+S/v6KOPGx+0HPsC+l+fbuXosXXqPXLvUs4DvzlUWO18dAIe
2jK4Zl0cOf/4NIoRbEa5mGWDbkrKbKKH9uiM2M+tZ66ZU5d+RSRcXy5oWyjl8ShttbnTjAfwvRHD
+SCWjIU4jL4nYE2Mvaq7xDPRKK/XHGpAmYhz16dfI/AJRT4YozWKtrUX2s6SsF+08m/d10bK7RhS
DoFgE0WgvU25VVEkKxUN5spQJfPwteBBbElmWcUmrTiQUWuKO0Hhkipt6ItoAYM8m25KUjviPZZT
i97XgzmcEWiWfPvu1Mc8u+EQGxJxvoDz6UzOhq2prCrrM+jOU+Wn/MJG+UHjlcqrhA+SGYw9M0+1
facevgh5okHJjrFmK4WjJh8ELtIFzgkGa3y3P0PwXM/QRRMopKiJmUTuY58XVZ3Bp95uiNX1+kmO
yMMyzs+3LE2WKhRycpM3ZCxqUF/wF3j+JjuhJo/h/Lk8InsyZ2vHfXW9TnCt4MRBFs74zLKulE1r
PnQ1XrlXp4UCMYCCRX7Tk+TSHC38gsYHfA86N0EztEQNcX/hYtYNuHETAsyPtxZggseTesfX4q7c
h0C5+Gi1Gjg7A0+7oRAT0fWNx67Sa+9iXyzA5C9tMTYYRvMHlOJ4W395YTFiJogISN6svMZDwKd0
R06YALcCI/oqXnUWwU+tKnnFEa6AVGhyKTZJaONm/HJdKjYAz2Ya5EDsviIMaV1pAdsy/YhxUit+
pUg+l2I+Q8XlT6tMsmC3uK5qaFiplLCTZIkDKJj4/yKHLc1ecaPwaixy4dfFqBa4qZQky3AmVXtT
DL2lUdZ9/f4GU87db77ieVXUNjFTDNpACtXFN3RZZZwNHukQ/g1ajWXFt1TIJmvIHLWXYJRkOak8
yuld1om0WlGziN1uMG0mkv1uEdHJzKRqOwnmQjks/3GEBqt+7EbkXTNUbNexI0kkvc0qui46su4h
cbS2etDOxuo+WPyh+FD2wwdKOe/XRT6HyPe71SPyG2iPIo/dSD/dkYeS3FH/n4Kt714hVzJKlpBN
MogB0+H/GykbOxQQ0v5M84FH2Nyfr+EAaAsRsNXW0TWhCFQYvV8K3MFPaL00goR+MbIZYGEiPs5F
TvKOYpV7LRbLwWXP61Qsq+SAEFoTXsZzlhTxfrTE/sGbQTLyja9I6hlIFKYk6dsCtgK8VnxjR5fG
OYmHJP1q+cBCu2pk2popeKRmHzbw98Kt4byeRyAea/nlwH3ALqB4ktEKg29Q1DSBPapffPuJW+lq
tpEC+AxgQoX8L7ZX8S2FxjytEborFY/gdfA1T8n/VLAjunCzI0hAd1C6Fw3hrWw1lzwPJu9XWlUZ
LFiMgDB1s/ZZZkDy4FoB8iC5zSdSJ/o45fUk18q6pQls2PtGyZH2OGZuyYkz8p+a1Q0y5FZASEP1
E8zCAfV+ba6N3A2Jt4ydPwUK0V0vvKwESxJedFFyK6XlWG4FK1vTo0RXr0I+areB9Cl8WDUQr6de
jpaJo9GpoBI9vB2Snv9jjGqGfPOD+GregDIgciMmlF+OhDTrjTYrAhX8WQBEtLjePe3BO2vF4i0v
dMOhZLHyx0Y5w7G7CaZE/AtBYPH80kVeetysV8oujzHOzIokcgb5NygHKUzZbP8/8iQgpZb6fFeW
6hJNNd/O6Amyakww1us1Cu+6hHg9DrDjEgdiGBIt7ZDHAC6usqnKQgBFXjGI+hoQKo1UnmPv0Dar
TPRwzJ/GK9BwNdhgdVkn50qJmdvwIlWw503JQww7gFocgi51hMjSa1nxiobTQtbUxjGqNh+6PmvY
2e2rvxsKyrmE5bRlKr6ktYTz/722FHAZiBTVgzUYDOmcRLETjbTdKLpBnbBrQP9KDXHX8cNfZfdq
32TATTl9UyFncfwJX65d9uczvpOtwwJn2TSOumw0s1sqUQbxUJb8XhJny78UEs7WVW+7B/N1Ik8S
DEFmpXnl2CaIKgvyi6e9oe+agV13WI5gULvf1rKBJx27YBbu+SS9ba1kwLSuSr+7Tdv6mlXy7DVL
paRLUhvbBBcqBi3sO9Y4CQpabNE73kgLUUUGN/51ziJnlQRDnP5pXpDBf+iDhG+0nw96o/9hIZd/
DMiLXhM3dygzkk622xcE1zqb4FATK5ZG833XQYWB0Oe29W4XjcIwBACEDIScPZS6VVD+F/sLZtHH
DYjCBQuTDKYBF0UE9dB/8/DrpYvt2u2rqINN5F+2smWJLpigvK+Df+QPZ4DcNfEdG8KyZKDYE3yy
Se0f8bDlL5MppK4YWk+4nENeCGmVBH94Nb0ryTUib6olXTtp+Ja+UJuFcIqtAzgGpVVdrGV/sCSd
O+34ALmHe1GKUFs+SYZAuvF7ZiG5x94xc5PaZ5YMhYioW5CxRJnjSI4bWDR1FQF++chnk58bZveh
A0yoBgZEfnwHnEDnq5Q8vbe/xVwQY/uuEIxDJ4TGH/pMnRQBHOJj4FEADrnIV48piCIhmu1hIxlA
6f2kgvs6QEr9yp/93j3vwxy3Jn2hNlyhEu7W7uoD/7F//ueA8GvQcWAl81GVMYNH/577U1gYAbNf
FAt+4NwvEOUCPOF5wmhKIr4VnQyK9foWWGlEF5fUiyWgBIuvEZ5H22uCytgUYzgPbqoMgXtzqb12
3h0ozS/zSh259+GYo0xjGWjSZA5UTYDJbNqDgNNHIDh8Pl3D0wPPCRWHwVX58NrkN/Ip7uaoAxKx
mSo8s6cBnrdOa0uwVUXEej4pOgv7staBYGrTluRpebe59pxHq/w+dIWd54NSogfTNYeHjLuneHIj
11/+fCDxjcoCf00fIxqhWnIj569ZW0Sv5zCXUtgQ9KSjcJHgFHKlfb7dIt9Rl6WQaWlJwL02Mrph
jJh8xrsA6WMxlFKJe/JIUljvva4rgNWHVgNsDAqd/upPThUBlgEQFXC57InGVh7UcUWs/dtLGIMN
Z8Qvt7JehdKHoabhmgB6+RIVt+kZjy8MKDtjxNI9IOlSWkm3ZIY5klfGsU4+kd1yKkb4zURgx1iK
uBXRSkGtGpRwzZKIWYUTYirlCVpl323qG5mqVpjqZXSz08qTqcbPD+xOwQrEc4ehVFtPL3fBNKEc
4TJNugFOc2MhUFQeOk5qtavGrV4nPOHAKYnXZC4WoP9lJ/NpFNsbW8DVgw5Bo8j1EvlpkxSDWbIi
ZNZ3sfYJCgVqLxIbSZbrCRF8tnmmLfHdK6D1WefG8LoLx34NEu3qVYS4a7WsP1jivCJlD9nbGq4H
+/Hg7mJ1hbMgXo2A3iCkMPSTh6z/yVngnpW3TKKB9UpE9EYUKLYrY6OVcF9hcbH6HGOqeyt8qkWd
wH0iltP8xf5ZT02VOQamQjmE3helL0hUIryAQ05zJvhTX/yRyDP4e6bufianajU0tbJKoNNKKunH
+gZ1YhzJjvxodEBhTUSbriNDl00mso0og8ttZFzi+hkPhCCqhbNkU4RT25Ds0/hgEvkkek02EPHY
JgJzDE9gI/LzjavmKTi3qpsT+KReyuPzvj+AoX7XzjBIivtx3djQcOVV1r1cY5MIoWyBr38Jjw7W
YARYIbzpnHGOCDO8UejMeBr9/uVbZC+2j1P8BEE/DuCEGgyOF12kaJmYzLgGMh9Ouxcaqu/1HQaD
SbE7QnXIPpr4xcVc4RozuaLYiDSWeLZwei2up2Bn26oNLnXbFA+FpHr6MtJMlQZD6NNGtLYT7xB+
MElWarp+Jvg8cbh+LMgwFe2lKtqJXQXSKoQL82Z2VF10hw/Tv/wiRy/g4uscaRSQnEkdWokPyvHt
SAAJzjbuIek2Q9UhKdSQyKvB37r8q1T9Jyxz3cMau9vsOPS/OGU9QSMMVxlG50RZlx0Dcl5Kjnqi
L7BqSfI6VaNW7WQPYK0K29GL5w2VO5XNxPvlWXYkTF1y5UlbnwW9E600OpGxc3Wh6zpuvwDA+r+a
hXZ3UdBe5kG/6PEJUsGLL3OZBJgBpLOJsbEhqzAFYUa8+WHxr12+eT5oJnTP2MuMf07EP1EbWcjG
x47VZFYLZhCt8dcw61zypfIaB1xeq+Ouj9+i4AjuZeNZD0qJPq7yKx+Lr1p7vTFFbFM9CaLFDJpH
+IRCVr2kNsLbCsJVDsVnoYRGWdBn1qBjwD1Sa+7Q15/k3e7XveQ9SA3ebfVsIo8ZjqpJKkrbahdP
1I/ndxaPFaWesDtw019fH8fk1l9iRd0rBHYwnaGU5sMTJ1ndJVcob8iNpsa62AkZhCRIuNYv7FZR
Qyt51WOHEo6m3SthrYRBORpn+42viHpF44b9DBM+mOyiL+6bT9d3Ap0/OnC312Y19rGAQ2mQuuJ2
aaAfF0AgO9ogcoAkbPXUNpM7RjqgSUeANtr+yWOHlqE73rQ4lrtu0Gr2omYQMfkR6o7zovdJ9znZ
4gJpzJQAfvPP9NS7CFDrlUmxwkOExaznSpMc2+IPCMhI4kY6yMfiEJNZN+3RZEiVxUd/S6lTcr9I
1IAgT+FwpM9rRQqA0wDHwIjVai/9XoLLqNASdf5BzZM1S6+nttdn/D8NNXvOTnwfE3YNfj4vqHI8
dlbOYl3NOhBZWER1rjkaQX/kP+VO+YkOmFpPb/EbXtC8xduxN6xXyCsuxcH9ZHSH/gIJRUSOIDrK
1QJVvBqU2skCCCjGuWW67kA/CCz8+bqyiSYoTplVsSt4IXPmTLmzwHAPcvDK0w6XHJTnsIVBob5Q
TWXZqjlF7M2yjY1nuAGkfjR44C4Pk9qXUjfTEkSulb4fO+iRLIOtzdcKkDKFhpmP4hLNCEDQnb/t
TSlWcMyj1YIpuBlewIc/gDB3HXamgnT3vF/bdwRhroXq4+WRQUnt+x1mk6ruoj8g8cK6yr9azxk1
D+7LqHAi+HkijzVTtkVOdE0NqpBJMOMRRihgipQWnuvThPjCeQPr9rdW/loHFBzc9VckpEfp/8vc
D6E/Iuvl7u3PA+xUGlcHkFYabaEHjAa49/xdpmBLN0VlUt593UUedIKO1CV4i30IANfjbjPHRqPD
qXr68WxXesr4iswzxo2NrnSy+EBW/R+HOR8dvcgroM1HJTjCfMjUil7/q4UM+q6ovCzUwp4oA0xq
SzE32lVu0EB+oVEuzPwp8gc5j9mBPSo83yxSn6AfX75KRRVOS6MHGrmWefQfd7oI4o15WgM/0VaM
+UD8krK9LCblWZLujdTV67k73oZdd71DCj78+/2oepnBF72YJYJ+oLQbpHYvlj2WdTX62kzZ2PJQ
Ms1ii9AMSazcNEkYZghiVsfI6D5KvyXcQQMvaeUK8j4nYHtMK/ueppKMhoUJlzHcQSppQfKWWofH
yRTeW9Kd5ryH/1te9pK218gGPSjkyDkP3tUgwTefzspuszkEs7E+KbefXq6Xu4vVNrod09Yc0H4A
XVmnQ8piutvra4WNs4PpUbQgllsaFd3g0qqSkyKI8H6AZrfGdQvd4EEDnfLrLvt7QId+lx7rLoZU
WsSKRvXaxbeKxAhZkVJ28L0hxgC+DvjP1Q/yEU+qiCOm2flmpSzG7paM/nXZyw67waj2kJhArVDz
1/ode4SpMGoD8ofC5/RtFVnTDd1kp5oWlPYJ5rYft8fNOm1CWjgr+/xDUYCv9emHV6OibsR7mRF0
sktc4FJ8TKVuHISaYyEkp4yYnQG5ZXjrFZ0G96r1gpko7PBB1xZOlwZGDuNmxGUg9+aBl4w5cGmW
7/iLw6uApT//nQTxdtf7NCzYQVR4Np5pCuPerNACjBV44IBh7faSLzybLD6eH1XPFkf4ZHsAC74a
q/l2E79I1xaG4qPJOU1Iu9xgDvnd9jP7k+nsYT0wyYDZzL6zr9q3OJ2thMrPsKBaJCjO4+pC9eFF
YFS2ebOGNcI7kNRNtZf4zYmXoiS58dq3MNEwqAkSL8PooGk8xxTAXRpr0KGIAT4F9UWcYrTT6F5B
NheWG8//kGgXDJV09eCS3kZfWd62GVjyoVVWawzS/Hz4ScvUTxcUS7iiYBMi/QdAXmtaDU9CTb88
pqGvelsNo2qdxBvG3YqQb6kGJ/+w1Z39NItjrR6dyPV8D1eFcycbnXaFJ7SmSOywcj1meGGZ+iVE
yjtoQnC6ZHV/xzMWr+7F+tSEBJwIh6z6oEaJJyNLpQlTfY+3zq+Ok8dY4PRDx0CbXVBKeuTV23+2
hdMcOrEPZ/QAyFlH/E2kI9v8U0w9pnfjoxqLBOShmhVRtakV2zqHA2BTlTuKj+VlRMsObPMnSeW/
mHmW7rrqjEN1L+rgDUTg7PrtLi1Lve6QD4/AQaGsHqZ7Y19SQLA+czfL7DaKS5KNuKawtWB1Pw7T
quVBX3tNkHsTcNqTwG+TN+UeSsw8loNTivhzpnK34a+ORNqvYdjo7PLgub8l0Tf5Zn+UMTvB6aZI
BQ+ltwjlsOjej7BZy+yaXXeh0nxQ/gGoVLzHbi1x396uL/YZ9IfbcpjE4zPrPMwpe0FrLfdIdG0A
C+fqC62zH6sKJEfiZtoWogg2sRH1oMhprL4NjnaS/gyR5dc/pLYCq8Za9wEPpRaKIrJhe+va8raN
1k39ppV6ZgsbcZsRy2qU0IlvNXNYZQPHK0Cs3xUcOG+a4q9528zxK/5FE7oz/HvfrlYtN6w6QDNY
HGIxzkA1olmOcGjqZwNer+3/KbgR1A7iY7kusgY9ZnYh4DnaO8FyWwcsAODwHWd0izuInish0XKa
xov0xbmkWyfMzRuZiJEz67XgHnUyvoEdqHZSiAb8Js4TaqkRdR0KUE/gVe4Zz9cE9NDyr1gKtL5e
xuwxVuD9K2hswSa52r3erhFu7PXmCrnB2x0enJxA+Xat9+Dgc5GlpMStnINPDyv0oCb3C3Edw47Y
nQs/7wZ+BkqzdA44Xq3kzlQhvtJJR0QUvYtYQDzHQWuq0GLgWnRS7DcOQBusk5+8qt4xW7/YKGu8
QCxWsXovOicfkUJ+35NatQPDqEe1WbANaaMvMSTOJ7ZU0oOo9iEd26Wbr/ZuP70oZLF05/YWfFji
fHKOvftReoM4XuVFYSpTM6S27TexreqXi2P0W1yy07e7t2uxi6R4OwJweoCH1ftAGXAKxBcX4Wru
HUWi6WG/BkP7JX+cRMVRKXWiweq6aQQWZbkcQqMk4WJhOWSeS/nJnsJAdDMvIVIY51WlHmX317bQ
R0vheGTAtlRW3go3HQGBMXTPbO8fVbMzKid5ixDARtEOS/LODd+8arnZ8q/D8SAdI1Lg/b/l24BA
tHjS+k8NnL1TnUSTHE2dK7fEqfV5jPfN64BXJTLHXshdp8nArFEXEIk+THLaQSrzIKX75OMcXlt4
nLnyXIixH8SNTmI/4I0OlfHM3jRlriwHSoGrze6gugrFpu9OqRyQKRjntsn89r5a3wxXmmsz/pty
GAYnvbJA7wDx3w7pDsgpedCObVfKk0n1AHWLplG4dwTxZeLng4xOSz+0OytgzEvnd9IV9pb7z3on
qk1ni0iKaool3eJv1a6hs1Fn6gJmjgeKA/9yEsAwtSvn3OwbOcpvLnOvyFMyffrj48qWAthuaT17
xYwTnr1Hh8yJZ3cxuS9Wqa+8y2oQ/yLzX52rRNd8WYLkyeE9CsAT5U/GCev7aqZo1oieyZoidpA8
7K2a1j5h9DeUK9EsUywhZfQ148dyhNxcpsE9YN6iPI8Ra18MShcxX9rcHObBLHn169/iGbh98YuO
pE8bFZVLpTq7iHmVJoVM9uDfaQJpB7+f4a3p59i3oHKGdlxXC8JC3n0tm98d0HAlvcmUhcsVW/wK
lEdUu8ld1svo69NWimTunbe2PkxYVg41j714zqO3iTPQt/wUgqhmiqVyTHvJhIcB5DSmHm3AIANU
bJNd/TqQ+1R8EPOwNikI6eHfNtEdWJlVE/6SBtkXrVgDjpBk2koJwBLDI8Yloqjn9yP1kNamBdc0
F5g0xEwJqqETCpO3bjL2GM4E0Rd2A8lmLLCXO2AkdJQYvRg/HFnSC4Xa9BDibGvZj34nlygCI/OW
xzOHFXYPGU41GXmZtWHBHCBJs5qDmSvZwqSrRbCZfZwi/KblDMNothAv3QWXYIg4Q104rHVjAO8p
5LohPr3uNtAWy52RA+f112SPdRM+VwvXEGY7JRWcsUmBXLtPjfn/pNQBmAhZQCXeFY3xkM9FhqV7
9pr8LaE2gyvSi6klsGSFCVBtU/N0m/+SoT3SBWRv+au6l+buaS5mEavYktFmQVRx+7y0RAtcSnLp
uiS4MR4Kg5BYUz+ti7xSX1qGE/6cHnq+WSLTKqfXczP7XA+5pzpBn5nnpJ/Cbnk3poC0caiD9+PE
fVVtIkv4Kb6CvVkyVxXmb0wxs9n1BTrlJ+6w/CkVrO8DwYGytOKPcyxgHLXkyTk+Lsk0UdvgmzYN
6c6vjxOYtZyxervYstg6nI/l1rZm686vQz2T/Sv5EUgZ/KIwcEF9uzldtdfAN1U/LGQS1hCU2QIT
AinH2lGXgslPvsIv+FjSxEelfREkZWHOgrO016fyI3YdTN2oCEkzCWasZjAlE68/7WfYyp8P783i
5glWCL5ckV7WLCQVDRmnvV1KMU5U73ybKOzZuIJHqQdz+2a3KYUX57sgd0FJwPKOsmdbfMgIXsJS
i+Cq7gLjOu+BJiiB4ciFqiHxrNlTt6h+PwfgnnI2CsqYBPleMXvGyuK9/AeL3i/DTJN5Rukazyeo
+hfr3uhhSrF/kVv4HPoBkkEwYAz2z2WcSDpGONkypa6RxAkEPnk7hsCneTUbIjmpEymnuIcDPTgj
r+z2PlNWfdunHi1b5aTgDtK7P6ErNRpPx0hAOrAazlhhhwKZKiijVczhAa6ETqFsfW8TLDI2lh8/
odl1UC5UvlLW1OD95MO9Q2tf2FCOqtN9esZWMYvDBYSRzCJ2cnTNjzYBpQoqxd0NB6XqM42lU9rd
jaNfjZAwpaShC/LPRl8D/3bG3Z3Har2X/Z9VIwezXf7a4y28vGhA8paHJh3cMlJD+ixeRnzne5w4
QK0wafKtiuY+Sa4d8qM/RRO1Ium0r1xHrx4lJKKfVxrQ5fuMijq0Xj4YJQODOeWgRJs7z+/lKLD2
Qzal0+EckLrJhrGy3azf/pg65XK2MDQD9m387LGIJLoKkmDIEVRNSXFB5C1cDOvRo79hE57z6gcn
MTCV7h9sKm8m3zaZLAeabqkaKG77SG/3cxHj1wfktkj3TdNEvuGTq5EiLSqo9oddgnHGKBHDXvLU
/Ihi4Rc7OZQcdraAi8XUvZvIfA8/tBexjCLxbb098SSp/ZcUqwlumUw6L+EdtEZoX3REZv8X20Ox
nf2p+vquDWEzDct9W9/vjphtHOXwy0VIAKJMdyOrmw4IyS8ak2zq4WGtVlyQhKF7FIs7FO39vTKQ
VtZFDHGy58nU3MmfQJZYcuUROPyZD7J9eHxpKKffcUZ8K96lyXE9iT2v0hGT9/f5t+UGGHwKUdco
xYnHCzkn0r1jEVmvC1gqJ+RDU4j/vInF62cjXXpneBne+Met3nvSLPrsTGwGOrUkDdhrI3LsViF2
cbj+pYLVYRoZ0uK5IBkPk85tHRjpzRFgKpJlc673W32L3QvNCBsvRz9tF9oy1OxugvRXFVHVbHfR
A4mh9RBTjdOWOojxjYH69+zt68wxSvcCsjwCrF/MI7c8HaVMG48RL1WOHvErStcByX2RXFBaUXxk
vmbYj7DZCNc2SdvATIlQdAUj+QHTVu/6HIpbPIJFtgpC8obuAYHo6ed1b1gc1mN05RjaVJZD1eLe
pnb/4JElaW97jr2/7AKft2TjECoMkiygWHDBJLLZzMDjF6BQQvBfQqrOTUPO51KiY3PHoGuNPBvf
JxJIgN6cG7AbNm1RP2+7Dgnl7jcBQ+VJkcXb6BXpAxUdXgMrHa7p6cJhDdwtUyk+XfB3QLLEy0Ct
RPgsjTvfGlrDh2aeu7pUZscH/hsHGuYplMqt3WUyFVI3evxfh8eJHXq/7rrgyaz/Y5Uu6HeHTug/
mOZsvUt99ScHu5PddLCk3KJ06ht/+Td+XTHpI85gLJc74MdEnF7mSJcUeHeNoksDnP8hvARXvKat
nq9PALuB9BG3yrYm6Ro8+761ljdeOY1jsN4TESXjv6GM+udWBhPU5eZIBPMb3JyXixcp1FtnA8IL
W/Er2kdcEQM7+QxNY5M5ldPKi/EqArQ+McX4TjM+P66O1beY4I9lrywvtqKQ/dHf7aYhTNIrWrOb
nvp8uDJeqB/LLVKL1kZ7GVpPO5d5J6QVFteh/t6BFRL8o81VDnJtUuPrtPeDwA+2wbUrDCvh1t5i
GPwg2kmyc8dZ7s/dC91rT9kUQHj9WE0eTitZ1KbW2IptY3syOlgO3drwvFmVxmczKYDZ+DJs4+L1
f5ztQxa+fO5jIHSa1J1a0ADTp1REnNe95TX3Wq+Kt/AZBOLxjchS/RbITclf3bJrxijyoI26y9Io
WuaVI85U6488Z7HPF6iWRUjmKRR4jwqaexWdHzK1sPO9qqkqWFlSpbve1hQOBJgILsCaBNrUF2uO
bG2PRmDcty7hQdr7mkWB6p6n1NzN/1hhp9b1iSK9qiZ8qf4x1cEiVvCiSWrbCgJHWV4bC0E2lG/q
jVXojfNRXOcFgvVVED8rZNAYPZXoExDCPXuy3h1IDh74hJAE91r5I1opWx0DlPrDaOwb4avn5BN3
5znO2dFcJN0JLlMnqWAfYzsZSZE5oRE9729sHwaDwZvboz7V5JP6zRfLdDd2/a44l8lyNUqSxuEC
nxurw18e3zPJx7y/8F+79zhNDHCsiRbPdCoYlTxKjUC654DEGH1oUSGWWq7nKekyuvqn7mBm0Ebc
mu8GVSUpCbsP+0GDglftNLoOX8jzHDy1UKeaRvLGDKzaH92NGyiqWtyK7Vh5ZXG1vv67AhyU4xKY
iTSG70XgiT8kvWG6+CWJFmbG5LXid/x28jRl6YvNxbdeFoDwL8JPk4RiltY8DK/29MQLLMoVO+30
u6sy7oMy/89O6/LGwzuCmdr7SXtp3QtY292oIhSSsHAp0P75BIrVvj6aPRLYVQsbcJWWU8JM4fEB
aQcTXqRd/AUUTXBGfhK7icczRNPCtBmAEbTG+FXBwlgnBb/YRVDaLmZ0LENMi8R8cJ6ygu4fXJZj
701QoXhG5EN/FiS9KDl0M767zdhVlTxsoxChYD1y8toIZyRKRn28MHEk8ScJ/utQNvitRGwy51Gn
JBRAxgIATebJviXng4PF9rVOvmnb2a7W3VccUMs3QCRPuXh5dKyg+QTOnp6vVk3vAvcqkfWIIUnV
E4GPw1EZM/g1bv4FZh7Yhs/XS+F+Z36LuRNK26WKZRS0geXPzl80DYlv9wrvwwEBaLFOREugZ4X6
fZ1tpBqhLi0COFezesvPcQayT9mJBK+FiHkqd8KHqanzFRQ7DoyzPGuyv4aSQk8Kth+EEgXdB6+G
FCcgiZWiSldn1cwwfEFfLZQ0RUTqPte40R8tkiloCx07DVtWKMEyClr8KfbMHJTiD7ko5VgebySz
kLNfkBGAv5xKBIpP6qF43+TNfDYE0wBbNrz4Rj0mke/8/V80lIumQfwEYqe22Fxm1p7dQP33XasT
gL04HALJgtDt7PszbBFsX/NtXuffm5+SWW1fHgGFWowN3os9Lu98c8nLsEEFpZ6hdbJWkS2gvgJe
UMzOxV7rhHQ32Fv9arecZxOm6wYNDkBMvg1egR02wZmrAidMw5r6iJNX6YdkkqeXwK1OkSE4H/rq
tuA9UfpeJKaOdn1QdR9VkFtHqUzjjVCpJyxBUnR4lI47RklObnR1wWe8mAhIIueyEmekTnB4GUs1
mVMqvwphggWI5T2qCwQML1AhY9+5TZPRfTSR7q1WVmqujdLfulRR1gpCCc2EhQDnNBy2wu4akenZ
63AArSGMFEp6AuB1HQZxkshPmJMva3nUndmKDmN5cna0GfiQdZzyE/Siw0O0fJJKYwkexDocyPZv
NAcg+0s6nGvR1iJ4NS4JMvCdOWrXMtiH1nZvMfMcIKeCG94PAJGgWhgkYEHCdUqZXqRIHzFxul5t
sq46vAEBjU9hehc+j4T9YfoGMh1JsvltQTp1+naSwhDRhDSwpQUydA5SHlPGi4+Gxw510skhsFkA
rM6+WL35ztS10BX5WhRPQM0DSpRyt35NuZoivx5SOqIcDOddsIAlKz9hyEMQn4zP6ArlJSJDYq3+
Wue0nvnbMl1TBusO8xg/s17eFx891bBVpaEX6xKw2Wt4hAwVFpKx7Mq1nMxIiz6Sz4poDVraEM19
S1bZordwZSYkorsKOy4EBG99xtBrIl/dcyBVPMSpTzxf0hELKTWgAq+BeBsfNt0Hqt77vr5o7vBI
zBYZdlDOi7QiqAHYVQ4snvUCMBNYp7va3LYJubzPia+IpdRsn7XB/fG5kNFwixIkQ0EWDt8v1YXq
ltIBgtTel9pCoKNEE9p56PmraolSZZPc+etpifzZyRHLjQ85bK10+Bg/nxaKeNjoI2MvfZQOnd9F
t7XRrWgYfieWVohgG+xWUpPds03csrcfYkNMBmi6niscpfQk6paJ5Er0h5131DkYkguc0jBcf61F
ZMcjEIIrRGchKYvCZjPqLXfwJ+OQXVvZ53IyqC0oVGfSl40/xg57jnb0sysIFUeMGV76z+g36acS
m8vZOC11iMCsiFUftpxInyABLdQHmzJbkIiJIladyAWu5/nz9aadUTU0UR+e7QcdJLfISVN6GVgN
s4kf6ZRGFkajFnT3tddOA09BN8gWsH94yY0jQzy4mMVJYesdrd8+xRWfFHNYJFHwZWJzwArav+Sy
Y2U64qlGf4V3XAt/XhsOFEePNIZEjiI8/rx/Ycb11kAMUIRx6ToEtBWyjAhmV57/zPkkcwgoW1YC
W8f1LFFf//hrCEH6I2OQa0rVgRClxa/1vY5B7iTd8xFDkZay2B6X9h+wRjMpkAwuBmntTuyRba0b
PAuFEGxQ5nd4ilQe9TMCS7oV2yF7XgO5mltmxHRL7PzZDi/3hIS40DRH8p1bqoTzCVyf8OFj0tWh
7mAkL7wGeYnIRo93tXGY3CmcTwajFeFsEOQs1XOofTMsp2TQLZDBtW6kSL616zVKN3+DzbDjVhb5
Nd/2BJ1jILZM3bKtYAyoA9kb7MHZrF7d1NagM64lH7GJbQwv/pCzXO9j1EA2kL/XZ8Dbs/W6ANHN
fvCJWKl2/jzBDQVWCJfSWz0PE1dNrR83PtM7tmZMBsMudBTxhT+axBvF4XlEkUJTo0Dd2m0hpChr
Z2H2dRbCJRjXJ2a8b06P3RbGvkmMmxcmn7ThwILZSqRu3PhHs+pAEWjtnJB4YpUXEnLTVFOLlTAX
VvRFfULEnYaEoiZmsLwgsd7sHNpBMWvG+eknD4WWO0u9606Fcef4NO3bfBCXhJNcZmh+M5zQ9NoT
4Ga4Ls6vu/21OC4Bf+TCywby/YbW9okWWjW70k82JtdDjgutKxBNggCEWgFc+8B+NY0vh/Ok0Var
D15/EkyJF4cy2B09RkqKdo2iTGuoEckjchocfS++Fl1dyNjthswVDQaFGHZFTZi2fkDbqQG2+bky
mHc2KF8U5q4U4+lzbcbhOQFgIhYgCLSGlC2HWbZR9xq7QfHvpCD1mjRR2WsF4I+UyZEI1Kbtd+Za
0pPZATmwqkqD+qUwj3f8cRALUQTPhb2emHV4iIRN5hQYmK+AeXpvoBKs7jr+6MS8yfrNDqrCICRP
jdpW2zhnR276kYkVM/Z4kxI3zCSHxaYwHuF1I0dSMcWimJKaFYFQElTDY9eRuLYzmRJ5EQERY2Fk
oWgGdx8uoQwE4XJdXl4KKuuUqp8cPAvYDX7UMH2e2yrkPLpmF+iaH/NIH9gqf0WudlB0fPMZbEq7
8bUaBs8b3xbue1/qMbCk9Q4/HCZlV+iTqMsPPOjoITS531Y7xESknjd5kqPs9HIUgZ2cdMDPAhM1
hGitVi0DRCsUcuEXximELD8WI5ygODtn1zdU5ccYnRX6eOH+atSoatH/Pawn8IBQeXoC8FEHa5T4
in0IO0DhHA3WH+TgNw6dlw9CftALMfzXYk9hdWA0bdwCvyQ3Aqnt4BW3SqJeLC9f3qPcPrib2y3Q
yf6yHeto+RHN8oeil7stHbktqVJ9I8llFyN4SVd3LbFFQXyspgx2ZYSn1U5Fcu2Fnom7i+2GKTI0
gluBObxRNklQXyZvh50QM1v/Kl5itnz0A3+6zyLc3o9fUIzVlzflnBaplB3paCe+1uw9b6UsVQlE
eWXN8dwhQhZIzPf/vNGEP019pNaRsodGcyl2PVDYCACHJFpCTKGLxbIAhkAJ5G5LjuQwWN2oTTY0
aPEdDhjALWYzaC3VuQ145kC9OCDXL9vNDOefJn97fin3jYOS4ak4SBNQL5JKPIBT+DtM6pMeWbGD
M83UdRQHY6gO4xVyCDMso9GEw7fV+juI7V/BCmHchFLgPGk2vHBZYsi8K3/jXHzI67DjkE+2uACE
iIiG2ehvkkbrZBB92xPBc14W7tWemBouiEQiXPgJpLDkeLC3yVB5n3Hbo5YMxFSXPemEGhT13iS5
pIZXHqD501b0n/9jXj/TB/g6uAjI9olD89tVfm5eBY989gROddQdjhlH+wfr7SDUEVMaogcWviJT
OddUoGOmhu5dynOK6Bo8Hy+Npn2dQjP7RV7PUNqCUYaqN+4PCWJY4rVkZznbZwWdAOHZM5L0pO+k
vpXZXrX5OwgdfVq3xsLtWC6n2TdT6rhKPF4qeY1qf4flISwS0zffjUK6u62KwkSthuBigHscIEA+
VpPAEMR0SGH+cSYuunm4NtKp7mJaZxPJxmYsSiWrLgPCb73ut1rM1Od4/e7nkKDD7RB1hezhVoEJ
zaF36sFmGhoqWV8O2pVKRLCZkqjJdrGWJ1KM8N7MzLMKAmgcbDYCuZNoqJICFW6hcTR24H4AdLb9
Jm5JTmnBiZIjgZ5c+zty8aAnHPvCdFDI6Se266jZXwIyGAtRTSWQBF2YCNtqtFJTp68NA9IBPHVh
bi2w1ShrzYgUwMhKLcnPXUrR4hjg4NSYTjHbwyn5hP9+h76NJmQfO4zHl9l+Qd336kXHHli0Jr8d
DWzbMajz6ITwK8QXyZ0KDdDThmh7BhznPUOSJLTeUldIlcJJGMHw91E+w4i9J3Cng03cu3JBXjGr
FCzw3mLvS4eR5TGQ8UmzJD9As5U8C9bCP2L8uE+tPY5br4WUCktLDLtaVqF2+pQe6HAt524bonM+
n+VUBS2Q/BBu3cJD7mDiyO+KCOiFd//UqAE01Z8Vq9F0cYbVYug+UlB3FN1BT3JZl9S6VA8wAfHb
BB7ZfcbQBk/6GVkBA55Mtyi5LiLZD1yDwR3cDhoFn3tWooFXtlSsWHKOQLkXUvt3KLLcNX8VkTit
4kJRFvksXIi8BE6BvWeq35B51qvTBsEwd0NEvCkULiAB/ApbTVIKWC7aZaZeoHnOdX9651dP3au+
Pl+BAan572YBfFqoU05lrRLcymbZCUJqEdMJCzoo9LS3Wq7Jwaq7RtFBKSWtF8RTNHuKGsZ0X+np
P2xBzvmF3ujkwTW+tubVrcADxDmjVjrCCiEHYw9bH92P6S/NT+4QRH2HbmV0ZfhbsGkwXJLMTVpc
W9JN0BRreUCVPdhcSUKlFnHpE6T1MhoCSgrsaUIe170rCUxIvXbEKO5hxUd0BSSawX+eJuT3urlg
8H1T5vk0Xl3PACKn/Hw6OSQlEPevV8Cj+9kchKh/mo0Mxm0ePUsxPEMbKcV2spF9IHu08MNgsyq1
9xGGYvChrVZFTnDlGbVThBshKu7TJzXIwL2XUF2gbSX50wZjOB3quJzYGKFVnWW+Oz+PWoeBH/sS
go3RMiWLhO3lRypSyAn4iedRkxOotR/gtKNynKegAlgKIAhXpPvCBWxhiN/zEFzxy7/ki0djZDBF
2UXRCwXPS/WGliHzXNE7gcU/V09x4EfzoDHLSEar7pIixMNS+1PpwFN/S9MgdSklVhq+CFDzMcw9
8K1c/n9lOtFE2+UGRzyi/69lTQnL+JIIaUcGV+qRU3zXXnNRd+OCiCXYNbntWFgoh51vkFi2Q8B/
p+KjVjvOkpLUJwpooxQe1IqzUw2bmlEHIYYx6NEO2eSu0v7QwmMTyuG7g3b7lbOhVMCBCzYKaTu+
1VVGojNCiO3SXBbKD56JlpDJ41D6ZVBTdf87ulQTpeUsLIEmRJ59vAtZD9LysQ+UUHix6k5k5f7z
mpWVQ5B5pTScwSlG+g1BnuSqNkQeYjI+lCjDwS/l53L/K+NMJjKOZz+O+20hEoP7gZgO1p5rzjal
mM55+6nouAS+uLYcDu/z/nVr5MoAkgn+2l3+8/fMoF/KIoRgeO7/aba4ZDFDpk4fBzjwiAx/NHJf
rajlQdDAYiqCzdpv3qiiIozm0gIcnbLEYio9zKdzS4aTAS3JfF0BnOZWv7lkPCHbEG72g3tRh32l
GiF2G2Vos2ihhFKv7woVGEB1kvNHkzhZUXzyVC5o3wmB8dt2FfaOUPgv2k8mu89TMwtaJahSv1B7
53QXjKP+w3K55FdVDD8gUiP23CHLpcfhTYzhNf9DcmaBCgQc/o92HDiqjSJkwJRu1a30jyPtJIBl
Q/T6VyElbq7KxEGN0vZ/fMUyRDzQ+U101N+Jetgqw57bnT5ZvKe7FOww+u6hpGiM9jYL1XEWKhVO
9s0og4YBJjZfIEDwZl8GqyA68SXFmvUsW/Xw8XT3aUt8W4F2wkhbLZr/YTUoix7YfRKrBXxJquEG
sr62drYiM4vIGsdmCTw7AWboGT47ihGbflUWQQ9dqYieZl70LJHwK0SsvU8jSpIayUZ8P9ZAVoYK
eHw7NjE7WwYg/KhaTRobCe7aV8cFmIN80JvG2QE0gp6R/jyETZa5Y+0H29dHUVldr3pGYHnKBUlO
MMlYLKq49KoAF1AamjJHp+XpD/RDf/nxFp4xRqf0QCfd83HbLbramiQA0Cz9Zqw9C1j7XUbAtgb/
AkNlb0XmXWgnj7clmFhFHOwVn1tXsz3U39yA2b3AL9OoUIZgeTbXyKhIuTXExbiU544nEVZX4Sxh
HtZXW7NYQ8rdOyO7Gnzld0XhhHfZd7glYUSSo6oHo2yMbKgkO89O1PcSPkCDiTroGyrpj+hoXOMj
DD6mjmxSDbxds/+OGKefJQ3cxFmfzpWCEniyEKcV7/HusZvKfVYXb630q1lqdKDennUeZkUxOxTZ
kI1IOvfIdicG79uRgGw0eyodMpMBTdadlU/UbWQFknlvEA164XZ1vuMc2bI+I/gdKLTKJtaRYGip
gs8LdAkm6Vu7kG9Jl6etOQVwdSaK3kuzPvHhjzxTutchJDkEFPZZ3HJM8mvjDIy17NIhmkOe/nas
Aq18LirWZG94qHmn8jiSdnwnzR3Cb0SdXeQvyBY2QMd1z5Mlm1sQjX3SKR2sKj50lI6AnirYPKQL
qA7mETG2x2UY/y+1c9WlcLWUtHTHXLDSREukdZnjBw4Yb5YqEXv0lQhqFQKpu5xYgRGmVS3Q0H6X
qYnEM1KGgE37qqGypvP6wOL01Mc+XLo1h27fsvfJdfc+MnEEw9zySYKuhsjk7L5NnZBUlUcojIA8
DDDaY47XLXiMEBxLrU+6BXPlt38tDhmAZ98bZp8wDsms7ltR/Z0e9sXO6VnMafIAxMU0vJTiwf/E
3p4cxLfAYBmkHMMZBdA44318t6JVF00wEqjVSCHhuMqxhxXOpkRMqDOgMC0O6H6zoCKyjuqrlFWM
A4RYpbEM42/2AF5OtEONhmQTuxWoaIE8NafW1/By3SbvSk7NatOd0VSVt7VehK0sxz6o6xfSSwhl
v7LIya15Mfh/FHn1G3HNLqhoL1XdsnQJ7/bXTQ0+AfFSGaYpkLYz/+Iwc1OefmTlMag9Nhrsu0ed
OEaWQlV/EF52aiAzoAPYh9Y78S8WkMNapRjrIIXit4YB1Sx+kNzEIX8Pl77rEBGkeqrTzWylVkKr
tuggBtjXF4p7E3kW0Iz2B4fHjUwdXFMNdrt1Mw7J7AiU7V1HZWK2Wx3csGMXEHtqFYR9VftALUpa
x9yeurjUbCcHXFPc+uAAeJY9A6bzEHSigtENIlT+R4+OnvlMck1Lf8ZNI/7juqcrAXptp5ZkySq0
WZxm/TyTQyrF6R1p/CqmgAaiTp63hYx0CDNmSSLhrCHjdkbLLc1NCG9wz+xNub2PlGkVgT6A6yWz
TM2tWYuco3JvjCdSRrh3Z0Qe+o0DjTMUD6mcV8y05QZx++sGNPuLwjq8wWwiIOKMIYlwrSJV2JaY
jLlOl2Q97ThIKQOmaR1VFgtlLeeA+Cwv+B/8R9g2+TF7Z67fRGbm9pG3BO6Hv3HROqxKVSBGvy6E
2lT8uAfMOjyVhNpNie8X4IOkCYOft+Ucia3/uPRaxJqa2biuSjG8HkQujy0k5PMzGUT++Ih+kmKD
zrAUX2rKAovuJQq4OelI3ZGbipEeTYDgiNSOpsbE9yYohphUt1AJMBiE2g461pgg6HfNiGAW8uvv
AQSA48INUKk8/xwn9OU6MV5kbWFAXnmAJISEUtMINuoR3646aDwVhcspY0TuACKUlmUIucw6XD/P
gkyXAppNz0tazb8DXRW7WYqCMVn9wtYvFcZAV9lZGb8/9R/kBfCa+ldrQWXOC1HI+FlP9F+YuaDG
G8mZfDCTYtHo88A+5LSt9IAATedpYch/yaEjLU7HTKZ+7KObbWt5vEJCKf05hCKNZC+/fpGBLzbL
nZug5avn7JG8Fue/NWl1b9p3/UHatsI9JEFqJTbjp4cFnG7NOsa5kJIYt41+IjPuZFYpOrV7j4u7
Ej8toDswisClObHjzcsOspd5W8qo5ntGGTkUn+cNeyDV+6Dz++YXazM7k59oFz+wH5Rr3WejPn7g
MZatYTE9ltgCcQlihH55KkYqOkM995DRD1VdiL9k1w1W7h3lGz5c3QRztlKI9Xe/p7v4bEz4aXd8
ykYwBMeAEYbPF2xhS7gNXRPn42D+7hyCAyHdyCvVhX+AYpR0SN8pictxNtemFSTMX1JFr1PP7pXe
toPa+TD4GssBJhbWFmqHSdBrPpuCfn+cBxuvYvtsX25Rxckq0cGoML/Cb0gbpaybIdQHiDkB7pRK
FhEag/+NJq7VHiA/ARYxF86g0VFjHsZYfRKcP0FIw23Z974nLZxKaQ/3twyXXQXtZMO2iROS/qoq
FLA5jPfSFgws9JghWVuyoWX9qmXkJP+A3TeETt/eV964bA4TX/LAmcYZs/cyAD0HTk+OsdgI1H8+
y9WgSh2v3mR3IHsFkYrk1tcWOURTc/8zED5/bQoXkfeAoyuUQEnF+T6Rj9DiHE2uZTWP3D5PcrRK
Cj32f3wnZcusCW2zclzS0DaR7nXp94PVoXVooj6l9IJckDo4/AYGfq41T5edTGAqFEzb5vZEYsuR
sd0bZaUNSw7SA71Ly1V4B08LmX5dtiBcaONCtulT7tt/r8RWHmrsKWvu8oNE9e7Y3/Rosm2dV1e2
htL9hFAOrUwDTl1hxoXfGwiWO5vZH8C/dvHwqmZXidIyAB/pBWg0VD2H8AM8BKpVpNyjfsFRFTwQ
Kbqyi0v6SlKBhTev98qTaXzCg9GGWCYPS3Eyq8nll566xh7q/qZL4xwaEnR7omzmre7Q6YvFYI8Q
MfoMwgmrlzQ89JGf3sxab/EhPD+WLqlHyvA+apc5GI1t+5fQRIZWAdw03yA7vS0XVuXW4QRWCcKY
a4wKCQQLVFo9JWVV2U5vj/ejWj6eAfc9P+hCS9rYExGXYdZOg3BS/5ar7+8PcHIGUxI7o3XdMKsL
I6IKCCMN24wr5pmTeUG0R92sMFQG063yMECIKylFIvZiKQ+LDydmtnBWvoS6AZGmRru8lnUZAHXc
v5vM0yOSvOAc3rT7ZoqNrBDVeiMVjLiAB/Gp/SoRDMAUbxnVwRYHMNGQcA0EjtmjPB5ddQOEN/tZ
VIVsMAQwMLWK360sG53Hxa0WMCgpnmC/sNipFLaYu/NpgRsN0XuQsXg/cjUCJ5f/sAeWljcb6CFT
MJZoVFZ4Ai0ByOgA2w5H4V+DCfYw55ciCzZ5bMotm2OC9uDlPBELL1pS72tv0ck2eMpVhUuGGy+/
uUjVNMLtP9HHvSVORAMCSqOdYWe1wI5zJwnG4LgIQCGPeGSvYKGVZ2bmMxbgynU583C7NpCcIV0Y
0f8kT28tqsOrlLp3ZMPMw1IUqRnk1uAPIh+ZU4AIHRN93fQJmQkhMYOsOjQDmEqjkkQzS20FOFgX
YXNGabPEzP7Gn11jEuPAQiQmJeA0r60z8clk4l1Vs5DHVroK1+qErSQ00rNUTJTCzKmuvOYoAzyZ
42xOPc+2lWqTaMDDbwz6F3+rMRt/G4qRorPoABPfxRvQxvqNEZ2b/HbGOF7c+8Y67KAYLVt1CyN2
91MktJCDVSuu2GZ31NdRTs02FrpIPAGX9HeGgd4EOTN/FzeHQZIIUSLON/wjivYsxgIMWUX5ahHJ
ktL3YZ9rICI0+zpisc7hA00BFW7yzu9jDykFiHS/2kJMXDIudPqNiX/+s5chAh6AJkU9t+/tia+w
8GV/rD1iJgac7s5ZCfqFlRL8nQf3TcBweZH5UdcMKpXIeRsg9tiphLT28fGDySElL1cPLCNSZlhp
ARl/UF9idjZMNRb3bbsyI5n0zqrrsu+TnKuVZnRwDMf5ACik71q0aJOBBJxZE5AZnicaXkBFlUFC
d7Ce7NUDkSuKm8ubCJdPBYoDaG3kGe8AMfznaOyGexEpBO/j6EyQu4Yq28cl/2C2bYifhEsgeqe2
SXEOKWjwO0JbgVsqH1HXsIFICLjlt7jDoqzeRgBN777sOeY+wGN0EdogsxXzwPply//6OohHScIs
SW2lpeqzafe2lAZRoVVcVF13NWURlx0ZvJQklHfSt3z+KEkkW3PZfYzFYUOUGdQv6GgzezhhLdtb
vID6DOM58WPz1vZJbkF6n9O2KJws9r7AWI9Msz2KIkpc5Poa5Bc/6u8o+TQbASL3rYx5okURpGBO
eX1Uy/4XfLnU0scy/2yNdtRKtsj4imCHfgmwK3ylXQ/+BQX99Kbkj4XO9u14wwZ3/D6gzFRFSZYq
46BNh1++5cz07lgAzdg+y73vCL1IdAz/yq0+Jv+S3VooVGIzfbdz7S/ewGNLl7XiRZjBctNdzMLU
VZVTKMmH4ps5aVAgf5VhwL0PBGFIURqAYySTcKN+teMtAb0aUY+HTatLdouYm4qFATBmU9Pcqiy6
Xz3ZZ/1dpLClsjyYxdha04ZH/fhPW/Z9/tIes/XAo1CU8SVboBcuPn/OF/wMn7MjvRsqxst6qUh7
OVZ9AtLotp2EB/9YLdePQmCvVcRdATcRLj7K11K28Fc5AXRa5B03ZTgHDa/g3p2ya0oaVYrGLFLT
XKeArCInOgcnNU7r3Akp58DM38aS4zP/DDP7LNgRNXZ0SOAxXClR61jh0JRtiYMT7RRqgo0iWsHK
JGw8X6LmIP3CJpWmsw9GKD4mrFAZhRobF2QJCcn964BMqbG1WomaYPhAZaYJpRQs0jPqDkGCOnjZ
rAzYHKMVWY/96+yvkq/+5QIVN7tSEEy08OjtIu4/fOQXTTPdYI4R0/5temNuEeP6lXmUWt7PzHZd
0kUlgDFpj3c/2FfvFm4BMuGbS19VT5Pyyfev0zKXRNVYpeTRSqH/Yzod2D7Pr0gEcHFwa0yqY8ck
L+SSJJevj9PrLbEYo/3kuCn7uwOe/B1tHAWySzz8GWdJ/2ssfsAqIgqlDAgBz63clyi/UkLqvuIs
DagM/Ecd9JQlTVHbPPV/vAtIMRoNWS5MwsVa2I0XwS6U8MzX8GmqrF+JGCEenY9LcBWr11G1/yXN
Dn49ItKUhbTLrxByInS2OEjCa26IQpT4z0lI+uIkI1YTLk8QkM0AjPCjWFz6+PkypXFZUTjropvP
ECIORTgahUxkz65dxDhIQubBkVmIAHshbq0tVonf06BT/JSffPagGUg7IcOVs7FPaQSIxfDc7Ugy
37zZbBPyNo1gB34LpxjzgSfKESfSmCh/7rePPHen3YQpK8If0SJJZ5aA66T4S6JZODJcbs4ZA/26
rrrVl0Ncxw7kYfpTHLVIN1LMD2XwHki5Pewsoxy87HtZpv9yJDjJkwQEoVkWZxqjXbXfiomQt3SC
wg/tKGuli9bEeHC8/wqPyECOiZgxc7T7bTFkx7fEqIAvMRjfJ6ALl150cQ7bSVrpn9vv1tmfQsE+
/+GQCXk9Bpr3U3Cu8EpCiUR6hlFd6ASHTZbWBKU9DOjnrCcB4hxLKyCtOsRG+hY6AbLFqURWde6E
snCp9wTh2zeVeIKpe3pVID6D4UvDfNedm2ODp9UQ4RIvWroWdKuma4SKB7KxzqOH+0mKU5gaXJAm
QZbEJIEg6Fp86xovZgA3gyJiBOPrQzesjL8VHuNXumkylZjlT1RKdEUGwKM28oHEhVKSyfQszsmw
blLYwfaUujsiJlrvQWx6yUlUQ9VTDNT1Du4HWARPNpEQProbUOqVgAsncEX5VkQBk4m7vBkDeaFR
nyRTttezPFHxccYL9btWqmHm+8q8IYZSG0kWZtdX6KPAvnCu7ZV/6QeaPGr9pFIo7AqeRGOzje9z
bchjie/FLfzLvgL9Y+Nmm/5ueeX8uzA9F967MvHzgFZc3RQcRfHZtVI/5dxRr9yfs6b5YQL8p7Qc
+hNvPbZb/LwGrO8Fa/OTVWY1zqgeKehGEwfb6Fw1qhKFaGX6Yt3fEtQMDZCvCGSn8rgRvSalT3s3
kl38xwl4/KPKx4jQw8rVGSykFVwwfIa1qobYvrsuv/nHY01OJdQEY2d7T0EMqbxl64auBTRnsHou
LCmoP7TTRl0SWIpxgD9fqVBInbmTrruZtT2M+2+cI/lWbsB80IESxpAQcgGWz1SG/5739O0ZtHj7
n0Kl3SNS2amryHe0lCnpHsRHL7c7bBCoAUHBt44ZVv+ldGOHLn6VG8iKpkRVsGNF3Oq2pRS5717J
OVbqCwBsL3eAEOqaBY0GYHtBMgpVMiD31l3+gY26CJulOqj2CuQ/KisZYmiPjeY5/6SDTKpzO/5u
HDSxdIpxaRyfKRRmFltbSzOqKkgDv0yKHDokzQS+9yp4VFeccSVFdPP8OB1G0rbuuShhV/YZZFBA
g+GEIRIoetnVF/mSg0RCFHpCmzbREuphs7q+954OxMq+5+mgDVqf6m1yuyaacQJBOwWaA6qhOZY9
/yUtKjwYyip3xlfliiIqo6T6jtfTMoFYmuBWIyB30IPYZIpuKB/0JK3XlnCZXG25tLcfoPRKRc13
HfDXkD+Q51qE1d2Ed7sUAS56cSWJWkXY9Nh2Kj79DA4pXMLKTzhYKyCNnOhodNE5808YTfZ90p99
tTeWbXWVbMdXFU7biqRLHRgERmWF8DKxRvhGS8i2bO4bKmfuQmBKcN0ZSlGNcOlC28dzvKkh5Ui1
OePw6rxbUwmNukTgGGu0X1f7L28che29Sm9xQqHly3+fAcXo+vPagvvRVWGAIaxzP9R5Xy5f+AJb
4qY0LbgLgi0DHFdSuxvzbzoij4S1cllUGgB63rJ4paytChYBnrE4S9JK5TmYxX8D3jyio5G48Swf
6WzcWd4ObLTzL8T5MN9ccgkwZP00SbFMXe9KIn9CSDOjWX0tWVdZ/tnmpCARLVlZ2lMhvGoT0cTK
qWaPNjwAzC4xZLWAmSTRR1foCger8hew0mIkABj3bQb/fCuYTh2544OanE5ex5qx3CNbW2CN+7tT
UThcEWcDlSfnmQNK0Wt2HBB1EXsB3gQTfT2O2mH7U9hEc+6e1OTs3U7kn2zYFBXRBY4quDbsKLhr
sUYzLlbtbEM7YUK1mZMmC8bBSCmsLSvbHBm0Nn+bi8fMzIVhhqOatgO7GfC9yAuOcUnLqIw3PWmp
kzZgbfJk7BfRn6deAhtJpazSRLxX4Lp2RNfR+F36++otLttuJ4D2NQVItuaDc4D+TNs/7xOuDzGX
LlBSyU9xidijDOFM4GforOSxA8siC8gERZQJ1O833rS6lDjw1A6rCIQXW8uj+57TY7aqkW/QnZO+
Cumzcd8g0litOwt+MqSJr7q6ISHRHYUJGfj//y8MAQpdGnKW5VU3IWKbdRUjNGSmlAVLTe7Uw58z
bbXTqBVaZ/Wgqxw/t7diVNLrtcoOLq0ZdIbfVN1KBpywlQRtYgF53cn3teHnOJZ1kJTG5M8wtjnX
070MetC9hkU7ElmnA5sbatygkSSGjVTpYfcAH+Khu4K0XzoidWZog0rg7IqPUOoW36TxeR5ACGAP
qQsImnMlDtYjez+0RNEvkX0uCPrMosNMGNDAswNuiFcDtrz0N9/zg3GBEbAhvSV66fRc9TpmMoS8
N0kJX/2k0dZ5Ks0G1znDE8825ELMCd/ut/u4kbR9KoFAOxAQgdVYmRd+x+ipIOYDZ8ZKj9I7SzcS
59f8/SUvT22PsvXAapqk1rk7FRURxX3Oy+/tIvDCHChzMMOZmwHAgPFgcwuFuf1rSSu1jRHWNiHD
JJ2DpBPvh1FRvKH6S6Ujj1/4p67isogDnAWAg/bBhkqZ504WwkOlDu5wFR2ewLgV+SXDqotPTzW/
tmrrenXJNH2qGxZeZMh3e8QQlvIM4JA4x1Xhm1uhc9P6frnw5+Z+mM8mlvGnLLe+OtVAAPJA9IKF
F3kzDW66xWtrf+CkDu79HVr0Nefa3vWu6BqSZv0DPAMxMpN+9vLRC0ubqGUerVhe7CrG6KRLe9F/
UIq/b6YYeLTLE6VktJ1qntuT4MFw1KfBhbRHCafQq64KICVhTUJhY1IzXYiU/AyqO4dxFmzL8cJP
nekBZjhNycQfQkrrBpUmEv0zk9rYd+S451YuIzqCCC0p9IFnPaUBfdkkq+4MFf6CNzLiClHLKkLc
zjXjWEuXh8OMDCT8SLH6YPCd2Sve1h6J7TLR9q970uZokGk2lWhxMCfRiqaWZ4UjnQJqwBA35Rz5
WwO/j/7TfEJGZxheTcrZitHRH4hCtLtiOz/ZNduyNhKNbxSrVywRc6fLicSBDQEMuuh22HZ4pIjd
VhAVB9DRBIIVdK8TR+OE5xKv1eUUq+du8FjTl6tyA2TbnGdRFwhtC8dPEU8aT97G2jtpmi9kUIBy
dNNG72L4afh1pCHWGXaFFAYuukkf6+ZB/sf3fbn1cZYPCKd/aSBvqanLg/pFLysvUSZ8Or0jo5pv
HX85COaGvE1BLRZz5DvuAqV4d7B2oeHV+JrYWJuOnqeOpYxSYkol67C1z0Kf0dqCV/l3x9GOu3sH
fwso58NPQnlJ/LdUOEbai8u0FR7cXMiuN/Xz3uJrX8v8fUiwsqsXaUUEtqAKXSk6XlyWod4+cz/h
KRx0mWqICOqB5JPXam7zL5NDMTJXCZsUEVFRW62yUcNh2n0WTFbmF9xK1cAkZeglvEqPI8Zd+tzH
e8925G3v81Yjk2bxcMr4wiymizekYGDEy3AInrOi8XHJVyVueIBhuqxufbBEULNV98zvI9N5BPZw
0rw/dklRSvpAe5iPmiVYIj+ODY1ctrjtF+vmAsyX4PSg2rA+thLIn7QKP+HsrQ+V2H+sP8/+8VDn
lbPkWeuu2gFrLaF++nW3aVD460B15pDHvqDKZdJrKKH7wLCnXUJtWiG4jy1s+wxv3C1NJuFJMBS8
aX9qK7iNUIikgezny6wXrMHnEBR/OE97ZGmcwOTTe4eCke0qaRk3YAZoh6lwxoqRSR/f7lqbdAC2
W7BRcnWjVhWXAcbM0NhycL+QzvF7mVwdIDpbhwh5AcuWKd//AZubJ/nohS9jIa2ouEuIxXBTLX4o
vMih0wo+NN0dKJQqOTuRQz8yPRPIOREG9WXBfs8kddY0TnEioG4ilPJiWO0zyM6cBY4MlulYaord
TZVD8dDdHZSgpZ4z+FkOIQCRP+E6uDH80PGJfF+93z4kjAmhybSvqH1AOeTuCHI8bnqocJlYD1DL
Esk8C2dsmEX4GArGqs5LqnFeYp1AF9QcJBzlkPW5KP9PW+F9T2uiVgt8Sh1zDNMd2gdc6m99C4uf
+t+Tz4P1Z/z+I/u8ZfgWeQazP9a05Z6Vra9K+rcWYO2fPCIKxd9COufkYOA9O/f+pzsmjJsHMjse
7cgYFrktiSpyeyKbgMohu3rdm/pu+VYnAI4/Sk4jSPmZw8TOSpAxKWyerUlHnlanZpCkKHB3q/EU
YaPBlnU/e6+vOzlmYlMYkWAuGeCQqDi67Z2KwWFf4SWvVNOzdgTy61uZ5NbErhoXZvyeTMgRW19u
BRrX+UH11Z/Q4Kzd97vnlSd1sD28FrWqUm1Kx+3j+gFUplmBAn6c2CEJtO8LtgEun0+0jCADtgLF
2k+yPSCpUVxtDLfOkXQHwby7M4Z9ue7DeDsVvMedcowCTFcEztz9rdm80C4EEGBLaGoQdlXVsaue
++eDUdLOXGh6F3024Igv3kHc9Si4qv9PWN7Znr/geBFSJ7ia/26/eIR9p+qS65/yhOFVFNGR/KPz
1mzHpzc3/s//SC5Z5X6i56n+nf7iZMmOlLE0uB0+D6UD54cWp4DJ+8RvPFYrnv714BRh4BbJaEt5
JxDZtd19vO/h2/P+lFPa1tdVmrmtTLYL0WkuCpJTyyWv4SfBZLiXhc1IuA7e6de6r7GaEZVDqf/f
SqPfy3H56zwibGFnEfbfnLofOoZBAxK1eE6Fd/V21+msc+DLjanQVYB5EladTGkNmxx45PQKm0ad
bAO1WwG4/zlhu8TQAwgMm6eKVcuO63flNCjPgJIiESQoMgW1Y7tCpGWE2r9OZWwNfS8VN3wflGhz
Vd8CAaS1dXA/zfIM6OGBLXGPCZz6svL2IYh49LdJohzZ1Adehsm3txV6N7aVgocDMIUiZdCer2uB
QbUFQVmXyMun4zZAQaDjHc04z9N7Cc/GMe6CLzqj0UAuCfWYbpIiZwIoit5FuySsczmcm38x3upL
Qc4JLsos0CJ1I5nugnSvjLPNC0PvzyMn602D1uDBfOchR+KNiR/5zopeQuMPU3kKLf8QPi/FgsDW
tSPSIW4Wbrlx0QFN+W1jU8lsmupef0JnjyH28CLJuQMDgwLvt6bYE4U2nFutETKToPm3D1o+u23Y
D4IcWXofAosE1A1o0zT7vU+YbmquEVkcyTrquGGyQdLVjG2rod0EJ/zSR5vhfAgFSr31fAn6Z/Qe
CglPHY1CtyEexLlEgIQUI+MqpErY9RwmnOOgqrIunFKQUps6dF79JiHzA/DMf42Mqf+ePXzV1ebQ
eu6t0Mh0QIBS1ZFFPb8Sp5DRNkbFJJ9pF+QLDujgwOEc+VzPeaPnAeLeIHERC+ZY1MJ2hohc5dxP
9Tgn2bo13kBALgLECk79yJ7mKIsHhuWzmmE7hbIG01XH1RjPbouskCebAPbsSYOGdf8uwcY4NQR3
aR580vceVwtZqI6fAZHujKXPG17smu9Hwy7SX+s083tQ7SDw/W+FT/i0orrVpKxs7GnuifmJmoNf
yyIRLkfAHboBebca/CWDXW+uAq9Psc9iPZ6KldHjc2RAU2hXWeR0Ry/lTpAylzm8SSWlJbuwYuGm
rETaM/BDsdpJ+2o8aAKZ8Z2JEw9ztI76+ypRRnLfLbGmpD8j7TSF30QoyEHmm8Aj98XFJ/YQ2cTq
sptI9b/qHwDQqs7ylJK424oQUy8i9TdbNey2vcE1GZX+/P7cSKY8+2xGBWuM/lK0rjROFuP1crRI
RhlfYcqF9hcv+je2YhfJ/zoaH/lw0IviXGfwBYB6Zuji/Ib2lZCPdffdd27k/U/fXkYXF7VC9DwJ
wb4iDP1osratlL3qIEpLfNbSoCWW+/xXRTtCypwtytghscuys9n4LemsEF1g7EDOL5jGmOISBC9F
bkUzReuRqeK6J+4HpqCTc9FqxS3vRdY3I8B+HM+eUj+M5tidx6u7Ubml48MtiYAD/mRDmtpjb1Nr
e+68+SVu1EjayV+Bc0OmewtzmJCZScoucu1SWIvWQHajegGfPQfIWr8xeCFWb/VsHyHnflYmepXL
i6C7jOnUzvnUlGaElGj16/cSyotgNEDNScSAc8EdjPKq34uwqZuv9QxwzQ7Km0Gis2Yhkz+Yn/Dz
56L5qf9GEcjItGYgnIglfMfgzy1izxNir+LX/6yirahYNFQ30j2n6XpSC74wyLeq9aQ87Kup33/E
J8OSgh+RA/TWOkzYlkbNgGmoM8Rpo3Tv4iExogta00hl18rAx+dm6qZaBU9/6xnlVDOM1095E9p6
ErYqED9aLZKck1bn7EL+1U2PN7hN4kDp3MxO4RAp3kYa7bcMN0K2ezMxD3MC3QX70MnZRM84sxgf
Sn6pdS0woNKB2lQQ6J2wrY+hTksY5yLTFuUdm4HhHC86CUin7t16M5dfDu/wKOBTixGDjOMnvW5u
vMsMjPFw7BraHA/4KMzkmfTA6zyIrOGrz8bGZPV9aRPUWGYfdscuiiGvKKY9ByNNuxkZB/mDXFvm
nqVOWNuVFGn0j5zYdetYLBo4jq4MqaoxXpQ30ZPergrpLl+P8F2XVPpiC3lkm/2+Ri4Kigjp3pBK
bUZqktjABmHBNT6CParhH//LSx7t3t8ErXEDKSVoITGtVkKl+w4zrrU5jujyazmafVx5RxQ3p1OY
p6tf3thJJgRSk6Gjcm/IWVinH1HACKJVE47+HebgzcS/bbNH++WN0efMTjoNlDJxvdxcy0Pj8vAL
CoD5NSzuTYmfBCxNOiKIsAfOP6VB7eMwkVB7Lvrd5J0/6i00zOelVwevEIe5yuNBgE0dbShyIstq
2XJSOC24kUt3jhcFAMW0TBJsCfFgysQjRJYYZlVhmobM8Bqy62piExI6ASR0gzyQ7mc8Z2/XnmaD
HecFLxcLhCLbScMk8Bo0BUmo3xQ3o4mcjjCD4OMu5/mwCsYJJ5gtFwZL1F9uhEXmCplAxSFDvpia
WJbOHUhWjWkFRXQbBYW7Hy/UMIwJZeg+8qKkpDuaeQkTfSgG/M/5vcI5DKzvJit0q80ucAvPFrhF
dvWkdKsfnpQJbRQQK8wGzDopz4Sruw7ICWuGbD1QhsIo30lS1h2L5Hi1WHyvGoTyDGCZqjYRGaTe
Klk6++VGlJw+zB+eaPMrxG3Bvxm/ZgI59Ak4KB5JTHaFdaDJ3F89iZ++MzWtfHiAYk1TkS9EZrlG
jRb2Z6nAo12AepwTILiF90986AhnL2xloS1hYow2JGefOJabGp/bvuBWb0YrPBF0ewsGiTIXNmB4
vbei0t/IOJRee7Lvus7ORN/B1WGpL5pdxjn80cK0URq7JhQiJsJJsaO2ckKuLPr8I87UaGZ8xDd5
9vuT7HPHbikU07et0nkP2pLfRwQ7Mkdw5ZmZXGiZmjN8HvxMwduqeWPvoOJq2uapdzfusSxXy25H
SBsblxxK6SGRQkb0H3Wl+Zihn+4AS6f7qxSswPDUaek0seRoL2dbbQCviCmOCmABA/aOL/49JBLn
xc/z1VgWI+WnLqAmw0hWdQsKRShluR+OYBuncfFxKr3q11avAIkCt0UaL9b/7m8eEhxNfZVpm4vX
G+9md5TvcfixQksW27po0OjfCfHstpAgATUIU89quOTPrL1CWR1m4RTnDUpqQ/AMaS9dfxwfF/6K
+A6mTL1cKQDzIuChhE7bgVS8CnKwjINFXgvoz1RvpMoKWiv6qiVmC3DYsxIgsYEGAnClHyMmrO5s
/hAhQ73y5t+fWxOOXnMdHv/qhv+9yOQGS0ApyASgLO+zMw7q9aroVi4gZIWA5BWRxRgysdfV0LXz
awos0B2vv3pU2qJrPOPK/Dk30ayAlQW1rNDmAiKcyPP505D7mHelxsH4dJr8t61o+fVnn7OANspd
mutc6wbLbTlgBG0cEbfN+9Lf4mMTh+JH0DFFEFgTkoiJ6geZu+g6Y2t6VwcogMELkS6eeKM9hZOb
CMekuyRekolrG1El0fl1vt0QjiErMqpv9muNPxSEkyt4roNfbWi/xKDQ8TLseS14Dc8Huu5eRdaB
hci86x3XkKrQ7pWDXQT1oOKglcCcnBJYUTkTKLKkDj+MHEMxFXrqsx61LSbP2oG4PS8USo3sj8g0
jk705/IrnxWg5DHkQaXK0iIqcW6laaEwBEJWxVBodjZJrZJt8WkEXFQZ0iAsaipkLylo2T0pyZ2W
OvonoQ4V2qpkA9u6FoH17/npD9yxyGxI3TWA3cWaOYOlXB4g1eDrAispoHyZy4l7Kq8PxAYH47fT
RXKtUu++m25pZ9z4TcGM1Ve+c5JYRpZIhqlSvuOHlNGFOnlv46t8QSr88Bu4Qt1UUnFZmF6oCzm/
AMH8HiQ55O/6pKOk7jr+sKZAa2Ke6itx9Xvfg7R1EHIM13LpPqLKtVPWuC6Sncffym/n9HVmtCeD
Ccn+KUSKdlo9HPKA6PEafRAuM6E3Qjc0WR3sSq880bUi9XQCR6MEk94aZziq1gUB5Jb9/L8MjUkP
qVIgfUMkrpK/B8d/Emp/V9UuRRzNiX1B76Lkw7UK2299RZzRyJQlWOkrreeOxIPx8nkGm4jIh5s6
hkhtbiq3cvJQwxRn9YVU6LWRfFdsoeVHeXlXHjz7FO5g7ry00HqNIDKXgkS0f2U0A50jq/Gi4Xi3
DQF58RcFokNh1Fws8DSQgZimwfFf7gr5zMoj8d0I618tpaC0SZRVaVKlKno4ZNX25hYz39TbK/X6
/+1rNdpkxbdqsjRZgFe6IcOxVbTFUJg+/5GC6iMY7ieDY91xd2pJHAOgRQ0AftiVQAHW6iYEWDoQ
A4i2HmMIifd06J6v4WsY7VsCuIhMwLiXXRvxwsCN9BVkf3xXhjr8/3gqGGtnsid74lcG1IW+iylz
vX0qxHbqBQfbgUtCIrhCbMSdLHHE3GxHQrqk+wLn2uRe/kiin7/4wIV0/LI4xqKaS2Ajm5xcbxxg
nZJ6BDQu50NQwq9drDcMEzqw6p/d2BY8BUelonYfeoSym2GQ9Vx8QpKeczfTRoUToJvLHGhdyJyA
NmHTaQApu9rUpw5XS0nL9z6U+FWtFEehXu9w2PnE9lO0UhbiIZmOgE1Sl3xNtMnMt2cGAVmluQmI
l4Qc1AwXulAZJv9TDFWx7i21n7OAVUEUOEO16OA4kt15IgziKl7OXw3YOA++MoA8uOkLyBGDVJ9m
y48t/gaytrBOJNEOlvJUJzdMasP/drdkUdczKmj9sPAu19CDA08IaNcxKinJ/bi+M0GVVH8mX4Vn
J58/Vy+s0B5vCuk9D+mtuvh9K/Vy4JY1wYoXsRxIWFBztuXBeHg0jQvFCiM+V+nvIjz/C8HysBeb
DtNZvGF/lvms3DC61MVWyjhnpXVrcmgJwXefy4UMR0FJklg2TWsAMe0Ch5AuO/YMsx21qWg+RQv9
830rMs2Sxy7FJO9b6BrjSNS7pvswMglFVijCCRXaWwNiYQ+tdvGxpJOfjsixFjMWgGk/Mhpncge3
Yeke1ksRqX0IEn+hEkZIzlzJ0WXSubHZVzBoEulO4R0AqFlZjs/tipzrbjKH0OthyDDzUyqmI/Qt
5dIxHcw0ooLVY3YjiCxBOBv292JGCIjBNj/VJWyrTp+TPAvkobtfldr3k3n9f6LK5gmIh7Mu0MQX
PWskVvTi3y6ZxbCboHA3B2UaHG6PtomKTixHdCGZkc69XYs3vMyal4jw6mJWXBCiewaARI9GfOvm
AusELE0+P4oVsn3X35Wey7TO0g66iNW+EMPQdHDU7k63frxKYGR1Dc44tSQGXidgubGnG/3WAUzy
kacOEXzqu5/RPe/Z2f1GMuRgxftjSa8vTWE5xs/q1rWAYfd2sYe0ijax3XC+aWolabvQRCydDNgB
hZVoADgGmy1EN7K+xwT8b5r+jla45tbtJntSwo9+ILOyUfkWfqWvY/RmqUMWnt4U7o9aIllq7p99
Zzl8h2fadr7QkulAZpihcDf2YkXflPTNQQceqHgedsXZca9fMc/L07KKWcUBG9rGN1kGmz1/vGmg
SLkonv1mDhCTMJbiGVuMRSpyL700IjslNsov7dEAU8TwBUWXIE5fxhZcV+UEYCDC4E2lShLWB/J6
9tLO6wdpxTGbGCx/aU5tPcszThv39e3Ptn9v9uvwK5fABgFXopD0kwbZscMB5YDwJXSXmRolBXsx
hqWsnk+6qjpZ5Ki2JkFzRXknbYRHlc8C4xUNK0j5a5Xcg341DyVmOkojDiHOuCMv6vdxKDjm5oPb
cvoBOAgxyCbzUBMTci76s4UeuymCtyUMNWvJE2xxGPK313GubjPCzytVgudLFH5iMQz/kQYAnQw1
pyKDReGoYxXASVAbhNHRclEMnqTS3Cf8JGbzOjpCKob74pwmztmy4cNZqPNcduI2CzKy9wbOzMyd
yEes6QW3mAS0cTvvZ2iLv0HOqZI+d8RcSmIBsbhZCFRj0VVsvWUoRoqZCRJZh4rgIx3SjATIOC98
Kq+QRKJqDbA+irJyfveDjJuemNbxSBm0/jQw0/bUBH/iaMLYdYbMA8lrW33w7IV/5My6DJl4dLg6
F9cF5NIswXO5CW1o/VFQgltdCwyih6sqAJA/O6lXXl7BAWb6CP+J9AAB4HYC/30hdaey4a4CQIm7
9f7cCA25jv+u0Gh5DvJ+/aAaImbZOx7VvHbMyU/0ts874CNDsY5OjKe0J+eW8dytD+G6zAcBWo9P
fADE05nCXoxrkArhJ0upp2+pF5Si0OQKPKhT0M5N/pZ+B/Sj2OnkSeU2Owsg+S2HyGKcY2KQioCx
LC4VGqBPXdlqFMWaobogYZ+kRezdN4sjQtPB+M2e2NEkNBqsIbt/C8ox7/6UPIFLbDBqxTRreAvA
u2g4yscZyVMLUPYK/ZaXj/ANCQtk/O+jiJm9uBKmBB6a305z/nGAj7j69ydpR2CLox4qgfIkcoMk
EdPUJRKESUBmxiZV6uX3eR/ql/9M/fnc9Z7nCGxfoCs8KqPJQCOQWMP4+60wYcsAY7CLjQG+RQcN
+ib225PlkclIgqH09qkZbcBUWQBxyhyThQVRujJeyGhQmfump/1di63dZxeRETc2cVqYcIvKgUu9
iwzt6MgseUQCBTqUo+yx9TPLxHCE1zE7J4VnVTPDwxxTQVgZUHNdVjCEg4H1RMKAM9xh2uuWnqaJ
rJg9FAMxJypWC+amFyJ7v1rdRpxDfr3srPJdCdYbN4QIRJSKrZ7IHJba6QMlzMuBnvJDWawAdwE5
wQYOEQKUwBB9LRAsLR2Kw+nkcxV8fsV2ZdzyLoaHube47GFa5MldFx7NIjGck+qj3QjkP46gRLF3
Mtm63eMEfcy4AWHvM2+8RcPc7GHAmvzdUGoN4SJ+UTRrsGIhGgMUFCYjNrwi+IWqm4BDfobnPjRs
lpa1NaU4wUvd1lEaj1623+jfuUPIexAOBZwSY1wAiOqgsesIxjxjrGpqh+CGKESQ1JKkSvQ1RieH
Zob7vmfqxt+StXuz8O6cewPCQrdu0tYFyS5FtI4nIR+0xmGlLV6NL26+TZSRzqI9hKdZhio4sZp4
I+jSuJsaK7N5CjY+ngCydWk4Y7F2u60V5zuWRASPJUxy8NsFJHlOuny7zmGf+b24+Rvz6Wd2wfyy
nh1oi85v84cJL3Mjuc2SlzaPGEQ4J/eBzoFfZZZ6i8lMOEtSJXvCpMmy5QlOUJtPBNteBBW9AHgL
KgGiOyvEXsouiIKGlAGZ1MwcK5dWJ4Jw85IsjSPquXY0ofk82+87yHpbmPF9kiaQpfUWZjIYcP+y
ConaLY9BAU+d4Vxko4oL7J/6KHXCce9KWzfphzJI4bmKjQRCaM8Ce504uL+pncpXjPDEIeeWwWrY
nUdQD+MLsTlWs7GSAgk8YKzJAv3fmJufIDs8CyR09lurkOX0Ri8UMBa3P9DPG+sNGwNI2Pu8GF3v
qqokmA2lf5HrfmnLNT3uXfX8/u8paaEktijQG0MMMJkUX1vs4p/OYlR3K6DkKiCwpmBHvvw2KRJQ
9q52vKYC6Q0Q5zhC+ql8f/XzSg8SrXCrx9ra/big5ZfsdJj0s9HiK4UKwrFF3Im3OrStiT0IsViT
m7L9mMxTynqsc57in5iqtaa5lrq2aoEj9c4LdeX39Ws8blkBI+5RQEHYoB81r55TOsk9/o9UBJqW
rDJottAGf6UapE+e+XtLG4DL9F/wDbGwreVHQqvHIynigIyUWgJ73AeWZOmkeBoXzwF1MJmpxyY2
N8ReWXsgQy9M0PIxEyfcMQcMMFugxx4lNAvdXbtOAr37uom1dcenkkydmyvEDwGTILyheW/aw/Xa
dsVBmxygJQxCE4lOtXF7eKTCoUxQ3a6d+4KI0CrOpMDGmhvDsAxD9kaai0KdkxvSRvAkDKnMaGP4
uaB7yS8EcQLjq2wwlwU0cGZS/6N0EEQ4qMcRHBsJiQY/ijptlcmoIjoudFKjD+5vq1waikBxtdTZ
2Ye+ac3avk+HjgxqOo1qS/J2G33vdtyqV0wjYLazNXLm8ZRpbb1HPLWUDdp81pSlq7/pYKihDef2
5wsFeD4y4dV+hCmgoK8eiqSEX793Wattr4powRof20i6F+jKxYAR3zywWxTjQjJ2Tu4/Qp4KIcZa
auw9svLMHJxlXTY0ecTi
`protect end_protected

