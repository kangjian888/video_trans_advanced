

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SFpyA3WDAkH/h6gENMNzEC70V+GWX/AuJRjC9uuhJRzuSJx7LjCfMePfd14YnV5eJpUmzZ71W3kb
9tnOI6KXTg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FappTG7uNGFdZRwaHkH1xaFvi8BC2aKkPLd6PQ4xkTkeceiv05HkyC3+B1zcjatywH/Tgp5My5jL
RzYpXDHCiS+WLEnVqDpcElLtP6A/XLl3ajXqKvZhmMUVZsEI6d4wI3wE8drV6caY5dK99YnGiCxy
c/wD5JKxsx7IEFSu4qs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LRNAkwpKrud10Lp0Eq/NqP5B49JnJU8WkULh5UDIksixm1tOfz3iui+8sx8gHS1R0x2iJMsSndD1
7xzPuxZn4a1eVkZa4n4EghKA1iQCL4jIUagjOF/A226osIvTkxPBVZ56YpbMiMwMMgRLER5z0xet
LPBfedO96PfexivUiLv1asz99hmC5fi5UUap1VwJdrnsIHsC0bEW3N+9FFvOSldno8glOl5txGSe
hOwrv3syYadhoBtySSxq9fjTH5UTCT6nikZqZkVb5yhHF7eaz/U8CnmNnm4+vrB5n+GG7KIVkI6G
7PqaCstXyxVZ0I0FOvUz/cqAZvJcffVN4NdFGA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
u1B6Vk0Eso+5EvY7kmrlz1476LggIIsaO8lHvFGJ+HKHly0lYN/LsIll2vy/lYtCwxTSlrDsJgNk
NtsXioC5DfcQQ4kEDu1f339J7HYisXvM7Lhemt1gBNgHhAmdUioIYx0fpzcnzuhwqs4zH51jdAXH
PU3S8K0B/J5Gty8ttFjVJwRIoxIqhWdYqBDiUuGzr/SoWf0A03jx+7IJtD5tY/voAJ5g3LhC8YQt
AWy8nfe7i7XNQN6Y3WxajBwMrXsrAH821hCM6aadbQ0v9Rva24HNcIHmfKUDspzFekOzU9yGfpW0
fWulISNFKBsu0+/BoJRhSZ+oJMcibfGGrXXNCQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ufS+qjgKdn2oE3oh7EcYzivo13DkHjOXZdvg+7gUZzbjFQGb+M3QU6lNcH0LrOEXll22KbI2ohfG
TzYR0mnCNIzsPfjq3uw6taFIWJM74+oLYtSXEeuY6ANmuCGlqaVPg2smc7PFDAPdH082wsWirRmd
5thR9q4u83J5L0asBhDI9ZTgri+q5MwrlbJ05yQiFPUliJgl6amNWt26C09sTCAwIMPW69iBKeeW
4vt5DSJ6XyglFS9MDI6DvF+Cy8vysZSNzc8P7lm9H64JZqo1p7yTgGY0TjifISAPXC1fHwrwfQXY
BsZz6suWdJqjyzpfb60JVTQ+/k5D70Xj1MXLQA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TI2B3m1FrAeKaU6k30ykyHfDnWZXVLw3GYVFmPwE7PU79Tu2R5dzZ8wRPsdfoPSTye6ipaIAsPtr
CwCMHFOrInoC4tES+00nqn8BAlNtkgIns4JutCAsylfO0tbo1jdQM1s3ZfLRmzO8TErqp7qh34cJ
cDScSpPoqwYzQG0FgIs=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pRy8ixMxliZyP9cGiEmLhkLpE8BPUs0NUJLS9EUfKEgqPIYh3TC0iGkIkNMUl3FvP77e0IxaktFA
/jqS+a9b+rZb/lQQUSJMP1pPdZyeKNO5EYTlJkeq4M/QPt/jHeYrB9fa/fTRWFaLSO4suMctHSMB
vZbG6s1wo4stlPecixWiLDS8vMBqt9xY7MLA6d9rFSok/TUkwwve+vf4FZtQpUFEhypIh+/V1Yj2
bwgtk5lfZpX3tS8eSCYcpYqNluL129jpVqEYjJIDkcuxvvuRJPiKMpRwiViOhJULCVRU7pAOu9+4
kiLxod5VBhsHJGbgGwc1XTZvGawHjedADbu7Tg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 124208)
`protect data_block
4qLsf70AAADIqX1+vAIAACWLzurTVZw6+eOqL1c1/26coegfc2j6bsmpx/88TZaPphQaMDaH8Vjj
ztJcpJG4X0iWM1Nfev+CVCFG9yGrYU22vR99/4gcZ3A/sH//uQgyhguAgBbIhe64f+0B+sFog9L9
Ndv4F0iintPSkU19sIXXiiHX5MypMT6U/kJrpf2L2A2tMm24r62rpoTmouo9TuLDwXmPtOjOp4Tq
pbi5+0ufo3UU5HMeqsNrz1o3FhhDzJt5latXD3mdKznietj53uO6UswILmLM9HxNsYsIX+77eqtK
o1/KIvobfUHkNrpRG3YbaGa4Ngo8cCMDTlaA/FapmvfSLdSKzMO5njJGmf+OQEI4Xe8p9SR2oLCr
c/u5imioZnzMU46NTcPjMFROUxDh0tYzfTBhH4SasVOV/xrMzgNf4lMzbqtFkr8DdVvkZy0C01IX
HTyU2Ta4KHksZPzJgIWwNLmxlNIdt/YnkCJ/nRriCM3xZKRFMqHOU2ID+wnEC/k2ODjRZ1JW9bL8
QiEbliY0BiSN97jd0kvpNGLjwjx28sl8BWgg819n3KSdcNp/yAXxNC34Su0peWuqa7KKih2h27kW
Hp/o/B/I7ZwyPYGUcxLz+erftsOa33WHQBqK5drQ9IHFyodGSOIS+FNcebtJL7BckVqBK/CTnj3G
S0+YnmJ1JnV6gDDfyyVkkvqj0J5j/OVXiV8aMOVUupdG7GzNzMAGoJ0uJj7/v3ZaWAObqerIE3ap
+okiqEp4bv/LaAA6MMK+booOLm56T0ard0wFAB3/hPCQlvateFfCHwbGcq609Zp5k+ON+7F6TUD5
YfelFyCB9WJCYkJaRQCZ4nQwh4N3dH5OwWNEXSoS6QLvJ0nH4bCxrEws2JJ2z+XyWbHAySiwpQWU
xs5d4rHjpaO7d6e2EkguYFEwESqg7d1fdvD0xGFETgxyfd5eGBMZTtP2c/6WQanb+R1dVpRfqQsl
GVR8eu4fHYgxci1LKyppFPlP8zDD8oPkww3XcF7oRltqPm/4dTgTOkk/WQmAXhTR0pVVAXxrcCqk
VyMXasnrGZR8T0/f5mqXE9endV0hpazFxQ0P58/2I5cWBuoCzLrEIbQcnX2/5CqGeDJf89L0nbFJ
vcxYYs7dRBAThaoAPDCovqzNihQJYlb2ULLO138TxDnkU9DDJGoaYndHD23Xo86M+gEnzeRBA5qc
xV6tVokDHw4ezT9nDZwzgMRNqD0Ir8CQYQ28D67sONIYQOtXepJBDuM7XZ2nYfiA/5zgScCEK//t
d89HnMZgTqt4LI5YGgOtiWy0w8JMaTW8/f4I0Zbp6rKn4ind2C1bQtXk0CP4NaDTatKWrosxAxmX
WMFyGh6n0aY5q7v8zOMWc+1XFrYJwWlPOTMNnPjZyH4UZ/mTi4FbWdf9Ai/LGyYD28a745t8SFav
7NyIwtnDFK11z7HuplhPU8JpjkRvVROm42Q02XR0+1034pN7VlHxEYdfDi5CFqQDwnLJVMRiE3kx
GDcTKyDFxr+tImX4//fmC/z3aOwzRBEq5BanLeO8MrEVkzkEsvbWEYHszR6WQta7xzD9AVs8vlBk
jkpKytsEL75KKTTb/C+/IiN7WqTCP1+F+hggnPY7zJGqJ8pz+APgulOIc5K8X2TGOjnx0osA6zjV
QbPpt4GcKn7FBf2IhzJe+d9pwQcFGadoJL4XqTIW90dAxO9REnBabm3C3ly0NiAHZJqS90ky+Y0d
JHqKmUGocRg7be2nHzqT2o9vbH3OTaCL66u4fRjoTIQYhzMPwNxMcA80UMubvwOHw6bx+RgQmPyI
bg0RpNtCGVT+iW+WYS1BrtsCAOx8nAfxypbebCMJXTGniS18fqHzP1sHU3dqqRQCJkvIGMOkri3I
Sbxq2cPUm+9AofzDE5UDJZEdwczC/WWe2hs672gl+8vruoiBZeUVpgEQLfPY6LSMTuzubriNqKBN
xPUCV4Q5mfIJPAXqIRmVjSDbcruYGsITXEVGe80gfrh6OZi1yBjvC4d6NNcPEVyAJoUj8A3fQ9fH
LjGybL94rSeyjrVjZGoN2wjx84QPuTJJmDg+KyeXuDWyBeC4vHA5UtoGC4pTMJOCTrTB2mkZAC0M
RKm3pLYwcsPr7ylq7YUlVfuV8i3TKTojbBElwnXAnGnDMbjpHuw4sQmw8yK1IYUBIXHT9D1b2zi1
fTh5Y2x4Sm+KCu1GYPGINMIxLBsKYY9z481Q1HiYQcgnlcNy07wGIlqX5SjdItqGnNwSgFLmFgd4
2uetFegC7zDyhoIV/SaLeiGRVD6Q5ARIakD1ynOdNFcjeh2wtngdUEtqk9vn/1wwB9udNG4GN9Sd
patBQFVUbR/2ELKR4t7T4BZYKqTGQ/AR+EVs6Prtb1UiT1dEBDvsnjAr/n1zbUytasdaTwkOAwfF
hludB4GbCPQpAiQzLLYqUxvlaydZoUfVRRjTZbLveBA51EMU1oy6Qg2FaMY+aUQ8EL8cWpuW7DSS
nd20w4V+rkELltucSFJ6etO9EEV5WW+Ysytthldjt1sDkICfjnN/OVMSloLJutoppmXsUgIwy9Rd
JDOnOBgQX3tyRCGEiEhoyBRZj0T4bbOgl4fugQoOn1uD8GSF83tye/2wFMApVf+RvZZ9eTokOpDF
72EEZYv43RJ4n88/lZwDCifBuJarSHBnk7P9wCBvoWKvooiICpRGn8bnuGg9MiEetFJ5RLAIN5EK
ui3CgeT324/3VjiXlN4WQxo5TPbyCR/2+0OAshTZMlrdHUFCz1TFzfHVM9fxR8XfiudkOJA2Scgc
snYcIU7cguxJgd8UMDxBZ2lOqp+KcZD2RpgBFjl1mzHpN3P6g6rtISRfQjt7tsH0PAcAZExpUGeL
0QTIBbIweIGymmDyNVII0kISAV2XeuhsTJMqMMxKfDkxx+rk6yGSh1Q6/PLoRVJ9P8AXj3d7tYY8
9vfxWXy44yjM/+X7/nq2yoXAL3jv0qkbfpRfgex73AURP3+uR2Yfs2u5GFbFEd9Zm7RJuLDIwk4f
mEpuTcQ/v5RE7xGDvN8WiVD+slfCFNnrfWnFft7/weYerVNtdbuK0/q1idrPO3e6IezhGuYzZdM9
BGwNi9s9ZNEaDiPVBe57z2RAmasCqeSESfILlPowcgBHndL0lQBMGh4293huTpzGi0oYOLqTYVuZ
in1cY0c48pD5xLHfB0EY6iTybG3z/5BDzskFhxSaNZyTrHCNCYPIYMbVaL/iNqBBZ31/ZCpMJys5
gCRgx7qwOcLgtW2StKDQUXf4FOkSb7SHixTfBK8GA62hUAXIsuunvf2dmsVWT1FN/DwW7llQ5k3x
iyG+Utf5myP0N/F/sHOyDzivda4g0qrICwlJr2joWeMlhiruVh2sQFQxllJN3OerB5dBW4X3tsgs
JmkOs/SsFIbjeac3VDF6Kr77jYWaULpYaJxesFq+qcbKLhQZKpa4ASzV/eh5icf7tQT7mi5fehvT
hf8g0zI6FwYmkM5tUCVdtxGcqMtp5YoVZyiEdJWIbm3mYwWuOQ4LRn2uWZCADQpigcX9kRybauRn
DuN3mIOFG666nITB3cwSox3Ju9+qm3ePcU+U0WIMz1qiIkQdIWQKIzPBxP8YJm+Mn9RCR6YGhuhO
coJhahAxKNXmflD2UFdmH+DmoFDwcUgeG+SLngCnJ68B9ZSdz2KpI9yicjHEMOaa4gRbMo0JMkaI
5AML25Zc9xg8M6OocuLztdkO7cwV/fSLToxyOggybbBCsgOdMrMXHUeJv90f6io0CvDNeBO8iPuA
uVNJDzRV85U8M0HMfnjdJNI6D0gqUymh67VPQfUQbBYk2AQnL9YkytZrjso2Ibx333vNmxg3uMR7
10lNTzQVK7kfSvLWwfkZdqCMZVMg7uKI1pMZbX8naxAhwYsse/mOdLf+qdF5ur41TyIVN5PsXYQI
g+HpVqxv+Sr5shVxqHJnFN6XrIbtDk8ojDAKy9JviICEfjvB92BiEdrdlB6gnaPJDHPRdjwY0+7H
udkYIjAie1Au1Z5eJitDI37Mbu1epwYfDw4dXFG4FTohJpXFFt+mnaJhPjJJKpYY7UXVvEA7C/d4
1F6aFopbk/IBzOhnuWc2Wpsuc1fT/LCe0A/UWkxVo0zCjz1rT+qVRPOWWYKiu3FfanJhu5zRXmbF
S5Ql3IcvklKTUb1f68ljNakbLA/mYtleL2nt/d5kPsKaHAfd6gbUJCUNulJONbqO9uMmi3Icu0VC
Nf2OG/DV542iuYzQHYvItHpgBp4ORAmnJuEyptArf6bIRKsuTU2DrlvFF+BeuvXPR0jq+IqZ0ywS
YdDxa/VZSOvLWQJcW9h478dvnXjMfwQvjpFC0ylhMdHK2P6AxT+bkrI5eJdcdGQq2RceCJUkyUs9
ONYLdMsqJ07pBUp/c4+v12+guXnyxxXzPSoMsjicUTmP9lKqVOWfyb2MNUzbAo460tXymbLoaUKu
prXV18O3oVpUXhgQHnNGbokTIVEGg7i8Weigeu7nKuyWvGr7flWiEgPFlSsyu3+IVskqw9STqZQc
vdtKTVFgoeRRmMMIIa32Etb+fzrbUHW+8zxAc+KEijdLnnSSvzRqn/VURbVm3Z4cDuCg7SgHQI+/
45aqa4QcQmGQAGOK20ErMWLqxbhdqfBtJHgOZM6kTBlpIwUlJ5j4ZL3sm6GqMTqZU9lIObpGF5mg
7cDW8ebEgnzMQMKsScqcmAXSUWiuTB5Nc9PNFxqqNvDxDOX83XKQuNEsWJ3aDTqjSIzODnid/uxf
YB0nSoUdebT5VCmrDDaYfMWZ+tN92uyzB6uZWS/AWLzMgya7UyRBFHLROPO5wZ1hb33L2+VZj4QG
vmnz7jcb/mYpoK+cu0zgS38EedCufWIsc+l/OUDKvo17s9rtYNQSdCDTaD0O+yZGnaXSncIlrKg+
NMJEIDjfFsArcSU9LQPzx2ictkpiT2rrxEXX44hqlnN6PAoP6ywz053O7vQh/2DMgFteniPPkYqp
/bGjo8u00HoiC2VDJ2jvnY2uv4zsZBBeNdvJWT/4mo9ayrjR15GRU8sjrgrWU2XNo5RrVzFcJ7PF
aZs+4bpC9Zo+Gl7dixxXrpb2J5hXfmZr/PBlAqENWKDLkvaqeVCbpxZT80y52qHp1HrCHINMzAhA
qZzWLWJZJO7bVULdru2NDjV3ttCMLLAHHnWtS9gSK1VWKieuXDpEUMCZijKFDW7wqqJ04mKE3Hnk
9UPu5B/nQpwtoHLnXSXxGXuTdT7FNcE/RM42eP0+TA+RD8GXLio1Aw18KqBXdtYX929cgFnwivRC
7n7qwEy8TsjikIUgRUqDXXPvSYV1qJrwohcEhCX5Yn/z1D+yXBJ5V98cgBf3HJHTglOlJ4C8G/pt
q3/wiJFAbieIJmmtXWyDk5ZOoY+KXoX0ZkzbqzHqse8U05D66IAaf95mnsBnUezuzAf67AG4Bwkh
aMsg+z8r/gOCvx6R6MGKh0UrlqdUFVibr9KQGqaSpctybsXcY3r7ZlaO/tbAAYyV6btq6epu+G+O
GcF7kVP/I5bMntQP1IFt927oPvXsMNbOhQo1Nm/6rZv2UhcH6zpolVL/GstNr6zTSLeJQ4QS3Mxi
gn8wx+jlGu55VYdelEk6wCrQ7CmZORVvu8kp54X83dm+64ZI3wrR2HYPiVtoyUxnyKZkWfqNAxQE
7jMgzs8rFGLfkUIhk/QeFO3Y2z9veonm8r5LL3btAjPCpl3MPE3QCHdczTG6JNmpbfAzB9YObo0i
pC+oQ5x/sNoBG39orQja2q+PlnSdtMdiFNZSqsLs5gndhququyXHME/MceCwcUliNbHODBmJCg3D
jz91P+hbI42OF9+slryPQs3+g0RxAgKN7XdqHIp+K/JOF0aRdSZ6oxWNzcNV42R5wiIl0I/0hg9/
1/dyhHPH0o76cHCKWG9b+EA6PfwjwAb3nmEPRLO+EXdhKIv/m4tPdWjO1BTTEal50WD5GQ5UkOYG
yLCccgM3VBllf/VZNfCD+isCdX+/NhvczFOgyrt+Tie4KeJVw/sQMb/RfBHOSb8MPBwnZNHbxf1M
S/aEHSa3OzGb0klnEQHyaD62yM6biXSN5axP4HQhXyYba8x1+/ikMu2ag4rNMDIVgBWMlXT+CMbC
shwW/RMsmQ4QMaITMtKZD1O8pQduCzMyjnZ2V0TK2pxli4x/IaLr24ATvjxR6vvXKEclRF77l8Qa
h2lxWOUFRlkZxm/8wQj55hvy7XSiuO8H7JdJXBzVrCrDbrIfODuLLQKJj125lplLDcmLjEtixWl8
TSrSgExoE0MzE+8PlxtgStlmyHWEr7hziaOHpt2+BNvg2O96kA+fs5HoX9ralS/hk7vKCDC9fWmN
VtoklMlGYxRH+7t71kTBZq0BePAA9NBGpucR6NADTJMTDukxG3fiPMYJhQTECgLbr4B79YeA3ssc
0GuIe5U8OADT+QOkBkN1wFur8u6zdCpkOKBqNjmp+SEDJaZM9uLoWO/Qj0Ju+f9dzlQxUI4pq1Yp
D/MGsMez2wyu0IaFWMjxhOOYQWQrDTi0NMkyfFAVkRvvvSFhbhii1SYF686Aw+++IqOLTOKmcgXM
uBhga6elY50Qone8shwmcMvzObZMN3wyX6cq6Vuwf+veIBt4I3nDOmceiyqXtdamQDg8xKAccB4h
9htFlEAzCn5P14fPJ9xFzKKZu0gu8PFOQFfbouCiYQQe4NWDfbZMCE3s8inS+jHRH5DIgnM/Hj/T
1z4aqVtvIha9N/S3aW/YHTz/WmrtdfGJ5vYjXo47TsYbtFH6BmOGY8Ydyt/iOogzJiRNOTBU8PLP
RtncMOSQfGqw24VIql1p3WdxyXFuX1kkTkZ0LFTOMlc1GHjmW3PynkauVgXkabB9c6Noq5147IH3
gFtUG47BGmTuZGjdDCaMA0MQQqcd62eKDsHU0OFeHw84Qpv/Af08lH60T+5n/sco1Msjhgq72nT7
DqT+LlWeEuGu5W9bwP1dtQIo/CQoRe9AIgaDFqAnLRS23atBitL2IR/DzIVaudH67RWrieWBjEo7
hBF+Kqjy1vOrdBbMRb40qf5Ltse7thDf9vnzASrcAbUhszNtH1aLN0bhhAJj5XgKyrl1FFHphQ1J
3FCV5iY1e4MyKUU/xBV97NOPwWbC+fUgWvrFzbybHjC6uuXGfvQ7h5fbRJZ6Hi3M3q/6jKZWHWpu
5YRFJf3LMmK+yHWlnaulUUh7XUjeWhdVCeHl6QWQ3jmepKgVSLggTHdz8pE3BpEj8a/xrh6QCPQn
F77CWYt7Cp2sQ4JvX9lJk/pG3nXe+VCg8YgmuhDAKEBN5jJ6yiplayVS0bHTpmf5A3Rd0o9GdyYT
Y+JprX4UD4x/HE/nc3+qbHqiQ5A13VMGuvt4BCdy0ureE4Xxq44GMusSzt5jwDwzLUMuQ1LmDFCe
YejjiChtT4wi4+NqVJ4LaGUlV/fML9KXGZGzynBex7K6u9LIq7Reon02cRY35DPsdkXjE6bmCfT1
d/hUwBEgw4PzDxoANMis3vSngaSA+VVUIuk9JHGu1SmkJVUUfzKde3rzeIaulnSyFSog7KbO/HaI
fzdCdeYmslhnvq2nPojognvSOnBiUBni5HtB3dKEEI+whR2n9x54O2pj2E7dpUWiLo6NAAodK1RU
kUNGBDChz9EQXlpzO/j52qhdcOpsZJakr1xrTFcKSmfERrQ1pS1TQoD5zhnaZe+lMvqcFfkUg3uN
jnOGrhf317kDivU90ArozNVIEGQ0NSukcFthysua0/oo47THX7DN7VHvNrQJJr+/+64Bil/DAlk1
G4FeaEW719UlfF4EtXzPxwYzDvvgbntz+hqZ3NUPzuXNjf/6dXpuSiQ4w1LOpFeiEcoxpPcZABq/
RVKTvPNWOSxZqyTrRsBcyJF2gNoxKQYAi1QQO3UQTPdMzglatsvl3pARFjVrZeOWKZ1Jkx+nZYSe
MpDpxvKbXc6SUGNLjwdW8rn7Zqea5iV8i/h6036GHFnCO2a42mzJu/Tff6YjQIK5wdL2h739TB4G
JNsYIklJ1opPp1PlX9cn3K6fN9zES1ptjfy14yFyZ/ywda1vgaJ7peMNdAiRs/b8eQkP3qZja4UM
BN+lenb3QU/Gvb18PBI6Y/pFyojAj7vb/hGvbAMa2Qavi5iN1Jtg+OH4bZLsW9P0IoXfl3tTLClT
X4ev6mjpg/zcMIrAm+FyaShJungr9qSWF+uW0ndOiuU8XelHvbw+h0MWXhgZbbTi4uhTprBkxH1+
ekERaiORwllyf9e/S0VsHO5WAHPlwFzzPEl/8VhUf/rqdbN/XiutAN8vfHOmz4Pcc7WYCyfV3M9W
OAqmf9ZMAetf/wU7v5yrS+lv3V830pB1dJPqMbt1AwyeI5V+TScTruFQ/KOt/Y2tpcnP2WkUW43l
ongpspDuP0giGOvL6QTMx1E3OyoDPDLytH9GHPZW8U5IKhmgr3QjYkTalGDHF1mtKDViGPaY9SU0
5piHrRLPC1xoIwwUv/OgECWHrt7X/7k4WlOieyi7xY7mH11JpNp2UcHsliv/7Z6Y69gIAD0NWAyh
R2glifgu7C3x7oH4SWtz4Tp25RjSS9Tppfs50VIhDLGCsXGxQDKO0KbHLlmmR4ddqJrMBVeVHbja
Ir7aX7a9MIp1Nb33nPEGkNSfKxWzysOKqPM3kcIqp0Rdnpn0m+eV2ZeQhfbA5aL3IkLHTJytRtIx
VA/GBJNMNq1Uu5cTxdARbC6eAcBlltRNHtRaMi/mZYd+MzOPclA3OinQvfQArNdLsqvv2DrIVpNy
HMY0YnIrXu63Vcr0QYbLl7MwEWAF1VX7K9yTO7LuVGgsZE58JT2yRkLwadhdK3AHAWmkw3yEFA64
NWofdNgbZ2XGT7sUdcvqYbhioTTpGhThJOGTOpHUEOXGGeZrKdZ4LV569KfR51aqi71d6MR28iK1
tWLb3Qho3VueYyx6KIbevXv6OkrAnmGfzlRV3OMLOod0KQ1YG0DqdQ+Sb4KMPtVddx3KMZhG04nD
aUlj8Tr+K7kRJfhmXD0XtPjpRp6ykMK3UFY1CBsEOcbAh6FXGv+ysiojAourRNQ5SaMCXqxnAx3Z
h5BxIVmuSBx3jjAWApvmamNoT54yhTyJIqdScTeVliAfHwDB3GN0J1BG0s+iokLpbETSJZ0Q/ffc
qALIjhoOb62NsDS5j34kuq3uEnJgwJ51CiNA3WcxkkYqr9W7DizH9oKeLC7pBCxrx25lQAVD17FK
7Fi5qgMTTa9el4NjMB/lGK+lnnU0sRcF7ntWpceUnSHiNaz9+LuZQpCElk9zm2Vg3BESwNlBDUTs
q2ry1oUJpNVd6PmgTjD0es5gQ5RDp4z13WapdAZBAEMmW/fqbhVfpNGMcsaljj3mdVrA6Lrj+RiR
A4v9V6IXEEmYDxMAXZwQzqXD0jswoomcXTSOtlyR8OYnmuMlSZXSYD7RN7JOu+JIspTKEc6e15N6
hll7V4e8VKvAFlcgVaSmWQtuxmLlbzuQj65fEtUQgdn9Gf8s4K0KuUBq2nsHV5T4B4tOZNQUjyXW
1MyMkCAzJGXJ0pWcAjSON7DG/j0UDQoKzzAKiSf9UeNvH0Y5mHws8MzANw1TNo0P4m0H2Jzgzjve
6lxs5JGYilf2OcSAlozjbxc2gLkQURRY+GIxqkA2WftTHBmcKfKJZXAE6PlkD8qkMahJi7qsGdCx
zz0NirfjBoatkILUwbiJHDBgjTvX8OAzrq7unBTbh+tXEz5G3HBSclkA82682xL5+/hNmTQJk1SA
YHQ7HcH8BmLFtmphLU/s4jx1FhAqJdgIBuAcapL6Et8nx1qw63YnlwkLx3FBPAaZf6qpTWRbDuBy
F4LY2SRef3sn6cDe1INOQ6WuyTp8r94lKH1v4tl81KrtI27MZroihesP2vF6eUK89Mto326Zj1am
gVLr4ypv2/GWoVTILp5ejhnrKsHgdSZcRDpCwdJC3ZOU8LRZ1DsXhdpp9Ghq1kfd5ao2YWIKg3Vx
5ujn0LDemoituPZYe4o/P/KXIJzERlbxCE1nsnRvmYDfr+mcA+8o6xsOXazNBzMk3EaD2Clx3Yuc
1ShVUnKxOqIJCSBegZMKE9ZCHUaTYDGZE3upyvlT7lPKc6c83VdSB6OE/JBulf52V0CpICN8s4xv
ODRlzu1ikrQF+PSoTixVziXAS2XcpmNmO1WUCwnSRVZbjqylLffd1U+1G1eQ8ybAwesvG9EmvET5
S4qeg8qQLaXquUW6p1P53UOdoLqxs3DghhAHa6COEpFtCmMYdvZMnxNGAteynZAjTEMdEN910xd3
Nlb2fyNAry+JTRVszEZJ3I8nLOjKzWryu4Kh64fu7LCJCpZIOcJnSgOIjwMuM+/ZQ3iNeUsP9kcP
ymOa2LrHaTngznQ5jIIF+F4gnE12e8jUJuIlbnr39s7uLRGehpya0VNW6j+n8btNkayBgJUv/nYX
PjT7o6KLTv+6AI1HFhZp9/pzPCqRhKSskU6vgS8qhfh58KMMqsDrQghrtBHzE6xYnjr676yHVoiZ
kej+C7VDqhZwlPazXKO6rIIEYdNCdpJzc/S/CD9FMl9BtEI4lmlit3PXZRhbjAVTcXuNQwmOSm34
tHXj2hn3KWuFnrDtYBJG+XDjMy8sCA3238fEvyYB30zZZbqBWPOb649Ok6PneQAlBmfO/mpwIxRZ
0k6u4AUaW6VfhJT5MyewrUBbSzwFPzptbcnyBt5O+OpDyUkSmGwd+jPI6h8R+/+O0CdGDY6/C0+4
L5nxfFzNdPigRTY7WdZD9psxVhWWFuBvE6tPbMht+GiFXaSWhK02awyJxUb4zlfG1FlzqTQZDiX8
or+Zz0fHj+1DXDGvtD60PrOACWA6Or3elsBFnb+y8oPrE4smCFwWYWzj9WU9vpCjPknzJ2juFi/V
kh4XGkdKTYsXPxxhxjU70LLYhNB6wrtc5ivEFJw5CbNVENSmpzRx6p6kARE2kM1LY8mdFBbB8Ewi
9KdRGK+YxhW0Hk5Iw9VBC6xLeNnMpPVkyxKCP1S2QuoSAcmJmWi2bWbAkNTonEdrGQeGdbilVs9w
rfXAHpbncru+UTVHSIMLsOFQpKrcpUKQITOwPg7nEaqHbZxE7p3JJliftEYqg1N62zvVwFCng9aT
PmUm4lu6ODNnomlU9Zshv5TqIi0N1KEgBaRqypEnyEOcdwsokgtA7VxjKBLHeY9gnjwtNigs7Cny
zOgMwKsY+vB4bNggvVpSKZUe0Mc4xr6NKL3hbre7o6WMadEPTSA0FVAZaN2LIkIJaSDHDJyYcfKq
hxKysOoPnfl3wuA+lndN6vrxfy8B4DlGMJX+V4arfkFxCaHm/EBPH4JxETOE/sWkWxi5I+euJKu1
vWrg1Z/ucjsF7LKRAkd6BbIZdY2RpBGX0O0378y919WQIT3kMB66pF0ATbj16LDG4ANVgg5Zs1dX
S6NHhe3dpSyQrXX2im0i57KdvzP2G7/pWj2oasa/5z5Vloyh9BtlVhr5mghp6Pvs0xb+xeazwXcU
o5iXwaHn9Qx9BPkd1u7I2eK6WceyUf3Zww7IvRxqta57U6jF57alwa4lJ8oXPyJ/ML3TTUDmWN5U
NTLLyeSMwllydkWstAIvH+NuOEuqnGUtwrS2R6vAUQbdgf/S32KU2suHYNLbsM1CLYUbL0veT6Iw
cIS6b2ypZGbJ02oc3GeKbzGSK9MxSPK4adE5ydom54S0mognbBraB6YIb2actjEot/gugc+7PYYx
jCF99EWvaOk9xyzlG6A+6KbSxN3vMypXnMy5aeqpOYbqebd4Ybck7FnXdCqTt6Fb1Yst4WUWZJyX
eW/VPB6Me9fvOymNxFTOgnYUNAbGZ0NQgUt/564z0OZ/0w0oEfv1tauE3lipr8p5U465teChMjht
zaEFFDIQPqjuqAuuh2rNW8XhENw4mLuRFDrKXKcjBGz9UWF8UEHAN+WiY1xVYMsDPX+7Z99Af01S
NWXrqMp+l9NRYUHv/ZIewLRb12OxojQ4TXh4EC6/X7pOpzNLtElQ/HxS7cIcK31BiBv5JeGBBO5I
+9YSVbm/1Tbe1NGqRXiToDEd1v7za4piRW0JGjk9eRfRiGoIauAnwPhuWsIrZmJHVo3HHcelVvin
Sln5gLbAEjhhc3ZNzNPJkADSXQEcbI0bO3DozLlxNaWaIwBwao4gs7Q7K9FeIEXacEOsg2CqjB5j
2mkQlSrdAi5rMeLAheUEgdSvCt+wFOl/yXuNlPSUwBUXOK/5UMj+eKQ8RasDAlVQwulfVrIEHIjW
dXpVGRfiGUaug12rJ7TuwdomOew3IUQmIFXyp+fbIVHnixmD8SHGGqV1rkYxR5p8QbUkm0dkMA4+
zapstqplssqMvQzUJkhWXQp0MObrGuEZ0q91Fxnkac9SIwiw6/iOEDR/OgN2iA/h9A34ainE6RlI
4NPfj1mFk4T3QzX2d/3GxEDEij59h5OkcFkttP0BY1z+amcf7Y5fiiPlrNAs8HEO5l8LQnXcU+7y
XSCiXHEScBALe+imAyhg0e25tYVrzGAH9dRILJKGSCRL+E/axDobprUuFTh+H2hd+4IdjHSKyQJK
0IsI/YUT6Kjt0/StUa0oVJb1BqRWh9DCnHjMBoQWkNgIJ3Yzub6FYHQGWplnO/VpU17BRytRKSFJ
2KQbvWyuxclGh8KDF3Q3HtTDoGK2U/WPnH/CFH80DIMakF7CGJNi9VOvDceYmn795EQCZebWlVQf
q5xs/cHDz/qU9VF/vTE6//ULOX43w8Mf3V+sNDAYW6/D9h2+RFawC0GhNz9WzfQXyJ7WVbAUeNNA
lQeJ2j5cTMUUa4GxX5vTsk3fpMvi9zkGgjqkwerpVTJGq5Ne/nZ4W+/tg0vYRDM1Yqa6Yj2gwwdc
YJyiFmNTRDMjb+6jybuXmgJf2J28E3jBB0PWGPFVcj+yW2EI0z6FmpIM1s55C3PER98vKE2XqyL4
TCIscL/fAFtGK7tT0yzaC+vdBWADA1CjwSs+Z6r0oftlOxKLPiFv67l5vkBWyyOMVtAOBHHUgNUm
deo6b61566gNEv7C1bZwT85/SHry/47nmWG/5EIlL4Zmz4MkWjlWzcBnNU4EuzU30Or66c/cP174
tDBV6iBpbiMupVibFbZ8+HcA/8vqgo5DFhCk8wSWOxB9Cl/IE3Vsrv2WMk8hFC0Im51f1JuegrIb
iRgXGscFy6qIN+XeZ/ZHFJ9n/TxcIC/dLBc3OGguJGYKP+os2TeA9aRfBZooTCa1852i7aaG/GsQ
ap4K3NSFbXbLL9QFLGJH3yBnkhMk4FCL3T6XNS+oihtjUTnpTEibB17vqeHC0PsgnOzmBfCBUTgw
iaYBJ/HMZpgCJ5PDYeA9ypEBJL7rThaveP5gINjZWnRQbhEa4boVpQoiIyHJ7IHAw1yXCXNGy8WH
HiUxHwB2B5973HSXj7VR9qVtLRCDHZqdMyyFUnRZ0yUYVGSb9mIEIlGhvgzQK73dlVsdpIXLddZE
1sGI0IahoUCJA/YQ4X465FsqIUDAcDJRKWphe1+P49YCTxH9h/Osc89g02XXG/FPaCDIdWzm281n
zDFjkVWBgWVPEMsIM2O2sPQFbp+HokvqJRHdgM0FFIzZKXoJpAuc2/FQBgj2gFZCbEQRDvlNIS3i
dROAdiO5BVRSObrpbenTlWNeMVvsz1xLa6vmeSD+X/aq7ajnZDiHHD0X2PvanagxOhkzgU6wG1Mj
Lv/wSPoMcCp++02PKrWrfD7ZamEWw/IEH9Zz7bc4+fsFukrfnagU27UgSbRUJ4FSy0Hu9yXUTil5
9lPe/YEow9vI8gv73IFrjsOogXFKHqRqRKAaxTJtjeveUwJc+uLKhcbvBMKw0a6DDhf9uPsGJIfV
ZNy4AOqwvPnwfND2ERbralJI64wUVmYwbN6QlJdpj/FgIWo+TS6YPuLmeJJRQRjf8OKtFl9Nh2vq
xc5WxQtBKWvJsFjqZJzgdzqLZ6KxZBq9hy+8N2Vfc72yErD85k34FOGvzqGcLqsdGle5NXBd9o73
TGM8tGTeWZDz9A6kST20k8r15SkvHawJoa7a/M+O9NWY5Q66WnHE/YZFnTgnF4Y2GgHOMwhzKq+T
1kkTnfMcdiEv3kBCP/F35JxRr5YcjhHnSaoeNn9TymBydwwoXzvbbjfYccGIvLloFQ/C4G16kPkq
idpqJGSWl9DdA41QGLZf1TTn1okS9Cc/8FzKaMIgE1rcTLB/9c3BCmjucl65cDr5s4jFyc/wfyxQ
2YyamGhAj9YBGMflbFWeRjvLKCcOgJaA/O2CqyqHyDA/E6ci87kibOGeEPbTKzPN5xLTx4RmPfPf
q3c/VYo0sH4unDpuDJE7/kBBBe9IvVx6cCcLznpv5Rd2RG+JhW6b6/ILfrv7igk8eled8zEwFHIS
Uc1U1VTBcLROu8+ZuTLzn2lLPif5ImCJkZ9Vq3+F1x4QnvlyQRz6opchdzfk8RKfVdZYEfNAFss6
K8PwzrokhtmnTtJztxfJJigtribGU1j1L/0V0yta7QDzG+wAke71NfGsweS19ggyzUBbg3K9ilo8
Hpmg+8tuPU8heu9dxUaV/Ulifuw7zLjyZyKUrvdd55wb4WR6Lb3p6LefIBpiY4P8GCgp8purwoZh
2Fas3y9U67JBujAk7O0voqOs+J0QYM2WLOZXxvQQ/w0IzajlYN0/13QYZFOHKaPnZqi74G5mvXrG
c1ZwGbChau12G3l0HO31iB3SQ2q/NwjFk74Ji8Dx/UXXfY1EOK6Z5dLwOKEc1RYyCvRODjzW123X
5wZisDNpzFMX4X47vzCk+KkJw+u9ZOnDYMPxerbGWE8PpQm4rco7qFQg3bNwz7KVGTq66P6wE6At
92uLhToHu1YhMRyGGRtQLJ+TFLZMGfFtlYhuYz5m5ghZr7Ghchy+GYK3bp1XZaU/kpjVyP/Sdwax
Nhh/3T/a1QEKLrrJIlg3cf2kFJ9t8MhiWnTtU+mfOQ2d3f2tRMN87X/6rl22PsFVV0A7o6bHgAkA
zPwCa/lvsK6Pdv1A7aFCUZbMlhmKnaOpXP3dB7A4Dgpwgj9YerTc80KwMRUAt2KJXiQLn99USZR4
2yzEebUH9Q+FSvRthjcWPHU7Odydj7mneTGgkQG2ieD5p6iJVlG8mWmmNswvU3U7e5OoPdiIGKAs
CEFpPfVbA8srnff0fUWeSwqF5nPEyOI92k1kcuqmgG7SngbmFL7ebLmO2GtG6lVPTmiFc263t08o
CQ5WZnztRwAGfsJrQytqD4ZxIolcEG+sq21bLKCU7qC+Car6ulWHu7/8eV2zu95eHg5QX3nRFVaJ
zkJZC0Jk7TdMYiQz4V3cPRryen79h/EsF00Wn0WgyOfT1xLDG2WVaB/cOYoqAqPB4JezD915Xrum
OsdO/ayH07IpJjumkTdSS0gNOYsOXAOsbeSor4cjgBOA0fDKDWax+6qYD5SQ+avVkzi6M6uQSs+U
vzQbB7gXVYSV+1CgVGmhtPmZQfqkdTFzUiJuOxE2zL9hbXdgeHRVlXo8Soz7i9wqyYYhge/QeiS4
/AV/kmsdwyejjUbPoMiAR3phaE8YPr7Sjoqi8hWtFGHpdcnpYB2GnuV4j8fyFwFdEeX2N0L3G4Y4
2UR3nd4PhLIcI9XLSjr/kKFTh6laBn4huAgvKizjtAVbvgJ3dlikm/I+JlD6DyNfhDl/3e8E+c6Y
Y5wmclBZnOOsacBvsS0iEtX1uIySdcqWAhieoCxAOB/wf+pgL6LKu+ag6EzHCU0jYUMYOsckay9f
YL9BVib0/kv0EAm0E+7kcEMO9vqJ3gW0Kv65ewKigQyuXlJXUiKLB8XGO1LYZ/QhocjHaFMSfoG9
ERAEmXc5WzdV+3GwVgiI8rxt11d7Dyz6QxGfEJRaoz3MYfzn14Z5CBmgwVkReQ3cPoCR7jaE3oC2
YeiCMbz6pet5QkoO/wHtMWEijxox1aijI/qJ312a3dkkNkjA8vuImRP4DAZWuNk5/SGkVX8YoG3x
Yncjx5PT8aIYPXgw60Zd/akiHkmcN2edwQTbeg8DFi20KcjNo+Y+ydXbeH65xD2QKataslkarPyf
ybM5C7yTRN7ORNnaFVfiJLpln13yOIFAi94lwFeDQfr4/Q9xGBnfMMoeDkjjxXFDvB67eHCt61PR
+ABAE7k31QH2h48XnVtTue1tXFDBqc+EZon+TYPTDOXN7gIbxlSlB6ocH9qkInBBk427W+5bd8+/
pc1Q6qV6ONwQDzB2W5+w3sSeJKQ7Agedea6c6QXu+tsIpnFAL/VWnatpFKM3E6EbPfsOMIEWowP1
7E+QRGfTQ2vSwbheUdE3Mw2F5agqZBBaZdag3YuUg1p91d4oStmCIbizZJ6ZSIwu5046/mvkfTOf
QNf2CgVCbj63dQyu0tyh2d/2BiBCfKDBrCTNvva7SqfxqAn1wp7J16coXFVzlgZ+At8xxGCgPNoX
OFPWWQNsc+0JoCF7R4giekUjU7yl5G5ziZ+MEeAkmDhOs0WgjETkskAtO7s2xayAi/QgoMMFxL7M
B49QioOJxi4sQ3QPZHCbHuTsFeLuIShaFVaJYrmbtEaQ/HLR5ZDT3k3nX/X/n0UoNdq7sFbEjise
IAQm8f7fpUXLWwhpVMyqSRGphdKtlPkMIVeBkxbhlWeHRo7YEB3OS/9Y0AOnVlU1tg5N5ORkOG99
luJJgUcEj00UQw1PCiciF354xN1T8aL56uCqiLOS5LeAjTngTtefUktK65m8HOP75hl0iumB9MUV
+cUuIGNZOU1RGI0bM+cAeSW9xAW6bb1C7j+UR0A+WZMFy9/6/DIyDA+fi1USmMJAwYal6M2XRs6V
GX7S2/KuWInn089QAvqwq1vWj0Dp9gXoajIyCWdrV6995kXRm0/DDlP4EKb9oCkyYl4olTQs3iUL
yLvjkwe6fmBDa9j4jG3JptdTHeWfuKyz1k0NEX0shW90TePxdbGd2te95NMI6Z9CQXLPjJ0r9HwX
kGkdWgK0bQUstACKewjinkz2Wp5LvgGTiC8w2K07Yk12kiWktwcaCExK4reD7XxkHKMoRdxhgo/j
lXAkyKfFh8INX9xrQwt7oo6DFX/QmwupJ4EpV6pIde5y1ZJQmqcmSxc4/h9q+MOBPvO1fbMnciZx
3OJC+LgsqYAXiWf9ghpTUiHk43BG2vtmSvfTZuCGwZQQmDqgAiouJZEGi4nAiBsql1bt2o2zGWeF
mYbQ3GQt441mkHSbvd56CyRYQs42NYzearyOc39gmQuD6crMQf47wGk89zsBB7AYXiGkMgxgJL8/
uNH8Z9227D15tqgWgOobc41Aj8QkutXsJ0K6DkqchGw3WO/Gz8WDEB4rZ0DAiKwgvPttpCq6f2r7
lD8+I1gOy0LNZaJtFl1zuVVSCF0MbL7/48EfeHih2iQQHMEqRop0no17KioaCdtvsxOcmkadL/R7
J0sntIrFkMiuGJbRfLDhprgwoo9kANbioBUlGk39VpVfdtbBt53dZODHAsEjyieVgv5UoPOFIRD/
bhT+Pu/nbth6EvEprq33Fl1/Kcg7SUt0Lj9I5ruMKVvC3KwAg4gj0hU10zR6Exlgwyl9bcnTQwnS
bIOieeBVMae9mwj9c2APWV4n+OYEZWr14Y7F+8oCsotD78CdpFjkYxyN1nBhlPRHJhjyAyzbWwd1
ApyHWWd7MH5Op01tAv723F/I2R2OFqj45xIZXG4IyVnlzo21MVIjNlD6RBiBNbGobXtKanlgZELa
NrBTjlLWBmqczngrdEfa2+u7J3rtEBozauBa4thPLOLb7hRjT+9NwnD59o0MUAL6LXG/O0c+i5Gt
gUHugQMwsaSVphh72IIaj4zLadjRnm2x648G/jiBa8+R1q3Ch14d9QtfWqnWXIUn10e3pe0eadN2
yVbYCIPS80wZr5D51wUUnuqAzwWF7emKge6VbIte9SbdwCcnUZJDcjE3CctLttQMv/EF7ghSzBfB
durms8uxUmfwioKt/wPUFYwUGbO1ZakJy6YVpx0icJyvquywcyEiCt8BTSUe7sLRqtjIPMibSx1N
ccbLkwrT+ZDLeqNafWkUP+HjfWKTRo4Z/R5NpN+eKPrlyCAiafb8eGSDgrkt3aq35u8lB1LC8fIN
mjSmMWgvKJUYiNPNU2Rwj4geXkLkV4y8kbCEE9XyhynFCIfWaA+Iqp+gUYar8U5FwzKdskzUzSp0
ZbWVziM66xWxqZgQi3Vdh6jabSkwMNKVnfpuxVwp1kt071KLJhVDFIqSw46X91iDav3gkCY5FQa6
2DVfje9f7OMqEDiEElSMZxjyx0/Zdj2WNjxz+aAO+TiJ01c3ps7zSLoMmxe54tYU6hjVRfVeeK3W
h6ojCehI7Hx9HYNj58XQqhY9EW2urHbTxrgONFBwf7mb+y20U2hXM2/y685S2ykUY37wuQ4R+v86
vTimD9bQEu2AR40r0f1a/tY4KfuZIZdbEylctM0eMc8+78HOoD5umWkkDCv8qypC4klILBidqVBE
hG036mFCMJ8DYTR7W1bRE40ZEoCE4bTWU9MJMbdhKqWkm4OKvVS6FOOmWgmCDg+7FpfxEn5c6IjQ
nBnkBu8BrgVNnofsqDPlwBVahtc4U7K7DUQ3aUGFMEPgQaFsD+2VveYamqJ6xQ/0AFtgjOIw97Co
6iYrKOa6wQ9ELVq3n/TAwpV6t0E5khmVLVCy85Xo3xXi0i1H3XlutEzu248+p1qlWAuy9k169W/m
1B8u3/mDh+EXBuJv13Cfqc5bjxsRTRf9BkxGegfmZbf+/pOETgUmEJVsJ3ln1sqbc04h2c4CIu1m
1APF5VqxJhDabsINM2gsGR65TU9C2rE7n8ZqmaxOCj9gBHrw7EFlgjLjrjvMfp+ALa9EuOl2ieFM
LWy8SlI/R5lIoS8+lpKWUlr0FvwK3BeavOM/h8R298rDfBLk4Np38Ro6VLNC7QZq3SUkgCHY9lJ2
8ytxcy/N4H0wuTc6pIAZKuN/POFDCClfifo1It3wI8eIy2wi5rGACh6FTcGSQf1Gd0/uxQPFZ1Wj
BefyDUq4PtjwDqVNMIxNdpMKC3spScSmFeSN5+aMIOaodLWMe5YfYrhTxABFElZ2sxi3TL038in1
69SJ3jNspQtcsI6pShPHZMBr74GqEjOeFzZaQ11TfHGFxH7HoyJaM/pbb0UI3fICbgLDI1lsi59G
gSP39yYAeEoBd0LyTIb5SALVrd6FO6bvl8qEHXsr0D3fzs2Fnjy62o1Z0Qkd+mgxjS218gDAJ3si
WyC9/uPoscaiQ0Y8Tz1iexOoxgMOWbQNDbURk6WJ+qFLthMx+J3Bi8k3PkGOJ/38J8JIebn6lQwi
jC2CrL9Hnk6XPZNPFMkYnmVwvmPotXGEs5SJHijtM9f83O3oWZCHXquIlaSs0SlmaMiq9zv881IQ
Uq0DrTpjUmZVYQOTqlYFq1EMYl4kHasX1pASuz3UnLEnq/7DCLWlv+UoiFmPogv3qQ/haxIDIJ1z
g/lD2gmJnvamu9ShLrtCp/g96ESIWpx1Z5l+Klxrm3mLlIEe5QjVWgWwRSRVakXsOpTpoAZVDSjn
jb0zTCq0zbADNDrwpEqP33UKKQZmr4EOERhmbYwWT9C9mvqAt3QtIYKab8EnpZmkI1GTJz7bS39o
yEMavMlXioJWRIJthsdlPknaHIF7jaVcsy63uum8Iq2VFiWZnW+PZG+MJ4eypOId99Z4XUOc6Zx3
vHPTYzFMmwGdN/ulg38ad/9OVTTXR3X3HdKBzFCLFSLiw50ln2x5azBqyIWBCBdNiuxR5Xk7CEmS
Puepl4N0w9+vSAggTYpfISJzKHucU6P/KAww1UVKaGl3okAKebdY9ghyxQGy0aGphF82ozh4Pb5+
82wvABFcy8QoHOz0ponK2nCt3jlXS8rhphbhitESPY7ZlYpipj4ILbGUg6Oct1MWOovwdk9ZrwhH
zIi+rfp1PHCcchRokBVFiDETOyO5W7cGqoReXD52wcvV0CEVqFNqZp88sNMsIcZFZqeKTM53l5Dg
U/fj0mRpPi3S7ik5/GuXV5N3Eu17w/dOR09ZrN+5r6DxKtz6oW2LR8MxqRAVxWyzwDypSTrlprFw
mLg8LXySq0ct5nZvYCErASx9FODhhJ/Rcv6HiSY/RBkPlvU/CulIgbyIXXowjagB9O/e9UTl7nqd
Tn3G8jm6FZ+0slFzhaidP6BkFERkeNBfY2X4UHvRaP88ydV8n/izY+9dcG41Cltr3JQZmDqnj/Bo
ooJ86ENjsRNtk0G4qc5e11VByBGAfEfJk/80D5wZOKfcN5qseed3nsBtUHLfRSE4c8W4Gztqifo+
fjX0Fm6eSsWLZ98kYQN6p2lu3Y53YcDT2Q2K017Fu6DsM0FuDsm7uOdvg/NH1sueAssvZ3YAM7R7
fVLt7Lb/YIdFZafqjVFKRt+NDTcq84ftwmvZqD+8fQrv22IIACkZ8187U4dsvUbBGm8jCVhr2ALl
y8QeK1FZk/dhX3ZqSlJ11evyKjDafUc0uu5eAaS0JH0j9L9607b6BDqBRXHeUhfSISGW/Hi1cUAJ
NZZU2OuZSaZTWe832cEygKlf6QVSKTnaHYYeNosyWU3xiFoUPQ76qPSmFqTtoW4dNlTyLwwTYH23
VZNIQC3HMMa9sMkYtDdQ3Jqh6O7/ElB2MwiG4lOMRq4BrW0CVi+55ekWL1BK1dsqBjBM3VbvghSA
0ju8zTa6FnD11bavdsnDZD42NyhYSpAuVeJzHQc3XZxCb+THG2XoZe/kxxQHdUqLG2ZjHBmFYDjy
7Ek3qoVcLJMGQVw2sDjL4crA/ZUGZ7C3PCKKJVXK4+HtYbvA/d6dy3fTwggnSO1aJ/BHZpXL7TRu
4N1fA5WKD4LvpHHdvWtR0k+Xe+btw0TOAtbVE0L0GTXIMb8ZFYdrJZBV+iqgO/GecBUSKmYpCTgO
astzh3QBXzxkJ+Vgurr8x3KT9kvoHN8d7gx+0FV0usla4Dk3pmeLtbYmuggVrIkXWHNYqHeRrR57
1qPZJJ7K+lnsC3cIMHUlaGwT1UwNnyd+0C89AmXvSsVn333EVtDpuf/6QL0vMON7eJKS799XyVtg
iMOcO8tldJKMAsrUFvfwhpFTKeGvebl8OTrXy/fC7BjxKmCZQr68OQQ184I46dSXfJT8R1vfNh+1
t8j7qgqHNXZbMMUwJOLbOGEgFZumatIc+E9JDb5xIp35kzn/F4FnJj9Nvzb6YTlYHALr9Z0zPUTZ
ML1xOuny5Mz1wBX1Ur7uhn0WvXm1ZCZTkTA1OskdCOIRA55vn5RnbctK4op/UvdaLCWt+5Q6pYw2
WWX6dIdP8bw8JnlSsFT/fhUxckMlxoFEeQBfUtIuwRSqMM4eLHUTgE1rlgPwX1yDtdLrtXNFzZur
EPxov6yYkyU0MI42fERG/R2xlXR/KvPHyNYMUJgaQzKe9gnRhzF8Aw8I0yDicQF4T1skt/exdZzj
a29FuKZuiddlS34u0W8SzxLvoPuAXKcarC6elUlFZrmu4fsn3YXGQYXvoaotl1/OrC6g0l6VOoc1
QH3Z3w5a8/Tru9Tga1EDd5ou5X+3XhXf8N06F+7vvJNU1yy+pkCamJYvTluigC2vPcbLuubS8oZT
pyyiAR+3G5zPqVr3XrwtddbCfB+XJpRVtUab53hTlr3SVG99O3wRwzg3rWufAamRPFYCdgt4lqGy
LCwbEAHC30hnt67tzGcJrPtOqJ8bC1fkZsWoeR/xi7pSJA+26HHNb2dR0LIaFaqN6S0gcqyLYRVO
9aE9bW1wlxT21S+D4I19jQQzWtMGDuXgQFu55c6CUKAmoBxTuzsHjrX57WI5tu6BPMYlq4wymOhC
t4jb80Uw4JJ5LHzBTrAU8np4C2DXtpnZ2P4WXa4TY4/m3xuJMXVEC38i8MnbaODijuyhXiDkqXcY
IsoM80Jxrme70Qe6CScmpGbDbw3EPAfEOLW38DjhHwa5+dP1pnYPGSnVzjjt99LrURGtLCkraAsm
I6RZrVVRu0QK3W/uNszMJEayyr1JvjTP3+aTNxtS4Aiio6/s3L0QlES7TMUKoUSUTOu6xAfFMyWp
pbNsfYC+NaXHXcC49Nr2+4CESQNQPWbz/2LCGJKXR5r8Do9TgNJcxQf6VN49vwbMs5n3bqlI+mZq
v9eZSkHMpmIfofty31Xb4CBmK86Pme17zodLmHWINtENY07zFimQrc17W7mSh0auA6Ar+jn5BsHI
HrVyRJQFriCZTdW4FP+RmNmg1SC6nMYbvIUnj27lc3W380ctl6jT/IliZG69+jsDBZo9NJyXe5ua
xdYbFrD+Dr5zSIK0xUHn6VuoNVRjD51TSOtQl8m+zA3t5D+Z+1UpYTp2Y8ImplSyZ3EIqcYv6sm3
i5pVauuexeIfe4iiWQiztNOIhHAzOdyEYFFfc/tvRXTGIImAsK7qvZAKgNX5ruK493Ap6Ec2IOOI
uMzMQ0X8L4/aYENuBmivVsaaoAsGHsEDAq0kWJzVb4gtZ6Y7u4kWniv2xmvqNz9lKePohtgY6KPZ
cpv5WXXrRMmSYPuI+9bwGT4Er5sdMzEw6RnJHt8hkpILeeLlZViIFwr8e73XaiSuOuJzKv8fpDc1
mhivMQDJM7ttoFEHtmnx2wYi6LSIIRa0Wb7sbHH4p6vD67ZZKp7NxF3AaLFzO0MXCKT7I2Oi9Gcx
ILEjsp0HQAGLnTCxX3pv+sMJOh4OLPtq2mnW6ou2rYEzsrThbb3DaMvo1NT2P9L6R4W/qr6YBBw4
SzDbbw8Pz2fpxCbRn02ot4Mm5VXVjfnf8TGqQCduX38Id53FFvw2Ee4KKXORj8mC/svDIeZxulw4
SXa/n2pVv/uukcWYlJ7m8lHw5rtukNmvXG3YeVw5+oeq7gj5JDX8c6pvx4HSACCO70Mf29KA0Xsw
HTBsSlQy3o18fOSrlZOkYVV27orJCkLdKDLp0fxxzwqgriyz7CncTGHsVEGlEUhJ5daHwhJizoo0
dEcJjtWy/Urh56n1QWUbMYX/nhSHzMjo8EhYLwfDbDY2dGECj2WPV3GZLvKflSfeQQmOKwKy8fox
XLdIQJkg2pWbdqjJ6aak8zEJX/0I8cxJKfLD1wi9Y2fjXtIr6Em23QyJ9sVTQzYwM+nTWXbhE1fE
Zk5Kfd2jzRVRO0cGCmHSIWtlVFD5hConbV8KMpouYumPthV28lQxCa1Sv3bl3IFY6+BFYKv29vXO
cl5M2TPap4wGSKVeWIC6+6EV5XM5Pq05x88XGOQW0uCESWexGy/3Veid6mOMsHCsauPZ9lYivJG8
1qwbOdJnBIOAUFVVdoidk9bTVtSgjteHuuCqxIiYLa28pLYksl5higfHxfCCkBctFC7Z7iyf0S8x
y86MRzeGi7blKPPrVu+QwjgvPWvfXE17XmajB/JfZ8aQod4PBxcnT+QGNf3Z44tASgID7iqrrtcG
xc96bV3H+209jrBy3JnEOlDnjqxt/MGmLScoPRW/zTrBJuLXpCQYlDMvp74iA+YJWK8/hy5gl+SA
zUh3OYzTgYveFIkqwFVgLM8HHcRnu59aWTtBlR36eg8Ah/sR0Py8CAMLbZWmwL/icdqVKFJnoz/0
OFsb7am2LY0h53Y+jsashfYLBZfN5CkEQCgT5Wo8LH2iRvysGTg9p8Mu79ljgH1I/QWmkegHx46y
Kvx7Avd81mYK79VYzr9e/ypWKl53zA+RwVuL11yTByHJGr95RlMSI9wIjxrsd3fdmOD3f0BsBldf
3Fhkfw9O4hsFmYBYYNaB1Jwb+AJQEWOtu3MW44xcPo+7qTt0KBQeWP1HPzFam+4c0XoECeXKEZ+X
/ruxBgtqqJGzJx8WFxse+GYucxTp/xflIz/Wh0hvif7EVVuLI+Ak/wFpuk0Eo1mkTjTj99yBrqny
O30mpm72mmEEInFlGWTVaksxP9e86jhcUbcwVTY5YHEbinOlr2jS0bno8SKzYkwh8tOTrsPKR+Sp
/38YNyaJJ2AaMJYp5XBXPXLp2/6xXaQb7l36MLhq5Ed9EYJBGUHZ4DsyZFLk7qxJe9Nj1wqgxslS
PvjWakw/rQ0DhyFmFjpwgTAsFDhTtQ+esNB1eIl9OUCLrNoriicmKGqGeF8k5hoXb8v2WnHu5dwD
BbMVwPlNpYMaCH3hpCSm26AUaMstmyY9IbNujX8Gghbw42+SGux5TiVclNai5Yqkw/BjA+LoAutU
uncyeB+e1fRmVSU86bH1OLOpTeX0xlspvlL0fIGDmxv1mMpZuyBcpoxYekFsCzVIWIMSOtXCng4k
1FfwSGOPgt4lAHY82xONh+NJm9Ci5/HFPIJfnPUClifFqcajPPNku0SrSDoYikx/0rYkAMvA7T53
a/fI3Fu7GnFi5vvLl0XydTkwit8dzWy0ajVxjAt4wn6TeXgBU+mzbrX6qmePeW1W7VQItF8YxGT4
1s/Lfcv5eEQ+T5Qn0jFpHpCQ8dll8WRjhGIr63CS6XRgBxJ3kvaQgOwG+hzfc44c+Q0Db1O562m8
qFDPLubUbnwF7yDR4tEpTyqnCQVRhs+MdkVA9BPh+mJEjOhjIgIZWVENmwo+uSUgXiQRdVCBKM+S
GdnWOMvHDx4qM+QQ/pLbDYJLVGxC+XsZzl4kDhwddkPT3QfzwWYDZ8pmbJbcFPnz7oybGqb+O8VG
GmUaLBunXgTZLZxz7eYZw4MCj26TlLP6xN2xEekuUJNGh1mApJWrNz/JhM6H8vNnYChKBxLLDv47
2Z0DNOMPXrDuTvxXyxsM2XGXseUDxiDPqeJbWYpcaYZU7qApm+z7835oZ2qfsRNQ+akDoJ4++V9p
qelquSP4FW4SuN97s4l+1afyU0Flh8zk2RhhxiZVwki/9cDuQmrI1E8UcYjrLrDKZGvDXED+60Dy
BHRce6HWbbsDL/2L7kyh1jL3kYZ6S32CVHbDx6OjtXmimUoV1wPq71FYM1uOp0L9SFKsLGsKYKvC
KvgqcfWF9eG4fsUk9JbpSFX+OkK1DNNQQVF4ewLuBpQTlvtCetBxwtWVmHMOYQd4zSSdzi8/qfR5
50X0Ppl0CCvb/FTzPou63pk8WpkXAKkYY1GnySivINw8QdfZehHCuf0tsSQ94obNg1Cd1+4SGjAw
5b9rr0IlH9wngmENfb5K1YXRJW1mryjzZ9UoqGDRwEBGDYMcum9NhI+PacTBKRsroD5uFM7+/LNa
dCTrCt5mZrL92mc/2w/JotrM1sfgziHpiYi8tmbRo0jFZEGK9qHSsxiX7Wmko4fuJ4v3Au1qVvsw
m0/qgcBFwy3HCEcxq4lyvdkh1Lwni0fRCFLa7MdGOFAiS5y5IHl/K5PL7MyOIcJ5IsuyKiHXO6Hm
CNBW/gAIsOQFDPzLUYOu+sX4LiZtwWoEo2sFxBTtte5RXUlBWaSsWkx9KcIwdAA7C02vvN7YHWdi
7qrFUkPDFZKcceaWPiKTvzennUzO3fMO+0rHwdRwb7TfmjzkOxyOHFcxcBzYuZ+MHPDzRqH8Av0B
2vHp6bJDB1648qD/qyMDGYu5rAFnTDDaP8WzGkp7jXwdYMS7JOyZObALDbo9M9QvKrhZKLE7jT5B
beLv4QzkzSfVhq0ceR3Oc0ZJPFu12BhoGLVWmRzEWKa+vIIxbLc/VWWk8yUJq03tLyheVdbtEEEr
g3zl3ya+MUHNi6TA1tN2gH62+l53MMLIAeZO+TQZ/TsnRqyzzIUiNnCNhFUWaTA/FRXKD/m3g2md
KkttNzjTVIgW765lLBgh196UMxDY/03r7BX4qAXuerX7f0w1My27lnvP4RlAoQ2SWI/Oi/iNdv6u
nUFBi7L8CcHxyj6KrWGmPDxLq3FRnpyzwE52v9XiWxfCrnLQ7HVY7BcfJqZVjoBD6KtoTFMVof3B
MtvrG48bV6B7xf6VZciN+ZXbxee9jpENh6A35hXcYhgol4J7MMv2FBv0FO83j16I5EYAzyGICfrX
RSXrvrJS0zzqfhfb9CKe/PwT/FMdDEG8YpQvBypxU2r/QubqXTaPQsy2yIdIlRt3f0clI+v2BOe4
pMFM1USiMLNXBVuJDlhS6XQh5VsGyRdbytZQQmcApUZpqu0gojIOJCExB3Vof8zEHTGoHd8z3nND
AmJRXRpBpZdvo7b4BUXwrdDU2/2dArLvpC259xpB2AyjgM4b4NGycNXiqIfmpHLdZo0dsxdb5lvG
Cax0WlCcSMa0MW5i0J4sznEy06AFlcCXXyAaiAykYjfaJyWBcHmNfiOGIwhl55Y43wC1LB+BLJor
hf31bBF99PvBDijJ1YB9tnJtqv+hp28+DkKR/DaTFngVbd7T5M1lg9tskI2Iu7s85IO9oe7lEo40
idp7xrYZPQ6WAOmXnazbEUdNMI18sUJHSwa57vdplES23CBgFJ3zR813XQVRnE71KGkZAndda+4k
bDB5vvAaAjJmLWrdSprK0poz9UFG8JRHQi4g+fhGyC/Ln6pkJFdbupsay95r0X6tFhKVUVodqGC1
M3KfHqhB/wl6EeBUGHxnolHkl7VALoHdBCdlzOwFob6nf6rUiGwyGU5FIAuyrawuwLy9UJy4CkOY
EpRIq6x1IeOMIrgM7oAlg/QB/HQCqpE+xV25fYe9xAFO9TLdOdNkDbOHvrryZxphFvhzqUcG6eEy
N/d4LRl+FIjpL0xDeTisXKyRbEjWYXU5NkX6xjelaWRZG5X6mczQYU9GIxMOepRSRZYbchdYejLb
VmwjbXAgeqNawvN9i1O895UZ2iRm9zdzjpUIGYKoeIyqtAXJMyGA8sYEGe2hIA6XkM9O8Vs9dW98
BxWJWRYxs1+eTZoeN2gm2K2qbMhi/3OHindzvBbelJuVnmv/L5vAFj17axkWVVpxLBytH1YjAYng
Hl27KjnVfMkS/c+HT1EYlvXBOaTiumPqH5iDv19FFOxa8G9Vse+6pwXHrKAiVskEnCkNTwI38Lqm
StYgSDAZQwd+Z8PibhQ6R4XmI/PFYyGOg61/gZ3S7lhnlfJWIk/bSYTKW711VDpn+DlV48IXwmeL
xoKm9U/QoarBfmq0Xs3AFZgBHWYVPoH3AFK/sgQFw8LMJFqwrN4OUlE+sURSnZx6xAzXoIcyO5bT
5ChLHJDJK1TSUtMK69lLuwEeUTUcAeN12himrCiskLamOqDN1j0gHLnN9xp8q7QfdVv8DMOfHAZ6
SVSrY8s/0eYLbtLk1t5FLJo2R9v++iXwCLuGkhUI53loOPX96t46N8PBsiFC/MzDEqJgkVZhLDmD
G15kPVE/AU8Sg2avUgqnYz+E5EY8KNT1koJXSbGToujsGD5HQjPAoAcecrMRHE7IwY4vjHWdIuub
ADZW7ES2jO/GDjJYOhlL+s7++FqcOv3BGadf/ks2t1WNfLPhAYz1HVeZ/bm+cyuBwAb/e8/+nb9B
ELKq6AOTBZDbMgVhaxmZ99vxP536RbKWJnSNsXHTrr76exwuT3DJfPicySaJC1K9FQ0uWUR8oaig
7rDXT21V1ulviK82yOdPkIgz5Ym9o+r5ZRfJrZUyYoYxHlaPb+4DlfEpSnNlPwapwmJdyZmjKiAg
tCniSiOggilG4keBWKPc6q97NRrHfGH568ZMVsjYBZF/EOZ4g/L/oGGKCceD2am62V0bx2xw0dRy
y1wpsUOWVlbleyVfnGAo577ELUQF3pjhRHuE2+BzrLmI6d/XsPl4ZMOaS33dNo2/vqYHOwllsQdM
MjBg3SURYBLr6d70X1jnBfTw5OpisroyqYwQFmPUlE11jW4r9GF9Ljy6RvAVD51gbKwPMZhjH5C/
yBRlAkwh05bCYe4MIOg74I8EXFlhVmhpMjOK8mUVdrZjc9jYNoFxuSk31yFmkJHMWgcURtJcb9oZ
jwl/M45eb3hMqiWGA9aPnxBXaEKvGN09fDUjTL947M+K3CeZknl/Z5Q2PYHIeXYMgs/GYO1Gq+hU
h9L8ffSgtKkp0CEotC3EqKqwDvrGxLmrp1hqxl/PzaLIkoHYuuPj+dHGLENlhrpYOxN6QyLbegcu
PFlr0Hgm/I8ohXewHu+zKBZqEei8xIvKrr089mQM/BOomjPOfudH+lzDtCv0lVkYpYkQ41OMAhut
PRlBaGBqsIBqGt8sw/9h6z/ByJeCArdLKeAR1ZGUP6/tolh4TyXoAHFim+wrtc4CGzq5HGxKKoxV
KfoS1O/sEY5aPN5s3zrGVDQxVuExBxdZdWHep2OkVB012NwXhAzdg30wpS3bwZw7gAddTiLXuCxj
3xqsou8FbN5aIq2ikUoCYu9SrGIeQ6FctmNIRxVcGYJzGY+rsfXjhQioQt19ShQfvTHGOBMdYbWY
gpcGudVisG6n3F/rEjEVGnSbQoR8hUuQoRB8Lf04ETVB2aO8NF1p579WljFf0quTxHgK5xFRF/A7
y52D7g5socJOVWcpFHnlEUYadrLDNuZQpo8DSty+VIavMLDX4meIxsjanedP014Fqhfw4DJF21Jt
L4xBYGNbo3LVTJMrKknOXQUYcRXdp/PH0ZQT+5q3uQDGyHjsSQMfmgyQBazP5nxNCTdu2OmoscJe
YlLYKDzZSISYsQnRXoCwOziqmYYPLswbMF2h47c6iak/Gsw3FzzV+EVsFDl7fMUZazPvGgWnA0/X
TrhW+kHgGtDjq5yAGtAp9D/6OYxgtEWhek3Xk3WYW9brEB2ndVT7rSSv9h8S0hxuwVbSOQHniBoK
TwmuZ2Jj7fJd/5RJxcT00SewbEhPy0ekxXgMVRW/S8zIzKFZLugVnl9owfV6LggGXjETyhhPFL6L
yTZtUd9Dhfl3gpFUY9uDM49V+VF2sEb1kI6LC4Bpeq072PeCtmkzT4E3hB7M6Cz/UOmYY8H1tuEq
OjvrfWXLFN+/DK7L4Tt/Cjexbgwh0AprNTQedeV4l4efM+w35LCnTbBAozCMFfDutmUSRFyiT3l7
aC2f/cwgH3PKs0zTl2fPA7vck67Dw5KhCcu4XR+2RKldElpswSx47/yIlp4J355k0WPzfefFk5PR
C/mEYyZ8e3IVquaMQL6ybd/C62sIF/I38A4uPjtNcSbNKUvGiAradF6TNrTD0m1GMQBcIHuFDhUJ
i6IMvfHeGqqFFZpGnkcO+hgqpcqyBwAy1O4gO17yo1GD1wTzy1Xxya7ijUCZYpqb5IrPdV5lUpfa
qQ8IrUUyU97dJjDJjFa2JI80BNH4ZLfF+fNzItT+DnIGZG+ub6KRfP4PMZGWOi37tDXDiTZ5hsp8
wNwS7XkcrvOBfmDQdXJ9EQ+wmjvFdyCEgrZDvZZvQpXUry++sjgNRRgkPIFWJAv8nPShPeE9jEFd
s15gWTE4OmVo1b3Wr+M4dpWEQTlAr0f5vulYs5s/Bji/dPxh/ny4aEEr0nz5laHpCF9AJQkWGP/j
7A/cERZI5IJrKoGOaTU/nhfxhgQ8UY2Nh5tFQqXa0eP1PFLIpv3PLKx+GXpDr2si939LqcOvyQPe
JKStMsfvF1lVfw4zWL7JFZ6jomRoemnaql88L9dkgnQOG095UWAQWLEGmzBrNdYOdpZ6T+qNSH2D
Tvg4h/G8Aj2yiz6aPaJJp0sNC9ZrrC6wm+G+WBxPTuuSG16QykxbUzG2tt1PODtfitzPM/9styhz
uEjC4jce4W67l0TH4/nSKmyuclDr8gkZkhMP5nRD3Ds48rM0HSNlAJQpSGsujFtHhCObGbC0waZO
k/JUe7m/rAgoqO9I9kKZWGD/1OoO1jz+RqKImv6mIImkUwa+WFAPrQDnNsxt000vQ66TpUGGpA6s
eOz+ZImn+cEhHiwjNaEfEhi0m9Q3AwVYPSM3FKuqN3xdfFhK0jwlHhsU7UfbA3y3nj40JeB+tlIt
5eJearIlN6DJijKh0oRnzmD+1LXnBm/gVeoqtHA1DGZr6oleAPi7Vgb2IBfHkigDqkgPz5pFF3xJ
iFslS7gDO84GUlKpw3XAEjf+kSEsnygLK1n7CYEpjL1KyAch3id4cTEO5odVl+WNYrSAbs5vFOhk
L+oUv6ES7zDGkdGDaiyx+VfErfsqMuMYDKpjYn6vcaCQdfKck3ptXhyQDbOgpn/8OJu7C/IBg5ys
3w9alOd2vUnIPruh4xRpDWWt+9HPdFjEcmWZaiAVx90loAOD8N9amJU6clBf3hE9kxVg4q6S+UgW
iYasOXzwPDeLBYooj/drJj/Jysn32TO2wZrYzHdjXbfKY3zdwQBT2W0/3Q3BAsIWxeTNwcFCWEPM
Q/wUsXdbHKcJ/Ywl0SiRN/G1LLS6t8IQv/Ljp8JGr6zM310eHjydsPCumy1v7hQAXWcB0qNnRfew
2VOUsTwa9DEL39mmJ+bhjCcJ4ZIrUxrkGUlUkqGJCeZrS+VWnoiscgSLOm6Skayrnc9zU0ijiHiX
Deg+ekZR+TWpMZ+/Jx/RvRqd6lxqTMGjGQDbr9Qjveuqwetxua80AHPJ+pEyUVKaJmiwOWqPl/rf
lqSt1JPb/3hq6kWmFrZCaIeD6/jp++3uJeIfOLCeKx/VKyFtx1W/H1DyICh18OYG93/1XKV2gNtg
fm+f+NMQm+8ytuZfuAcIfoA9/5iPKfaWbmTRSlsY2J1AyfFBflB8gU9GfhUaufWft7OI6kdKsm6p
BHULN2KQSDNbL0Hp0nAIROyrS7YwAYUb5bYj8ML33h0uE4sPyVJa651rZQPqByr809+ty7pDKX2j
Phg4hOgNgi0k2jkJEwDXrIikMisgv5KFUVh34UoU8vNY46uHA8sCHBBUKa2Hhsa/1yMRCiwsjNlF
DrK55P+LuZPgNsrIVm0mHKkxxCUmOeN108HB1rg2GEDiZYzMX17b7Qm2G7obKh0gF/FtqT6zXlF8
uzYQ560QEvFakQ+i2izhL0uncJEiXE+1sEsJocFvo+fHzd8rnpiUkQyV/ORuRi2zdz2LTYflUprF
T4w7wUA67SWXKOWOCWOELoFUCmorQUhAvklcDfR/GL1SOwcLSkDbefx1UfNA3b20J/+hVSNf1IPb
zSJXyra8wLFkQPaBUDNaQQtMDOITbokKw0/BoHthpQh42OR/HRVPsA8XExgHnlS7XFqdsv/G19++
RW2XplASHviD2zZZ5euHMbCGY4nb1x5A64DiiHEvmd0VU1aKzdz4z1joTlUaxa0ZpFcbkrnHnfCM
8zpKi++hoX7IHSNjlvmkg1ke20EHtCPihr8cC64HjOxChl0hMWybIW0Q2Vi6aHtwy+FmlMHhQeL/
m6ygxAqsvNlPAyJOR8JTQMwv27Lr4KbwmtL8FzSSHxw7yN2Ooo32DnbOjhGbBFBoPKB4NvkMVGGQ
gK/aXYR+ZgfJx0DZryDS64evKrJYFsg7rnGwFvv/akTyOJ5eNz6C6D0VffNhievO2oc49VGW3Xgn
6K05CNv0lhhAyOfbmLssilHvMgrBa9GuOMjsCONWtTrpOURcL+qrfa5B7Q68katqbvnm5LfIjJLG
ZDGRZgua5IWzulgtV8FGNTgWwNK0AbvrbU4sQZXtOS5vqkbIJCE6ihNQVHtHqeU2OlN34DBGChRP
mL5UH8/CjdV+p+ZUJ92yc2p660BOdjdojJCT25qgo8/C29jEZQfJg+22I3voNetDtsMAxe2A5Npv
Ck8BZxTQ+edB7Sv7rqpzMoXXTfSuvI+JqLlI46G0NWBBqasGw9A1CWCtEbu1d4hZv8iabCGEwgjw
9LZ6TAa+2OMa7GuAlLKYnbQorx+v3uZfblqYJE24P6G5wUS9e1WToXOSeIMR/9xj0owwPECn95Pm
6IcA7vMIXPE42japaQbc9MZhKp0jHn+d5z6ke42vPPMFVbHb3HQswA5Hk3qr4WDp6nfgbheom+J3
LOQFKspBiv34bfpfrWkceNDoNk6gM6RylMtdGUrIcxZkjZisQtDzQnsF6EitXX/FMBRMn8LF43vO
C/QNx9/AgZSnH29ngl6ltM/RTFSP0fDzIAccUiFZImVv1lKoFMEJesSSlO1Si5wkNrJhl4et4PeR
7yrqHCezBK25nLX7ppXAv6cg5qMLL3aOoAPkMPqIypKY2FwROIWFOW/5rJhGE5Pi8FUx7fpzGRF/
CNsePMfL9J5pi+RwfZCvK1FrVFuETZFXNLqUzEc/LOErNfC28GNsjG0nk2tbZuUAUWYsVCQ7BS+E
Z+KDQ/W2e/hBZd9fmzXyKPiSn7Z/erYoDzDoERxV4fPzcLK7bS7NNZ5VQUabtrxDHtYxBg2CGyLi
uDE5FkjuzS+m9GyGGLiXgRMh04OvlwFt+zbjRMpqj/2GwWgpX6pabGbrWztync8aMIg8edfbv5uY
4+Tzze0OFMsdH2JpSMqQ3j/wgm30VxspSD9gNp9+c9+qkDsuKcTswDTPOLl41VYyVwkJNTZXS4P2
HKEL5Pfp+bXaSmCgHEyxLEs0JZOc0Okw8dzheKIELR/9kA6cGJxgoE33JO7EljQzkqtYEQCTAbKA
gvO8a3FbE932lfDz0s6ivTtLTuMgbjgA1oTebBS5LS2aNSWMqPt5LJHpj3VKELc7WZ7ylAAs5Nkf
qLocQZqVZfzUaYM2/c0MBaItaVzDLc7L3TBhPI1hLRh2J8y6IJw8+/I61gRz8NXQAXXa8X/LfBTP
OjCvAd1NlmbIt0vGWF17ypGHQU7g4fEAoCDxArh/F9wAic6v9xdRkIKLto4msdSwooBwAXLinfPP
h3zRoQLvKet0CgZc6x1QfhEl5Bkthmkkjsvqzwmxld5WNjUGqeUnbk6NoblYWzsyI5kPhc6xnafd
U2YdmIINstvcwFBEco0gyHkpjPbiWASe5Aads+vQkSYR1tYjoLETdvQJlPQKD/e4+XeBMJWOg8qm
t1D4hU3qqADah+Eze7iy+HoeAygeeKPmCGkT3QNA8z1+sr5ev5rJ3Bl21eYC9rWAqi0+uDu/7KEV
dTsXHuxl1Qxk6LQ1GXka7SOloVFoxflTNlybMMJGlibK8BBJhUdQH8OIXUlbzTg5UFuuBe+yZ5o4
OpRGbkZcivU6+nnsVIzjOvaakqleb3chR9vV+7/whGeMvjVa7y5eXS+a8bgG1W3/v0fZydA2gx/3
xS2A/9fvLk1Tbi3/3rnswkCkOSlBkq99bQpaVX5MdDZi2yPngxXojUQG1hrKnom8JZtOj5XIbAKJ
5KHHhHX6nQDsXyYmhk4djUSLI8/KbfMP/NY5OsLPvYnEaic//MwQTfA3EHonIi+ddAa4xVDjcjLF
x4yAUT8aXQqY8MPX4qHHD+Tnm2JhYB1WZxDCk+NeEVtTwTMe1ng1Oepr0DvuDqUkACs85RMSjLkm
jRbvK6T9yRj+rQKj/Ho9MAKluqFuAJCckdE3pi0T+9p0EP6i+E93IpQJdxoGnbz37jsLswDqqE9g
/Se1VRyzGqOab6acJWTji++bMhQGFtLUkyeOM0lTNb3Bf6UMrBxdwhofq8GuAWDUyJl7TF5N9Yf2
HUUbbgX7f4RQFoLY0Sk1LIsJlnqWSJApxFI2fNsHqJ99cd55w53Dksfg7nZyDfDWbV+FKuyU2bYa
7vrLPmANqbDRadmScrXwHuquW37h5bS+VcbSl9xlVWPwaMWYTCyjPUBvP/BfMg3h+V7Fob1mUxbq
fXEdZHOji0y4alfSxymRul0CFQqbgquBS+mCNK6qNpAJqDzX8674EXNznvZWRJh9P6vBzNrt+xmU
XstWC3vKX22je92QnCt02KOKxhCm0ceVnHA9BQzo8L1L8n1vStbYHJ0rzUwmxNdso1Wx7I+6Ua4D
umGIw5xr7u3Q33lUzC+H8MXe3hPmnHYGfCsYf0n6V3wssZHFUNuhWY2V6MkDUkCU2Hd3K28d8ero
ChnU1BQpeSQsSefHwNE3HBj0skGYxoTlk0JTBvQQGwJu/a3HJ8ZX8ETFwllEnfUsqdOJRaNHJVDE
SYpUTU1Y+NltsI3jRWnRmd5i5jMa/G2XxXikT+eXG6wuaKlf+DhXzoR+X9tUYFIojtp4+1kOV18z
Dm5YANCv895xMxnUWp+g5DivMKTTLw0plHxc7as21R9ztgU15DbwIf+LzkntoVVCND8yTGW61XrW
7JCIbHa38fzblZMmu41Xdq+0JY8cNAj2RfMC9kVGJ0JZo9ry490geenW0XL063Dfk0mgmZhN3CTw
F7Z+LBvyV1IJXAegb/Ofo+P0B04puiVmIg+ez210Ol4YXjtfLj3dJEZlOXzx5HQLzY03akuze7sL
Hzg75ibAUh/5ZSMOw/pvpYdVGxO5jKBMK09MxKu0kz5j3gkZzdem7tjOqsHjKp64wd99Nnfx1zbO
clrT1gaPKSATEGZnbzTH56ZNADgf9dg8EQO5LLEwVx37k5Mbo83zEM+nEKOaYnNOSfbymL3OD2zS
Zq9kOVKJDHDgF4wyKHlL8XtttTSTvWkSTFHE3rwVGWlGg0nC0ryDdpruBwfdsydDzwHdfzfwnhU7
rXAIFHWcSIza3qhx6aqTlKblCWmkAtWrFzkMW6Lbgtj527G0jwjK9I1no9rgeg2vOS+zJElZb94C
8cwJMZpa4QeWId47ZAT6rJjdAC+0Z57gGYzvxFqHXO6FsNP2kV62W830z+D/6ZqK+9V0LaQWC56D
0hlc52ttVwmmJAhLP0QAOHuEbGlZJvcMMoviZDGyUq3fgaaVjQAmEyEhiZFeQ9PL+7YpB7xfNiRC
ox4hE0shI92oONABioOMDNN6LMpssHuRKPZF6W8PBo8vQcM3hGRHhCGLQ9J9nT0DX1VAT0Fex0+Y
XJMNa0uE/mMmmJ3AZDgsTW0FxFMteqVKw372vWMyekHZ3dKWxWZeWBg0W90Kt6+Bz+bQCp2Z4ZfV
SP5ePpNixLwpjLbPdFp9tdYNsGtlPYfqak4ZulvnFIqN39ExgxWi/Mt90IeQOGNyGBtmrYQI/TvK
Hg1cNqFIuyrkBixScSqPXnq0p6WBBC/zZIqFVJ42Q71O4qpjTCoam/j6/6dAB2SGZRYmzFO23yJO
TFVIHcuR+Vzdmd8REGoebtIbHf8EmrEwKiBWbrZ5MssjfzsYPMoDabSuoB6LUI3XfW1VnDGp7Dyk
/BZNJN45cEiNvhBtYPANqxf/0p09Dkwc8PWbLMj82P/r57wk5SC6k/4VMZTp5P7n9Q/4MGCLbYXU
4jG2lmdiXmjnkMv/eG/urNnp+K38Qed7efw2S9X5CObioAO7ZmtHw0ETyAen4AUFR3DPgzcbpL1t
s+o+bY9LUNege1CSVm3Gq9AJxKF4qwBCMXj46KrA6B5hS5vIICfWwL58OiFnkc0nebbbYEbsz8Af
wpd7z6a08EFZ430/DkZzmFUIw5MGFg1lW3XAgcJ0oLzqg+umiAc77Qix/uM48sB+af8sl/9ko8fb
Nzc0umHMmY7sCvB/Du8jFO+PYX8/4GfuE7nGHe8ndbhGo+FD8hyBurFof76jycABgfo8ncN7etVZ
PKdmt+JRXSrPsZ7pOZjMJ77h/F8cK94qOzaWSN1bFvAn1x0ZWugEE9q9WLMZ8OEwbKNSpsEpYqM3
LmS9Wd17Y9wA8MewfWkknGL1qQkOfdANU5Bc44FI/FSQ+bN902CNoI2a9D7UPmxq1eTEDlVk2xe1
S5ep+Qhwiv3S61sAdNUqCIE4NyqWFgu/YcEWhpz/ZvjQ+AmfUaNQjRb43Vn9Vfb80qwyfIK3cZHc
0tt6iYXzmZwjFhi3QXHJf6qJZABJ2f+l8kBddXOqD1xTSEvCBNYO8dPef+FuPXP3ZZUM7pXB0h8J
PS4dgBhpcxJVKf/LANiIy+cnhAOGTLiJXD6PWkDmN3Q7cZrX2LocccV1/XhZ0kRWt88GSmFzzPxg
U7Faci0pHS/v/hcj8OZ44EldNJcs3hpGmmmhfp7QZMczT+Pdvb8b1HmXHUtbSp6oaVQcYfmdl2sP
es481Xm/NlKck1rvn7Kjq1KmJbDZYSLc+FfP+d8/uyWx6wVs21+E3F1fQKrY3ZYCv4H3GQKt3hqZ
fJx5YhKMXSc7O7FD487f+YaGkmrYnpincXfKLVIBrA+iOlXEgwtY+3EeZvrUXgns/ymxl48XFIK8
0nuKjz6ZA4EHpTXUlhZey9N6k02Su4BN4P60MJrcT+1ccHAJUYBIjVkaiWslIrJXgaXTqdLcyaJY
BofUsfP3Tv+TQCRsqQU4QCAcYTSlqrLkTXEM441I1l6v+Vn4bez8K5fSRKzat5lLGqjuDlr/BBzU
w+K84hZeCdKVhyVTpKdMyxDkM6iPF6sVmGC1sqhb6LuEAIMfcASkKK5uH5PZ8B8WNDC2aUcFJN+t
6mc3HshsjgnQe0y824NiRkHOHeamMnweyZP5sMvEML8F3XzrA5OOypwhdRZhtXeJixgUSysiSTgd
sFe3H+xTq7hDyi4/SwZj5UETG5yTQ2v7VJnaL/lJZ+6E/ptCIOF6krN7WU14z6xdejolv0eGGo7C
Afjwu0ZXXYQLrHIShDRp8W/WvHFy7IGSTaDBr8Kbii/QZqbXansVJl1MkO+KjsOBCAqOW/OthvOG
gCRRq38lv7tsUZqq6tIAw8GUdIMWLv7xrR9XqFaOYwviQm9rcs8uvWfTB/SEPbm73U63cLAKYBc7
/4SpzPTmt/DIxODqNQU77pdJMBvPzIxdok+mCuRY4GeGsIhukhOqfbkIucJmr564YZ57ScecSOCI
ywM0y5jd7a0dNSTDoFkT++zeBVYvTOGHAD41cynuwjKxCcss6ig6E25frwnXKCOjVO2Ed2H37i/Q
d4qgA5H48JuJ/FA2XcIv2bc/jRdhuKVyTP1xesBVlawaH4mWybJ2CxvEhE+oNgkytoMwbD073cjm
cDEoX/w85s42Ss9+03/8LqLnJ57I/bY4VKir83pVtxR77pKFoHg6F4F9wCq0IEMHVUjO1+EAxi/S
1EEyMeEUCGvvH0UVjO7JJVgrpDkIY78WXTbrrwv8pm65Qjk9HKrxwFIkmS2MH6eY/m2LnIJpIx3f
v0OybPw9QOSMOuKBIEq/U15y00mJosx95cnuU3s9AqAEhdCpf2EueDq602qEkTclMfxneYpjTfUM
5ntcD3SL5EgYcNxGADLOKihjd0ypaphsr0pLFDXrK5RxrNPUUtVOFPCu6yywDZIXPqKN3UZy1ONq
o5JFSALKrSsrgcpuYsvb8r/zOsADjxSTLGiLPZlW5ybCf5IDtZSUWXcEQJSlCYnwpIdhFJ4mo8vP
aSCEkQbi4yjO8xk+3HLdkS8FMqK5DuZno1d9ftbbsjdH4CPdkywGoZublFIRx0pLPSYu4eQtHl1b
q6AX3SHZj98uAdqmzfxQoBgNDx2M/7+0P3LZTfbDIxttnUJ3xYT7xm2T52ukdKhDouOwZ8t34eX6
B1T/QNudCyKdgnnsSjEW3Vm97RVBVls0KzXdUs63sY3WGIjqrG/9z8GmuyiP7uTaqeAhzMPXI2ob
Jb6yXLJvFyd05uOqv2dP55FTfrTsAgpAoyPiFbmkCjDodFLBoaHGjNS+bMoBZB+EbNO4J4EgGqDu
me1QY8rpzk+yvPNFuoQ+y6208CbRvCluloPN1CJ6Y8uAZWai+SEz5L+uyXEXDL0FsZV9baRB/mPU
6IGLdEdQuYGh3Id1sxQQM6NRhIy+cmRsIKSjyY8clfvn7amHyXrC0SM7K4cbE/efzgtqYfI+GcLZ
ZWDEwGP/zKhWMhlGg7/GCvJd38CzQHecuLxJqm4S5BIIO4o09uPNsUw0aeNXHZPJWD54M+5CrNGf
04h6mdHwQbdm9sPcnFf4xqiRmUA+nR95+ATr0ymbaZ9CyDbOk9kjqglpb/aHiHrhB/Z9iRVm/3tw
tQqT1mMW17EGQQNBi1HRr0H7SJc2HlmHEmyr4jtzALu5/urvMBXLdY5T1x8gFWSoEkiAmomIaZkQ
E2H0RGLsaYexS6b3R6Mq9YVkl0iLEa2W13EBCuNTFPfW3Dk/BXiB6gsDL+fWE6gU+EtEf2HGB/Vw
krIADk5Xiqp2AhBK7YWRXW0Yiff0IdeED1yeLKAig5jBIekU/66tIlwJFqDPfMnBEyOvFG/oKQLA
KP3+Mqq+whbar0LHthOeqrabDtwfYKB6Sxd9RSBK28vWO/JkUaV1z+lSyeEdD5fyPpFdrKAuTVlJ
ZAadVK4/7hvyN6xUztJbeiRayQnA4sn7/FI+IwXX9Scr/9yKdk49eNmC+q/KYFugtxt+qodczCUk
kE/5UftU78lWbBAVC3HwCygk5DLwcfAro/RI7dlSbzVxwU2hbz4ZAdYvs8NN/ugLXgAen5kBeC7z
GZ/joaSYpyGZkvruBa95e2/YIvxwXK//GwTUBQmTmMAd0RmCbAcZslKIOWp2k5bahIaq2aHNW2OV
rHSTD0S7AnAuoImnX92tHO0e+w49cnNOqdETDSFSwgF1lqhw6DNfdIhSl3xhwNUNYw4CXRxOX6ZE
wIklkvUbY8rT1HoektAfYmarhdpFX9P9TB+eXdSlfWZRontQEe44MHBz9lmQDoo1rzc+xEpjsnyl
Ex9gtlTMpfTnsv1PisIg4LTZDX+Fa7Cjpjr2XxHEvC4rSmGM3RsYnONuyHMdBmNQX0wekKibCsAE
qSmgu9SqJNzFmK4QV6BXZaI8X7JOLSl55BZcQQ7LR98ZdjYlxeHeld18MR96FQUh+zjzRKxuU6qm
5KteMFP3HzTk1vKT5lH1fimFUEOt5t2+ZmasNWRQDnRcFMefpupUzTQ8U+BVT9Y3TD+uaJewywXP
KxQrmcYXEFgdwV6F7DE9e4Sa3LisfdzmDqKsCaqjB3REWSb80WhYNkcqUdKiLw4Yy3+nnQNi59Ja
F5toUQ5jpQG+aFPD3AlmTZ9p2g/UNjbqofUE372Hyjoknw4Ipk5QAHQkVVtXnWB1idlJbTyIMtJk
gYOf/Pmoc72NS170lH/kGVralJOtkwUxImxUQB1GAK5xchFiaSrNvR5/tFUzh2tyCTUHYPK4u65J
E+TKWQ00llqsNmiu1d140G5y2Giz1VC6Q4NuUAHlmaKV4LjUa7rmwRv4130cek/J8lIRK85Xpv8T
SQQ1lAA9gnfGklAs9FS+Cpxyae5c+DsPa4yTJL2pIN90M2brs7r4j/74cJt1Nh3ts3JoInlTY8w5
tShrz5B+ZN5IIYPTlRn+ONTjFpkJJc8xh/pgX/OFHOiw66yG+G7pv52pIFvrKc4VW/E9AsJdlSjc
QwzHIuNA/0F/m1J7BoC1FFDUJrW71DQaOoequ5KZUOAlbk/1P52vRsJvr3MhdUblny1Hru366bIW
biyQUNlkgoRbX2BEmORpP3C1ZFLaQzXqKAbiR9Tj28N6hEh9pEzbfiexzaUS6/r0espBHKaCAean
2jkbJI5NDGClxWiv99PrLSZLpp16V+y8PxnoUtK6cDbTfKWt1yeZhpXMKUqk7kyl2Nj5z+xkVO1q
f4YJYKjUyJXWWeKB2lAFDWK5syzSiOsYCYp2YkJCtiKeVVrKvvKc24zPMquMAt6oz5SkoQJ/4Jxs
7nErOeVu+xAWq6F7/sUszrAq+C8T4R9/LnErehqJOuhNCx0X8r4YeVivFaZlhG/KCnaxNewDXloq
axDbhXv5jea0gfYwqXGU1yIckSo/KCQEss3T66c1opUY9+MGVmsv9onM5E+jyjIVskJUW+dU3fLk
zmLWF7t7jSCqJhOabJm16VCT+1uxINOTHMt4RZC4dkNa9hpu1NgTqhywwmzw9EntDBZfHtu0GY3L
66NlwUENDVCmNsq3H3110ccXPtVRxbe/pfc3BCESy5aFlXfug3j+2JOqzUHteja2nVA6U0OEe79M
OLXGNQFkQzlgLO4dS4cAyujxDu+4dxkg4Ooj3++9IXe04LiTiK9VsBw6PNh/ifOW2rLBbW50+hZg
s8UWDeIdXu3BVaf8zFnlolGSrMyTFrJCxW/iUh2JXNik25TqAkaRM1H4T5bvhRDkoxfPHRUBE4he
RMw9FZsdlsVdyda300vC/7mpGvNRbs06N3a4C9mhg361Rrq5pUV/eS0Is31nLLxxf6Z7JXHU5LPC
zL9QEPhuezOlYSNjcx96bOiHCrBu8mzfxj/G2fQVRsn8bM34vg1qUUbPixSKp/PCJS1qsbE7frNY
BIhjWQKbCtoR0Wqt7AeH6qmueXA79uwZ47iNOsCvuuFvc9RlkJgRmMbyjZg04ETMJGyUlhbU2y8G
1oP6XM5UdAUswrCd3Jk3xaRsWSDHsDFRKikR4IBVKYnXTG3EDorW51pg8igiDRu7TTEEwrPkLDEK
Oajud4yDygJbSXlv2JgqkpDApts4TP/8Msc12oAW8GKJ+SKB5vSXArFGy3b9s09k7i99HNds83/9
erOjwFt5RpQ/SM2Ri5clVhLyVSOSxGk71WIkB6OnRICiJg34040gV4NpLUJMvpvfAKwMbQM7mVvz
3MKJozKO/0SsAM4GZqGVjIOk+zDsdZMuExkZxRK8luikNyUm23oTArKGQn4RHbtkcnkDVEs6vZzS
MGa2Uoy6XG1Ht09VdLylL9In7Jdk/g7TAxw/a69Hhb0zMJNoL+lF9mlP6hC3W/MbxEPy+QAaLicn
w4c/YmRBHBTsDwqEK/Xqww+EKdrEgDlAX4Jydu4IIcDHmEijgQdz11aF6KtQqBjNuqAmAJHeK+JT
6wznPYOzqLWknMWWv2tPzd7NXO++cM+QxseyGBWNKxpGU7dOMSq274f7qgDi43m64KlqFjHBHLui
7hih61hYbCjRVoQSZ9C+SrucWNjtUKcngtSoypp0ntqNoK8ESKeqnD+/RbBA6/epRuei4YdyDbUi
CNse5dysRm23nORdnu+UDXLdXEIzc5asOSQf9Me+CxQa9pRRL3OqosGsOTUPASRRJHUpqWi3AmTW
pI7vkqeY7Kry7KnVrigc1eghBmsowauqmJN9iFogXHHu234W6I+tNZEMg0u4F6pzSUSLAmI/XbP8
JbIJiXEDxR8arGy8dN6g/EDmXxzd/+I+Mol+OmeMbuTfTCEkcrJfIaiAdzDhS2KhoJjM3qiNHQ21
hr26riNuQw7AMrZ1jAFRuky0f+jJGJMU5l2RY+ebLfEua2b0NJo/B4zl24j7S4+UYFuDa3kQV4u7
gGdWiCP3dAh1s7Wne+iDxpFvtcpcTopoqbWjzDDtyPKp7kPw/GwefYRKH7T54kovYyVPIGeUBDaA
6SaQ+vTGU1gNp6AYOSExPWrLiyoPIzY7uKOIFafBZ0RAO0dPnulyQlpVQbeaV1DK1crXAOPlUBRY
JClhDlORNOVpunKIRydhrHVg27q0o1MndBh+4ku6/IeheiBPj6JxdIaF/UE6+C1/Ao67XYLUnEwT
42DgbEv32qFTSb0iVWUvBVqXe6Mxga1sybThlfwYLLrepn2IpmamyQDpC/0KbQdnBffUnzdzcMvP
zPNpWACCl+wCFUlsrPxmPEbgnT6oo82WIq1EaX+2vDg7HG/dN5N+ykFEpX9HdWTwnZqWWo/zQAAZ
RQZUxRZtr6GyHsSIpl9u4q5M+XfgNiCr7p6d6bOmEVJTgLoEmsgPi5SY1ShJJMAoGl5VVDLj3Nun
9xj229sCeCDa6rulvxKR8aOo4aD/jmdOvzD9C/ZidOmB10gDnsbFn+W1Dsi5MwpD+QTdFsRhWN1Q
nFd8cn8gNj4yEz3/+IV91X79+gBSC45zyr3ARelfDmzNzM6xVL6Rdrbk3CVKeciih876acuZabC8
xiPmu3XLFeN2/CfwrfZLHtVNtqv3m3kDRUjx7P6DDZKPpEbxnMUhi2S5wVW6QU8EFYg1Q4scVxEQ
wjlF/rKSeNxwL3mIL63xCSimREQLwxe0yPgzKuZz4E7Qlo11xsONhw9cgefsfFFWwVBd+eOakuP/
ilCm7lJ90sD9ABSdQxZjKoLxZirFaeJKHn7RvcAz4xEBgXtfgT+rRDvzkiB/t7bJebgXxGcdVJE+
qM//yxah9xf15X8Av1OnrS/Fc6n1F0cheN7fRH2yR5NLnP/j+2w7eylqZo1bfnOXgSB+c+DBkQ4a
4eXIzs/rhGVZRbpeQ39Qw6waEqOQhKy9Kw4POQ/tWYCVJRA9xW7Bzj45Thj/SZOqwoSfxIVO2ecj
ytOSn0DvlX1mJPSo8d0hqY8QOSLAWidbjkbhMCt8JHuPR5vC2DANMOOJQ3TD6ahk0rlElhF+6dnA
s8LAImyw6jSGwu9wY4l2Y1+okrMo2/F6G9/qiDJ8mu3yUmQEwJAYoRwj+D8Ntk6ImcmYZRXdkKyA
Gb385rRb1+8D7V4OmLCB0GCax2HCoSaPfYgr9CUG3VnFo0jhiSw2bDvaan8wlIbY7rmyzzucWFkM
49CqpkEw4Tev6FCYcGPBxBmSucpEYclpx/bKDsbHx45LkbJJbTn2DtoY1MCG5mfoy2uE5B2l2XoG
F03ikX6i5Ha1AlqKdzYb8oNJqq6iAOkKl1k67+4E5GfCDvWgQkTBdV+4BpKX9BdfR6Ca2+K5IHHc
yjinUVmubgEqdnEBkR72ioFyyhBGg5oI3YsAILPZClb9J3RzMwCv9gq1oufsDrS4JN/6Kua4B69a
4MmjgjRhDxmBWvtMRCno4GzEgmRHwpjnavsk2Yc5pBX+HGnRrxwEoVGCQ0gH+p3h3MSSVF6CO+DY
sYRLqtx/7kweR8FaI7vbcMZMgtvy37D0ng5rUiFG536VKJKvoYlbJ8Mse1Z3+BPpxRQ68z/KLQu2
KdVYxIbCUiVwO7xbgo+4xOJ4yIyIUBnVmQX0Zzmbui0y9WfZR2kmEwb0iRdaREHxzw+BUu26EHav
j9TnBPSVPUTT1UWE4gL489nNOSNbE1UfqAoXviVCIuzi7olJtEIeRdNcTGQnVxNCqGu1R/ARPMFx
gBVZW1aN1HhsZGTP0UcnwP2BEHDRSI2UFzqvmpJiSxg5lyMIMB95syCKAUVCprJNrkCI8TBH8cW2
JFdr3GzSLsloen09d2XLb4KxKI56JeqCCru86g1/Q+T1hx2Dmp57iKyQuAG9S9+aqfkUrqYi5Zej
F+AeA9mNrIMu/y/XJtukMqxCiEKq9iSF+8k2V/TeD7FzOXR7bFao0SXZW/I6X+g5bQFLNtz14i2k
Ph+0SfdXqEH3mxUqZYY00RoGRywZixJAZRmlzF4j9WYH8H0qtovpyEXYF2abdc//PbeGPQ+5EQe7
N6eY+z52+H3GoO5Cj7u24yDigiW469KMVKOQZTrbW0KqdNRU6xkKMxXq12rRqyBeuhk5T+hfDwfq
tTSVwyzbE6cc7V9RzZVYx/C4JtNrg+xDSkjiGQyZF8sqgPXzmPABdb9FdwS/+rL+s6rv45XWdb1F
sumBdFjGNgTpdlTMHsKzsc7TV2LbeLdXvVCk968woLe+lUirpGgsOWPzdwHEmF2aOl4wiNz22mme
lnHFqFaFaaqm+2Z6nqtpkfAtNu0ykwN+A9Q2p4HQWK1qcZZteqb6/vEk/9+ixhH+wv8LqTnc9Oa/
WXg8aMmVBXH3HRvzBkM/1cD1R1pyHgwdnJskJ+IY2Euk/7UN3mqHDGwQEqE2ICTBDJSYBn+WjfKk
00rPYb431ml6tcH+6yQYOlWM78W3W5rRXh7Y0aUevfJLUGdPIfiXNjpYJ8Qv3OY0Tr1oq61GDKFL
GhLDNlwRXRmoiPeEnAxqjSWdhb6C2y/DN8/HUh+lS7SXNDSq69+k4tx00NDV/I0pcggMwCp3msWp
6L0kJeCoSWqnI2Z17hbEWLr5T1Tt8vhctBuPU8ujIurkbDnB9KAx3tqi3VOHcAOkEH/WPCjCrS2U
Gt2hja8GL+tMx9fAWN6wIavvOnhJSMEY5qhAhsSn4d6Wfwjgtggwy/G3kswyLXIUaMeui8qf5wsl
GLESLZWjOvGoi3hEKkkzwjL8LRQbzimQmti5f63zikMw0rKhR9fsrDSIsXylfk+ZlpR7VZYImyCB
TU9IhqctOQNU8FRQWC7psFuAZjentgGsznQJY9GxKwragjgSX5s4wImCSBBQ6zXAadAsjTvAq/cA
qZLD/QEt/F/oEJvx7u++V+IR5rUVvTB2Z+oiO0zBw6eTeB74fqPZ5nEZZ2Gl8ZyBRss5efWLfUdy
S9liJ0D/Mq4Zs8CczhWIT/dQp+fJriT7bVDHR7qF8t5Gjqh75mb+wwmU/R5/L/t/LR0U9a4D1wTF
oA0Auz04SIgXwbxIfI+APJQXQu71Ta0Xd1RIZM9plPfJugJo5T7s8J1zMLK2J6FhAJqA+tET2cKw
uWAgmN+poyXYZKiNnw4ewEG3hJil2Hd1B2dXA2NU2ZQU94jmoi3ti3k7ffFFC9yZqP/m7K9M0hjT
8wuDdzddQPh3Ix+b5cK5sYmq8qqDBhFqKiP8ObesEiPUpsAaj7wiG0OV4F6pY1lT5zB8STLSrjDx
BBCLVKDP70JcxSD3qFJOQ5/xgUDE3u4Lq0++9EpXUJyYTAVPNGurAXLkV6jiWHMlDoSlXeYFoKD5
QNkMFN5ZImsjXgPbBmhbDQL6UBp+krBrxLDCIPZxaNrtibcj6jsVl1az19YKLmzhcxM/kuiO6yWp
pXzxQd30BPWXjeHRpn9MTqkAGZV2sHUWyLaHmFRze4wiFBvRyhXtv6wZQBrFjBGunLNTAFrS2M17
uVMQfTwQV5xF+A2dBkf79ll1D+7jd4WJnVnQfdKQQ1Hh7uDfd8Ahz/SYK5rAF7op+6QDr67GLDXL
A/Z1hc9LC35MYrpfYB2IOf5XCqhNCoBCdJyM0Zw2HtOclzPmxEqQb2nSVfmHw/h1vf0iq8l1TIB9
/v7FXeEUwLoAzpPxboADQp46qOa3NcmtaoFlz2Q8GKBAAdN61caYmrxR1Bq/FqzQFBMOlTwF5aqs
5pTJ7bagE/h8NC+5BRlF/PvbWWBh7m9DInLo8xYncIhlBqD6JlzR+Ru+v2AtpLlyryO2G7+WI4A3
x45o+ji9zTInLU8Jvndp8rXLDaZ7cut+sjsFmP/t8JK3bzxKDcWgqY5+iZFvma9wfKdJ1vWCXpdj
KKoyZpLb+ncOL6rX548K475R8vEnWTYjt/7KCgKPsdQyBClc1v2JDucRbRtYgGPXidrviiQZ9ye4
Wm/lMAoCC8AKmYccAKTzcBl25mqkPTFCBWBbbGPh+ToHFEh7hKzvjHdUnEkBl+ub+i7lfGDfNl5E
Xfq2CjDAddcvccEjxibyQON1+PFkERSaU7xWlwffwQ3ykzSExUFOMy4VttNLl3NxrTxsqdTH3CwY
XgQv3LL5wgleZDUteWyW9SXOAI3R1NOx8ERgYiqPsSUm+jd7NzccUKh5TvRFwvwoWuPg1GineFtl
JcOTvMOP0pBrxZlsSR2jJZTDCKSy32rxkx6u2qIat6xmPWt7ryBfcZLUdGYPxpw3HbVMXnVj03Xx
Y7bOg+LgT3Q8CfODG2ujJ4+OElUfgekBKmlG+W1TwqOHxmmArmsUtRpYTU8XlXMJVWox2MHQbfyK
PU5LX6T60aIW+pwU1fIC9F4a8pu9J5VWPHs+n/Tev3oVM19+4pQG7xlpCPv4oUTkSws6hPs6yLyv
VEUeu3/oyqi9jsPJJnWU9QngG+mjzyvhJ0GXENO3dG3xpIxJVE4zOVcl9hFVgMIiAzxbGDb99hOe
zYIOyXsQajZ2q/SSq3/8iAVl11cZ03PpUo4VgVJ5ioQ1bRD75DEU03QZSJlB29XEmmHFHmu1R/vd
ufHDLIj4/h4VV6BvgJB0V9441pbUmc++2KwJh+WzkFzxuHbPrpgcS7gxd7+WMsxh5w2A5ynJ9yml
lBmJ8RDkQ8Bc/PcdTI82vSPOph56bBpRSLh5vyznyxpdrgCiW1v9lHO1xiAZozsMIe9d+uqe35Ex
g3C/04M6Ua/S7A2B4i6lf65bSAxECREe+Jd3ThhnP7ryphyUVFWLzp0dwqIea2zAk57y8cQv+tBU
IM5fbOvoMEEI/QAMNg7c7GdBr3Ngl6cN8xBwwOwAkVjLPl+UZnXh5WQP70luWjlEQvn8wblpnaEj
84CG5lMDUVXYqX2v61PMIoZdb+sdTl9YsGqO8eviAGMH0GBzeU7fe/vhlEvaOK6MutuuX/vwwuCI
Upm3Q1KwiIlHgkkMwacJjH6HAArLlEGddsHV0digCMLSjVni3MHazJZgIyFMNR30t7OOIrMl/S/O
GTNegywOKIGA1OQzgmhg4859f53hH/ZCYkFJTJm1Z2R9VodDumuICNR81qxdUCnkj1sPG0t5Thof
/5qvhgLVo/WHpRIIB1EqXgmYbhmXUHwCN82ZNyqDDvmjGvURQna8l3EC3yy2XXWOynGBVPkNU/PR
ELheL3lh0hckR0KcP8ddI8nj1lLkOq4bN2wtujC4qlnp5OjFC2+o+xpTSm2bBNvKWbWp/xCLn5jP
b6wMFqD0aoicdvL1ycva4tyqvZNN1rjUHb7cu8pP+bnTriINbHQxRbyT0+TQz+fml10E+g6UmS+J
4t/rpEFGpjDfes/VLICK1RD6zrUWVydGvwQxjF44QDi+s+EVVBKaUfgz8hbM/tIdI8C2kefWQ34g
OSoEQuW1wU2UzQzJV/64r6OKnq7ef8RoLUBU5PQ+H9qREDaq8UhaH1fn9OYCLOFg9FQQpCdKv734
1okjtoFasK5XXVBBmkuMM5Syo6o3nvGNKIEcp3Y0/DJ+eAllkLvjFEKNelF2O601PAPMOGuznNrt
qkWDBHkM7W2ePAV5CnJ8arPQ9ElfDRe+sPmB3JlodSlbZkThswtT/vhErlOPQkj4zJZyj2tSWLzS
2CI5zWwo6aVHRZmTK98DVVc1Z5/pXOF4hCsDgc0XmKDA8L1we0WOIgKZ5F7Uzk53PUZzUpq1SzNE
1GWfngw+/dex2jHRqlApKmzH63bE+gAzjKX1auVU3gYOHIUW1p/sVE7PikLkXYNOoiuI7JwNtaLM
bLeqUJm7xpmudENUp7HNsSCCUJNgocz9ECb09CGhkMzmBR5y4Lcc0lQIVusG4nzB1jjB9DCo4Avs
ZKkhcrqHpQznmtyCGRjWYoL23PNrhIKkuyeekIkbRaR6OnJf8kCJDlchSih7EPdVKFvAucLwL5Ml
Do7dY4u2cyZlhFyfb6MERtNGS3nXYxmrb9MVYXCz6FkyrTiscLNQPwkQJ4qZXsYwaXr++m84Wka4
ApkB9vFvXE7eoznbDvmgTxaaILENe8GtI+ZAh+kPQkiiRgd5d5bD1jzFuf0AQIvAeZiMWEP5YjMA
90LM7TCOZXgoI5RggUeTn/g1KphD99D5BBC3w/HIJyQcvS9JFj9yHx0R1MaSefWBrmYfvdligAIG
bBTiWbnhVohcMz1NUBllbowSZa5eLqkgkNBv3JWesETSFXhrEFwks79vmV/knQFCrSt+GMFDJnKI
dDQhahionsIH1jZ+Z9ES2cIY2Jtp0ljVXb1AnaW5+aVKM1pCB04QYmENClmklxH467RbqweLjdRy
lGtQbjOHUcCY8vFH0W09IxuEch8+fvu6Y4trvllaS3prF8JWGbN2cdt/POK3ves2UCrNReBxcVoD
RIRelUNpuQT4PMQnEdUcrD4OUKM+0tu2AwEx/Haq9+WdJOtaUjSWWiHBj9Jp34j/OKOVoVqIPKkW
5pUdq2L60A3N5pmdi+jyxYWl0+xIQYrUCZOPDwvBs4zR444BRlwKMcpNyGMY4LUx0wE5YtIhWYti
q2cX1Rr0gli1CjOxo5U0CalG2xnTBRzcLnEgAKAt8ssFuy3LYmiMsgtZiihta4DayITMlqznlrYz
XyEoSLB2w9ujUv4/t+hYa7o4XF/7ZSc3XSasx+HRmHf7qCYJktYvg2yHX01nfME6VlsbPuQzGfa8
Q3oa0Mdr27YOjX36offT/9hn79tMzPlVGG1xQtYFguUs2RusljV6HtCUkeQ4GK9F1oKBedGUtPAW
Q8YW+ubYo1S/35w9qZ0hpFgbLAMCUOMrZFatkZoTZTQWx0jbRBmiRa1P3ity64d/lyZw2TGIKmCU
Gk7JxAJtgV0hM+qEGz+AZFsB6X3agcA8yp9EarvyemAvOUGBkBdcsswdCW5lffOfUyQKm+NPn44a
h1j0FE5NOynvJ2vHiZCXjIu6LDYJ5pGjS7djusF7RyPvZUYgzqdhQ/W7QlMMTX1A39upGYgRGtfl
JPyg5BjgnMLqDJiOWqvvvELzRiaZQwWbtpOMuAfVlv66g/Qhgbc9bIX06AHpBcU/1YZKBNZXcNw3
MG8wK7znr9PnP4HG5cDAuo26npPYEn6Jkv/1UokWce5s9MwzFnH3KL6MaZ/3Y4zJIE2OA2CRnCvT
IQSvgKctXUUEDwFD1NM0uHxUvXotXa9N2d6xwtn6iFS9uZBMeL7IvweG4W20bbGTSp+u740O88nj
XUzuqjPCopRyqg2dB0eNXXjhLfM7EhL3Uw6CwdgW9bTPYVob7y6F1acSPRjd3P5GpeGf/nWlWD2q
IWWc5/7vIEJ2Hneo0jUprk4SGNVZYwkuyJcyn+D+UenfVA3oy3JP0cPFYFkHHBJu96tiKugUQCeB
QAA5qdivns0fomT4vYgYvq8N8hE+pnNy98KW8+GD0M6mDb/y5n9c2Bse3SGa/A1xkfq8b/OaLVJP
KOhzFd04BzQBkAvmjzPTj2LkHFq3fVl5acHUA8YKiGsbiatYk91swKt0FNIbrNiiXSWW4VsBXu5/
ycy0EOunSlZI89zXAjJEBQ3miO4hHtGrv09xWWhg2cL9QsL+5LAS+SN2Ck2UKdfXhO5CD38vLzda
8qoZX5lrOqVVjMe+htOyal1S/dEZ8EBUyi3Uu2ys2wDyO5NnP9zccUHv8E8AV9I5zarDZT2oISWp
cOwYldbPK1pHtFs2cDrmYsZaIhVbNGDBk0UcEj9EMvkBp7PNSxNNUapaUcXvpeloIVzT4nGi7oCm
Nzaicdh9UTKrnaKQsnLwvpWHslW9YnFZfHH8U0UiDIZ0mY/aJYMZAyYyYCWLevX35r472+ka3tK5
CD2Arb9zT5aEgiK5cFyUSbBUeZRddWFwIWOs5k013qA77hoDyJbZ63GwMAxJWWNoqUhC4dTZC1jD
tgddOyAljudOCah8W3cVdSm5jcV6TZpsyqsFzsD/QiJY6nHZb+UcOCqF8S4WbpILwkRUIbH4/VIQ
/S9Y2X1/V/4dJOmePDz1/G6q2jl8iFcvg5IZhzv5Vhoz+Dap+d/EKupQgfA2ImzN/wKkhGdil3rZ
CtEqSL2NbmrF4TT5j0JCntjK5bF7l7zNRKHp4uzwc54KBy2BGw+gUtdGh3e1GxRLTREu5nOmuLx8
F+g4DdyZqSnZEgWx2IunCSEn+8i7AHG43S9COM26f5rfhN02qt0+0YXBqgn69dpHTkY+cVlU3Dwx
TTwzgRwRsTL3AA4xEbakw12I+r36fIgQT5KB911K2+MGOCIoithi6VYYh1/RzveOY7OJuzO4fkOH
nXddaLLELqqFFboGnK87/5c2eYjkmLeegLEEQO8DHilFpVyFFuxj4eck/jtCqjbhV0fIEnUINSAe
vxmlehubgu9ee4pNcIxHntrLwNoIBhA0fpSuQRd3NsVQt8nJAGlrGUyjuch+MVJo/mofBxBuUUmt
w23D/t8c51vaQHcjSMp29DxtWJVb3tU/libPZOU226tZqshbXLbYrHfvkjsU0J07UsKcY8TF/oLp
2gwQ7sl+1gnwgIQu+q6RUDfXblIfmoqQNeOfagHvtxjRWuyAgngLsDFpZvvaS2RX7Sx1ybfQ7Gcz
PG0qVA89dX6HHrCA6ZhyQ9ARtXAwELLLJX/d1jK0CnLEZkQbYxJdGlfUQgh6idcKhSpnp92WXuZy
lU1wh861gPARrQvm9iJD2mc00GfL9zVfOkbDSx5H3w0bAgvRA8jE1NvmSMTIYIot5bmznbjqNnwU
+IOVzeENkHyPRJh38uEWOO2/ijk7rcMMCZlvCKmkeKo6x0N2WjeHgZcbfA+eYhcfVDVedxOcOoci
5/DFQDVAMrLyrxaha5Kp+HTygGQQfkeavD2y2A8LBwhqXxobo/mZLudZmwgFBr9st1XnzaxE/AY0
0LzVDILSK6T869FPkkVtwpMHS7hlwMq/g50DJt0IHuQ3R5vPVY6+kIcpycZa5EHRWz+8W8A/LkwN
qqxR0chBVBfk9fbWEwfY2LtUjxGIyUDg3RvWtYCAWwjojVLGj+SVp3Cb74YrjgtzNCTrxDP4ep2G
DtC9NybQ00+rw/mkVh5QF7U8zXhJqFAQQNppBCHZajMvdTfR+iZXdqT6FULAnLZ1zoWcYxX9di9W
cREBioB+qv5fJyAp7ZCNz/xX9P9aoSvHOcZjodH8BK02jDtUDShNtzXr/PcuZCJyKvRXc0PGUJhq
4umYGh4fvTogqFo2PjB3ufwhxWcZUQ3xJeq2C7lra3wEO1zLvR0cdvU5G7sFbEvVz1dkyZ5ZgtRz
/VWdWDJjimh9d/Y70ZK3Kn32PxJ3hNGPUwsir6qvyvO4Jd17Cwd2grmhBhdXrT885mLHX8JUEu5L
SojRG4hn3/MI5l+Rd/Kx3gQ++Ho0mC7CekcWYSoqADfteOBBaU0lrJCdi5Hp7ynspNrrzzMfcoWX
3eYHNGFA6DLm4Kk2CkhI1y5mTwFzfM4Q3EpVRUYwbzOw1Qm/lgpIht3d7PoLYgrDuPq8Lnwy7J3F
oIkW6288hRYs/t7Ao//ri5rGv0OPSS61eSSQM+8nvFJM9G0McFTgnijsA2NiFHHvRPM70Jh9j4tk
7053nXaTlKMLGA+EcWQFjnAtaBP86eV8jiASc7qiyZzhbm8oiuqoaRY9CUAq8zWMY+fd6BIEbqlm
3JFHGvSv7jZrkAc7z7pLvz7Ubt9gETZyn6vqaGlat8gcvN2GBWgwKw9Bn+42zbOA/82WyoN5kzXV
VY4y7gFg6P8tX1zXRBGKQ0dkrvyeffMxGv1zAbIo4oVSLI7nwuAgNAWC9iTYrBd3cw41NijqaZMQ
bJ217ABWyFazNSpXYVsqKuEJvATQW1FXwDP+oNsxaZUsYg8B+JyYWTX6r8fqbcdpyC8rZbYjsQU+
7sVW0ENXlmLFkHQ4zggEokS/S97e1th1Cy+8tjxirdjqhsDQa6+vJHwd/S5S/HcSe+rt+XPi3RHH
tiTdqKMEqClJTiaklOhBEq6bWETKQ/Zv/P0984jA1y5AW39UMkBvUKaFNhN1LytZ1wtXOxToYJX1
VPY8mg2F0A0ycKkFmCsG1bqZAVElx2Hbp7jirs3GvGG4uNHRvNmT9uUn7ZksD9qHwjFY8iXbVAZ4
q2fUq27+o4l9+I3xKeMi83jfFSxaseq3Y/j5oYOlJpOV06otNNE+jlu8qHBbOaJz10wd0M57eWP2
1rKijFpSK2IPJcRDR/oh6+2E19ShK/CPAZ+eruOt31y7D7jnBHp4D+nIjtZ1uM83m67oC0Ns0qnx
QyWkGLRk7SuSOfVhX8JTC0BW8W52HHD0by+y99+AjZVhI93OI+uWN7w/0jjF/vBACPV03Ea9j8za
ejASSxqfldOZG1MVK5LvvmlLiabO6Wu/LNqMxBGE0ks7RyjG2hpH6CANsJD/+qaXz18/8tnSkWWu
iCwmXHUdNu8W2+9w/tGogtDKe1ARJfgUBCMxLpkCguSd4uegxYA+8RjvfmfMfVkAXJnvkUCDNdQS
oMu6INUj3C1myf+WX0goO0JfWyt2sDXzzNQg/gY+Mj8fEJOG1minkMlwvvMr2CRn+sh6amihy1BP
NyPWwEjWczEAlBxki45/rh/hPt5kp5XO6LSGxzklyOpYrc6deu9CN2xNYKoFSjRvlwNBNb/hJ1+1
rlKjubROxaWGJPQVlRa4HN7ylnjZBWLlbo6l35376ayK/ZTXwBEu8+aZpAceKZMIsIB6SK3MwXp9
nYQMIk8VQxDKZaj3vBn9yYT5rWTibQyHSwYOwj5xlRnXNXm9r7REjFmJOIsAALXAgQ3xmaCMX+y1
ycCKvpqVR2BQQ9Ql1AzS2dXS21W0+aJBiTGASw0i7qQ7XCXARZLBi9Mi1nEEhsnV8oDZSGVgG/rv
zeyFOnVIamvMNUi2KJKQ0G4owWTXv5CyUffD7HDkShCg5PRLdnM6uehVXb5pkmdVEa0DVRdQYlxx
NwSdy7YPBdWGmAqMoWCt0BYLr8OrfXK6GqC1Pvy4q2B8D1s2kevJQeUQz82eLkK6jMZKu0MI3J2G
VCYPvotfBFCYUBcrDznJOwdqyAdOR2hvsLIlJ0N4TQ0hRnLVu1xBlA7XLyFal76SfArnhIpl4AX0
PE6PJpQorhVFivLPZeAHQ4dWTwXS1UMy9ArHr1jwudriZErQl3qmxZISSXecgN1/pL8tz2vjz5qA
sKfHW0y0nGhvkjkuwDoEsu5qsOlzOq9wvOyy1qDtAX5oorGpxr+dSffsNhxmL3TSV/g+e1K67ppC
bdAIc4PFYHq6Brl808emyoKlMPuaR6XdwnKoyEHFwpqmECpvqXEMI4216jE4Wve74DgTkC9EO6su
ms+2//DOcXxNbMIUXLr4kIcCSrkLpW0DL8xSJ/n2Fi58Yt1QXpxKb56MHrFWJCrL7xECmvlQEKOn
VCvcZsXeCHwAPSnvrgboWptpNx9yCTHZffnMhq8zSkQgQHfDmHVpHbuEFilN0PQrhg9deKImjaip
Ldgo/zM2Pd3gWulVaBSME1dSiCU22lhk35T7l2d/BMPzOyu/QC54chsK38UOONm052iG2m3cJq0j
qazu64i2K48zByONoAFdhW3j1+hesInXRPoJhwhgvJsmwy9PAXkJRKgNw7qOJAQcixiokuJzCVoK
97QAo1Fp6s3TDra4Zb/zgsT5YL31kh2evtuDuGVPIGlp0MgRWJMVRxdtWLa6lJnKhzBmQiAQ2Fzb
1Rg1o4CsUhjOnIME1Rf13XcqAzNyrSXu+e6YKQ8JEnltxDQF2FPs37ZYqTQnv3QdnhvIzhOZWHM3
D44AsZrw1p9fKoPa4wbr0x1M0MOpHPa0o4xzn31uZS0E8QPJl09j6KK1YvffpJ0TnJbCXVRZFCMr
CoNP5GK7Q562grR2vlNXnYBWIhvYlVd2+s3zOLUf7miHrZQWN4GsiL8137WO3enu7cKVCLs8utKj
02krkwczyr+2X3TYl3NSsAdmnRC3EaN5eKRfEgUQtTE1q31QmYmF952WHDeMcwJ0RCs7ntirPn0Y
RJBtpWe8E9d90C4jQNLwJNF0RMHCjTCqFAcG1VbAJXwzZ7AMrNCfIkwhif+t/XSmoDsW5sivXLjd
WJhxRrimwEbyZ8ZlHT2VgRuuwRUlTbT6lPWJ/l8XMhS75c6h/9Jb0OYVn2+qGFkg6qeCO6PHogzE
mi/gNhS9aYz+3NI1shtJZj/DFP7I7lgZ8oFkAf3Pxy2rAdBCrOEPEHOi/jRE5xz4OoLatn+Mnl7i
nEuI4Ry/NuSMBCGtlI5pCoQVsyKV8f0UVhDaM7Ef7Xl12qMWFLlFcomZncTkwGfootNQ6fwooNQM
m2GEaH5+Qv13GV9xmarKoA++08rtGIyYk2aBSEBVFn769AOvH+8EwMkV/IPWI32fc2CMim3K7BQB
dPiuV9Bpv6oQEoeoycE1Xkz9d5oeG+K2qh1b3Fnt9sKZkZwb+BgX67Y5TWfZZcReO5+xLSqy4f0E
IZuCS78n0uKDuxaYC5nfkB9xNfk+5weP8zOtK5m8ChXEPXIzx9ZXpwaPrvT0oXYCCKD4K4rg0HbA
hmtiJfGEoKUy4s43047Df//Zh0iF+1eFjmNS3x8XrFaLxM8kBJ1dnHonoGrXl9RoX3AZfgO0eWXw
yRxZ3VrgQ0cATy7Q8B5Q0gPuMFWJDkAN4+QGs3Ds75JC/7RimHLeay9gubMqTtdBg35H1s+lprvr
caxFDIhkBMu7IjCuRoAw0yGdoFhP9fp5lN7u90hOw8gEOWEHq01vJuCikvB8fx3+fP1x+M90gDTA
xfr49HSvxodalI3BPUR7MFKFSgEdry8Hcp8xzLgDcoj8W1t3GSkVpVO6QS13WDKyewb7dzxxYX3N
7knzv1kw7mUrWl8e5KLMYDT5WTzsM9dZ3O2MF5c0x9fOt6VK8Sxx1P7BAq1dOTAFMq+fxi8Kt43u
hS7dX3zr/E1t0lNg47Lj+zdRDzqpTKLCMWmgxZ5OgncylK4xogB1GJD0rclnO33m5WNsFMQLoMl5
CUFwNJIjBB/rAAezeEN+iuJ+FUsmz3jhuX+V6hWFx9p+KqysfMqGuQYCABeEpnJOHbiC6fYgR+At
goTb9jQleBZmVyDZknX00eTlUtoCiOq6hrRkxfxpHiygzUTHTbgthlQfNIf2qoZnaKH1rh7pZXnW
7E9pHUuvE3i10I6mGkuli+hIN9Z4xtQLswguumuPsrALB96bNlOvoIxsSdtTNQe7P9NfKjtk6/0N
NLdcr1y4BnXwHfdMtkb2VhHLDpKLVQq/c74yk3V/xTyvd+8EuF1R1QehldOYW421gFd9ES22CLcF
arjSOZK1AQChh3uKRFUa1j2wdgAEEaApoNsvzot8J8qbNLBlh5hmKkZRYiDN6MSPiXgQwPPjMY4F
1Nb1K3t+ElbaUP9kOi56/sORShtCKy8RlBbzncY8MbizJwe+/l23SMFT5EIf1C010K2xLhZ12qO3
0Can6bUFdgGlF+qOqQtfxpm6C1gLV/xENSr/1qatYVQjNDZBqF0+wSl3Oo8DiewNit0oHhN4dnXN
uh08Xb9sI8SJXLiyUfDSsd8P6AR8D1WesBQZpWFvYruvDRsqYZl3231imrO0Qrn+Oxh5oiPlH3N2
onVumWtPcg7aun3/G99JV0C1yA7vgW/ksw/2Q7i2NHoahA3u1iJ3SCFAuAG9Pc0mjtLQuCI+7RJc
YdEG9yXlQ0ihbzmZW0cnQNwkISELqNg7jrWeXk3ZT3j6Ztc2Oo+jY80lfGUr6mRbSeGrr8pLGz/K
HRcmyZxyjhQjtaVyq7XiZ2wuTtv1Jw24ch76t/6UAj4/MHa+RRpysVVx8F0ih/ixk6ERzT3ARKLB
/fNgZjtKTIGuZWkbriuYH97yWWGaNGXoXygRgNLfAzGkO5RuwVzrcrPKyZ99GrSfQJguxCZWKHbw
c4+S5ix+Kfdhku6BLrsdlP3Eyv9A7Pw6yeH1AwwPq6pg5piG+Xe3avP5wCee2YJct3CsMxsCSblW
igdf4azqXRxrQtQwG4SztqAKIBnbex5YWN9jXShXcZVPH07Y2AExqc8QDgKEdrt8tYHdCES4OQjF
5vhEz7A9hGnfO4D+8X3y7b36FoSW0eK7tBel+I8+4JS0dJUsFBx5CyN+iCGYPOaxCKGy/a4IeJ/t
ON0uqBdbMkTpviap/p4wec/olhYrF6Dy6K0nu2948Jsg5YDKBOMANNcoT2OR1VpifTVG/WRxcFww
eNcjGgamp2VB8+oQWzqCBDmiZzW4zh/aHOY91jFiVCwJ1Xtzn84trbRuVA9swSZuyJYE+gTAHpTU
qu0iC7qme775mCk8q/H0DzSMsqhyUB1yYbdu8+vu8GcFcLf2+8eGiGpXCOHbb2obojx4vkKwErPY
vUSW5Olj1Zp9b3BDQR0bQ/Mn71WxAaYXHPn0XTMve+OvDJQYMGrwRTF3AGwGuQP1DnL1wXy7mAeq
mz2kPoY4TU14cJebJ/rZGBkrodbD4gWdyl4e+YwySFSHatSCAl+MTVSAMDovBc3/e06/RGaOarSI
WJeEoQI5ubEi4Kmc4jZCl7QwrBCr5Eqsq1MVLWD0zrabf56HeUrf3hye3RcA6tYP2T3oTgFEDHpI
lvhC2IniIKSZkGHBs5AofprvexCw+5AdYEo8iHAqMAFiYBSA4WcLb9OD2xNqAZmilpjTGkA9Sb2s
HJ+XuQFYhKWAfaAX7eBrSjUonqCV2a4hBkWaV2zGTJ7KqsWK740+QZINR8CsFrTJg5/6lKiRFQlf
T/Rl2re5Fq3QbsDdZfEtzocxLm/OZaZcad4doXBfU8TmCVXu4Q89ae9wZPnZJqv5lVVy2+vFxu3i
NO1JJfOLNUz/ijcYgXIFv46MmbzMa5SBHVGi+krScSKvNjOpqvzEKdrvV5wld7DVZmad84ZiHxbu
+9PlVb+qYXZ1H0aIOA0yMm6WhjI2iutP9KWz9mEMi2Zvt/SEaVuv+QicHBWNf59EiUWSMCQ03xrl
VKCEomgp2v6aa0f87lbjlpBS6DSYFTDD0u+J6PKZKo+KrhPFGpptOsyM4qVfetpH8VxjUYUCu91I
fDsW16P8L/2rW12EfpWFrq/u61o4+dcaFekRl9DRBEKuHHgNUiaNUJWB3pcSbEza5GFCBJJmvQKy
FweHUNHBiw/RjkZ15F+0QrziiM8xLkwD4T1itoD4Cf8VwelJ5p4zA8Yh9VT7Lr/bA1gBCqz2Nicm
of+VVPFqwWXuW9FL7qf4r7vX7HvAF2/fZlL668IxZL7+Qy5ongux76u/QBkU8wNsTzAcaauDkpH3
eRkZGXUjqXtkKs+4s3vUiYMut6UNFbQogRmlzP6qVrz2CY3l5+4uR5nPXqlf4TsuBCSXVJUyjFAF
ZfJKyffEfWFWei24XojrckYquTeGIgLjY0TlIGKBPus/7ytL1JrNs8jQz+Zu7uwrDrn6mi/CGjub
S+q3DDTlmo++FH4qja3f8TdNTYFkIkhm5OfZ1ZqpMbfAZMNIQ3+9iWqWT+M5lKB+dM6yUysVdVO/
5X+cADFnad9rHi4M41MRM4jNBQ1nugOLOK4vSXO9L/wCpEMlLq1hCA3M+FqzTeEOfO5JhaYmz94A
BUWB4x68VpNOFU8Yx2DqUz42XmpG+mT7a8cSXMOqkCL+G8NTSSVevdidSLF9o+4WvQVczQ1MzzVw
nUoJeWNzGwX1v491vmCEao9uSrMip06DsXCBeBe8/bKyH/bQ3qn0MMd/bsclZfysFxdQiC0qWcLO
G9e9abPD77drqmdxeR7w2uEqde3J31acJN3TTEJ1iiaP1tOQmwGZT5cvHMP42WoUY99EkOEV2P3f
CgOd9TcJT++LOFMPwL7QJgFaqMZkspBmwx9Yce9wSxQX96GoDhXv6auGg0lRKNaMU6FJokFYyhDW
qciMxHAwJBYrJsZIgXTavPnd/9Z9wbA0vtFOus6Wt4v1pH2bS6/fvQuPUkA0Ry4iwW7qNMqGwMH7
ny7uUhXNkBbcpUyiaxHk7Z5k2Ib92xWJ4+li5e5LMbGCbrd6e+wu6bpMkrRBwYLIXEOIqh2ejraa
KXIr0SfOCiSrXpO1iSm7CPf5cO9M7VcHL2+fqfSqLvhxwMgDK3W0F+wSiJrV6fNW9cmCTlKJy96+
GZHfufWtBOJQ5T+/8wPQsw0fllNB4E+oQpOc0zBpAZAweDGCwldNt8QWNcRkuxvWCGiZe411dZ/7
sVr+Kz/tKJ2mJ2io6Qx1l9oEJjDxHAhHOlEu8CS0HlOf9OLTAunzGn0pf0/yqS+FtNH6Lz1BD+NZ
dg34AoVpmDS8b8TZfQCsYvqLczf32w3MV5toQSnTeblxi4HOsXMa2gP9cQCwdnHkpjwB/QTkzUcH
LDxoMJBDjevxHNyBWhNACOdaA+I7eIv+hoPJkx/lxnwjFM7r0Yh5FS9p+tThSCtoPU1QZNq1862B
XZOt+gkwwdzkmbL+8pBBeubP4X7pkH9FXKE5txrhHgxpLNkQgiKb3v0kmrlRhpOJEoRs10qFKdaT
Qqj/PvXVISuROKbnvGVPrvX6pbJyjQYdDeoC0bt1WHURVwHKBNMnpn3XQ8As3MpBM7vMcRhZ1PcK
bJPbDLMmj2msC8xU9HbAwNTV2W5EEo2JuK63g1tiNCGvcNhULmzW5CD5ebVMUk5MHnm78Ula/fCU
Kos5BnfNy42dqeZ/L7guJab1h4qxs9u28OXyZqli6OWW1bc/q6oxNqT/g67rZcj0P/JbQzhwWFal
KzLZV2gp5gaTOVh5k0dPtCOK4vzp/e0n+8/LszSZKUAxLdZG641rnANy+DOiD7Mzx3mfcfxlKzXP
RlP+QwyRdc+Z92lcP9FloLWxXlTVfM9/oh61Ozt1WNIn6Xv2kRmDsnl9qGawICgUlBVYf/jjwRb7
5f8B4YgUXjqMMjmONOzQ3Ou8yUdYQ56NGhH/ZKB6CNsOHGQmDjv7YFaEZZ9u1ykxeg259tou2T6m
MiuqZdzKExFHvoc7vUi5t+BrK2sAZIWAp3BYEY+3zYBjny667rmljAMz+U7gv149lJLQOyQ3SPj/
8XkzJsPdXBs+Yz7zg4XtDByWkbOOU2UW48uJ8btew4AeaeUWAkUW2AmnVZRF+FqfB5I69QxlKaGq
oZCHjaZwpQbR4+BaURSoL4RLtwa7RpME23f5CdPJNlw7VtIrrXA9p1H7KuC2SIR5Y4D7UHrHcbgc
ACDrX6b/V9wSlw3hxIhYY96UwITfp0LoLcX06D9GXF2OtVmR9OzMCYunFKTIeVmd7TlvhbuPPxyV
qj9ku9u6XZesOazvr/7eK87k05ZYiI7R1NmQ1DYxSi/IEV1m2d+ieetTtYhjPla6NnXd3ORwA/z0
g9WnHUhW8qAbg/hjfjayiLMOQj2dsjcw+Ct9SA6+SOrQW0EY0yfMUyARlT6ovvJrzQ2MKyI1s/p5
k1yvDbQYDxlgf48o0TDD2MY0ixBlLJftWZM2aMKOfx9GTvYzbJvuP1yyKXNntUMiX3ANAEhS4MZi
BgpcuUUpMmAVftlOS22aSpnxdNZomhUzpYmWvs6VmDQVhSjekn+QIhFJtjQxyodOX8ZRCQttWCDa
eBF4UrGqQacQoKrxQ+eNxKxvYYroonfuH3A6gKbKliYBPnI2ynOHpQ+yIZsFNRYcGmS9EyedWHRA
SSLnwdEqQE6Ep0/9dfpa2chFtatQeKi6GiFKer3hyEA1etf9/CvheEqtEqcVAZu2LkLFwPbiCD+l
IEEoKFhhaYEX7/owDs3H1As8NZV8fv950ZV8T8ulpq54/K6d+ZDptECbgy22uoYzW0G3BiHpqI7v
moTim3Lz3aUcTbi4OeUYrzZcc7kFAcf6rz92kxHsHMimdjIsoYX+yMz7yqlrCuZ9aoGrS42wpHGf
dAUphtG5pMpkB+jYaNk2fOTGp/6gbya2cZmFBjX/el+3CmepcmeEQ6KpDN8/md17wQsM5trvzNSW
t77Fy1NKNJIvCbqezlrE6aDWzLl6BVK6Zp1Xq0t9+WbXjbq/pZDWIDp8AiAfuHlT0m5MOYQ5zGyb
iHW0NWkE1kDVXWW89oRdlShy1cdKp3bJhsj9Vbnu+NU53c51J3aTKZek8rd7faLIG8bj2IgiDbIz
LF7tUvZQIVJpMVk7NDZ4lhADsgxvnNrKk1lC3xFbCw90R0j7Ocb9/WESu6rXdrS+2dOYORMT6vaW
Z9HSqR8TvNZEfWFATum/8vdAlcA1O/VF7thkt1FXeb+DcgzwkOzfQJxDmOP6PTp2tTo82nfSUocX
f78wOYQ7X0XCZ4ycePP9Wv/VoWGcPA3BvFGkByGwCWXIhPVBH7cw1OSS6jVPEc6WOBJr8BrbWC8k
+QJxmc+oR7KzaPEL/hLQRNSQg7r6cpC0/dV29ZlUykmJVg5gw7uBzlnX1mGDx55wxOkHn1bvRzk9
/c7/zEHPnkTQ+OlLY50pRX+zESXy28H/+2IncajpGQjn9pJ9fHrylc21CZr4noHQz1xkutjJ15F9
Mpkz1BXNcwevEEEKQv5k2lFe9ey0dtKlyPg4jpb/STp8jhQDn4r75ieMBz+/+eSz9UhyrJaE1+RP
+1z8mgAgFsP7pynErwoGzgwZLlzogW6V8Z99aDMxoHTQrKcO35FoR7yB1j1IPtkt4umHoVmnxcel
2j16L2HAGoLq4JoScfNorY4CCzz0WxjABLkLzxqHvuHyyLSg0TGdRdWkDmFXOv6jKN1p+TEBSZoE
UOrrCJh/gI0qv20ufpsJlx6ieVUSw71VE1e0qegj1+28CNFSlDSEJ7RsWec4NUYBCeCPYwT7E7Hj
y+RCu7Zkx3XuIOyGe/QzWgSHiSc3jguOqXNbJ37hcfx/NUYpkAFqkE6R0Wo6+hN9pP+PX2tFPyFL
qnRxsZ8cxnaAWhLkbM3KXO0aTDO0F4/XBbW5kCNSJQo8UAqnAIoFtLz2QF/YEE2c5QUDV6Wo98xm
EWMZAF1mSFybp8oIfMuebp5d+U0oWDggXaEyz5Y+qukXM/ISdpXSZDtxvm8btriz+jWsKZuoPA4V
lvyof0zqXHRRhF5neQqAC4V1vVSjjESoWt1DyVxNpfhPKJ/TiPNn3OsCI7eXNE1+JzLRFTgJnldg
3BXPstHsBJelHvtaBzhO6OJ7BDpku6fkefCJHpe0hNfNhv4/4oAlBS1loJQYMaPEs0SWrw/T7d+W
KjWWNPHJV5W0C5Z6uMG9/sxlO9vtoLVPigjGuzaKRXoJ3NHS9YdmJdDNSB/9f8kh8lo1VgFEvFxc
nsS68UZ8bDzNHVm/18JaLyQcnOCIDM5Otquk8Z3K54Eq0ZBQaAhTDZLnso0f7wYPK/AM/fjQoC+f
3oGnqNzAbvLdpoeVYivACKZJCLUYvbTp30s8DADd5ki7ths0rUk2Xs+oBhwQYd4AWAkQnHiWmGZI
piHiI3R9ATX8E6IQYSsSnO0P2W1xmuWR97OeqCYICP7qPU4o/WocsQS2YLmxCCpofkIi3GK0Nrtt
QRLMtvyyVqdXS/cF7keOzNanMfkUTL1ySSyNKRcC43H1alF74UJQ6ZcMvCYJHGU2NC8H5mGC2zPO
Sfg2/Y6++DFRxSmLPAHnlD+4PujGZdee1DQfiG6nKHlMHt07mNiaGxFQ3LyouEoO+7PXHDjmboXZ
H5YDU3UooLymnlH4L6Kwir+S/fGNHSNcPpg0XekS8PcVLcPxHIlStjN8Oh//Mnh8UQ9aaGvpN/o4
4Dc7SlUJYWDg3i4yB5LPtPe9aYAV66xAMuYIPL7RCIoocOtrMXK5APca41hujkgQ1NSUURrNcfkf
9A08mi7A2cB6qI2/TT+q5rJWDxiHB0UFA5OX+rUG46itz/2uT0XVOPgSK0Mj/aOGFIcCJmJCcm4r
prh2pgxRyUMOBTsXXjFggMf2JJb4Wk9JcIddxSU+0uAeULVr7hM3IuQln4ThoxNA8H/rjLyo1coZ
0GUH/rBI2TPsDY0J+gqtexlMl/csDsC5unfgimcPRBo81H70ErIsyIP2hbL0f2Bc/Wst5A7H+X+S
e7T8RWf2nA30GS62Z2VoD5pKhXk6pMJZsPtsK7I4WSLgzev0y72oKwf0rSgeIxP5IAhTSqIfuABp
7AmsQGhwWgArMDcaOC2mWq1FurZXl0LJsdLQ3Lq1Np6qB/GF3Xg2qQUIlztrWA04OQFKENd718i9
iX+myDxTHsF0pwKOptANG2ZBQrGa1d531SAjkZBEhDQ9retkjVNUFPJTNk5e4xiHx6RctNDqKtwL
Rkz0oFfuH7AQgiKuhb6h+O4Wn1iVcPuRz6Y7sxPSrSGa2NVWpL7ES8O0U+blKUFkTM79r2tyVzxs
extS8J/Hr+Jf7GQMdHzrbPk6C8H2LHHt9xfxblyq0QBajVvGLx/hi5nEcR1uptLbGPPI/w3p8H8Z
jDDClQ+BYBMu4Q7yAmlKLl/UnGSYvAC6KBqqw0n9vbXlzFZ51j3eLechQv0WXo3qiiSRiQOo/2sa
n2gode4pVHtz6vFyiRSKoOHoIkyUnqLRGasQzXcdDVoKAJbqSnNQLFS918dS6OUpaymhcUwEVOeb
MsZzufjXRBNvUwZ2iRrCsWZdw+kP5UJqGnKghipb0yE65ciRY4lPcqJiRi9aMRXWSreD87k2L4Yz
sj1rXYrbHGKWX2Isq84MqKFmcp/vxuM6LqKC+bY7g6WgPHZZ2zi9AcjsCNqFd4hS9mErJSBixiAg
94HmNTcB6a5VQ8rfwgv9GM76dKXGeqbYIgUtemHR2FWP9UTIWgdBSrKYok1CzWNuKuhcQxwZWAZA
uS/TJ+7ykfnnpSPcqUa5npUedbvmniDH3dD66Dj3PhDuPClkLU12YLsTqv2P/EVQX/hSZ/YjzlW/
/dNzEj3TWsMdxgwRfK+Tadcgxi+0mixfm4pEuNJqyNQ2LmWy0kQMeUEj15VEryYflZ8Z0W7CR6Mr
sKSVobFsjz+XGj24bJot549Y1eWiv/7Vqa6RmXGdWdg38ESp852z9d8oeoZshHe2KYXPnMY/q9MQ
R+rp+QmEdcmIyNCova7v/gOKLovMhxax8TQj2H0glnjRY5ayfQfyLNuq6IkgE4bJSaIOBoHGKCQQ
ok6y/WOlmEkHOLvGS2LH5QkeXcDmbep4SlYp/ztzgrdeQmT1opVuvA2HzSyG+2ekir1Pu8natRhj
ZPEnKCXPzfGBPUwHnyLxBt8rfQoGLKU97Yu1HZJfzsFfyH4Efr2HpP9ca8uUmTUCcTLYx2mcYdOH
WtcSSw8RYvuXXaSzReCK24j/5JwNZ0WlADOLZ7+0hDerkvjYJX1IXplh5cHaDL/XY6Qfm2PEOKfW
xbv81FGE3ffhvAfN3DlLqXiC3BgEVtVopJAe+vzpZtqlqNy8iBXLJILODEQL7KR3bADlmN5Egmu4
ezVrjoSHhSI1hrt8uz2X5IAVT3twe8R12kdeMI9uXCqlJksA3hb1A37KSY5r37Nh9NOWCRCBc7UB
dqMsomvI3rCCKLELzOFrJPVmV87HtqNcWznas3r6//rPSDk4BTIYBEv7yxGK34hIqSI0VOB47cnD
PAbykE9mkWHdgkv60YPsr0DX6Zk0Vq4ufGN/ynzGZmQwIU4AfwtndbiMdce7NOgWpiF1gb+Kcrwx
4xtsKZy6/159fEm5fKckMjM6Hebthallm0ubZN0tQ0uJsWikg/i6pTpblNBO0j5e89ghIUZsqZO4
n9ABtdmr6ZS3Hg3hOCFAsn5XKqVEilB1uZO4OK3GQ5HZr87C1sAnNJQ8iVs36IlbnuBnq/lmxPFP
23T1TK/uGGf6GAxHJ0hCGxeGaggHf7rNcPnBBa2arrfUrtp9nHwecqLsiVrDRSbE6ScHR/iC+igJ
0RjnKWiR6QHnlJctoDoD7UV5THzAUXmP7Tj4WXbQ/xh0TMbzXsQDxodYBkIKtaWBRx4CqbbATrzz
6SrTDA7DxjVJxn8vkNSMvelMkwyqZOtugo8ffRaIjP4OjJsVCP/dXU68IpI4/5sSnkdiT8MZ2hDC
yuo7KsBMnEhYckiTuKDtsNZHCsjs/whW0pfNpxKNZeY032491VZNDoN8O7J1W+ROUEHNePD9shvU
3xxFEqeQLjFgp0uVJmiVptuD/9h25lgcUmEcvgVecxp79daQhjUW1yX2HaEKlhIbBYIdj470/mkc
Y2dcJ5ZcaOLgKW9FQehTbvueWO/dJUSGY6vM+hVK3yewZ3U73VZCGVOWIbHqUWWK2/vzi9NFa68E
bcn51gx64AprqKrKwGw+i47wxft6GTTugJB5/aQyLmJClaNt1rboYiTGoOccmfiOArUlIfjAqpg8
PxDYRbSpKl1I3Gg1XzBnwgwy4eTsne/bKkEgAa7J7TRyFepUvylWfFzK7+YHWeMUrLczQUHQ/wIM
2Ffb6sM+5yjEsOib5bYYYl3kMpOBr48bhhZr0eQv0dfToowCiD+Ea/N7dPShp6GXO+F8ak2MIsEs
240K3Emng7BVB2pNVUxTXNHJOvxanUi41+dWBY6kYKgsM7n7fjCwQl+vElx//cqlfsKRnOuSEmfi
udQXgGLFiSnxGRitNZwig0jyFTHDjyad64ZNiEdx0L3wZ8C0yi7Eay/aHXW3iEoo2JqnFGcvtQcu
O2cVhGFj3HD5P6wsUAbLJqzxTm6xNUYTbWn1sQ170tiB9MXrwdcGTpgQxarFyKiNbv3bVpnsrT6A
DmVoAB86hIkizqGjR+kmLj2JI0Hb/wYIHu1nlLO2Z/GFFWXDL107VbnEkLFNTl8YUXRECM5qxnzK
RziwGPJBqOX9b95lSpiet5dbLNLFQN2k5IjOQp+/TAn/+lh8KMLO7wEAnmIBozFgi0T6eD2KRAFB
S+Rrsg7L4ThC9mlsfwwM3ZTo7Grn45mt8gc00vCYKpIg+A3LSdRh/xJXmRLq303Zn77mr1P7hwR0
iRW2SXtXWxE7RHOiakXJYiyScdIagZKdjGNlJXWGlCb8sBw/elXbygB4pdICHlOYgZGlvjRb4uA8
YJGlxtlgB1bkqIT8ELSM7BkrcRF1w2EIY18J0NaB9g9NOY1XZpU5Vw1wkl+D+o8GshG7+adqsSf8
QOqLTBl0tlGPRrsv56g0ssRsK8CBpiBy1kTANwaKi/6T0K2gX/3EudzBwk9VdZa19qDxicUXoVpy
OAWOPb8IcKY3AJKNUrhh14+/F0FE2ltYTZcAz8iXvDtgfu1UOcQXaD8skZ8NnNxzu+Jb0JH4kmAi
MmH3UQ9WVMo1DojRVwSVV+yT3GAXobRtZzmUSQw3k1HLjtld0LomGGWzQ4DPye8lhZTagujOEAO+
anDbk6Mta2K0OW1w7R66NShx4UXOGU8Q6h8H1NTEs+Snem8qLzDuGyq8FgHy9j93fUm8QF6F0Z0J
1MVpUB73Wt0MFG0h9Mj0+y2THXTFWw0UUbz3szp51APdrWJuvDFr/rSZeDiJGqq46wUeO1XKYjcn
SkGEJSP8C7f4IyfWNJRh+ROgBb6UyTqw+Kpe/4HedIXJaXF6vlcMwOeK+mt/S2kteHfUSIKqFHSW
ru/BLOCs5O/icJi36ucQaGHZWKQMOnHu/JJn2YYASHRyIHKJZdv9q5DZrnRTBGwnYYZvbNS54NTZ
ydCpeztzXRwZ42GDjO0vcj3xpgd6c5GC4Is4GdjAbwPvlE8ldQKJcDO3DP5Gi8cNgvx9pGEOq3dp
XJ2dnVwJA6gl33xGYT+KlZJkUnCdU2d5l7QiJxyNQj/QSX2qvp51NpOSvV/7loZNGsFePR5SrsCX
OpbsSxd5G8C62NXWlAf8r+X3tNEJnPm/1hFmPlc8T0WQjSw47v/87EMZqXtGs09jb547zXuZf8CD
mQOdbM5ijPrLXxlnepIDScIpFS8GBgXbItujU2PjpnfrA42LxZjbLlRsloBDaQu3DsY5f82DOmAa
X5uzUFJp7jb8rzTxRo/M7xFpnmjzJfGeNIs4/hXXjIAgbDOpRcJ4LgC+EqJHaEZok5P2SThwB8gc
seJKWKaIaY4zGmmcCX2Sz4FoccIJzjAr1a6IOxdf5U7VnaG4i3QSXiL6JEV8XxnsgwBT9U8HiX7H
5Z0Q8nrUOSQ7aNkKgNXHrRHw67EI66Zpkq8aGULjZJU54beOzD18hAYIR94i//d4IOqdr3epMF9L
aMuk5/CBM0X6bol3PwYhEj8coACMlZgPKcAQ07P45S7DUjXv2ZSKF9bWsD79w4nHqMtcTAxg3jVe
LMEJMxHqUkQPYfWmhWZOqGc4tu6Wonk8V1COTWfMfbvT99rPHiCws5yB9iArID/c58k0OlKipbwl
E/2qR7qH5YdzqFcH2Tmz6VLZ8wFlQEWOfsremEYI/tG1IgXcpGcxiKWeHYn1Ddvq10aFPG9j+9R0
SJzaez3eI08TvrLST3ToGEWqcKsTzodZlzhaIIfSBziEBnU7Xjeou6ceth8rWc1hjcquAH9QicrO
BQPzv7zsMI6V8NIS4PSO99PgGoquyHXnihWrdn+yFJa3/vYNxr6HN/gIrCUln7nKghqC3hqQgStu
vWxtCaGHY7EPXfkexXD9EhMpEnwHzkmSwVHITyzg8SNj3THchU+HJSPCg5NiN4/zdxCc9vEHEln1
xme3bzT9qZmO27zxK6L6VU+8fwCPeCVDMYzl3uJz0MvwSXa1gdnJmXHzk7ZmePgfLDTVrzSixH6e
k74h2RYD3YVvYt5nvijd3Vz9ycknBkbjYVHSm+6kXcxhV/iFbv8X/QUkacybIFkDIU38DI88gPmV
YXVOA8QJKmbwgjHOhT50EJxb7Jth2GC52LJROZFzBDH2JAv7g9XaB2xUWpzRryvkdMZjcbXO8rTr
2rVFHDN2Pa+3gT5pkZZEVriSdv3XDG5sln9BWuOwUQ/AW2rZoyP3hY6doH6NBuKjVlg2guQZgRHK
sWKFZrHEX4CoL7zMMEeFbxmL2ckHydYN0RSUleleYS4wQvwAaJUTXMCM1rx5rb5GEc95oQqg3QTJ
GKTbahLa1eFZDoFUzeVpN1lY1hoVRuBs2hAnJYZ62MSCkaARudqazv2kwveQAXsQOdlwMrhYq6FR
3MBmdpB1m6y+w9pMlaaolUAPbHZFbeWsHHPM9kFkxs1rFLIIAzlsbKqpG5pLhyYp5KiT6qJDgHQB
xzVKARDhO2jIxrQmUVFzzcSi9Minj0/1/hMw/LMQrllcm/f6ChJLkF7RQ/QUAxYqWEUhhmkbexb4
VBKVXFMkQ05BAboXLAFvSN7w04gJeWXaxfwY0yU3epZPiJyZZWPvxzweDwayWVG2x+oo0J35DRIb
RN8nY30qpBHnlpfB7274xb2ZhMeU6POPvt2Bg9Ja++Tl08UQ+AmcV0Lzi/Sx8sJcXsq5aV0X3h+7
jX+um6ggT3wyVusXVuVKB2LkL7ZuLBIH7aFw53Q7eKNDfMcv/KodAvWEoJjLmjWwL/iqZPwuMsmb
fYyw+nYptx/pfxK3Ne5ShcW1hj+aPctINUPFZRial/gdcLalmUH2+OLy8+GbKtuVP5rwnMBC4+HF
ZWEQaBgOrekvoGpVMcbt4YgMq5X91GG4+ne0sVotsDtW9pE2f86miEGzEbmjNmkJXc2HVlN8yS+u
pxsL26zldOcn/d+bq3ZBhl6KHzp0bs/KNt+736jvk0OX3pJ+awRIO2+WunWvzG0X61CCI/uWwFfX
6RgcQ2UUnpzZq/llT1hEfwUxvItBFxt58FKrCrThqBxf37r5y6jy5KpPhOp313I3/Xpa9MsvtGK8
g9uZblm9yoHQdS7k8JsscOXQaLtHA+JTSWJWC0IrO04uQlg9OpjCvQTDe0EIbHY0yrrRukwMAGpQ
wgHwQgzAplSEa/XU+jZE8MmXGVHw2GqHX402VmdLxapKQSyleKNc2ccTVfYfUsbYvlUuegZCXQEA
EF9cDv48azZenR83d+qRb0X45p6ZamTt1c/P+Q0EzEv8MLwlgb8syRpcVFhF8fihjheF4X4mGA1k
Cvtb7YDuudD2RVTmhiVM9NYlJO+Uo2x0Z992imPKBMDHMYmZX1tlO8x04fLl2uUJisIHwrlkr3gF
DTrqnIh9iHMWBtO1rCCMdkatscR2i6wkMcgqE6mJxvF+6PyoKHLdCCtAzPhiejPjlB6lk31zVILc
IZU+dEMYmrrPXKemab9GRNAR79e04Rh88GshH6YASYIKgNIfIrcOZqCiO32+y+JJ0tvVhXtQIqWB
vVlhkbreN3jPn5n/Wwnhpp9KwuPSfMxm8ObJGH4sxkoVAZEM+CvHsG1UIEDRypiOWCO3kZRqubVL
+Hnu94VlLZYUxmD9iWFVRwzlGNrZT8vwBvPHEWYplOq0gkfCRMAnPeZztEwRWXLOQ66Ml67a4axU
mVoNBidy740lBFqWXLXjsrgOTqR2+vFKuVsGTUGq/e09ExVh13iz9s8miaji/d1bD+eavgJFbWmQ
HnMM3x8E4hEWukE4VIGaV2LAaIkPq8YimSVlMyLAarUmfgCIBGyY3JuR2PnVi2YSUtSvrhFLBVIW
23x2xIKXI7vrOI/KowTqL3T6+HEGqUibSLUQeyWwiVfDaoVo89lnjM9v6wRB6zGpiKRDJOiRkMlD
0ZmYfh+rcmmYx7MkulYttRyD8K0h5NFYRzm/FeJwMRUGcKfbz1sueoKuzMPH/dL7mO0hil4m608/
Vn4Bng3e9GNQGtAE1SDmBUOEoq9vRqMrCmlAOwDkjLAmjzxcnGX22qloKng+9LG4BbiPQCk+y3Oi
PYgGBfc09kQ1cYxckLZOQrqHe74rxzCBamxmSpvkqvzh6Tw6JmAibA4qditBJrTYdIN2lKjODjgT
Gu0uw0POl3AWZzPKlq2fc+kRO1bN4u3I05PH3YMGDeBBBT2IN83RJ1azhCVMdf3pcWUagwToDOQI
g/B0XNjqF5w3TsacdPsTiPNSYRG2yf74W0mWZe+xQ/fzbmGeWJFyzQAdTiKC1B7FQh29iOA7lhoF
j7PQsab8shIasF0iF7yr8oErt0yzxxnlMXn2S3am8AlaCypuMKN1ntTzJmOAn0NtyptK0DEYDWeA
BnHvJNAUnyc3oQObDqP4TZM1A2Eo3z59WbjETlK7Ek3567yRZWTYXY5p+xJLGh9mCEpCR56xgLRL
JqG/DtiWFtgMeVdo24cK4Q08MJfQoPE2MKu6fbrnlbwge7CqgUWlwEd4swHG+6qC8q+i0m+Y57yb
W+a3K6zk+t00DC8Ho6JewRMKcHVxjhYbDKyd/p2HnWdy9Uv7zsQVDP4fSCWBSiBD4QtAKNhZrOrS
LTbcMDNg97dekorXPFZQRGio9AD/8ozF8OF0YR5ALE9AhSOBu988WKLDbflmLyCUxZwji29ma3+9
u49MlnOW7wQ7+nSNjZo545PXm01L3HZhGZT66gy2Qi9Y5wLmRE/jMbHIhmsf8Vfka/E1AtrTRLy6
KhhswMEmQIxW7QDcP392ylea462HmitGJuP4oLaBC2NMLxZNqx8OqMe1ilDSKWSKgyb0rhKk8Egx
EGRySxil4Cg5PDOGZXF+qEoS48t0D9i+usdjLdNEPMQYlwjrw6/JrQJRfsPx2+k6AD3Io+jUnr8r
G35F5zKwegCjrVie3feIfEfqnO2QW26ZucVuCl44DrxhrAjtETRWncf2eipdfN9mFA4XNETDYssd
I0NweWmVwcYqhf646YqxkcoHXq8spzmg0Eml7umK0hVbLv77mJvwwPZ30vf2TiFRD4OWzDgHPr6u
aF3ofsqJDcR1XzH15aktPLgUQtNgJQvRD1J+2f/l0X4H25MEk+1pHjRbIjlpZMLDtfjKojf5Ocq1
lBvaCEg2eo4TNDDa0vQ0U79oqCD79ZTwtkdeBEVpTKbRP7plrwV8vV/vcVn53c1MpFSCv69/ty4J
w1/whOxgTqrjb1FEX1D1QxmmngT/KNwhL/tVbP44DVqxDXMQWbEn6QAjPjPmiUlYG5igtJRpxbYU
wS0dEqXUKcEdP8iPEAB4tH2kwBYUymXauh/+oUJ5Tz8/uMj1FsnvExSFOrFqlN57kokpwq0YYx6F
BHUF3OVmzWAsjgP65d19X6sI2+a1+kGDMqbT0PHwy4g9jmhAyUKtH070xUi0YZWdewWYI8YrC+s6
tYMoNFubIIn8M324tSUj83J5DM2OHqabr1Wv/ckgTLwTpFKJcRW7d9cjHCm/XartC+4mRTz68Rbg
Xa4q4c9EVxIoq+ZmHHYwdUfAm6hHP/3SpzHojQuYQAQ3fklocSo0zjLz/ozRIg3T15zZ7WVdi97c
XvOGcuUoEA8+FvOMRxs9KzbOXW/y5p5kunRGsypJMElijG5zHkbmlPV646JGyf8LzYgnW+5EDsz+
eozkuhPlmvIGTVkDgpAT6ajVYi0QcN8sLZCGYMLJuJ/o+7aqXWTGtwocDBzwePi7KNLgzvJvE6ua
0Y7M0HFDoLBbhaHD7al/mLiyyPSckKhk26uolkPtiW/x1eW5q5mIQrwUKCGe7+DXxoXXd8RHJrVu
s2amgGigDFoihuGbDmtayze8pOzKeixHv4eVQRN6c4OYatgZbEOWmT1MW3w8ZfEXEm/ehmnE3l8e
JTEqbjDLDCI7hmQf46tAhzZmq6NHWorWiZRQhf+/Zw0ptNrk+21M2b9jcjgl6xEffCpfFHAEodos
wQEdCq7ittlMrp7BrDw2mz/Sum0UV+7OOUkqoTGqvWBZyXJLqneyLEpt+ZWNSoQ5fjR4haX3CvDC
XbHH8ouDQ6sWnIwAZ40X0v6I9FIRK8OpWXCH8NTjWzAmZgwN/cvn/IJ8QAvUlY7xfd2/iNtKf1/d
jQk7toFI2dOdntmi9D6dlxIn62TSSyqHjH4/SnyabCsTu+QtHxRQ+3Szy3veHcavtedJkX53Zm88
xJQcJ5lyCZV8fp8SWViBtz2tJ4VyRVAYCYf1CZjSg9iyiUCvPmgDKVhhfTCYHZt0Ug1RmA+1y1ZL
m9176fmy8jv1NYumkXE0Jm4ykmxAXspJF6u2SI4CCZxDUfIg52NF799Ehw64+w/e226/hiLQpIeK
CgAPRc9K6SYxTDdHjqlePmH1vOXBmcJjI3JgRWQ0AbUxN2ZBeBenlgw1M1tJYrSbe9hYKH/upKjf
0FWzBP5PdGwlqi5cJbgiSGfQdnjGH4B6v8IJtMnBDEhuN2OOI4tCKmN4vErYEe/Q0Rx1RU8fB2eM
tF7A6zbGKN9B16TMniCd0MBs/5oq3VMClnK34rw8e8EOvXhp3/Fc2zYXHJCn8/h3lde4mbwz8LTH
eavUlJUaC+7Fn9BETwmziXofS4vCXnm5R6P9QmgLKY2CId2Dlo6UIXVVYTrYD1feJV9M6FpBsxHX
Kl38y1DWFHFLlkrlDoUJjlk7TvSAhbfCtGk2iPS1BV/UzH9fXejadjdxbMRFU516exDLU2Rdstly
tPUdyoiVM5xU1DOWjWHw3hije/KATGxn8kaGPWkNKo8dbu2aVAstk7npbwQsh1IhClkpFQFKSTFm
K4c62XlIVhU8JoX9RKG0MuIbn0wg7M2gY/+8S4Bjr69vojj3UZihMPwH9ZTEjBC3yEu9K0QE4ypk
KHDahWACR476vhhi4FbvmXGObiDI0YBy2BAkxxS64Bdvp6TjqvvAa6q7ndJeP42rMcD143iSR8bV
PfmkNQy1yv6uit70EO+u0QXfI0orUB20Tp0pczhbn3im1WvOqWOAklzPZDbZI1DaC8tTkaaeJ0ZC
WjRVsE9BAyMyMOuCzaBA86VI+nisTgSGV71UfFaJG/OT8pXmpBg6xH3VJZ6Qzmc8VstnR+0dkqKs
EFSddxfGd78Sjfrvkiwo0FpxQB1HllBSk7/kaiTnkUw66hGflBw961DJRHQcfHKhBcIPqN+O9nFW
4ZdDBpEbMhheGrrRZjjMs9wKx/qP3BXq4JGGEcz46WfwTXbRvsZPL4UjYO6bArtL0M9etNiTMqV4
K9gN8UQSG+WiaQyLxWvB8xF4IJChGFxivWuLYWCTBP3g/hiLXKimp9TOuFIQAg6Yjge2c2MkoO+5
cCv+JTz+1KORyNdjAewNqPhzqoDgif7bbD/Wip+5ohFL9hO3GnUIrgFiE0/lMQfgYI/yJ5J6mxqs
j5OZCNyFurcHun7wOuTq458+iI2M85JbGr8UrAL/j3LFeTiRi3qtZVYKqCrLDYGA+FO1BZ5Anmj/
qrYJDMYCfWZbBTP6KD2Z0BcGduWFN2ajvOjfOAPVR8I7PoKeWhuAGEKHChngxg4X38z+VWMTyxEM
LB8/4tBbcLKd5TxaDuJns7y48HiOrnJpjLB2n3EJvQJiOb5AYNtgb5hvpE7LYiDkbeQuvaQTkR9E
/zrmqhOBcgzL93zccEXsm3jVcYNSdL+Kjmqb2lJReSE5JGc3MhBZK03lbjQ4+ZgzpZhU/UJ6ApKx
gqv9Kc+Jh3V/yX2kzRvZTZ0LStwcbW2oANNWIqQTrlnX7xXqfoD3yTymHadp4jKrm4LiK96m4ZOZ
txEIhLcG0ymS0SpmwMk8I8wmHN7gnbhl1n3d33r3HY6EAeEdXaz+QswGzw8fABgtrhAwzER7M6Qb
qiIvJmFnPECdBMMdSJ8OO5H3wXkvBwoReZOZtXJ85338ZuPw8On7kBQLucHZippMpBqa3MKTUTZO
tn3EOpq14pwpRMkzSBgFdgVaRdY7iIsD6HXrqRtFFjwtUnOp/UII0oW4QGjLHW99wwxq4mMMwAzC
DGf9k8FC2LYpUuiGjsMShoL/r9RSsoCDihxE+hqiKsaGiWuIW1LUSDTj9W9b140XxdU8ko78x8ni
lQuSy9duE2mwxcIZkRKkBMinXkGexuO0wHbsyKa++YSWtfSeFff1jXmXn3YKKDJD6x6FzaDLTYEm
4Ry8LCruT9Erp5956JUusCPrtYR96jzTGSpJh3YqPIwOzo7FoY948X63TsmhoszMHw3HxG7Vw2Eg
Ab5SryVzAvvqB8L1Yz+kOaxCX0/p4KnhKbBbE4GOi2Zc3SzBhuJs2VpR5fLfMjVu9DLwIipTetY7
Hr8W7TU07CU4XyoO40aUIFefsyyW1Upfcyi2QWLSBaH2HmgahqW8ODorBFirBqpCDvZsGpXNSWIr
b+b1Tu7ELdUc5bdtIsJpGctm4a1iw9S5B+hQz8TEw5l5rquHdm0sFjqoR+SsI7oJ76jNZkU1cltl
qShyP8N7Kp8XJojVc6u4S6ajUoXxwAiH2NjCS/tKmgtkzuRr+wYtFtbCROYq0ChwIeSWw0pEHbWI
NhE9NWy/xojptu0p4qUJL4yyy+6ZlVq2baXlZbOntwnvgcmG12zh2Er2S9AjoYm+YaL20GANYhuI
Hg2kZlw//GnLCBXV3s0s/MzpZ4UexXyLeeVwvlgYHrsfzRNY/+8d6FIq0EuLjPKBTcAYGyzK25mE
618oyvkGsMO+P6YzpVLmT4pJhvjyu6zXmSdhEAcTSjjDcXNalk6puGJa5c+GSuhcuPOfEIYDyUvs
t7VEM/v+KXshS9qD+cnNA1PUmIZzX5oqBD4emygluacU6M4dFCy48Wd2bVyTueK4V1B2AiTf/9LT
4/YNNIMUTV9IUxti6yrG1LATfmeJYuwG/oc2q8pfcJq3G0u5hP9hIL/PKKRFE0uOQAzlo2AQzEx0
ouC94dBRYqlPNcCNiJahwzJbNsY9ANF0PQN9LkY4ApL+GjRqhcA+m+g6smWcIW/clmN001X9lYgL
Yi0T9cmElE7jTEi7Bg6NhCbzopc9SV+UsN7MHiP14rgYry2oxeis4lX21HspXRYLl8+7hCfB/10Q
fuaOlSNAqpCrQHbYSJ9BWtDXyYvqLJcPBunCmcS8UtCKRV9Z+1fEj20e4QRub+5WmM+keRM6Sj1I
EPe2d9Jcg8U1FAhwwF/c2Qyj6HVVSPCC2SC+YcmQ40RBGJXRciCuiz6FEqRW8M1f8+jXnZXrsuqs
N5vSqAeolNa2sGF4OYYDZG5gUpz3uJ36m1Vsk37MKSLrcSnYQeEHm1Y2FpBZi30zFDQ6fg+HBJjZ
/jDv6jZ8oIrX5BUQ0pBd6LF80C8iS+4tDUjeuxd8hMLEVX7McFRuN/mI/GkBV/2/AFEYn6w3Uul1
nKEt4R5hb9NRT2HW4vWaU2EAdTjFE/9yc6BRhlVtFXGTnqzQ8MKi+5akNbACBbYLLCmGTC7uez2X
FlXfJ+wEuZ4Dg/S26Rf5VzGIrDwy+lUvLy7QAnKx2IbqIYHfpoqg+XHULB8KzGDxo5pi06klcThz
ltfZ5oQ0OMcumUSPgeZ4gnt4rUQtVxrlobjyYQN4ODXCcdc6/BzgX3bJC4vbx01F4K6cZZ3lqyRT
ZjQBfmEbd1FYGRdUi+SqAF2G3p5CcbmVuqLMH2CgNI28cWRU3iqk7mcM7FIBXbbp97G1HwY6b0Ab
qrNIJm01ZgN+QjeP/L+xqdlECuP6zZoyJ6/Qj458ymjASHUT05x7xrxTQx1gn0BFw503D4gj9iFn
zQ3nyJNdrahdY19BZ6CpEWNRZMRzC6GYcb4zBW8cBGieI6ZmSR2NRylkaGN9qlbsL/9GI9YjSCy1
y4Sw0iJSBuKLplO2/BdffpTqC0aEEimAbzN5PpzE30+R/ZW0xbMVzroXQ/Ly3rfJeDCipzn6aqdx
4c8xtjujOiHr2CSVHG0Wo5BQwRodonesboLw18CKEB0y1qdH3rVRMydAfKzWuBBypsAUZNgxMDFP
SOXX8shXHazn/EtaNeQgQxS4KDzqQzAequyEkNbYG7kcR6Vj+1Aqlo28x0ImfiHUCuzFxL1aB+9q
51nGbLPrLBj1e0LadzLsQrZCm8NAcc/NUDLdzOFwTrz9cUe1ok+ZHf3v3/N4fEmQy7PdIS9dGwUP
/WuTDTk36zJR1yMdUta0k1q5wSpim/FtHHpJxrsWEQT0lx4sLhZ0zz78Ucn5mEmOmDuqgU1g1ro/
imOnq184ef0Fh+/jXAGUmSuopZ1gnG7EDoWBFZcFlAascFwAdHnQeb9+RD/8LfNdZjBlKzDFA7FP
jGHEFXBliEOzpe1n89csJtUmH7ZCZElNp0jMCkZb7HUebPB6Go51yMR6K42V6810VwaCv224pwil
xNLyoXcZg7C0HoHZNY1YHI8x/ayS7IXM1QYfiP5H6oKqTQESy93Wu/s4puG4aYd2Zu/zWioNr7oG
xe/XV3roQaQ1JmQL1vQ/zXFxqhNs1PMtMTqu4W+NCQQoC71JGWwdJvk47x4Ivcb7NwbzeKNY1+Qw
mz4GyT1LBHy5w18+TzzxA4mY+6JexQ640HpCugVkfSeeatrCFYIbw2Bc6xLs2s6L7p+KuIOnVRB1
/dldYQLKtno39HbMKIRKBCP2tQUAW/UrZmN5es0SfkeBJTNFmapxdFBcaJmS2JFUQVhVRqgNP2f8
+UeQMWNCcKIi6a+YbWbKbTRf2r5pzQXzU2gASN7ir7n1Ka6kqPcOmbiIbNa7tHQNVArIgi9fqw//
TcyCqBU1HIceQ5IvtV3MCzQBAtrztMmieo0B3VyT7L7Z6C2eWyHYw3r47FPw5FhYMfy88Oh+CSul
GNdm2brw06ZXTkjwj4dQ8CgxN3wMsO8nUnxBZOkeVe1nBPRkIDb9p/MeOoSlQKEAc6vBvLtfBwJx
M3VjwqcNJw1QOV+cqO+VVAmwESXaHFJQnFaFBsEo2SZpLYdUHcUL62xeWVSzC3jXrvJh1QGt4isq
pOgUbEZeCi7+0c5ZU6MEA7SGnYOHvdv1jmeKVvr95SSJMAmVE2CBJFEvZ8aVOq2u6hJ3R1heQIGh
1AL5qchtzVe9Hy6ZR/o9FAla8VG82d6HbyCl8U4ij2pUg55CtZNV6aCeB+roe6MD3mmK/hUPSs6F
8g4wvVaT1/lnpt8wQryhEHqAIml8eaB/DyhKw5rulntrbvBNn2S75nhJoBNu5OvoNq+Q/C304vtg
cLWzeRaIyjkpu6r5oBPJwf9QuDQc2pCDqiW4z5a7FS/fJkg5KHpQJ1iPSbCVPAoYJmYr6v5ZRha2
7nVXp9r+ugOBTL3g7j/grzd8XtuSknARNv8NP61wELxXWgHCDnLc4Bd2GVVqZSs3k+KI1H0zpYIT
zguVmxl4VaJFJgnIy39+sYYUNMfVbI6GU6f+45BR0F+CRddyfx4aR425Cn8cPLL+dZ88hSWlhHGW
z6DM2VafsKwAKS1HJuAH44jVUnS17YuE4uOLeSrj4j6BNjlBP5WryMnegL+aI/MgCjXPTsYNzzc4
fVxfrzwa+Ka27HcDnB89Ht9m5S7wcyEi9bVHFIchxotY0gNrKfxgJImkk82Tpl66+yrZ/NoTq5Rf
Q8K2na2AD4UPlHASoMMNXqUZHtVKZiweydggebt0jt0Y41VHgIkRdWN694HZvZjL7OsV31LtOdE1
rW1CiAGgPpfDC/A6xB6/EEMooWb0+v7kO3AUc8Lqa8pQi9+bCEqOvAPEzE7cmPpZE80xz5hFvEw+
ErrQCw4RGffAUOi110BEkQWaHh1qfRGYxbTMMnIvcNBR5XK4xt3tY0/BLMTgjiL4Tv38XzOJtPIh
HJ5Hk4mlZOa6mhrIkRivrXUCgiSd14njFGqgfH4BkNqJr4CsEPRKfeo0zN3PeooOsnCxqu3/Es6N
o+Bskj3kLzbMUUO948P18An5XQEWGorUK1wI7CXbcrxzhtX036dfcMXZqXRPtmJB0kq78XkI7CxJ
VAyzIaxDW4JszGtaBIAkAAWmrxQIIUN2brnFnEbj5/Ch/4yrGv25BpRAWfrT9rGxRaMhjDzRJUhb
rXG5n1XIgziCoeaQ97NYnz2PDyyigacvag8bKLxW5ejYfBTUEBP8MXxOSHNzGnxqEG3M37bQE7zR
KdvjQDxdNiaXAT1JbbHTIYP8ghi/8Nf1QHZU0zppJXIcW18MYvC+E0kb4Bb/4EFXiSQcGinPxEsl
1xsVWRs9giRuQoyi6p8L13spYVoe31q3g1Yzzn5WzjVd/wjG9xu8lIDZNehPOCYMwdwBNEpxuH2w
mMBYQ2yMaQPbUJ2iMmgsng6mAwnUg73tfpI9DvCoOU9GMCIm4unBh5Nhbb96csyGU8kHGA83iD7/
R26msbb8RtG4uBTYagC+xqheKXT+oZwGkrvhP2sOCScCuqckOuvUAYbLN5UuWxkFW8gKe5ggiqVA
b2QjFX9MH9VY6IJI3lDh834KzMrdLt1TiVlkwKhAxy8IvLGlPSbesKrok/0HNoUo67dZHeDCzyLn
jML/vfh6/YOa16l+sNvPwOLFQGvYGgUvb4MD0qN9L5pP853haAlT1akb2mhq59Y9gr4NhZzDtHFa
8ucACfQplM1x23tJK9qw5jlvWd3Pc9mSd60SnvBG6AVgdqJIFbZ1P5hQjkTEd479K3wYoTmmWC98
3D+jvky5d+F8PXdV30FKAuOpTL+IeezyMyR9htFD6S26jFqbkDwYdOoMxtEt9CUAY/3RDIVuX7DM
2LGs5kuSs5ub7PrPyljxDk5tLft8/JLRbz/3c8sLUcsyYQ7E7tvRz9uJyA6VZynfTUNkgImwle89
1oaFXOwyWd9BhrWROWY1Sfl2Pm03xuNHBZVcZW7PT9n/eqXPKNajUsTHa4DtsmFngLQKgVx4iBaa
5OuNDDU0cxmqKG/cc0lswaAoFWGQrEV1WKO7XkYoWE40qozj1/vFjgrZAK5YKTi0S1ZXFaum9mhU
0Oe6L4PeN7v1GjsrBurdS2r8668FzST0QJwBpQL83/B4YCudM9wA9O9p3AwKtZm0NHmc+2ZA9Sji
lT5dVBFs02x3/sH/63KdvRmHHrtmfaZ7Oi6ImMBgiWYmLSvmvDVLpRei0broJL9IHkU/vY01Usqh
XOunkLjU0gRg1E30adncVmcwIFt+XqK994ASI5YHVZP2Is51oN9iwUuG6vqd4gjlLSRENI3wBItU
S83FkNtAiq7DB3/0MRZiDUzIChV1pvPlk7uypR9goW/f6R9/wBMCIPj+ouqcmsotYRKUVzksC1Al
x5ArrIIZQZMoRUIzG+xV6DS/ItE4+XkPJi376Ku6SLh45Z+37EGWOmCEbtYMavg65ybEF78A/n4V
9nXtKlYUinyV+XQ9DaQqvMuYoTuGj/hwLdQ4jUseCtWDPAgTy4LCWGTwHo9Er05EPww9hqnbPT9R
rnMtbl3LiYIB5WIPeovtU4QYMsmyFKow/ZmV2Jw/nSXqgueyfpCWn65rwI9+zSSMY1rnoMT4xUvo
PKV0nYBjM+Rql2eiEFlDFWN3fBWS88kNZ9gtOJSTCKEmZw/tLcVWVbTVYtqqEbsPwQHllGhCTOtH
j1eJ6vQEaA4cIM3MLo9gVnVTdMvJO2gqy2Zz8kiizsWMMGIIkoxUvo27meQ91kK04RsCsNvoC7VF
3kagfMl/f8hrXBQwzdiArQyTvxvZOau32aUohVHbxlpNtr32GosmLp+V/ibdIqrtLkKpn/0fXyjy
MBojKwNarRWYij0hbbzz5lk46kx4eIKTgHi9bmn9AdZyKg1gzYUgqI3psE5vqU+0amNIELEAoa4Q
JEmt5M5otyogzioozggLI+Sd+Ik6Lp6YnJwOnZYYUzlAeZPxdbW88EYjVsm7T58+2/1DfLkFL/Ui
okHvca1Qo5Ynmm771khQhq6ZK3T2mLmHL+ts/ABipoQxnsY5C7ubiDqhfB+tbbS1x5XjZiQkV+mY
kgmYUqBk2KJRj+fE563gJCGaOyoMkhldtUXqk9MihHrrKKONXVS+1K2gs1RkyKhQKBMSfy0mxKFt
sCil3j8y6A3scefxlYz1VeIucNrqSxsqCNsDJ9CbNlAfdKijZv1by8ulkicj+VC3emX0lZwH4g0O
Tt9RVQ3tvg30exuLxvcUnw7i7ywmigkLSdbKFjX8kaLeYolEpZXAcwjlv0OYcvkxzOD5zlxlPJ8L
240hH1KMe3Ezt8kHcEKTmkHuMBy7pULUneTgpDWwFP0n080rLzyvAgAZPN/XB65MmrbpkIVDuD1Z
kq0s2XO7KALztX/cpAk9DxBCzXRgONJLqFCaYd4BSTxpu+mbQacphbNa0puEtwdvDvFLzaS9MOpv
m2YOugHN4EdHEj68rD1jENClJ3fwrlRN+vrjaCDk8ot7JM+cGCbtkk+TT1xA4b0qwiZGp8D6hz6i
97NtXxp5EeFjhARn1aAwAfueoYg1bKRHLMoLhggJSB4f9mHTohErB/5j4ltKL4BYrQlYPkN4TqY5
26a1PqmVee+GGQY7uz5/dIqoTyserd+7jP+RnguBdeYKVrs/jDxsDeNGed3at+IOC4m0rpIdJ6dU
iCIjJ7MKgMspC8bU9dtHu9JzGGKBh/EVL/xmEdEx1+u+p8R8fEFuhQXMZgaRSOxUHmqMEmvmFI8v
QX6FXhEgYryYe4OFsHtgTGx4m52K71mfgMMeE4eU73sOY42TEdWDRpcYiF12sDonViwk05VL+daZ
CSVlwBdCYDbYtYqM67HdePQxxknJPQf13BcF5ZN4NqEunYEMsLT7zp8jX5WcU6ne/n0nqTN+2sQl
pHJptSjp2Lnh6dpGUK6fqj7+dTSy56kG9gaqTHqQTE1MMX5krrFdtgK5ieP89vo2VVYbKyRm3eDX
KSUj7wbZ2pEkPsV/NuLX3+Ozf2Rxcx8MF0G9yFLPYP1idsbnSekonggMYCObUtoNonXXypZBJU8r
sE5uaXSdgczNzSjWjex0GfdA4lkelsQGdhCU9LKhIytBfWmHKICq6gOPXcu4C/ARbkhq0sk7KMNp
D8UhIk682sbWDCN3woNjwhSRtHqZERpiwd4QfykSCr8MRiBKkBUsgPsh4/Owh6z64Bt9GhWM0yUc
5iSQnFTNhylcVAkGnTaF86XETRSmCwIUYp9ni9D1aXxo7ovkmWiLWY0Phdb2eIZMRIZ9AxtQ/245
LI14RRsxbPhUpAAsQvz7nP3NfsvrOyTK4/7ZKSevxLnCokPKIkdCUDJkbxtv5Jhc1wWCQTJAobdm
6Qs+p0uBj9QEKt4Zp8P1OtS169d2IfYbe4pDpmHyYSLEnouad3A+fN0XVOY8A4fIFJbysDVUERZe
6apdPKT7zpMKUpLyjCHNDZ3uCT0hS3tAh70zisM/yl5Xa/L5Kc/DrVoU1z+FSmoCF833ofLB45Bu
t1De9Q3BwWAK6SzSDMpagBFALUISzU22uQ7kCMjgxCgH1zm6JRLAldp58fCApPhD/Aqtb+xCiX08
kB11rO4bhsanYahzeylq2uTlrTOiCvuLaI6Ae9KH1Cl/kLsSfsPUzc3rs7QE/MLhUYEoywwEWD42
NhpJ0qxD65Ho6XtY9vXrS0EiFjqITxtH68gTG+YY53WACKFGx1tQzrC4zNP3suBK8NQUut6D7L+o
9ZZuWoGg9gGndKOp9dRYxtDo7lhHHZeWORIhq3J/PCqIoRqpBcgdz5P7bBuF/SeaxYEwRyHM8XHU
qST/T1Lz1PImnhd7/kDm9LJvnAviHF500g9hRa7gdf//LsWLl2fcU8uXjONgJoW/DM19T3ePH7VT
xRZtxQGofvsgoAIg4MKqrZnsfLK8235huetW5r/CaG0WATMxABqvLYPeYFPTqEsqMjL4maQ2v+9n
Z+73PHhOl8a6U5JAzEW8OtG8ImhZQ23jS0yBlKMOo2BMVtPgq4Z3hDO8/1ewTCuAv1W4O3/Qctzb
TT+d7E3EilomheaBYTfrWpVvYLMdq0Pn/t7B+Bw3aitl6mjLoPsUHqpIOwI8zcfqffS8mvleCzev
VNKE63SJ5lIU7Nz0GlZI98LjPnuZTUTs+6IAA7QM1Pxm1JJf2ccrVJ7voonmJbwbv7vgBqAIkbRo
r9LC1nocvOdWcJwPhfGzceB3qaHuWvun51QBthiBhdKddrfSy4eq2uVEir2p6/CHW5UOIVTEXLrn
Hm6GqrMUi60c5NKyEzGZToUJTX+h4cQdy6K5h6J5rcxODR9iwcW5E39sMF5gp9tEPc8/TLhLeXOQ
BpoqhIwvL+HX5SL2D1uFtfNHIG8ey1qmaflRTCGGM19AuLkIyqmKmuMCB9oY49CglfGZ7crbvZU2
RxmA7cWRzUwe9HfZh1kVYcBn2/eLT0yuwPhQBmRumaQniNRkZVx77l0QOQgbDgqW2bZD3xqY+RFR
GtEz12caUmAIX/zpSl8sP1luCX7718OcE+HWC73jF+7PeDnmBfSJ6jjU58T9cgK8TLrnfTFJ70+O
cvSGQaFM0cVRkOnSRHcIiapRAceRC6Fghx5YGvjPbREtZFbjhM6jYuINo6Vr4JP1zHCz2f37gGFf
0LXDHo13DYUIriwLKBQcYn0CdZloqjJcx8icepabeI0AnnQGfwpPz7ccA5JymiwQ6ncpiSLoYBB6
o2RUmwc7wQWQcMYgB4psYHclozzvXM3r+U0QyTKM9ubG8opO+i2ZqNEfXW5mNN7qLMiFu/CI/Shw
GwZ+pNDDiDSNBiA5QCDdi2oALz3hV2kUV8qYL6bdCMtFv3ouKjJsH2JMZY+UvhbX+57ZRABycVpH
QJ7S+J3WcZIz6nVPD1yasVqylVnr9HpLrPVny96DvtFLqpOen8DYsL4Y16DYfvjauwOl1Sdx1co7
+lS1Q5Xx8nsENAiGQ97k+bRvfp7lO9hqNo87jhJK6RlWkIuOWukw0Co1c1vTo1lHWw5rEaPuwSFV
sQuS5QfQi29yHCJDYRZ3xIteFYCtCm7NVW34T4DR1MRY51TlT5SRKfm7tAo06X+N83NJrvcr3R+h
P8rkDYFW+jxieZymmDkmZQTKjp39Gs5bt4j9TQ67XJpjfdOGMTzRSDubWrzOTZvGR3g8GFdJNozG
oGsT8Coki1faCZkg8FuwLZBHSHILqgz5+XArPBWTiz3g1qyv1x1CN5B7BCtcRR35BfJ7d0WvhNjN
loy8/lXoYu7sj/jjjiunf/8W7zkeytnRg2BcAdNt46knbCftL8Dk5bYEUtdJJx9xbtHaCRIGvdfs
/Yk93B5H3XdgKfeC6AX2nw+xqBc8zY/bZ8OFOBJZRnMfvId0pkH1X2rivp61z8NCU1cgFbWZbgEW
1bUefsK1vejVWpoA3jlaUOfnMsJuG77ilAZifcbWeQYozwihZYN77t9ZHR9vsQpsu//RCujMr08G
VjOLxoi9TwDPM4cK1HKklJ4CExl/bWbuK8rNeHrnTAhFTYOzBGt58QJUhH6qXVmQafYxxECXj5k1
e+3FMjHrhnX6bt6ajZKbYkKkA6iWkO5wLis+GEnOaqFZ9zYCWpbXc/05jFTcxWsHPqkOZyAMBfQy
7PvxcW/4XUeXGOBruVZMRMpnVUj91HCG87aqBeAmHn4UtaxyiNgutMvkkBRtfB4019f9YuMM10ax
tbLJKO523js3TK6xa1I+s7BbZ7Mi2lg24xXAIYFM8znT7Dn6mlr4JfbbFThxUHKSHFxyicQMXay2
bMU7XB/Lllmbparv94uRgZs/j5VuFdwgxJ1SDTZVs8D9t9GNn6882UYtlHxl75/tpup9N9qLr64s
ul5s83e8HKcrLT80RlFWefbERTbeccIVXhLKpUgSFf+MHsvbigrlX87RjcpCiiMZt90QsfEsxjFz
rdM367riIIMCWzlGKBxFNk1ZNVqpzEs7cKlJkHDRPInZHYB8Ozqa8xLUoM0FUEoXqYVa0qJMMHPG
s1as3dRR8rWk2pT6EwlD5+mt8//prmttLoZTpDTulotfUMHod4xowMmL1N6nQRwD8tMzhv30ao43
sR+e5ORl3LGljiGXgsAmRuzwcQbw0LwRHBEz4JU5g314tGMgqwWBmhhibdeoEa8kVe7ddDRlR3dB
nG5QOgxc82m2OnGtNhWjxiVVbTlbabcziK0o77sRw6mRJVzT+INw2/KGzEwlz4IHrqz+0og6SWhy
GGQ8UZjiI5keZjW8+u0FsGAd1eomH1DkaGX6c3pUFw5dTo52FRli3VnSSKpyJoS2ogITZVfbP1t9
91qY6/PtAGgQt6cT5yVH61AIxy2hrm0a23piR5Ob4MJ9tJ/nNWJQEKr6mXnquXouf1wTWQk2nNOk
mDlrygo1iOVUL1gdk6wnz91cTWME6SBn+6Sdo3Pz6D/cLOaXIyQPBHkRTSAXtFc0BfoWQ9kHIu+r
Bc9PPksMsB/Mp+jVSMgEvW1wcVYvksjEPbo3HxRUmCbtgwtrEnIoDgspoGLm9Eyd4TeYhGxD+u3Z
d0AD/H4iqvZS3woOTnThbsE+d/mE2mS0rrwrIbm8z56CKyWgBpYF0XbgdMBPtNstbP9PYRjV1Blh
7Q2VYJkrx9Jy58xxk2z7vwiMsbzE+HvAoqBZxipGuYziPOWvEBjoK9CRWAZuFnQ4PDHfatVe8Sue
2YQSIOZ8QHN/ZA5kL/afHDmJSDFO8jQzzk+3Bdt0pAf5j883Gu7I5NzSWCpbTgxu11wZX4fIjKT8
o3hjWqmPQnBmeEjVYztlZMUN+1Bx5+Tw9m6oOijHsBWbnil3gJTmayXL2TpceubRJeHS2fcOHrcA
x9pml++QCjdWdfdail6pT8BEhk+exuMPb0bRj/Dnq85Xe+/sa9eBVhyAIJRhZsQYA/yhFUGzbDQu
ilk6cG5SxBvJX2YIXg+IY2ukQeGP7xLaD0RHuqCoQ8D6r4S4boMUbbY7BpMIKUTUAXZtJBbRwuhI
SSwctoPZEdm9PgBQnV/2ygqXZ7lIF8WqJQyjnLFzll03vBQaFLNvCDYRcPzBJ5lNiyKZ6ZcYBRer
afRqiCy3FZdHwpcdpts1FQGiVSAvxnfCTkgElKWXnVdcC3/aFQzcmYFk37odssMIUV617RvgS7BA
GBxexTpnMiY37rq9//g6Yr4B+og9YPLGLajQMM/QVWJj5P8/JDDMfoPJqYbZQqMdQm/zoyPAJ6P8
L+7JcAWuzj8SuzH4bPuHjjnS96iv7HIjcjVa7uA2M7Jn/lDpEKm/Dw09KH++wUozJrpFRRqPnm9E
7aAgFocyANKCMl7GL4Y5CjYH4KbtVjTt4Fgj7ykJxCnWi2zjfSKvJ2+uTLUS0zQP6HkNpPM8ykat
e5p5h0KbuSBZulkDsqSism3YaCo9F3KY42dKKT1fe+5zGHuywEwPnFuCpkYAf/dUQLLHOI3bYOpe
/WNqD7MhsY8dmR8tLlYSAqDGUZcYus3y8GGFX68FPEp6SEXt31yyl9Eq6/iKoBoDh6XtXz1216ds
nWO+g3X+wVA9nUtf5Lwbk/pvpo4i9eAJPAgwxu0DXcVz31tAEKgVdlvHX6a113jfUkQEcErktH9W
Qv0KxPU/7dhg9cQsPBCq+Um3A4vJzbHj+ztdg4olGDaz6E4aD+yCn6WTGiuhhYMwiv2XFtuEkSN+
XmnuFyHUAuKt9BMrW5rF9BlszaqzmB6CllRVR/pZNc4mI+vXuplobL2VuSlI2xFI/Yj7/s8HOnZr
w31OEBXfL/nRlY1FoGhuHZDhyQd8AB3IdlaBJdsNFK4DxexK66WgJbhXX2tnfXlSG6n6naVSfZfw
mSohdoscIq93NEAyS+RprK+i7e3FxkzDdZ/7/H58xi/832Nn5knvto9jh5GR2f7512epo5nGaGfO
FnnR5f1M1Bd/IuYZsG0G3v4BxJR7Pt0ijBuohw2f8/7S6MbIS2dJVWyG3bDNMCD2PjjYFfmrG7Cg
FIKOhaf/YSTwVwTgcJkueWPVIhS6y4rp1nVVf7V9rI036sDubSAaJq0I0cVxrLB8YwY5Qbngj5wn
Lk6NqdGgYMsxl2lncQCoEswO2X4W8eGZw4XDFmpjibYT6m9DDPoWTroayZDGWBajTHCjIM0DLp3R
EL353hZrpzEtBbEQkZBbCEMrQFm/pAGwgYYYU7arEqqcBx1P6ymdaB6+BOmly/Sa6ouGv4VL7hvs
tqdnhhUEK4OTISNM0/Qmwz5UVCA+u34TrwQAziyWYWnio8ZqJcEXg+nz8dt7kaB1T3V88Zc46tLM
GRgO1x12uC9Ra0H49gaW5h/gaSC2X0K3WIjy8DEXbda6SjcMWVmpohswza7QDYcSBWaJZg/eJASx
2uE64Cozx8pKg2R6iSxA+SkBEGAB7iSuif5eBmUBta5USR3uY1hqTcgscAD5xE/Kn12rYgKTV0ar
EG3elmNXkQCamG8rb/ZHpYrSBxE3ueDsyD98Hhdt/vzS+nKfj99kMnTo+vWMKxaLF81hUwYpJMEh
OM63U7muIcmZc3qS0QlvKu+uIVwNVbHGQDW14RtpQqlCPpuPLZUOLieOW0sA4pI8GRs+8iHFt0F/
Tjc+Fk0Rwes5WjmDg1WJNKUKOK0raQQDoeF5lr/BtGPoJQR36qVfP1ESQBBSVsjbQHLrv907B4VC
h9cmyzLhfw8utTbIOiOxS8KAYemBy6S+0PBDbeBhoNTxMEuVCn96s01juwfnmsJYU28kYj4ThohM
kszBvW1L2RX6BFwYwMqtar88KBcplAR9l9uGNvdMHIcTP9dhnZrkleYkhBsyVBGHsyQZ3JyAg+6l
aXTH4yBO62TWz4DKe1wmu2Xe+Q/FBYpw8fNipuPe5Vd9CJTnl4vmy/W8FSJt2bic9ii0IgMS20Xk
aj3DpwhiGB8yqUTZrP5V6clVvv3SpdHagUTIS4ay3HnU1Nnx7OV0ogHaEuW61UZhUkUd0EbQXJwh
qiCNg1820E6curftjce6dOAuLCkoag5ddthxezGuDNQD0CyKhggOiOMAkmGajIngQz02djG8/9lb
8H7U4Q29iCxUkfl0AS/cut2VSFyaZeEry5Nby7qznMxUt57WttFYYkilG9ChUVeUxdyeFbBhkaJu
fzF8KLv/AGRqmOmgBhEIm8v5g4GM0QLfQ06GcZ2B2NznKJtaTnYpYj1IYCAsZrxZG/bjhT+Llky4
DzabLTXnIMRBVd18yi22tAuLbH7z3MSLrGPAjGa75aRurOjKXTZuxWah3xjQ3emoStMgdDTdjte0
lrSpPDbs6ezTnLvj4xqktAxLS7j5fe0nUQHcuGeWqUAdv7mAj/OLADNQEnVN9jkWOrjWliWH7oMe
x4A7xIFTSK/mCHtQB1AK12snKo2l5Ahu7UnpR0H+EZ9jpMyUa05YLaKJ+1wBXIGcZ0PzxLBTPMRC
PpWl5qrPsguhtHwdp91u+9Yl5V4o+rFepYvyd/YrhFAPipt8/zliH2BiMDraPQ9uuqtA9RDDFgKm
n0bdj9xsXyS+cmTPAGNVrxy8GTMkUFKHFUVoNq/QEtzg4RwocefNiZRFxk48FypIXRdoK3SDMBRm
kUsJ0WWygwglQTLaNF4IKaqnlG++6zonj2TRRiS/uJnQQA4XT5IbyBAetr3SmPyZbEpAEAWtH+Tw
fIAde6t7y3CE5qhI/NVFjub94T8jLTRFQLS758WBLI95hbL094xRh7UaJyzV4I7qTGg4wnJnHaUF
wyYym1OkGJfcsK6ndZq39QC1/Psvo1sOykiShGhgwMBMKejvlCt/90LpmFqLyH0YDxMW6BvWPUs8
GookQFgMBHAj289Kwt9RaUe4eWEqeMgDVY2DGo8+ktGt0OPlfvQRuPZlsGavTwMDPEkI0gFydUgD
E4ZUvif95Ba/MyhQKEquoX8PV83DTttShk/dx5TvpYFHf2yWsu3XU0kC/nM94QbPZQO9dd0FPp8m
zMhK4PfZ4LkiYKPkPtHbPcPVJLlo2prWgAQb0jyZ/r6sMgF5L/7unLJA4E9ZiNHaI3ZPyWZKLzRL
3TOxb4nOYIz6wV3OajSFIJ5c7rhLvUfE2KG2elRXHioG3fpqb7EfVEhpV0cz2Fb1UQRCE22twgGJ
qnfGtZxrCnIB4a43gxP9cAGn6UqtC1pPrY2Ra0751E8rZrMLawLnCuulh0LrnB5bSoueD+bwtlDv
SxZzQHL/+SHEIoetYMOYZIvtOAvtWRGX0YeJ91HgWWYeNzGOF/MvKJvngq9EbR1LqXRiTZ4FKHzv
jLA3zC1CahMjJ1c2frGk+OpuaOweuGh+Zg+I52h/lmGQj4FNXvjFIMmOnYp9+ReXJKViyCh3AhyC
NKwAz9jUnT+1LdpUlDrL5H3dhKq/B9aLRVAr61K1PBtcJsynmiEC20nnPLgzUB9QFL385xYqhRi5
URq7OirmFDytjmG5zF8vN5Tdi+GprXm7bk4Px3UqUMf4MHesiuqZTHZXHiXigSwxnMvjDyddV+8q
IKTKCHTLAt+Q6T5R1kMuInECoouicsYQfhs8WK7N+TEtzuzaIOvFsmXNp1ZZCccGCMrjJNzFFrvt
YWBNxgbYQGiM/RJ8yeYqfFwVu84LeI7n5XWptDs2bc6cYpzk5PtNoMIA4D7dJ0lh+1bwY+NdYXtG
iVKXu2uH3fE//Kg8LZaVkZkZj4+gfR3LsQZYhqU0giR6h7igLDRnfCcQ5d55qOqc9k14Ljhw6tYS
WxbqQVdg1bCsoSv+C3cI0U5tJHy9IY0EnfWgEP4/jq5kZJNFoijnq9Yf3apu3ceQM/nog3csOLDG
WdAongURV/hd9JRsg0z1XRnaG7NcslE6Q23fX/MAdRvuxwzM1/yOeipbHjzmqFLRACm8E4McdkW+
ikh+CPvctQGTEIJdQtxmKC/EcCicEr3lRljfB23tQxS5zmGMNzYdwQ/say+iembwrGEiAJV2Nzug
T9e9rDnw6kcAorgqyRrKKfd5QXyyIX+dfk7t3zFB0ciSNk697Rd728w/K4/Qsf/p3PEHs/gOzuci
ZeCdKfzXZXi5EcSvIpeMYU7TLvzKW1ntG1jw5qru3vEBIWKv1Bz9U/bMU9z7MdG1FRXQiqnO6U74
qa29EELay5ty/UFjW1AFxnoW8naih2k299lmEUgCc9puEjrYeprnGBsrqhD7dRGCEZg/y207cHBV
xJP1E074Yx3sdfM+m3JU0fQJ/ZiMp0zZiRBKwEGX3mdv4xAnSsaPAyK/kIQTnPsGdL/M65E4jTlo
EOqFsELk4svZOukB49FxfkqSCLV8SDxOpsLBqgL+oZnUzkHW4K9FN7UjQ2SXNNEe1QMTm5E8qhko
ZzXC2TtitHadXXtW6wWoDXbZGKh3UvTUInws+E03pEKAG3iiwfiRl2ZRMaG/C5d+VjFkcw8/Uw7A
QAvg1JziqzU/XcRAwKL50K5lqVcKmAbGQkAom019GvfrTMgxe+nEdLJ5I/LTHzXEfx1Op/zylXm3
tj354g/iq/IQwVJiaX/0RYdceLcu0DY7TOkXX6csmj7uBvZcGUiElh9beBp/UGctlMkV/e4cjhMh
ImmqZF2pqPRnrCpT1O46JmNZqXbzN8RT5MTVHOECTs0qeF8F3XaIaTOxGi8E8zGMTZnlZYt1+I5r
bKRI01lZTCkfBj+uppbPX+sT0KbK33ah9NzOp5KGf30fe3/krSf/X3FAh4cXTHiJ0KE8GhZMjTqx
5OgiN4Oyg60n3Vb3fbdHsb1ccaOFsTjibeJ35hPnEEM0ShWhiK+w10XMDdnI/QSja1zUSkZL1Bxy
L8kQ16r9W5mSTXk2nt5hQgKNkiT1dQWwPd7OVX/5Y/AiWAuMuv18IEeANIyMSDDJ5rDPQoEGTA1+
yR6+X83EVlGSH9YOvhq/38YzfLoUgoDHnC+ACi3q4g1Pbv9W8PTrZYEmW9yxyVrc3IbgnmMkWyMQ
w+HZ8I63cGPAvTMhjHPBJgg68fmUdx/FSn3GRH26aL5ggwF9g/fc3lXY/oE7b8EznGXMQmBLqe57
Ua9tknoyjy6YeItjVjoC+8Nvc35R49XHQiJJSev1cnAzkVf2O0fUEiuR+zKVjP7iKVxe2gQwY91s
1HJ42kA6eppCUg5EE0E46r24zxDjF6gp2Frrcjz37EleHYPHU0zltza+JcF8WAxReWSyKQuwm5Jc
VivF8ZyzFsvTQNfYU6xD1f7XMMr8fwRxaMBwXBDUqup72E79jTlVORKcI/u3x7f4Li/WV61VwmSu
HSBVusAM3oqG9tvpWDIZTh6jSVGEnC2fCVUz6Q/+uLxRV6ch8N9uoaEQzlJNI5BZCeKM8LjL0h9m
/GI2MqSM/QTMrLoF8LptjpKzcJWQU5DGZIo0YFmgY4OKe8UZIcMJP4ZujnxVZouDqqAOCuNg6oCv
IgfMf0YNPZOiKTVNKd7HHB2GVp+JCJ3FR0++c+lkhgwhif4QL8/eEIzhe35OCc8JzvxMwtFE+WSu
a+JsyAJs7dhfRiqo/A6KIm7+m+k4ZErUfvtbzPP+MlUC65OofXFfxUnbK8bLZNqya7h2jeF86O87
IBoo/80DGU0Cp+mbANTcfOnyVYw965Xek1uV6pz/rwrAvqeeqKa/vGb4/M4wvVsuU1ZSW+3yxuNK
lI5E0YemTT7OvgOiXuvoCXLdQDR0HaMkw8yrbXNgyt6Cv26hpMifqaRetQD75ZK1DmJVWQ6kyx8y
rhAA4XA4T1o8j6P6sssgjOVPilDF5xHJQt3sZC4oZnrAT2xWgqUWPklYtNwbDHS3lb2W+L2eKzoR
aB/b0UjBIKi2H7pIspZk/TV7Am761NHhENXmjxQ/DzHB+zums+bjorddJxLoyckzgmVRANzttBrZ
bHExJM7YAz5516GtixnOuRKUIFmIu311cf9jzvLsbxtoZv1n+ZD+QBgxCYgxYfkz81OHRUPF1px0
blhjcxnEzlK95knbRF6Xz25Mh9NvwF9+OENh1ey+GGVHVw+zqxVSSQ6RZWy090/tS2u9vGe9XxKo
mwNNLgmP8w4ViDOa/1gmwzJrIF4fqM90AXL4qUEqrMGXV3szPJStn+RgkD/Dm6PT0l0NABd3fjqb
P3mFEz0c+U8borQMezRYndnx2B2GW7R0/x8oj9E2K420KFS29uALWGcbPMCtfYGQGCkyqSACPHL+
pbToow9tvLjBrRbjAel0VJL+7zI7SXmOmx5Cx1Hp+kCv/Euc3P+4Rwd1jOIwMHczz8EX/7pPI6mN
EYxa8rTUEds0IKeTKP3fbsp60n0OZ/UNKvAEJ/3sJmzS0uV1Od3Q6EYynh63xyX5i3TUIIx4DMxz
jWHrVKgkYX7c/AZxsq0xIQCxz1LZElPx83fxc0BbMbDUDJC2bqlqlQSV6OH/3iU85RUTyzuxCKGI
V1WpsXqlDMmBkhwRypYzf9Q9q2xCyFnfXCHm1tXUgkGWCYIZhBj9xi4C6Ckpq48c1Y5siBtcun+p
r2JGAhCHjfRvswBQaupj6ekbZSBqldD5uQ1S+EXjX+RWjoh+24d+xVKbvs6gd+zUwrRwa4KNTO0N
+dA3rTy32+pbUY978sqemeY6SSyEXGxztVh96oiKoYCwNSVl5j1LnyUzf6Z3Kf0EJQowzA2ZGD3g
GNLiNvRHgyFMWwBFfWh5TSX5tup/B10DG/wS6wFlxRapLjrIG7PnnjgiMEjDaaV51yoXljNV6Chr
rioan9mDFK8xRAat28EslQ+Ed7VMZGaLrDdiEBIJ8ffPsEXCUjotif7QeC5wQqTyLgVMeZn643Oh
aI+TIKTlONxi56+pa2BEbJ4hhseEJpupM4gAWXj7QPt6wLa1B8UGefCyVED1wIImHkqRmY7rM4AC
RdNSqL9701rELQexHpBv3oRQp/M0gAc7IO0WJP51kqlQ6/yg+35y1sDNGBGzbxCqPEqIKWMYgg/B
oK5q0EX6vawWG8fgN6mUOEsLiTgsS4WuSMhS7Fzi/tLLj86JlZkLFGz4apnthg7GYtDTezMLCerX
SoB36PoSdhqaFZHLjhnE8tSmvz8RMqN114F1+bKSYS8MUNGdiCbZYBwQ4lPhNd42C5orA9ryh0TG
37EXeAS0vAmt++dHFjsWD0ajCaTjUcw518oGCrqSzPGTwZQwuY2psWwB+goYw3xyF8GZ8mFpfkW7
jlto0UIyAbeHXc1LNxduWwn7FdjR4g0Pj2RA7H940Sq7+OWAICCn5bEiwthX/H1a6dKiYouUsPvf
FieJ//kw+Zn4h5hjmRHSm+mz9N5G8nTH/PbZK2bbKgNExE+2iuq5SQtM0emRLGJlc8X+9xlIH0Ra
XKdS3Pzr+Vkia2pp32F+2tVZWbcpihR5EM0F7A4te8eWqRthO8h7ms0Y+juFTU57e0Ex4E6B8S6W
kLYGRKQQdfxGBsLX4m1KONtre5lCYpkBimnfakiLp0HLoLs2RN4SjsGpblgYjbS5M/aooVDhs64m
uWmJNIWUiVUV3Vtvd3qc+BmX6cXNeCqmfFWdAFM0MnzGXVAbdZ2PTNr2RT7aI8KNJMci7Pd5wNv0
MWxK5ZZwF78TGmR0j+7fnwU5SzX/Zx8YHD7vuTFnI1aL0ydtcd976jp9zY1wKU/KM3ZB8E6nttST
s5C4hEFqQCPXlAYQecl2AD2VjbasdrcWFWH8p5rCdLy13J9fxj9soIctxpR5ynxcm503Z4Tpr4mn
PeCDVwzkgN5h2U9uyzX7ONTbHFg39XLJqsxcdoU//TuJW+MqgRBhtWsxmXwJCQY5aXVVEyodSYPF
6HOapeMbgOGUKYG45N4SBPy2CzGvmlZ9G1EoySP/OZYVvIDXlNQeEbvhR+lFGXXYELRw+SOtjflm
P11p0ux6V8WVo5rgfMter0XRmjl9BYV6Z1JSd6MrAWntGK0Q22Ei0uTmKxCi6qenYJcgBfX/Bv3Y
2eknjm70qziuz20RLp/8rbY8Omu65Ms0pPgySM48+cH/tkXxcrbEcjU4nfJ/bjBqciNElvV0u8x0
M6GE0Kh8gJovFrTYLqoeLABEzBdir+rmPnjbaCl+kiz3t2eST3xk2TpSFcWO31nTDkOwMDqrB4Jt
IXXYN3YhprceLqD/2hC7PMSWJ2bKBWGZj2wOnUBUs4DEfchFShts8cDItnH/tcUyWapjglX1h9Yp
u2TPLROu7ExveXNLME/ay2DlQWk1iS2tC9aY/57urC2jx+t4SlUBW/emu2iDEdAkrCi+AYBqQPjW
lw1/dDJg1ndcMCOkFKVIGMPDroFH31ol0j2BocBacLdkNlU9JFIRwjENBwtm0EL7mKMczThKkkSD
W3lkDSDUvRiOoiSeyxeqoeaUK3Yz/XRbKQirMaSHyvLGEnjNvFuXnQ9z8Wd0ffu6WrGgZHw0Hpfh
YCpcgkWXhq0I19Df8QBzx7iKq/BFzP0uLwdLkV4OWKS/UL6KlHUPCLl4bRiTlo0ykk/4oXesmZtG
2fG0cYZDmc2WfiM++FHSyJYRcSUTXJ9XTibKiV7S5v69fFB7BnSyfQnS728PXjQosZBy4UcFW8/W
s+BlxS+bkEJ9wuP4bXZ0Ck4maURmezBWGPSaAf+E6VwUPZ5rkiB72fVqCDE9ZftrA9bXqAOcdBp9
iWc0HDQoS/CRlWrQu/0qt50OX2u7fS5/8HsgAjE5Te8j+BNsRIR5p5H8wgdlwe3FucUKt+de52TC
D857JVYcJeWPlPcSX3tznfMEGYj4XTvg7Xj/njUAirDbiK+Df38xYDBIKxPCQMLRCF7IoFZk/0IR
a6kkveDCwSTeBAXi5/rCO7hryJuhGMZa+OQtSNgLVaZakcutdADH2x7KaRG1eogPy8o3BTmCBtwJ
ukx01zGyGZJ+OUYh7hgsm1nBDa91bBdp6nmk/Vi/2wukOfhApu0j9nDO+rZCn06TU213LD+2AcVe
WMKGNYv6t3qXr6JNqhdhsIHQad9Uo623UhsV8mserc0fU6spaY6gkaButCQ1K6YQm/ij4jP+Moc4
R6IprukEaEcJsc84OdNrKLQgsf70YRGmHn11XeXqJcgNU/xH1Vk20RLkYiQKEUL0xbFuhCc5Zv0q
yAoB0V6YZMmOoiLwbsA00HksbO8Ch21kFYCh2KW4VxgPpge1Y/XBUQF7+hrFOeWsRCdHrPgbcY0M
FYsFOHZVd30ioon+BYe60aNJqw7u/p4bAy0pxTrd0pxzhLrnWXaC25NOTwxFumBDALZDqvsGgyga
EK/WvTXf2PBTHe1Q+1M9ga0+JkrzXrYykWSLTA5fBvoFqAOUha7Pva9Dmkpp4wKoWfGRJE72ndS4
zpsyKzs2/cfl/7niwqN2lQHnYzWWdcK5DNJxSulGrXi+WoSJ8nCma+xe03oiiKWRxhbjg5ALX7N/
jPA4lIUPW+eO51S1Wkzqq0gR1G0uJMeGWuzG3ip4IFPbpuC9WId2NfjW0F/kenATLdjZkFifzicR
oO0+WXT9CoPK2YUZRuozv0EB6K4e03+nrIXj9IaL/lxCcNocyS0Ckox9o5SVCn5d/eiMANw2FgnS
sms2dzu8k1+b7rHddWr8dhrUXwyqm5+c5go1yxp35nQ9U+KV738fWg74x/TGdo84Hp4ljv4FirmR
O8QVb0jSZ/1i0QU0cbFKAuPxy3ARK1MSa6ZsJ5PW8qm3oHM+fNIOzR6m4HGoThrO7P1zI5cgwxbn
D7EhUwchW3qkJ3xzFeLylb3oGfJFRcuklD8eY5Iyze/jCmoIOcyd1c1OLKLM20Ill24YfrR2FZCI
uLTilv6HRqvtESMRe/WsZiy+hyWa7WMj+SfA6vzOmSy1WuDbRprWwW4IGRDIVj9PG7p7s2CaUpjj
U4ZTsLXyh+b2I6IrABHsqHg+DCvm8290Qg/oCSwiz//o7audk+hU5EhB95Dqci1ZdxMDA3XAn5q5
zBuLle4BG4lnHyQJJQYEVMwoEdW+8mmsPUQQgfNbkBJofNfbrgfr2GUI4tIjF+ZRELMedmPrd3Bc
+RGbNZmIFBLrdAM87RSmBYFB0kYI6XVMF2eHPQE6/zVn+G0oLhB1Er9woGO6EdNuHRrEMv+Kr04R
0/ZLjOZvZ2QGU9FVlOCQP962dn3bioEbk095JkQQRK0JRkyDLs8s0CEqbQ/NqhA6HxWDt2RCM/xb
JJUknHgSFtXlh1MMk7+FphDSx3Rn+g5LxDD/KCd8lgLhn2eyo9U1ki/R90GKa8gGgZBSCtRuPWUT
Pcs4B5KGeh85txyvIitdopr9NkNqjX/qYxG1ZuEZZTJB/VTg7nL79NwdSQcOBcEx36k4uaCEjhlZ
b6nIvHYT1UDkaE5WLa1c2gMOSAtHPeFjGG7Do0AnZ4CgLkmdbeBpHJlgA7D7PC1MsjPbLrt712OG
QZfzxtHg8+Os/+aVXuaWc+URsg77/GNDXvonMaxwRl4yJvegsekTMj2kBbpFALib7e7j8N7qINcF
EGELeW5IOtSJ1pHcD29IbczmddT3BwHSjlXBgiLGyLzr9RInABxtF/zE/HxPEYmjaT/QH+BdH6Pp
uq+hcXnv22ud94S9MlKaA+bCYAaOa+3skTbbb6rphfjgh5+QL03YsPx4WX46ar25I28vNdK86/MW
Wuw1Ec4qvV8jQs84qA6Dbg4aRj/MRPEiOF50pS3Sm4DPI/QdcQKkIpN6n9YUIQ1YqbCyem6wRlQ9
xZA8l0xYNPN8/EdAYjQBO/wNVpTBtI7JS3uPlz8Q3pQ11LneXYEPsEjlHrcRYBa2J98ZZe1XbigZ
9qIslJRDa6u54cYdKyn6uVDIYQF/P1idyH7RLMY54mFImJ0v57blI5++ONLQx3s5fmlc2z2sycsu
uFuBUw3YvfYHJMSWUDnQGdP7EpyHxoZOK8mXZNLfIWfja0Y+h3SjMkwWXdt8DQT9Ej2ZdRmlr4LZ
0BraMi989FPudSNkKZwLQhSDHfsd2BfY8+gE0aAaHT8TarppJ24PvQKjL36QrugyrckzOv/i8skX
IHW+7zAh5mc93Ll/Lxw8qguvLoFn8rZIhRvUMebnXzNl27LVJEuVXEXb1AVudMJApoEmlw0NgVyr
fvSj1djOYyc8A8k0eLXPmO4zH5g2VfAbt9N6zrrqLlseIovwlhGjT54iWYupz+3skalro30aor5S
m1ACnE/HG+qZKXp01cQtkvwqvzMaDoRlSxiBrc0ug7wmxNhK4y9ibMNTVNRah17rJyhXtz3rZo+0
kypVws3ahI3h0OTydVkS6xP1fBjIlWcDjJbUQkDU9fjtlvY8n6+wRL6s5XRrU8vKF2AIavmmJpUb
UbkTS9UeIj6ZVvvg83xWXW00KJhC24WMwPsMjZ82HuyDRhBpY2RHDeIwPmBr95Vpm5oL8SDQNslF
d8ujV/Kc4p8uAsfeLAps/rfUwwWpGF2G6A2xBbKi7IpjtYi6b1SJi/+pTvfntkWRLkTbR6CO5eAu
mzEnETw4itDgcmb2aBpcZSyLBRwJNZYh2F0t6RPBusdPA9OuR/5UOnCgMQ+Pg1EFVFFuTz859t/M
nLRPGKiThrHhkeMXMcJKFUZJOTnWDPeIUaCfGc3e3brzYp+GHUV0iY0PcrcT6mBgZfZLxgaaT9Uv
pkDeKbM7VtWUPKPxmh0a7Zo0lQ8VnWLwp7OIwlpY9jtOg9Lv/m0EPWJVLGyIsy0FtHHWJwqBW9pQ
1v6zFVeXQkFlEioO/eEycM7FJ3eTqrrVB6OkQh5H1t7VEiQ2UbeiXVokbVqUzF+IFYyx28+nkCuR
X+2ptfn6kg9tEcj2HiDjDFbV8v3D0hmTgTUdLTMDQY+CyHn5BWGlEbDcwiEAaDTA7N1FLB9T9IGj
OhMl+Y7FwZxxhVIMauad8ie1X9d6+tj+Dr1qg6gWEjGopjXes0S6BUJqLoSiniAaBWqHxLMbALGn
UjYDB3QUFV9otVdj3rO1CS2896snStpMMWr1MPQE4zdrAQP6o7ZaQ6710ubwGXCa3L3EtDOD+fix
JWSimvOOx3gmvFyqmpJksqSqqG+lm/Q/wYKI8OTVmQ8Yin+TeejTBPNxjYlWWNXH/3DYO3Al4an+
95B8a9LQvvsiOhRDm38QjBUNRGl65bFXjd1DOUVqchxw2ly0ysXPVzj0zeCMgQLv84XMI3AlSp52
47NWtjXbV2kc0T7s06xXiFGoQWB7vgdo1B45Uu3WBOQxXQ87ffUUdiHSXwiATju39R3XaehukJSk
biP0DoTIHs9L0t775D5iyR7oSnEpAzu8fvKIe90wZKfi33qNyAN1iGeRnXhi2wFSKPp4KLWGxA3J
lzuoaJdPIDEqfItgOvoq91t+AwlHQvMVL7UYAeNJoUczPclhhDVi3Hh4PC9mFEi79fF9RS/AnsEj
idZ88Gy3kHSaXhb5nvoKhqYH+y4SnFSeFqKVmwMr2bYqvyLsjwql6+07/s2v2ySxFuyb2UtEelzm
sf5WuqUkQl3fWNpUx9C42vBCfQZyzCPVY56Hn37V4MnIqPQGUQluiShKuJR7qqOvS6+IclcZfP3O
raoP8Tj+0nAfpEHknFYoMwRusGhz3ELd66Oqhon4FGvDkyaVLjzOidrY+kIVpD5PCi6lb0hFn0vz
GoHUMkWKbVuYFO/einrlFBVBeemPg4R9taUif77Hl9lyXC9HQz/oEoVcmWk1RRgbdtXwshh8y8wV
DQoVCBWCAvGOFUrH3n6ye8qgzvvoiUMwtJaWl57kgIIKODSHqIwEbdBFYuGacdesqEEfK9tuUDjo
llezjo7sL/EDl/Onz2wFXFVCJ/k1tGPpn8nA1cfSxapPtBrU/REHIk2Zpm1regz8O4RD+lmRl8Zc
spruxAx5fadmT+U2kYTt1B9yZ+fBhVn/xSmfxfrPT5g3hgXH3Af+UgHAN7+7hYMdubHUt1EG7mjn
/ZSqqXDEVB3+iPdt3KEtebE7PCA+2JyahCncalGiRPp/JJkxxWDGnSLVPyMB8WkqEnOi45x1+aK9
4wGJ1gSHX1NG9Z+cAyyNlhc+3IHAdVxyxKThA0hEznZFyeJfvcsgx2VfcAZgywy8LiZgMnPO1vDf
oKB4q1OTWBrF24pLlWfXPVUV+KbNewhk3q4ohhHKjXUkKyeQFPSS65KMuvs5AdzFCtKwT5Xu8Suh
7FTCt5DUW54yYB1ZlegKJ8r5yp5ddlJKzr2bvq2sBSL7dB/CpCevZCp5pHkbRspTO8VNg3z9CVng
oyfUD6jK54Z2+k+E5+3kP22X1uHGEVAu+/cN+L4ku2/H9/cxo44YYy1r+ip5vHydBxLsRAdGSXGE
WYi9Yu0hhPxZ25rVARWVOdvry5H/NNMpR6l3ZRYlOoctNlMkPtGQFdqxq/itOa4waPF840niuYVh
0uxLhIgiLTOxnQSBWWZdkGeuMAZHoDPEBM58HoXXaiVFZkQuTMhNmSBnfthRzLA5Vdrkc9yvKKPL
EfsApG8MOvY4uqQUQRUWb2SiuR6sp7ELoDfw6A/Ki22ejw+8LPotsYsqEZ6pe7xLNzXCxgfK4w+I
jWlxRBStrWtCXWoAsV05jccfZNpr5J7OM/GY2CMeCkYBgVSyr7sHIaP6feULYXewVrPGWbACFcEY
GkxUxkMY1nHJISsnqtlGT3URoR0krzQwcS61KLq5ECvm2BilWfMvaZzmIgnGaoiwZcPFwi7wNsvP
KLvC9sxccmBBSmnJGmpIYF1dhgNViekHRJVFQSIVuXFK7WklvnGdu1CsoZYgpwqDuQ2v9qlPOlft
Y8ql7DqpLHnwy6L9NOp9cduuzmYX9pP367u7OTinJcZnj6W7Ms/0+70BTxVEtbobvHsXmJeYE3Gm
EbeZHsqoESa9XFJL+FvVe7jsjY6CGGRujFZ6TrSPr8a5iWZszkkOkRoK5Kt620v1BSGL8zf01boJ
zW9r7sd7tkgBTknz1gL4Gwjw/Db+6LzuWBGV/WOFoIf47CAbsBvTHjvPv7pqCcMD7U4P5RKdDlRC
wBtMdvahEilORZQJLm1pGSpTLfmYs5UkgQSVyUicDm9XpRjj0buQn2SZtrGzH76T+09QpwDGKhIB
TOcZsfvfDgWZNw1h31b59E15EkcpDbEA2axrbzg9SkDaa+JqH1FYRUHGLqA+0fy2ctlsI2tCi39/
LL2uR10sXF5wqxnRgGPdzFiIL6XM5kfvDrIIsSv5ZKsagl27BHUqWhTvb/QfxPJUb5UCn8rlTx54
ym6l8/P2BVgQi2vnexncbwLRGECMySgKYS9zmfGjJrQgk214qevWZ04Jj8HoV37cVVl/gk6eyYSY
eMRDXeLqqTo69gxldooAU5lyPldFa0AwJn0RILagDlnmgEfNz8fA7s5AiMEGGcmQQoDhi6hk8Fkt
HWc1523fD78ETg9CudfSXZHtI+8Ffdws39JewWAaCwSOcWbL+Srz0fZk+M4iSkT7G577gBp5RaNN
IQTvFDYs2suelY46Kn183OYLemTlAORtIvSlN2rSL+eKNJwfbPQn5VwThUiyowreORhGkl5x94i3
Ep2XoSRB7Q2y0wQJMDLgo5tS0MSh2s4uSIlJJYGVX3De5ABCI+sAtujp6rPBFfjmcNt786dAcqux
+CJpDYnXxYQwI0FyhIVsKedchC7r1ll4qzvJC3Cm0OVBeeTwuETYisC5Qgx9mz75A02Aya5p7jzO
TIwRZQGbtNpLSTxKVwhPVCiSCheGJrChyBA88jj1n1LKlABXXY32aG4fRvrcKMTnLkYyCajfhMk4
FX+eKl0aDmDVz9POcP1jU2iWMJ/RTAOwFwmjruNYnjQrMmG7w/cP7HiXChrgbIdlHhur8X868q2G
slLvjv56lBuCqoq7MwzZqMINglHJmRm3E8BkLjYcYqNqQg8ML/D8sDq7bBxYvV++BMHJAn6gmn6d
rTbB67TNW31tRdsIr2RKhKZEHNn6dtVm3u0hnoh88C/kwJ4vh9n2aQi3Q7cLnCsznrNnTzXNFp4S
tUmY3cwJXuwn1b/QRExCK2VRsbx0Klq7CwKMyvH3hAydlOmotiYc/EBGB6zgJOc2SmiDmvDZIh/n
AaenSayhN6qod9g6dTMVJkJX5kF4H4dxVjnwe/JbN23gxGSU1VDiR77G9yiXB6YMHutPcHW/5qdh
k5JXudl+WJRpJzJRFsbe+ylg+HPKlSXTQfygSpbRpLIdPxhRTWfkhUmDg5K0jC4T1xLUvgWRLy9D
wgBrDehFMH02Jhi9occKCTV+ZPJGMQEccKMZi7J7S21SlntianIFG5Y0kepcjVWJff2QcPu9Lcgl
BxT1zbZLJ/8pp9K95q7s4tXypg74kuGqlFy5EfxzEjNULHyUgbwlSfwnpuYm2KOxUdeFZ9EO8ql3
c1sH+iVdcrkvEo7UxZvcSjExAgRJpb6tBFvyms8klPTB0Do5de21/8LyjIKfcjWSobdaTdFTDqQJ
7TzwR15NHvp4qZgfZhjpz2Yw93g+9QEmuozt+slQG4SeSC83xlYbexCAVHYq1H5UZxfmDJoqxPeu
wtIHA9kj47qROD4/11G7/yxsxojc/KFXC4b9aR08ApsUvl0AwmOu3l+6fdZgzruoOSkgjGXe8Zxb
nCzfzHTieKk3L8VK0QyE9QpjupzaVu2cMjH+c7C6WBVfkTXc0k+CytU8Aez59nZNBuAQKhOB672K
DHiJs+ZC3ssDBp/j/Rj4TU6QfPjwHOLAx3YhN/SkE2u6ySfGeB1VclsPYmKx3xFnc6OQXDAAEzfy
nnFLXFZin9bs4q0ZLJdmNRsts5ZkgRaF3is3tsj8dDQC1+inlez6802O6+w36rDq/ie41uaAL8Y+
cg2U8z+UljYT8wiNGXed/ucL79hdoMeU4m9OGuaKzgpGoHYZ3B+T6QXVHfZ5lVBDt9uELk6EDZlj
6eF3ST+z6k8JC133rQvb3aawYbUq/YISd09ucrV/v5cW1uisXEDCZAGG63/kTppcPLU4Uic7vnUr
rfWTqZUty3Qm8fYxv8rS3chb96bJnbvCAfgfq6W4uF1/+jmPwDjdunm7djW4t7uYzD6xNSF3yFse
/xXbRMZRxODHHvzeqhgSrGWN5JBqSOBAdrPhhKwOA/FGcea9XyJJfkOgyJTsp3lOoPi0o5wegjYr
L0cwD1Kj7gd7ECYmQL3M+oEL3J4ksvmvXwsN8nn7aVXZiQw101wGUAWsSJY/CynS4YcYjJ0Q2XZL
wejtG3rPU3nb9jMye/c5rIOZ+E8EvHpnP4Yp+M5LYi9jiRd0b8it/mHhmRvQSZuhIsT5LYk2bZKZ
qUeBWGlL0lHs/yQjiJEZxT3k8S/CMMMidC6rMb+XYZTEwzBhLaRBU7oDRtbJt0SpZMW007Amw3/T
kyoS6f5UBJSxlfYbSFFLM9tbej/ExE7gbIlrkWaVyukTfmzNq4JPWif4VtRW+XaxBgj2ATMoIm+X
qisJ8ZhEtGlHxZg62+y+yNa1mkxjQ2mvnZcvvd9nTGbAFit2h4OQxYPBW1wBSkCWOxcajzcV+juH
MbmOyH1XonRWpT2ghHcyXX/Hpb0ZtUmcEe9FHiXr7zdhtj2PkLyEzVgFrJXP1U+/XkdFOWjIH65+
p2bXyPbWXkIffDRSf7BpDjFAdqNjWRpzeR3GQbDe5djjJgF0lwDEIxeJLhFbtMTxuKvUd7ASNuaO
Nv1sZ4gRx6ntld5bHY3nZBU+4HR1hEL1WQkdp6YTlUan/9Da7soe8t47zOnFTtNoqLECa+Qb108X
Npcp3j13U6VbqpScL+COhHSRTjIECkx+Uq+T1lN8EWOneyGuq1ISH5/TCS6Y1v2HLqTY2l/N/uKA
M9yLRhil4ovPpw5Ikxb10SiYVQogRiJWM2qNW42ORlqWWDXfKQGU6ec5A8+zlBDSdWxbdjIjil8A
O5ErH7C+Ab6r1CjoJy7+5y44oMfVs2zC5Ve4g6x1xxABCpmc1plRmTYt4L9ADb1tFpfNabIilSwz
rbkDKUoyza4NCKQFPvxSD9C0b2lNOuMHUqPcdmpXYYFKt5InrvmvOZAX2+fJ3JOHr0ArkQLWGxwb
oo+2Sqod/jfv7iRO4twX95GFM8S495e1iv/PrWi+vvR4+Bh1BgFcde7SEOAZ9ywjWnrgmGRKuCAV
06oNlX9oxIv1yRVOMz6tm1S00c5JCPiY4H7CwJA3SDYxTTGMclTMaYujiz+bszlliRRpSISTeECF
7aXVJUp1wK7haOzQsIrw8agp/7fM/bmGTnwUVr3eBn0TJqzzSOnVyiXDj9SIBmsyRjVJSyNkGT2E
ET46W2OVDJ1+krTdswyGfJS1Bh1ECtPlVTMCsELsxriRjcjIe2KuX45US6PgL6U3NlrXAtvSBMfX
G8pZ2R0ZQoAtDcPYRMYIgMe0JfMrZ0xLUVyekaOYBxUBkC3yBnkcrMVhEdHpKwgXqMg8ZKZPWHiS
xytLXBvBEhPOHzVSOG5woEPnl9r6TDBg2J0fRbMhpDgqnlIwywJyB31u8VG8rWjH+JnQfVWKfra4
spw7mAS57E86jfOKrg3CTkuX844jC5Zz7xuQ/CxK18K0aTR7UwRiSn2P2AExF3toSqJsttd+/KVx
4c8B7SUg+hHbr9w7mvvoN4P9ueWNBEV5BINW7UJZNiLCRgM80eW+azEi9UEsOoukPpJwdS3w4MK4
wpUNAMjXxqfK2NOjzPioIqA50SPetiE21ZvYT7j4a5YFFg+8ONRB7xH8kGpxf+olbP710V97yb4z
ZQfjCqgGwtXsircnbxgGLjepDJ/nUVdLX/eNClNmz0v3rR2E3QxMtIy07nGgQxjcKIpcbqoU8S4a
K7RUhbfszTNTSJyydIDJOA1tbMJjYwTMhYAIml81WyVim43LEPI/EPp56heypSPl0zZqdBmUOvzP
1Jk4vo0ulGbTcU+IXMfF4QxLQ/NvxfNMXb/Xx2+8e2Ot6736K7ezLnb0ntEwJltnM+zHO0TT/kYe
ugfbpJt4D/subsGma1fuKG4+uez76lpyWvBDDFjHTEaHL1njixgZRsCoEDQenISnt89ew16oes01
nPZdjiH08jb72xagAxzRvikn6k8RG8rKPtEA1j5oK7maPTc33plmSTsAMn0MRTueH8WEccH0r9Cx
7cIB6fdOkCmB3+PUdr7CQ3fg0G8osf0u71abbvobiPlB2dm/Y1ICgnEt92niOUzuqGT5b8iPBcyh
Bs9xErnVfV5QGWm2n6FhaJ7e13S1Q4rlkyJv+8W7QUgEUfqJKQfQmD9gBYsg2p4TsrqF4lmoGnja
sY1ndgKWViCPbC42uYcLDzXJaVJftyWJKqeF0dQ3NuPmMdkARRuGtxCgFtAe+ULKg8KnNFBtKRjB
0JGVc8ysqcEgYl4ZkscaOdn3Y7UVEU7T9P5H1fvWKOcoG9e+k9Sh7WHqn1VLi7Ir9Idz819GN/27
Z6SODeUqlx5rbC63IzWGQAC//J3TcguSy7JyWXHBBqfd8wtejtcnQ/8psUkK4n3MCfAPg+BSId1Y
S1srYgSu2oTLx5zIEiOpTOMZwdLYjW6QN+tDpw/biOcEqWBZ6VR8E1HkXJcEIdJgz1XqvJhOv8jm
gA9rSgPVtoajP9KkTIPHBC4jhQW8SL/9rUHNpz8vvFiS0jqAWknx1Mg8RwwpiMztf2ES1ZIafbiO
JV9qXn450MU3MoDjqF1vBuisw5rXQ8w7QLrLwBMKGM7Ue/2UlpkIWry+fZiBcG/ZfDtNqT+04kG6
mEI6TBrKxGnx0mgetR1/a9A1FhaUD2ftmdrEQ8TWJBOfU9LytyozGEiYNMM2+uwYaOtPq3u2D+Mg
tZJK0fCb+jZg+sXrhPIZAt/8kRsHKwVYktPUgO3Uyge2VFup89ZGBdcZv2m5EhFtFPp8RLf4m6zW
8h0GPUqVPPS/SxHQn+7+c7GZkBAFTsspxhLf0orp1ORWTVX2fgW3a6aEioD762tqEjKNj2beTT/E
Gq6Ynr++g055VU8NE+Cq3g9lGNRvHqJ5ScPczLYjdHqqUYAG42BGmDPFl9c7ulMaOTsSot2kmcIh
WjiDcss6TnUoJl0JgXFI4GcS4DasfLW5Q6YAKbm14u12oryE0+qryIcb1g1z7j2rV/xuHWnrlWxI
tt7dTzJO7bPFnIRee36kzrG3Ee6DXPkW2G8BMflhibWv7p8bktKQOpfZo18pkjw/DEaIIDsrsNdz
EfsaR9NbKDGW05ZtTEuiytexYcaqthwwHQJ0udhD5Z2vid3t4Xz/8oErtwEjORM7ViK1GsdZkkjm
pZIVhXXoEq4ZLmVh6oAM2UyqRaQ6j3jx9oj8B6dsPRmPTUaM4qCqdLTePAuLDPAitTT9ENBOsywq
HvO8xMy0zYW2ybgbuuQQOIkHcSsMlt3QiY0uWrS2tO3y1XdfwzFHzk4Xc7fsdHkbp3xFk2HomXn8
6HrkDFEkbt7/tteQZxLBumUQaf+AD/gZDcCN8I7iYNykgbZ2EHrOPn64FZf0KcR8CBf8bX+akUiw
V9BsEBNSKceIPRJ7AiszLE8/kezpMkn8jMTgb36IvFDXP5q2+L8VYXF4xNqq3esy5TjG/XRSf8ta
JuPGo+y7GSkLquzFV+P9x3oOq+IlGcT0J47BfsukTv9zh8SVD4pVcr01ylkI7GBhaR4MU+K7gjvH
gkwixd3Oq4rAgV7w6qstDJvWlJKs7X8woZd9ihzsH9Dzy4kYkRJ0ZNbZ7cRIKPx4K5iv5bXHInCD
ySFf6jOW3OOVQgGu2UvPLu1z9JPMOQoSeRJYYzY3is6mmwk2BTj9XNHNLkEpXzIprjTS7v68WG3w
m+6+/aO1ij1WUUZhym9GjEh521mur5jGDX7gVnRCH1VrnveWtJ/kYXBaPtsXgCL7Tr4lw1QKRtZD
OpUtol3Rd//FOEXFbYWk1MiIUtZ+qh7SubxfrBZYVoRiORS2tKov51bxdGSLNMwVhyhSsG9OGmAJ
MpQ4hPVYdsQ+1wl0otIHvutemKctxkj222iffj1/G2gMgalQhSe4y+LRRsJG5vu3Lt8b6D2Bk7Pg
SOmIN2N9xw/wZmjL2eUl9QH3MUY6p39ZFyFxReU4S1TDaWBvVb58EjYn+wa1df0RGBQkBfnWEj5q
4V1a50tK8pXEbehFXcF1CIYekCpb4UFr4sg5dZtKSEJcyhJw0UU86qJ0zB/v37AkfKYOW0oirKBd
bvZT6s0ePUjXiyeOCERtA5Y4lhtmRUQ/2tF8f6Gr7Fkp45Cqvurr0OvCCLsHnN6gyxXUiTBs8ZHz
/Xqerp6nrrz+Z4YdVSiTH+hzTsHVdK1IcDfnDYE5nJ72zsLU6kOgmXmVgyhryIpUXZl3MZrEz6Oz
3jVSC+Hz728etVfLveJ8tTXPbtyVyJRL5hCHCiNZEFo/IR7KHbY80EanZhAJILEqyRRN0iMGZ6MS
Wcv6UTIykhRQeqnU/aB3r735QhCkx1A82QlC5G8XHuI9CJVWQ4lRyLzKt40tyYCWWHLFQm48MyqC
7Xj5Ysxs3q6mI7lMU3ag6gGCz/gyWC/YIYoVovkshUy2iyhR0L7BjQtpW7iHztmFlAalyLLP3pPt
Zb9NgDzgqM/BWN61afS245FEBQUg4zPnHROcNq8SWK4njQqCuSAZbn3IQ4zSXBHOJHjNjjHrelOe
ZAIqXXInmjtKFV5y8FKy9vmJ5EHbwEHcXCtLOr1Moo0LNMK1eJQzUZ5l/0jMU2LBMWc2F94GUqIn
MbOSVPeS2RTZVADXfARKIKegHQzbMdS3hWXRZIjKnQhIpFAZdopLH8j7bjAfAPj/s1NI9gG4VaYz
d8Q5vKNye7X3Zv8ExlLHTBRDA2QljBiqvrZhARWLAIRf9FUjAboWcek8/YySih7YgPfnoHPDdTOK
k7il0coA7p5ovIJB9kvi3Q89fS2yC7N8POj3hZcQIVHcbIzoxUhJ+jdz7+3ghirWWN3tUsBCTSEQ
Fm1O/9cBWU7SoSG1wQR0mJY1SFY9f+VTeHcAgUdm7Oge4TwVakOEaqb/MUgKmQMP0G4+FQtszWUO
kpnC0VU7mh7URZbBfbhbFNp9MCvzWir8KrRxPk409wPoOsupWiXAX5RA124//Kq1ESJV7nueOaSW
IDnk4hAbON5rtytCoXImn7DFGIk7v3YzjDKq1OUTrQhmUfAL8R/FTkFgDMv9OhXTz+5sbYhtP8ks
iXR887J0cevLm2t1WA/HH/+eHwJaOgyOcdo5qIc7Z5Ze5NKrWzdzu77++pq6j+ltXyxMjVP1dky0
VsWfWK9PaGVP+RtymaMQdncxt9aKPoLi/bZOypQMQKL5LuDI4OkF1hrhUkiFQkEv0XLvJmW0Lqcz
qCQlIHp13G86xESGvKALpnbRMUQIUUbz5ppwCgJaiiCIk/4m4/VFP0UGSmU2Z6etaTSwHbmBjK3i
vys2U3ApBjY5DhXpXTkDce8SomgmMl0LOQn7PLufLHi5pchvJm1JcqyLklLX33SrSmINNqv/9NDF
3NyET/33WglZJkfFY5CNMsz1ZHxZFoHX2tWT+cH9O9dwjLO0XkRgTiPnfHmJr5wQ6qkrwLIokiyj
eLqUmKcM6pkoS38dzVBrwMALQ8MCvs1AIAa5sON/xkt/Swdmgl9Si5uaDxcIY5iwvAoTNXxPVgC6
Xw4+w4fZN6sf7Dkz13g88dr+AeN3sc2wGrZk0oZrxd/3gnU++KD2Q9fUsnZDt6For8ekNB71Jqmm
2RScSp/lXnZXLVmF+/1Zg2aopJT+gGeoK/S4Y/sQ1zzfvEUlBwI7yFc3Nd0O1w0Bvyl5N3zBC2Zo
A3IgQoUtWRyOWzgx6E6pFznOSQEF4GzF7nJyOJ9fvy+nnPOSDj9vgPjVAiQdFsBHVs+AHhWOwDzp
RV5v/3bB42GcoAXgtYN+NeUjBp9wn129TYwNa91oj5DoWbxaqGkOYftlTVpuAJxlrS3sI+hEWOMp
b3DXDDWCmaw/ogo3JGXF3+iNsqE6Yvf98dIpYzZJh5nOmQOpQinXxNKjVGhCIiJwEGY90fo+FdI6
XpR/tuGWqQDMv9vxxvktUGR5HAbvR5WshCPGavalpwPLpghTjnHpRj9Q8yX9eBaBK67uTv+V1zDB
awLnvoLCxT4c63YrEAFp13imb76DG2comt87wLN9DP2E1juiZ1tLdN3QQGzdhTKbGBAUfWyHndRN
VtLmJUGLqAH9PFvgwsoExrFWGtK/3sL5r48U1ZJZuua/daCrnBKcrQ0tVR0kpsrJnub7CJMg91mU
VVn/uvPY+ETZmGoNiSfMNPM88G0TXq7hRjgv/YcDh+dr/xlqf4nTVUt9RL65JmMUWPBf35SRlQn1
cfQe0GMQAg1LsHfKAOR2lqwTr6YVz8n4dekyHJ5wUyjgqb8SA4Y4BnCBmgMffDzB1Da1eHIEWDrc
djYSDY9ecQVeObmeTyc2u/7gJTxyaiw1P1GMuIAAMauCOBvi1KHyCRdoxltElieUAyAuwmyAWnlZ
HPg+M/ci1sQ79cvbPnEQ8Vo+vs1S/is2WE/vrkzryaBgxRc8BlYUTvNV3VPL9N9+s+u15IozsN0z
n+3lvVXf+220QPGFYeU9Hz7r6xu+RN7Bs69BLLDBHZazX1mJ8s1Fiot0WnqiEZlfBdbd/auOXbjk
+GJM5B837fjZTAfQncC0ahY7lezq5I2QYbV3jWQyzQz0E2VZerHLNrZaIkJsqXXUFQzZpHXgOnpF
kFTDcHZlQhJLdfFpD5Yy0ex2pMDOf+CeZM5WolmpiOLSw83ni5UwRhigH5qWkFHrIE8RLd8FGNBw
bDDNwu5bUa289jLC1IhS2N3AKOe3TkdsmOe8rpIGKd6fGAAr2KnmhjsoBzxjkCpjPpDv13Qoxylp
Ak0LVK9Eg82E8WZpzJkrITt+c2M0Nj1m7OmS39U8PCjtnvutxz1LeQCmNohh3x5e3lAXmB9fTrES
dIU+PiXhCGqYGZS2wLUVEYiwW6h4XFn4ZDuxdcLZB2dXsJkzrR7b+fIakEhIjTbbeD4UxG8jZuif
DrFeTgMs5v2+BSn0k5yPKTmMqz55h3wYbYfyyNsWE2Tf4yb07wJHy5bBHXOIpTK6nFtdRzq4G0mV
2+SNcnz1ADLy7gAtXQJmiW7lUL86jtBft3ynuhUC0LsX4dLqyb7EXcq0nDjDX1qZ9/0yHvb+rCJO
dr1FNo8HGyh4XnpgssUsM1i45Yyigf0grdRySkv9i4uTRpuDE0JCrDDtZs/b1k6nqJutCN6eDy+X
zJGb3peaACMCKXPomYpjb/7AOXMeovHKczjmZ0Q5Q5H15sk7mHtWcJs9CokMvMf2GB+WfOqeESrA
jOuYjEKw+Wt+t2eTIcg2EEMBf92bcQdZ1pBrQnliqXnP259JuY1vvT5ltvduG4FXf6+K6jciGcVP
rFDz9ahvfHxL8vDedgr6+/zfoNU3xSw7prV2vTe5/RPNT7Z/XYx1IgBRV0ttBAJh1FCyiF7sgXP4
MnnK2uhAF5mc8zPmMCRZ0cRJsiW+9tPRCgNX9c2uRHEfFUc18psSRManD+EOC6Z5I5eWcSN04fim
MGBpD8jW+12qBlqCOhohpQggxkh0EGEVMsEcfGgjWbRar2gbG9r0X5LRhKPaQDaGl9chQPYZbDSd
K2zM/iy6gFjAGcoChIL7HAYm7yi0Gq0NIhSPp5OJH+NOdJK7mqbwY1GRxYwoYCMiXnSmIZSGa1zL
+du7mYmi4R4vzJefhh8hreRc7DNiFHokI3iwZIj50L13VRGWsKtp4fVoZ09RAidB/NrtPIYeYArC
l6Fkw3tTzf/nrMymGoONjgFaKExC44ZORSmnZGivFurWPh7Q4jhc9lOIDUTyl6fbynfpoDMOSvNR
R0LFEcaEIRUrgkTuCmQu+Qryu5aKMaByODZ3fuTjI4X/zMzchgxJBc1lY4Qb2H+TMWz0wjaJmna+
leteJSfQuo2vkUivOILqNinsrn9DKhPLLfCa+ujfT/DMJ4WGXOmcvQ7QCST2n8uRH0pxPEXtHPF+
Tl00RIprm/+96D9cy+cFyVLEAbpGQbpPvczUQvU8w11ScWSYXumKcEnOZQBzfnrzefNAaXzvgMLz
EjexbP2OyGNh2ysJL2/ITtykcI+FqQypwg+kkJH+VrvKg7VRvAyLjMJbackKLl1w97cDgy9a9YpT
QpoNSk7DUsfDiYO6vNTwgRvajjehMYgISY6Vb2i32bVxH/DW98xkqB6yfBRJ7i3Vzo8cRw1npIl3
RImmB16/uxICUJ+saJ1lbpE5AhCOL1eI9T62G/pjVvFuo2Ts+L5R77uWnaNwvxnPj00U80q70e/Z
RUZ51+sdPXq7HOhHCjXhNUUNq1WgnstV8mMPEmNC3HznpY/1WvFfXFlJjRgA5fZK0EFr4ay8veXT
6xMaD8WrErwH2xWw/nKshfE+rJcLuUOGHPe95z/5CBn0PAG/sraQrGubkGgMrwj0sbzoivDp9e2s
W6GvmjPEDGrMBK9aFpkx39tAeLCuLt4/cyWuF8/ajQRt3601RwZZcr8Ubh+dGT/DDnHFPYKhx2lF
v8tx0RVnKpp1xd07Igiz4ROIr5KQvcJNtFmwE2ZTxpNTguXR7Wc6cGnEj32Hll2ay7U4iYT+vnz4
GMd24kriGjI/gZJs+B2qC6qXjr7CIPraOkvaV2o56wMqIKxFu3wWGOvU2dLuHVEf060fVX2sfd9Z
iNTEe7G3j8bJ16V5h6Q4SswYZgSEy69p5lfYP6aH038+G1A9mLyYuuDClUFDngkuwUSckWPQ49kw
xT6iZ7XOW7oQ7n/ITvEFJQ7q/8vr1OQaKNTuQ/HGFyNXmeVVnIHwO3ulQ4IedJqMevJ87qbo3/8z
M/UW1sESz8gzya37cDKkWjOQncZkvjosOEqDiv4GqJd2Leyy4SB8NlJXfrrRT7ag83jHo9BODpFf
SD42rELNVhWVGpiPwtk97+pudAhAQ2oqAuAhDBCetk/TofafauumMup3XuNTMhu/ridbLK9MfCh4
JkWgOENaoqwvdxd48WnVw/XWkhM42yPRwgl+2kvE4BgnUVYaMrz/1YWSYtVJNQGwMHjPWK4PUX4y
Ew9TMubLpm8fMeDh11zw6FnUZyCbSJqjdiv12b6HUjpGKUJntdpXa7G9uRYQ/zZisxe/TaJcI/6O
CKb/4U+/od7D1Rv0jU6VSNg23y9jUL2fcV5/7hbvaqu22OxXXGQ/eIb3LGfrf2yNnZsynYqkBozU
c4umlT46WxK7Fdv4ffcQkuskefn/gKLIt5HWO3ZJAls60h6EmaUjisttKDpNmsLmm0INpoYy1cu0
jJjc1Jaygf7VI9kaywDEJFaSNY/hB/6xeT2tStJw3e+MBN7ZW2iMU1874m5ZN7FBqwoQgGj+2GqU
g2qN7EmgdTz8V32INuTdykrUbFsG5giEcM9k9jT2Fle7fBehuYH763jo3DaQQs9fCSbcd5hOxdgm
ct08UuZiED2J/Ff/LFdmsOkrXJuUZbegzUvdgrvskSmveZvYvyWEJYTFLvU6Ch8YXokSaf8vChqy
bbuyWsGCQfYX6CdRHxnV7akR8DE15+dZsCTqnP0oJrGc8vQmn15JtRZltjOAwGkE0eRojD3fifJg
Tzrylpb0GDqOEkYb3ZMC4/9ISAuXjbECf65Bz+xKcvBfDL9qs4holuLx/W+25JtXTyXf+Ph4rVUl
kcolfeb+n71r/r6s3xygD2QTjcDq3L9BmemeQGxW6yfoKTfQL+Fu76EDcu/s1GUqbObFk1jkyclM
x63wv7GhXKSaRWpbheGDyzs6mPDwPrhPnvLeqfeECJtiVdQ7VS1Fn8Tf7SsIprGirLa/+tKmVOzI
P9wS+1MrIgn0edlGu38BM9R4jeJSNP5Uoh5Dj0r4CFCEmcdLDlOt2BYtOmJwc5MDZ2SxrxWQJx72
grCQ8L3skHkwTxjFct5mEPBu2V/3O453X1qhjXnVQsrOoJ7xEQzUXnDjVNo+4VrqZcEccdzUVJh9
nupBxWKCoTaUOiVmx7woK0ePYaTB/1uFp1P7pRZgGysdflQZPnvKWaBPef9ckjmFWtrdiopnEGLx
LRdT0/dNfSqm6YI1WYIXRZ8xYfYIhOFrC6T5SU69xUiCS8sljQxqonhpk0tbkP7Wy6lp2qVqVhbO
STYLJKVlElXPeM30COAi6tjg09XhTKg4cYbF+rcKYPOx3TtMda/pSrhZBm3YPTVAubz2XG9Liuha
/bov8/QrHyyDXz3vCT6QK/xp/J6hDzFzph03UjYrJpNZRnW2x7lWadCN6s2ftcXvEQNA0RAF5lg1
4CR38JZ+W95J8iOjKeiPKJQPpPTTyVY477WJ7qpIj9GFbzf4UO/7mEeh9gR2y9SNkjYNRRbWhpbI
F3++3BJO+YaSREbBxevc1jcbuWcyFiQYlYobuw/MxNsvb4Gq4lDL/bJ0hOzkAqvzJCIQNVv9v46S
Njjty8e/9J7UD3RSf1r5rkcVxFaEAQYn+soghcCy83UIxmWFJHIkxGqOss+CyxiWdlhsE7XAl9F9
anSPFxe3Az+t01FNOmUKvj8SbDj5KFSoVABIj1ql3LFBThAmmjixvyCISwN0Qa/2dqgkfWlX3dyj
Bkr/6yx7nq7Z4Lwqu1dr9OWQowPJzAYxl4VY9KwtpuaHfyk+OgMHjD/ea76HHKApdwzW3AKVV8Ts
bvDfTa6PHN3ntofF2Lt7kkiMRlMea3yPhohUU/dcqtUaqBGfz2JaKhDWCBnP3AKlRv+T38AkTq4B
hL/ViEpOiN72F/r9du4sNela5RsHUmrPBSirBdXZWDanqNn4pdATMreBu7JHlrad7Hs750Ofm5Ny
mGEzPyM9LJ1t+siLf288qkO6+xq2mJ/AV/xcNIKnMEkvO3t/HTuO3RvqrJUWphwZu6H/KtBnted3
PQ2mUIiWrayEpSuPhvAMGPlKWKj8i/07V2u2RpVexIoz2pfq4irhtsfr3qPIGjudTsB47oTIKaZ9
o72Ci483dot3gA02Txb0J2VateXr5P1Zs9R8JZdH+1s+B8OLDW0KJYKnG8mJAL5M862rGtPz6Iiy
27LwaG953wHHhocLpLzuTyMHl6p4cL7gmtB7fnd4yuGxuPMMrPYmTzEunu28cFaNj7SOxUqfK2Ht
ODjR4MUscDBsxUy5RUbsA/dbs1yE9OFVigSGODBxJ5t7CtJNw6zaIvN4KJtyzQE/uOappGelmsFt
q2bH5d9VnHpfklYf8LX2Utnx8xfns5v2nnYJfuLCvW3P+mvXh+Mlylc/z/kx+xCX2GFKDODtKd//
aYowrE8b68tPfEmVrOwPKEdGq/Ck68MnB7fzLEpjwfIxCpmM8y8DPFJTA3OEUPbeBScx7JDWZyE+
lPAbeZGZlI8t5cMLSZNcpzNaXgFAnuA72Q0wEXpLaBsOKpSjrLz8LV85q+r9EbXeK2CjFUvbg+5x
AjV4qc0Yrc8T4a9qLef56Lz57F9UOKgg6NNdCqBd7AXtt5C0S2CDLSX6JwrJ3ll+ZJG1fiXGt9Vc
xrrViCb8ALsckck2o+BFA+Y04xFXbvlVmfFsOdZsZLJtZbigO8jnPYVnzSfZP1XcFCVOu6xinvrt
NGvUnoJJl7hlqXoVNVInzqGriXhj1x2kxVrkrYzZ43WStxz6wtrqXbOdtNdoINQr+qi8UtoRZyLZ
WlJB0XQs3bWJYVfnMVcb0WTiXtv5PFrynHlZ6Mo0iJTnD0Ujazs6yHq4OrGBfDI6KfOeBMgbO460
Kd64qiBXuNklcwFetv8NexLuXrW8cqqsAK7J9nK9OKurGhb0MkDVmsJgn/zZOhZLUNqdYTAg2n4k
bKhvZpGWGw4BfO3eF4mjbPjMXw/wRiY9qrCiJn89u3PmzKtLxPKqFoWBMYcaZtAjAlAtFs1ghQCH
COIGWUAPNTdEVR3w7dq2frC9TH9JoAICMpdQBeteXR80VsFBeUGt2Z4deGoUHIMimCLizrSwFkTV
xL+CfKWXcdqedTeV0JWDhpUBP/UguHEQBnIdMMhDwPHdOSGPTRHKuKIpRk0huEeyjL/4jTkUzkWz
IK56ew5xMA9t8G6l74Cagc9gvNwKSCvmG3r2a8YA0XWJ/1Gtq0C228Fzrp1jiRaDa9QCcQE8Ff2l
/S9xy/4ZgQmNwPpGGEQpLD9LFYgrjn6CbSowQAvA4czNJjGY32wTwJ/2A8Aoo260AuuGMUaml/29
MxfCZ7eR6M19G3x7XbV+12KOtWrobWYGhUHXWvkNk2LEjbOJjgAP2vDx3rp7nwrGvZyTXa1N1CRE
uJihY9gm9g/APs1WqpQfJV78mvOq2a6eOYCYEkM8ku7FGVaovl+8/42PRCYVJzh1MiSGlrNUCt8P
mK73NTyFiFGoQEpJIL3B6qHzjR8hzKQVLp9yqHJEOfNOG+L/qhq0zcLtBxS32gnNuiAumC5UTRFn
15sLInBBue2wPX6TshOJhERO8aJarsfG/E//RuIYkP1hiD+V9N4fFYvNNoNV8dV45GAd+gaDAQZa
vE2NEUq7Pa81FhMZ+Be4qwMZGI/0gkcPHhr+xw7tULBbCkw+gGxWbh7VBhYlgejmh46FQZBXIj5G
ngZ3yOqyG7Uom5McFMw3Mbj61U6Szz39BXWRgENKYdHo7oC8SoHDd+QbPvVOPOpdLnS5yZtt5Lhx
zL4647s93TJ2eaINl5vgCIMjZjsLXRXjHrb/DljTSgjBSsPuS3h3StZW+K6aFGXyEkegAeww0KQB
dOUIcmOG1QgbANvlUEJZEXZZ/ZPmSQsBbHYa74eShW1nH7tPf+Lc91rRHRY0FAuREh7sTYn7NOKO
xoeWRnHzgQAC8d5UyJ3B0t8rWV/KCHEC7z4G6cAXdALShdpRsO2vqLp5mBnjbuDwvtg9p1MJhMbU
rHXyx3S6OtZOaEkf/Uu0D6Mr3IbsNQKAF+YTIIU96Mvpw5nLwHKslEp13JbBG2stQJ0NNFN4ytCE
b/1+h/GHnTmuxqpkw4li9g8HvA8y04hwLijdMiPCyGTSIUgnT3wZHunk3OW+ug0M8xjvw8zGjZ3W
83Zo5Buiaa9bKHhWrM/n1/ExebNyDWlQMdcDhUG+PfX5Rejnzept/siDKxZgeg2yvLgNDyHvoeP/
MXrvTxAIipnIocUpo4GZowN416pNHqtEnJ27Q5aXuLWiY1ClGhbMU6tjGDqEC8Zvv6E2KJsEFQEU
Unks88KeATSxheoH8U/2RO4CskZqiB7QRbKMihhF0k7rgGiFec2VN9gwI1NtGQRdmqTnclRS/rZx
wW5NgSr269IZHPrAVKvB+zcJTCmE+TvfprankaSAsWNeSwCrPrlYA97sYh1+PKcd6yhU/c/WFj2x
jWpS9ombdBWic+UQm6xlYECy6lL74ZHXzHTZYYwEbNSa27+i0MYTLIFPEes4MsuGSFdO3dV5m6Kq
9hCGLyGtt48ZSvEog2DNQwnM5hRuJeboFSqx4LVFrrgXokh07PYpMRYatNzePnDr21NTfRtqkHRC
964sweIOY3bPrFzg00JQL91CSOjoJIbUkL4zfgH1DFQqfXBOnGFSwsU50x40K4Dk2lOCo8UTjYFK
ajYuoPUP4JtM3WgZHqmUkMK98S3SBlUbDcksUjzxtijyqj887DFuYUksWDzP7nUtoeB0MzPaQVml
bHPEgv6k9cwG3tSC3V8EQXWx6J8JHLfP8Dhr8kynGn2WpzfcvVZNDZ5ceNcAT0+/lHZvfNslYI6O
io5cwfV0/a3dY2K4/Xnr5LMqZ8z2XYhK7hW0a5OXZDZmAAspg1dkjk5u1ZWU5Ld2XW+Y6tYPsyja
48jTUw5kq8tSPpCqf7dm2XolmvTJINq1zRT1XP5Qe61vGKE116ARay7562nMn+EdvPayQXmULQfB
MyApucguqZ/Zx8cNJcVXfq0xLuVT4bjU0nktbLbwZasL76uX67UTi+M/Z+Mt1wwm3Xh7pold8wxH
mvYEGmuxTmvE2zhchBJ/45IjyKV4ibm2g7FmAqXtWBOjKnYNCvF+3g5HWjmA06IhRqRK1vV2D9eQ
kNpWqkEmdiiVnFT+w8U648f9V++sM9akxXnXw8+gXqv2kSNvKah5YDbU0I13Xj1ex8a64Y0sprn3
IAzvluQpGg9MFlDgdQPwcN/OfwxAka9OVVVS+sagF2HNCDjbsDBHLF8M4wCja2jRYJuFD7yhscwI
HcxvPxcVKecHX39BdaiKf7+SBK5XfeA7fCfRvbPDvkd+5iDMLX4mVTHXZ1d9xNi9OnhnxwOteGx8
RD5PU1DcVGo9T8rAhXJQG/0c02JNuhiJnxY5i5LVLS61DKFEgyXU6/ZZ36XAhpIMNxtq1tgWL9Vw
xesAVEiQqmYQK4TCdaBXbcMzc9BlPDZh6PPowysqnedBPzUwfyz+coWiW2vbslBzBEBOMt/b7sEt
kx9afhbrFsr+efGNH6xKqbl/i4jlhGyNmFEkEwBI1AFPa1F1s3lgi1qQOoRNIEqoRiPrR59JnzCv
P4r1Fzo4mx/MJL3wEDMsZ4oDNHc4DlrJ7R5MBippLMSbsU6/vHzz8j0srOY/IiXxsQRfCgKh67gm
sX1cCtwYd/AlJEGqTPqnFZcAyUQ+aO47asvM16vMzXSg6buqingpttNcrTt036s1GOvwUeWSwYe5
os/noATf5MFaCCuv3V1CQdY6+61C1Ko8dMp3QMV6snw76QAgwasF4hKahVnPe6wIyI/uKGdNefGu
FqzWWh18NPzfZQwG7exXsrx9rSSDvcQXkSwlOR3hu/Qff58rIqqkmY4hJOju4mmA9OqfHSYxucqI
YwDoSg7rGw6rDLz8tFY4Arg0+XnxHcfyne16/fP8VYbJtFdXjbdC7HBOotEVhXM+LnaKlYRPTZHx
nZBgucp2Z0fYJG0UxNeMQfUb3wVlYrAUszdS8eN+eh0N4wFQww+NCz3b+7Mi4QPggCpCFnoUS88r
T9Z+pPRaWhEN5ILCI4anoN257eUurricjrum8rClxtReyvFT/TeT3e4Hzzo1hCauAfj2vFSeex7K
goNwjnvxHnteCunUydQfRGlvKxHD4OcKLLjGPcM/2oV2a+dX7T2n9loTHUW9sl6DBn5R4/FgcGWN
Pz+gji24XWnANCOcpQlkcXdAy//RnjlEYn5T2r7r304lAc7MkmV5oT+hqwEr8uz6LgwkA05q8K4s
AJHQj9BR6tUa3yANimzPslTpmaSmoiWYjVOrixw4dmR3KaBDngDnj/KfvO9+FQuKbXy1RKXXmGRj
KQpFSPubzu7uh7yfZfnd859DQnZjovMe2FV6jv5uASHB5WoskhBaZT0EgHMuxVIxduk23bFiJzTn
+ZKb146oUwYT7pc24BJuFYtb8OylKFj6LJj3OYUAMEZKQvDugyQaStzPFoSvaI0lGKqfbhexBXTf
R9ipuGDBPWlNDVptWbnmXbIygETt7XY6wLEoMUGtqEAIoz4nmU+jF1GHOEOXGmlFsf7YXuY6e49d
uDpNuzL7gPLEi54kWQAhTuzIMN+kQbkw4P3gW7QcffcQdhlSiUNSlUcLtnqmoS2YgBQdwOkQvRfv
M486Gw8dmopegRG84Vq3+nL333DCSiNHluyzrdnkcrDpSUYOwK6wWzpcvBWWhqv42BKXWLySxegK
CLRpTW3ztVKSVrKanxSTLH5X3Bn1CC6mRxdJbIu8RiFLzrvPktPEQpyZJpvnrXlUQgRejHz7Ptta
5m9u04+a/af7xpy09JHOtNPNUsBKtM9BNQGb3IcwJDJOt6iHzSdTmc8pINF/vmsfhemJU6hTz0dm
jpcLASrPDpNYo90DNdkKwaZbJVZe3l0O78W6H1dTVbjf9xOYpTPe3bGL8MT32NevgwG3zajieaeR
4CQabpT5locJhYqh/0PYTzTEA/942kwUzMRxxTIWz9IgmDit1K/45rrDXkkjF6io1JOHwaH9+K81
ngWxp+iiwLS68UnMKyUQ8hnK4iHNRGyE3WOInh9UYgd/sOBskaN1qKeGQx9PrmFYUrxX7KRI9phF
4EtmZ6lOxxaEZTiTZ8THn7GosYIJmY3Jyqne9gMKqQkJAMxiprRvVHIlwXsHZX+cF/486zKKRG67
Yk9Wr6JpB5PJ15yj+yOrvDsZmfrBFa5lLgPR1rQ/pQN5tsUMazGXwmLpGRHvlaVCMmumokM3vnhn
SwS6i9smTAmuq8QzvYpyckPHi6yabmEjpPfdcucRVMMUqUt9t5VxFEXR1GHnyeqh84Q6Y/2Vgrg0
LAOpTFVCd/fKCIAJXwRzqObLEKpQJFUZVrMcWTu1qkOcf/bUoAYryu2HNgEhG1tmNPKcczDx4rYm
FqVNQEtkMngtDkuspAeoUPo2wwEoC2EHUcbgbphLDCuHL72eGS77tqlobni12PfJh75kR8xl3/Ly
wapPMlodwy7rw/DiaLtfTqzLUBVCvKqPYM4KtPcLBX3ax6osrIkfJXWiYp2RsMBEl5MrFT4nCfU+
yapPLUp+2lioVeIkr0tPOc+YsUAkcA45oilBK78s8ceqr/Ntf2m1lsOkTC3MF5wHBy5udLtpNM0s
kA5kqPuDJqN/vqfDjCx/wSp07F8yojiUSNPUbTPDsM4KroWOnYQOBWylG4HnKKpRDemmKOg7jNhE
OLd7iHp6hfbMnU9Mpkm2UNXEp91BWzR47UIbnshRY3AA36ug1MsvuJvUIw3qRDtFgs+/VrgbnJkr
Dv7HBR4hgapIzj+vcmW6C7r/WMjZaMcD9YkqVD9FAekf0hIexrOY4DLtyAa9V/A3AIGGLv8shvx0
DaYoZzYP2YbcyJq+rz3GjVpUavO4vKIWcv+y5XBnAtRKXYlsJkjTUrWJciGNia0ARUiTq1uLN8dy
CqfeDpXKL2molUD1K1KTfdFh3YOKc+zgClq27wb5s1VZru4sEi2NBR8ZEcXb2obMTkKeU5d/8vd6
b3w68W6Z4Lui7I+v85ZxftskoVCqE2FpzwS8YAzOeQrM06qbzX/1+JVccNIQs/dwr971MbrQYEq4
GSqlGZjeuOdNKDpUuR5fKWC3CrpriAwxtbhfL95Oy8FgUcPmKz5NJFYm4RtpaJnnpxuiL1S9d5xX
sjWlRgaGSImd93n4GnJxpas8uWGuHewaY4NOj7bAIyl/l+klqLlueNJYJsAXVmEYZ4zipEhVkg3M
3HrnZ6VNbcoZ4XyEzxcVwzhRPjIdkNBN7/jBKGbv6pDZMg7BDa+JJdt9aYE8z4o8O8/DcAd7Ic/+
UmeNC6Hq51XywN54Lx9oTIrep3MD+c3rEqDRlWwOit+sX7emlFFnG48LFVPk6g0fego7d5b5P1IQ
tbEHxgvN3u7Ueg2RM6XpbieR8A/LBhTOPHPNEQ9sMnGt3LVvrv0H+HBHVZrLcmbcbR0vois114dS
WwiLliCFJjlHIe2LEl4maHA0/5aXUgaV+Dis/y8Lyg+sLCKtsHXQ4uyzxCEvfOsI9Xy91uNaBTua
d4IYJPKp9Fz0ZFPKYppogUbcDGkhpv9YLmB88KvnYqQL1cq778op0i1XnhQxi02HCW/RhrK1s+Qp
EZwn73tnJfZ98j8z3zXWlLwIRZStQZw96x1XkdL+d6ofIQ4emjWRlD1EVCOT8R43UZVBmkd/Yweg
OnPXyxuCO7J1J2i7mreah3MN11Q93nuleCIlWykrQKgFHkw2jRXjVt80RAzK97oIqrq5Tqii4oiL
QM2jVHHcYlU270yI0x5Awy6e7LyiSET32glQKQf7IR2xm1c37cIvtKMVpGxXaFH2zGZQG8hn9Sze
gOE6AkyoSCSrYOaP5s74j2OUKYzQauO911S8mylI9o8NueIDbtZ02AWLcsNaqPPj553gtUS3IlzX
sMv0vvA99t6UVUP3Mc9buiRAAmA3UMK0zCH9oaKuwA1R22wnG80upydJq0CMY9VaihBp9D4+58u1
c/sgariBaPRkP5DHv3D0JF+3li6O7GpQpnhxgqlL44ro0bw/TugsBdckoiTW4keB/c/lTCD5Ayle
oGbd9BT8SZjy4aRD3Tovu1VCZzuTfWTdklUWd+GvBTlb+jbfiJ6xPXOEEbVsYklUb9P6qkRpVkZn
zeyrm+ghWZUreusM2WGrqqCvNWVeby2jG6q9zOfr9deV2mDeaBBg/oCzzKsXA4bEJO/P5HWtpqlN
iIQDy5apAXnmZkZPBGEKrpGmmupjnz9fSPSvlpYZpY03l9ue0GAFGgeeEtFcDhks2Gg2grdl7pWE
LIeZ5PrNu1yNcC/EqgFfI+DJBO6UjqYt8pwing4uuogyQ0p7YqmHsQ8AYqneUmiIM9o4TFV1oW6P
S190TvjYTeWAybJANk4+g1m4Uh6AZbuHgJBl4e1lA8z2AVNUYgAffbkcTolfwzcQ3y9AMjGOOFMj
qyeS/Z/wbGW2V4E4Y67ld2JwdPVFzz3oPzp+QGZyGJoYUagrcwseEIigNZ342bvgPORTibw9fpDn
2c6NNjkh0MwiZM3uKdzwoLc2PDDAoY8Ly73xg/SruNX2flHnDQbnDQj7ti3L33KFM7mRTNeE+Bsh
kDIjJU4pBn1QhficgnrstySjeGnQbxJjIOr0/mkB3koyQHRTJDH6M6fPK8hPgQinKI0aRSrCNInq
TXd7Pkr1PrU4kd7C/fN38/9zRaVIaYzGkPCKV9tegm2iZ8dSk3gz8lEyRaAV/7lTuHiyGN/0NHVb
yW5n5IPEa3K8xznnheEBJgMQGMp9G1uwjzmCMXsbqKPl5RphF87DNDlaC4O1Jildf6Fc1eFcELqq
i4hUvnvpE76EJfW5ccZwAY5IietY/8oM6p8UOPQ73oyXHQyjiUdgEtvP7TVFp+7hQSaFHJIjW8a5
L1/5y83QeCYwrOEIHeyPA9W5uBfDv2bhz8YrLNTzwGg8eJ/QfBnRTBnjqwexQjTqHQWr/SVBxzdr
hh8/xToX0f7CkuP82aGXaM9e6bp1vjs46Rv9OTmVM6Bp58mfx2wSY+JcvURPdXe7IG9Qi8voyMUN
Y9lqo5XNqsjM6UoffmpFNzeSft0AlBtTrYr9au23xM274a2WgrbeASyQbjXZO2E/+8IZPDo62ivy
FLeIdTC+y1YkQw1leUlruHHZFV1kF+aoHRvq05UR4DR7TDNz8Z9I69KcKo0SV7OejIrDA3fS1his
gzkh8l9q3GyhHiBdYfxF9FjhnkcCFaOHvyD/FdRg2NoA45Fzpt4nViHEn2aSjnzEK2O3yrHrtgbV
GYeinXSzV7/K/fX11npzQTRNidb3JSxFsKRxRaCvOp7ieoKL6z8kkcbWMu/No/ycwwrA6ZqcBCfq
8+ZNMFIsFeOQ0jHYqyTwr7lNXM4XgDL7tojq/ggzbcx1WfoKYg5CYUnM2dMVUKiRPljqgKkBiYeX
YA8R+ElDZoSqM3MdB5oOUeHtIzVcdkHSqyLoWImJh1Sf2Bro4lH0JjuFGbPy/63GRbrDmqDd0b8l
ElVYCV02b7ljMNPr3p3jgVeqQqrwbWc45tNDDIZXNOeqKFbkjxnbPqxHDzk0UPcGvj2uMzQAg7jW
x29/I8a4QoF+che8klyOxtB/2uz2YHjaLzpFKHVFJPycKhaZTiZcCKRtWuviZhlZtuG4dWlBLNWM
IiW4xOS9xaoSmhnKfO4ZAiQjCGcjm6QWGF/6tbfdeU36bgSt2TQUK6ToxYKvvWiu3rAEW7yr1px1
63+M+pPM2vdMwSU93b3JmtYJmHTgNLBkMBMVMMEDQAvtIEzLv4hv9MochO7yXs98XWJc5K+EG9P0
WuqZarGYQDXjpT2Qvm480+zYSKlUcNJI/PKxy94JsXu7HDwOM2kDZAoOENCabIs8dgvfM9UmhrlR
GXiWFgiiDSYtJgaCwnl89QTpSWXZ5N1Y3XSHeLW2ynm9gdhnkzukUDnOaALk0FmPyyrgUft63AeQ
k0TrTGPk1VYSzC6OxCM/s8Z25Illsygdstzr9LM1kGnSZPKTH00ngOg4zzZB636hwpVu9mxP1jm9
wejwWhWMRoHQEQTUHiC+sH74djXWJE7WhyePeKA4dTTID+YZJWat0X9X2H8KaNaxoF/8Z5tP+hHx
ToizbtlNnlM/dQtdq6KwfIZNrdjBg/CdS3DheJuq1gXab2LHQu3FR3h5HUh0Kxc9SSSx8fOyuXOL
ddyl7k+3z9OFulQFplM8VFkTUFJUTh6trdRRNRB6gWP2nk3NSsKSAgk4ojpmWY3CUNAY2KNOp5fg
lX7ea3KAHGICmWMk2WZ+FsrzwkKM5FWI1LGC+MYWYWvu32gJzMprABLtIfDsZW8auRlEQ94sI+3B
J47O2x2aphiGDoi3/J32dQpNDgTi6qGp7AXrFeotYqTJfWPiOhOCJsUNoggyKUtyClHeWeqNDg8U
vB+jnAlPaH2UmE86EMOD8BIy6DG1OvoBe1uigfXydbPncQMRMF41bg2w5cx9xrn8y+wjF8xvXaDQ
7K67y1OkA8P1YJtRaZ2u1iV8QL1h+Qxf5LZvMTSO4l8VN0qSVsTdX6hQz6E7tZQbjaWOOqGTAn3f
DQnR0pg/x9B+MJPXMNKJro+FahAbWSNjqvhCJ+NxAinmNUIcLnX2Fcr+Ew+4PwbarfxHL57uljs1
Fhez2gNh/K+DBQ1VJ7rgTGNICBEQ5JCHGnzlsN4eSY5J7Q8oXG8PJ/SEIw9NR2EH7mjSOWmQPect
K7R5qsq9HlVzHIFeF9+eaGzpmWrdMMP2fo1MPOicg+nZjkXahzdj0jJbGSr2uii12X1qiE92xSwS
I5VBQsoFw2neEnjKIT55Mjtass2pdZuom0BegfmB4fXnRqnb5HEa1+MmXnoZCOzRf/BBKynBuZp3
j4VpZGJ4dd6F+SXFsJNK11WozOjIjbdvav36YxXa06RVuu/fmhKSkEj5wpGwJxYy5TjE3SeUwtVF
0xT8buqTybj5G+8JoJ/fEbFuWyFUApdcEnneoZzU6HgYIPDRSkMARown+RI5cbzrCji2jrkpNhus
db8r2wwpqMlWJpkAJooxMSDmTAfUVjN40/+uw0RPiDq8xkvMrgXRTrcJArTT9EZBksbmndak0yXz
dSb0L5/mzg4HAw9JkLLz5VWdrdGD2UYB2XFnPdQ9jalu9lYCAnD3lXpvY2pgsptHh/6yhYsRnuYN
ysCtI3T9/bQCbI1wsh87CnF1FRaGfZ+OOEzGDsMBDq3THrQED2EcmugXVhLqODWFUgwES0pnbu0W
7npdhU6KsmBNy5v5veO2+XhnC24PWfS5QEdC+xY2C2E2uSiPPZYkutDjzDCOLEIE8miCqP8nFc6i
kntZOGNqcOXVw2zN1HtbW7mY7ObwYoBsGS2Wepp+2FBqRZ4sGhA/jxYXE315AlsxKHTLvBD6cAsZ
GJeyY/NKNbbACeeORhNxCe4M+FMkeJJZbYYQX8Q/WVZc9BNPNcJaNB8lAghMQQsh0i1eioBIigVJ
Hp7kmr+pMvO5Tj1sr1R4IsRh1aSJqZaIWDo2M1/aDEGBgPZOPPzvyosdLScTMfCLzUGFpAa7q1Rs
E6TCBcydCGl8TzsKEiIfBDIyDXhawxm3AZRlwNY+JmbDfkgvo5Dh8F/WKBg91B9cM6yxjyy/BmrE
b+fy08Kub9CnnD2seOxVn4Jyjkg/i6C4OgVN3BxKU/yv55dlEGzhp5vRXYfx8+UpuUaubgp7jMJT
rPo4OsC/PxkR0giEJoQ104pVGSAsujmCVQl2vuW9IXbzoRnRu0jb7BAe2YiLuRN5gvO4R/FpJrwy
w26NwKOhxffA92hl5blY41mrRuF05t7c0Qfw53M6R7QN8kzJmox44WVn8QLT3KvCAGPOrnEIVlK0
5ZNkEvDwuxq5czDxq9NgZEikR6q7+BZ+7HI4uYKxqpd9cqkESSqGXGtlM4ErqpENq7QWQ4tUunxV
yXIGgkpOcrFR+clSlDm2JDKeZHhVVeK4UOW9tUtB0XnliVuRc/o90vmdUi2CT804cKikt/G1IiQt
ur3bHjKm5ew9Ng3GZ4xIE41jPJlyqBPnDc+KcbPNU34c5QTZkTdOo++c+p9y16U2wLAkQ20PqAH5
kiSq+dZrHvON7yI0VAbhGne2gfdv/uHrquD8/1tgEdoT/wBRwEys7nojc7ENy89v1CT1WCyLcjad
lPr81FzHPRjS9cOb4PwGu/392a+A037/WHLqvVnGUie6pD0Hqs/UgPYI8VUEiZoDy/saQ81hM5TW
j8lvu6w+LpizOcrKA5RhsRs1Xxp1a5dnBBN4cyOJ+vb3wcsC39QTLh5jJS6Jd4iOU5CdcftWR9Di
iuo2WW47QacY1EXXQjr6idTWgEq7zbYyfTGHU0lyQAsJZ9QMQoWAxF8kzEFrbMYrAqxBAHEFrpl3
qiW8qcRYuGoAkoBk4FRFDvoQtEGJBhRp63rNxPRSLrq0uDn9p8BKIOKSWOfwqcgP0RUonBogezuR
kTUvrrvnPJJCqa79Bkba+eYB+H3PHSYPduxqyhcKgRZqQY0kSqxukhw9WGdMwYxXIUzI4FhlpUER
ew0L0IeMENqbC5L1XiWY8JwnkLIQHM8GP6T1afQ5kwAxFhbV/u5bLAOC648bwNYm5RLgKuMVSTbR
y+tFKR4GjwQ/2RSblP540odSH41o0tQhoPJ0KHWS2n+/mhAxE6ngr+OxhpNTtUoS9v7WZQOodazZ
QY3M7SL3w0ejOzxeVotVf1C014ZVs5dSgDd65az75bLJc5/zzPgtg8M+k+rFHmBn4a000+ZCyLb9
xhcMNDtMYqsHpX6T/8ZlkfJPTP5KLJcH+UQmwlcUFl3kgfZDF1WigYPcTUZZoPWMWqMe/+48XDTN
BGb03h2yCqnvfmhe9IQFYZUwogGFJuXUDOu8xyWeYPsz5mtmCecARG6Wmia/+9u1WDbgOXKSnfJN
xyn5yZG+ZSstSShNGINmyn45trV4XcrjmrhtUAEm89Em1rkU4Pj0AAH2Mpu3mzo1LBaMr4mkPD3z
yonJphIPkDSdG2aCKG+gaXH5/a6qiAFIUycW4kLPHzJKbnxeFXVXyWgWYvCnrPWmSNnupN+9qgwC
IJNq6abt0RPSueMnvxMsdNcB/Czt+GmHRguTP0GR/gveNe0IvaUZvriFIvbIXBFE0uF7RDcgn5fC
vLT9sAHzUhefQ18cz7tVD5BS34HafrimhDF8DsuhaCkPZO0KQPOKQ07JTdshwRy8UwrqBhDE9Uo4
lR3mka29+PmPMbgbxf+gakYnbBijhPib+kMvabbOaHMo1OG2KkcsJ+f7SuhEJPH+WDYGF+GbAfwJ
3pQYDHBFX3Vk8vz7j67g7/aB03Rzb37G1popY9Wc/wu0BQ3k2Cn1jU4SbANj3Vd3jGhUDJpA9wjG
XDreF3VJEiSumbF+VCCZt+Mwhqs63DDXSM4DgJD6CQUvKFY20qrVpaPnVLOZeZ4ZyCoy7S1DDS4v
0QXRIqbkn8BCJjCOYOi9Mev0I+N20lBm7XLyYIJ5ywJk1tBajk7nrgGHjBwgFxUoDN//hRS1Cjej
fw7g5cdHPREbOgzwglutiw08UcpJef4jPpYxPxFedqQc+wQtybxJ73ysiw8PGZTmZBcvc4KKnHTz
CmFobWLmxx+Edd2Likj4iZdenbeEQpTvNbtzr+pYZUYEVNYlraRNdTks5uP+gWV2dgZBkW2ToH7m
Ow5N0pIZil/7VKKJurqreVBy6TY7dh0fiR8Qp/5IeVP8mbRKftS/paT4Fex/+ZkvIPjY5/dZ80/b
YcIBy4nEzvteB+x9pSN3uCzFi9TaZG+qTai4yhhecqHdxWE8ylzMpfZkYvA7lXV4eJNtSpzukxQX
KWVKwgHP0Rq3Kac7tWCpv6dDWA2mFrLwSUJhJYYkSctveTcaIGHH5bA62DsMTy/z22++Vf7x2167
P3dN154jn8JY3jpjFOFLV9ZlVC8qdaP6QPYwzrvUI2LWXj6YubZRdmcvumyFfnSgtR4NVz69Prnx
ImODG7q2Wi5BUTQHxxjaYiHK2u34z3XAtwDPcqj7pnv2i7zdoA/soNUtYKrDx7pc1roRX1TJeJJ+
P4kJ5RxuzXIStEYs9tgVpO58Ft8XdDU92bYkpYftiEaq6dQMC6SM7SBsi8lVizfOfWqN9LN9ZfVm
3lcKNXyjK2aLnpJKTkjdC1/acqBqVLVW4zPfkLVNv8lASOy9llc+xiBM949lhbFgfdzfZXBoTmo7
jUThZw9a7IPJLuYdc39wxqxLDLHn8W6x9VbThyhTTR0GRSlVRTY+cL2iHSRTxqoDXW+Vjm0aM8rR
KllMIdHhbUd4NFxpsQJFqFnM1vjsOLdEVPC79G2/IPZPeNjEMEg9FiKGdQLL42sKAzN08lIrZ0Dc
Vwzyxzb959EHlVLRO4DoIq1o/CJb5B4bvChA2VoAuD/OP81j23PNzwfC397m4GK1ekHF4jCk5Mgh
zUrFWXx47IOzgCDzSudBk9tTRuSGPe8w60CRLJlkXJslITEwZpFldhKA24bCMhHkC5HcXDWESfUm
DbZGE1c6ox4grMbdabo6HuzaLFWoBKt0xICCTVPGnygjt/x+0XomRtUA4kdC0RilxcsTqjirtEbw
3mOTNHxbo9X1gpyhWbXKwxNkV9Tz1ggRPMid2/rnVm0nam7H+KZ79OY/G4J3hBp8cUUF4elnFx0i
ush3ooLgAcwRtMSg24UsTrMQmCMbrA6SUyW7MSqo6+YLFvgngLGX7EMUL8BBoSdB/XJsDAqmeKwj
Q+Pghd1zNAgzd7SGGx9+ibqp8oK1tJYVyjg4Y95JgLV0+UlZdmJ+wIcz4buGUvzN1JR2Vok1zxCF
AD+xBRbrWf2ZDkSpKhKFOX3LjJiz2TjrP8BNlUoDQSjiYzdaqcnAD47GSkLbN/9V0c5M49cOvLbX
2XroIafOMSsNXCCSoDAktISpGfDwcgFYXNKoNFMr++30FJM1NOD1GJaGzooGAy0KTI/qOvv8hQbx
+GWyMkcvejTO3Yb7Bv0L8oDrrT+2i3uolnowCkMSw9iXi8yfNM2OlnRh6MdghtRVNUHJmmCVC+/I
gizWvnwk4KLISjwsbMHYAQLT70Y1P1u2wFehaJ711K+JkZmNHQPboRWQf3pYadoXOYeTgc+g9R1S
crg3lLxRxgUgsljwvUVCuJ9mKIdwTaeLwWrEHIbLD+mOnrLng1AYEldogoYrjTFm7V+8GtsWRkYM
o3p/MMEggTAD8zvhvjfiDWR5BRIvcoC9pJUQjoFec9rDunez0FwU9syG5HHQEja+xKjBQmStbENg
58OQaLwEhKFkoD+1QPFJMzRk52IBubdCkdsLC3rdasT0et6PMuBmEDadAHAkyV7DW49zU/6/0UWt
OD8yHrqb/i1f0gDHzIMbFm4TX5ZpexrWc4A8tJ1wy3aA3xOtwlbNKTGYDYCVNYvFf884pu3DgZq0
mulSa6aMqCl+XDk+da02p0s32nzOlz4Th65U+LIgYHhkgOGJ+UKbMqdmwWcSs0pUrsGfjBPXwleI
BhM6y9aaBAp1FAF9l5flHvB/hl8nLz/KfQLKJxcZRSduGUMHy/wXwmaQEMYzW3DyhhyFLNIXT9v0
JUwU4oXdHmyCkUzee9CmyHYzajdW/Fqz9XsUnM5s5nLnoAxZedw/jDQAas5o/LirWoaFztExuN+m
zv5lwUeoub0H6PVme9WnPQURjhxUzG014yalNTIQwhjCqyZ/JwLiyU3Y1eY+Pa2Ts4troeD7kTgC
RcIJwfta48DH26lnMAFgB/1jjkf1HKuMOxrxdnrTwpCbbV2xiBMxmfPF3adQ9FlU4cBnbbTijmDn
pWlNGurZEBsJadcaWR/CUVCUVZGWNRao/zcMZMPM9HqoiWaSKmvcruqsecPdBPOf+XNPySASfvlD
vXhHGuJkN1kyBNpl9ihDX2d3UD/QfdcfNdVDVCZWogyVlOdTCT7xQxS3fJ4rh9FhDEUlXUFUceor
TQQ13x2CGfgbGoDpvGEAaiLV3Fb/atzsmC4PsvjFny/oAwtSUf3lhv5MRLYEeT9atObhjy+tRVIg
Ej+J3Sb7RDaAs+21CLRHLuUnE3I1d3bAZ6oUR4M6hGbbJ3W9owBd9kW5A5FxQeGdkOAUkcLuUkpJ
s8gmYbrqc/XYYO9CCg5wPUjvefNtW0fD/4DPB5gLGJheXGIJF3YLYMhEuYheR27AkHXfq65QPDUj
Of2qzv9bwrMjDI6DZiUkXn3uxFQsGMTrP7Rbo+shzjOuvDPmAwK9B+aMSXhannEsEP5Dm92NzJhx
lvKMJwoVkxvdQjSPwgqy2/1fwQs/tK9vGSr/67O82KinhouR6yLzR5LvApviYSXU55PQWucnpmcJ
lSPmXioPK5y54g6DitRdGHh4SPP4NjMf3CXOscKQkR2Y7FJEArmPwds32w2XagHW5/x+2wx94xsi
BLIbezLVY6azBAc1sKMJPAx0se2h0y2900Y3N+pFoKr3WYnxdKHulKuBd+GPmQ3wjd1UleExhm3B
Gd/jrLjfKAuXbIir2f5u2y8p52map9V+cZk+NdR44xWnOk6lLKFnNO9XOFxrxnwmnsnL7Dr6sNdH
STZ29DFpNmhkihycZwHk/yYeBf/4d5KTR638m8Fly/vBOJydSi4rYTQshuWDC0+SgPt6iMTpai8L
SBBEtE43P1KB9r8S2IuNrahjnTHMh9wZrtSqLmEG3LIWnGTOFBhcyAA4Pxvpf1rCBodPdpRe7np/
sjaXmWaeLuaDWVnuoePHIEZORH74h7GZuWivlj41Bc3vb6I7tkbMu5EF1MVe+97/XL83aM/x/Mrf
ircFowI9ES0Y5kVYplachB2YiJSOSmLeJgea9QK5uo78TPf6Dojp1uF+9b0brsZ0fRybH1n52XRM
EdOLFJetqTTljgZA1X9T+LprboL7ZXOpZZdgM68H0o9hvw2+XWvE29czyjOT9kpbugegYu73Wepn
MBiTJpl19rGAp9GXL3X3Q2KoKzth/srMP+UYgHe7fxHuoZS2O5YcpX7l27ENKh2iYcpTXD9qQrZW
dXEyULRDcITyumvTUa+6i8FgWyO3k3Fl3Xx9LSMzNDKw9VaxfIMQiJGfleyZNiBQTQ6aAB69Ki05
i9Z2gilH3ds3EWzfBVOzaXBqgmH3DcWcCWFtWgNwZhNXKfho+caGW3BqjFA+mRkqAQfncLJgrc/K
bjIiNjPYAlI+ep4ZOyeA60sYqKThXEGZBbMCJ3P9QmRpiVv4blujH35kB+UENY0HsNOzNAiN37BS
cPktU0av/Brx9DFoMNS+c5+HR3cK45a9I4S9wwOq9NlPhLT+jqAiv40aGOpTNGdNKQc+4HGUMpxP
rcfL8THh5DN0hJONKNJWC3TavXz7/TTRDPiEKAK2437bpQArM15gD+dMKU8gKZrgzOYmGF3vOWkA
WhpVgeNpAYQkitCH2YVvyCdLpTjKKDN1tIpXSgIwcn1Z8M94zt7YNaWC4TjLdDOoFLzl7KPzpHZG
Be/ykKb3Mng4oiUn4S15cpAC8MGDFReY/FxZLk9x5egp3LcJuYxlKCqd1egu/WF4gKV8NabDbdKI
At1X0ZPYENZU1EHpJ7LmqKYYG4mZXzZSBLX6PFPZfg5zREUMVKQhMS7Y8khyoOY9MLvj31/KxMGO
VNP/1BpVce4PbH30KoQ/MjvYNnG+h1UwhQ1WKi1h682Hh8ooj6wzmeJAeBO451faCVqZnvX4vxWA
c+XIMY4VxgWYU/ikLQyi7dUvS/IN9eWxcheed4WIssKoxwgyyFirrlzjJVrfDw5VI9Vnu37F0BNL
6MShyZYMWvrt6Gh0ZUf7n6+qimvWntmi8MXe0p7nw4SCUFCduMDMXaKGc18YYruB+Q9sajtNIxqL
tkK5lGDguVmy3RLlPhcK+towNdq5cz2fjJHVt2GvmqwOGn32Kc/68ap8cqBOC3ndAeILM7frizdI
YYtkqeR8kY5V0SsgJIiNsi/zlM0QFLuaHHu/k6kFhXCq9GVb/EZQb7gvP5PWHfdZ3QcpwGYtUpCV
tzochci0wInAVfgk0QWYlkfm6yj652WwHPvd0m707p1PJ2JCCD1uG64e/Ci8Xq3gbRRsRrPUmy/A
tM8wG2u25JukMM825fo0fdsAhx0O5g+oQsrH0cZ83qNfQgrDXvAd6Ssfo5r8MF0mWQVrNviTt+WV
vi/JElTdwrxsWl3Y+Fl0tfzBjBbKy6VLNpFX9jz2N7hC/6isuSk6Nt5SGtQY45T8oBoJn5UzI1Rl
fQSfh6hMWnCjgHaE6SulZZYjd3teWuIXj1qOb3EqLqyIVSmDbWd0wvrdt73+Dh9lyVJhXaafYUkq
CsNl/8gxVffcCk35gE3cU0zgfQr0achzfi+xy2vE8viOXJ7xgYZsXvATksp07wn/TJ4byqfpWJ6L
xo20pe3LfK78/MvfnVzaRjID0wYVvlhn7DDvdH81ccTIazEXq0VDONV/QfIJesFyGjsTm62oThHd
47HQxhC4vSjiXnMO/tc2qR61OVPa97L4xy8wIF8rWG4kFYjx78MTIDI9b+H3ua2VYQmiwC0a+tZc
qqEun83IWqq1q9RemgsZmzLUNY0VyxsDJrOmMEPU8Jz0Gbbxgbd7vkBaE56qXizzEO7y3Y089ipW
69yV2WgUEDRefzOF90sbcMjdgmK0ivNhOdsoHTmp3O+4vRMbMyirWWYiNdqOUGl5sfvDsEwTREmH
U2OxOpmXFjqJ5yU1AnA1fdKZiRmVg44FdwLKb/qrDUG97fkB66hlcnv2NrH70hVjv8VtD7GYELFj
/BFeX8VQ9siSrXO7MP8SaqxWoJ6M+/VLVxFwkdCGFvrAXT2y4PQNBfwccguFu8rQQlG5npF1kB8M
+rvvY6MquD5QBERu1dDmmhDuHd/CQA5MJe3l+o8gwBwPRbVgE32iJDPbqQTOIttC/9MLRqK4c3jt
CJdwy9aQkeUYvTK4AYezdF2jcyjMJiHqq+eHNTcWs8wK+buGzhitVvpa18cDKfUz6VWHaCvPBiZD
YAcKE+Vm9LDcsGLAZ2fD9a95+daR4EEUgbSf+KrEtEiPkgAlCmUa92b42BoaKB9qov6GHMBkiKS4
6BFKcXFB8qN33PJ1Br+hFgU8OcvWDuYIYpTP2N8weVXItEAJdMZZHCBSwBOI3XTyMnEbOP03STlE
2Q5AygOpjA7ewnw0ckeDYXLPztsZQK+6pOsspQJuMzC5VO4v4I3UJv+Bw/nWYOr2Q74j/XJ3Ql5d
joqsvB4vt+OH+MnENXtX6ZkSA0REgI078bBuLvuSXoTHxn4zHsJaTfvJ7B6jM4f1ARvOjxYwbHe6
CYfZrBXnD2/DJh6IvBQnS6y4d5t49M5d1N9EWu6KCkMJRC8QJcBspi90QMwzNTdki3d62jk5N+dO
KEvDeiWbl0QCldZEaoDRYLSFJB8dAQUGsa414t+Wh+c/r/l1NIX4RrUCj0cMzpK/Kany2QSj+Iuc
fIlsjDxsTcb6WpJA7pVMhPRKJFkGK2MbWAccWc5a9DIvIFpQvPJC8SU9ELUmsbApwR512DXyQTZa
jvLN1JxJrRCXt7XDOI7gEmlJQyL4K5WtxDaoDalbrM8aNZYN8CyxOeZ+ir0WQN58LT8OQAR1ITdM
uX3Q8f+KLAzr3L2rs1GknxgPM1uz0jr3RZHHC3TNLQ+y9xVMoe/LGycDltzfz0jIjvBaI6u0+Oqv
Bzam25JJFghtMV8k+vUjI4NeWmpWPR24GcATRm8Zsrwpy0hp1POkIqMMHJu70k3ITplPXN/GNOEd
t6AXRrEk4rv8yaWdZ9F6Jqz4hUQB4mqnHkKUcdPTrkoxkGl88d0tGzLmCMJAJs5YrYwMTZg6OXer
syDqj2kFoNEVIZ0nDaX+z9JGRvYVfzUr9Tlv+CnjqgtZpXjEMaFFY03U7Mwip3oIPIkFPsCPufoB
KeM9h35eFu7yXSzxcAmsT8SSQvRlnpQKVvE+goY4LL4waE/iCnej96i6gM9AmtPy7YgQflwCKcM2
cFRpnBuMxqVY3YlFCI7VZAxKozYcu+ZlqUsBFyWR6zOQI1ZZnDKcZ7GxzIU+hwEURNAIh18n8ySN
zQFFHc6cK6kZ+7ThQyldMsi9xoOJSSsVn9NNFziyf6tSL5T09BccgTC6go0LoCkkUbEq+oNGXq9G
PzOQPG3pSlLmugALgsnWKt2Zg9VrP/acK8VYwRYc8PBpBwMK/Fxq53nWN8IaH4ZrbfYK8rtIPZdI
n3uGz2oXcEHjAQm2hHGVss1D2py5m//byrAC3gaSzHl9dsEe3whrWOYCmVUgqSdtPvj4hvz9xMB4
9n6L2m81On1WGRRi0OqW8R3AE14DsSGatvN1TUX5xVt5d03HVDt/3LWn5YS4d35hi49M2JV4qc7j
KWqdLnROS7YgtZ8Un7QaZ0JacluKd5vrgN6PlYYOhpUBLN6x7VR4dcQiC1ACNz7ekotq96lxh1nP
qBkK+XM/sPLmSwcxsNTFCMCQLmB0TZK+JI8KgNw3/K/8UoWEXg6Kct9GoPVt6hCFdqR9zVX0QEJ+
rIhtyrN7aP7OifkopyfpBRVt9p7LMembcaUPsVYEvN1qpuaHPkUswlol4JT21+ALw3l7jOen39ZW
LckjpnJs2grQyQ9tGs5NdMqMxuxbB6BQ0JT8WGgOjK7gxATe+kBucKkgfMuPk4aWGV2MFOTP4auh
Maz5ecOrw/BFVhkwGTIO9D8Qy9FlXLfCcKrxUBnAyXM4pVkAFzMLGwL5fhBOprgZZh0YxQ0Y6DxT
qQC9VbpJpnnVCpZrsKylNSf+C9G/Jnye/1ifUvvVXr34fs2p9fcUYVaDGlS2U+boEX0ud4gBle5z
f/+cao0Y9mX/XwJSGJDC84XuaoN9lcfbxq/thxTjIPuN93c3cF6bJpSmevHovEXWhl+KUAHDlpCV
tg4aP8lPVeika/+37ksHZ/cmRu0H3TxcJRKSi1G2HbesylP9c+1VCSuJ0xSgEZYWvJQutnlaj0t2
cAiyKzrZokyfPCEH6Dy+jMSGUPjeg8ly5wBrD/03PyKZoBANzQ1lfPvALfJUpYtfXA0EXkHcWB+E
oqayVjlAl1ZLnLCW4mtD4bKrSrnBq203DYnKOwNF5NwDvOTDgFybB4ISTvqb1Lg3KH8zcuRgUrqL
zvBw0j5K37bgGV1yDEWc3j6kqVDeySm1GYyoUGdACtuBSQtdD8y3Y2U09CCUnnvQfxWv9rq1AHbM
iz0HlixnhUXghFOVzXr8W/y/mQj4ju7AuJaEoyfiDvuV/7dnWbgQMtvPN69FZuulguAgIwDwbe/+
Md7C+hILiQhDxJFVPySZRAZnK6Sl0F1dxCCFJbdXlWWRLI0NcJip0Zz7OOhuE3lKv2ly7OVh++Zr
N+vHSidqCpkjspMojBGJWv4Jt7mi+Ffxn+copDapSwT04pUM/b0sTyg+PJeLUyfnqz8+oj4DXaUl
Ff+Y4CuNFeBBvRNcJfN03qSHAD95eaB2KGTK7JFuWQh6LjM8/ZmPRRw1YEDrc0KQGfhcn8YEW67U
+zCVxNWzxKI3qn87at7oYe5nPQ/flHy90ZE3SP2RJTXHRPkzbUy5oewbClT6O0p8lezpP7qx/pGG
9ZF47dA4r7NEx217FCkoFPnI/WnnnZK/vdmz2m8FlSMVrCD0CSADMqDSUQ4DwmMsVnovLBctqyng
LhSiyJFw8gtp3qs/aevoBoSTai5iHdcZQzvLPYQE+p+hvjic0AtOfnX7X+sLCHF3SjmsdZQRoSGG
PaP7OV5cWqLajd6Z1wMZGj0utlpib9I9YU9rJaYS2A6hE5j9FnVuQt8OQCnia6sjqHQl68lLPZ9c
+Z8XqTPayjxWiPxBSNBS3sbYm2RchIvIMrq3AFXXwsh9crcciyJaVIt5BwK2NQ+xXhrz2ev/VQ9n
G7TFjDoau3mR/FPNiZb8Sm7MIYO4XyF8zC1dGdXEAzQ6IHq8ug/6DrTieRRUuAD4ZsSMxb9UFFGh
sgtiQPeUDJGHTi7pizZeeOpSF3c9AqV8x1EckFomh+fKd0pi9+uILfaPaZSlvq7R/S6tIZHB+8Pv
k4Fn3qLnIxNtTsxabV9joqDYfnm5prihiLOCRqBfN/x2XC7ToJeazqJFimp6yHCDeRCevd4mV99V
41DlQ4VobU1nnQ4cXqIpvHKX8rG1g9A0YOu9vpdxxtcDpKKM26Q3ORivlI2qFQSCESy5Olez4MS1
psQ1DgKBSshBkS6i2xIwVL2dgEhqDf5/GXislrGFLFKe2YvHhhnQIa+B1xOfs2izViwRat0+VSG3
rN6vA3a4LBMgkVgh0azGyOMbzzLEukJFFNsgmhDRUHfelgbsA3nVwnPlVMfPsgFFs6fyN+fO4NRo
uk0xVUvHVyAsGRxGAGSdWVF14ZK0DsAiAJnu/jTF7eTH6QJv8OuIskbdw0Uxc+QNMGRmyLKwldiK
2kQc59XgXxMubLz5LLhoYJIXrnJuWeq57bnpbXzIrTOV5YuHsMqokobdChJsyKb8vLEUB5yuhNDo
+GPHOjZ+KWJ6Pj/wvlfkhWrccgbDH6xDXRkmHCSZ4OwAKecyRO0x21KquPRyNfTbV6CYC+nWvdM8
DLY+JHnJ3ofAdyFZNbYPuFylodwhGruG/l/w1pf6uzboG+kOe3uex+JLbCKPrNQuFB9gADSeR9Xg
c6I28/aqj8c6cXSC4NOPfcMorxdYeyE+AQc/QwWBwI+MvGTxeYCT+cr5XSV6gE7qFuALY4R4ipCt
g8pyCIQ4cyfD5DtCTjJI+2kO09i4/gynJIpvhLUSO+PFUUz9UW619YWwzO1ERs6EcosY3AS/xm25
4Xucgn5rMWvcwvXiWzZbWzyzCHGIJmxUFfeNVuieeC/MIYIWP/KiMFm4gJKNNwcLaxqZSVPiu4NK
yUlLCXKnSbEctLTUg5Ci56k1kqlLczWzTPKuwBkDshfexBgi2/DhRTJ5ilitbQa10KI5ZkN0x3N/
tq/xhyy8nw1QfbUfLVmnT9RPO49u+25A0l/TtwSVOwzzjOkMZvgXkD9Wmx4u3iK+guufAB+lvwpe
yIl8VB+3GCB+wvZBmb6WpMVKWGMoMUaOmgkm5jjqN7iZZFPLEVSgCbDcDZVrLHGW6smD1cqCmETy
n5et9RiIy+3FLaK2X6/MShmv9k4LNp6Jq5rjA/IfUriYjmAd+jmCAWeA06nxXgeH0Y2SZBsYhfIt
9T5wao65r2RyX4ufBRWLU+fqZ5P8gEvL6rKod8opHRg/q0tn5nsDelIAH9Mz8OHjcXiOWiLomQal
u6Cui83KQEj8IuWMliBJj37ElCJjin4BYQzqUrXqgFRdEu0Qk74heijP8SxW9/UbwYfV2aTDLGXr
9bez5GFNz3CsRdUdDPHTG3lcfzbSJhjFGtyefbT+e5xclipQKEk8H9BQlWB0ybxMdS/M2Xe6iybr
5jF+XO559xtITnBu+CsdPt9FdR/dYr3aRNC/EGv/AXLUJequ59dbz9u/3C6Ok1ZS07MfM/0/5xDY
CkwxlNBTyFzT4Qoa0cOrk0dr5BCjnDJsUUMTrtXMwkojOrn00kU+0aklTriHJXzIBVm+WjvH1F6K
FMTAHMxYMLLA67iVRf08q7jLsTSvHBdwVyimnrTEOXEjKXwD+anDtIqXLVqDZ6cxhe6YlHcbwDVN
x5qyPPbtZQ7+UrRTlm5YzyU4jwwFTB2bH6GEgDFnnR7apYYCLMahkQtZNbEjcjgdNJG15lRTrUBy
aD/GdwzGtrAP+0zSyV31/bEvwAla7RikQIXewo4Kxm2RyQB2E4GpZfgsQg9b7HpieUJBwnTKzZbY
d5CnW3dMfmDyrBTUmn/1Tmorz7OQOTtHJUY2phGjkAR0U6l/yx21NEP9xf96jkX5o30V6QOu5Cg5
XU5l9+XY2UnQIvVFBye/ZUXopVmTZn8ywQOaS4cKePok52e7p/GcKiLxakppdCo3JhPTI6MP21qX
pZpDlNoy7qWhVGPXtAROngwDZ1wGtZENJ4YjZ/tb+1n9N+S+ZwMSGcE/4l3PjmVMowOdfxEiaLil
i3CRwfgbbJdWKjFz32y16g5rAAM+X1w0wjvzAQMINGhSKcrOeJtGn8RUpVIuTqqpyQQXzDAjnfo1
XX2+9DNcqsSlAfkkGseFYz3TCTblgaB4hwMz/1UOSBwVTQlhE3dX4rU3AXhG90KhpIDjHT3eMBsJ
fal12ISE48s8eo8/2jVMc8fiDlllMXfcwAo96tkVEG1d33JDC1P+FWvDS+V7FVsSfZ4Mga2Ega1V
uwOO7zW+P7pnYzmbdN5CeVqbb7zzT5LbhtDXDHbWpx9Sld9cs980dJzk3iJMQwwsviccpqB1oGAf
LqNAhjTgX5UbmVbduL6mfnPHBh9f9RL4rPCfq+nXn8bq0rj1ISjvgaYdPmbm8rMfvtkcXbSwVn04
572xK67IT5vtGdkySWzwed3b+Gt0a+gC9RcqZVTnTorMvG+HslXlEjlgYatBSBvXmzbxNglJ+rV/
zD0LLEhyYbxx0oXpccinTqxuS3VMGGtcSRVNbJWkwckytpzTlX1MUE0ZaBZ6ler5tlbgGBdaXYwF
BWryySQAUDGyphdfes04VlDelNEsttr2gtwPzjMSHdL+i7fzDaBY/VUeHh9N90E06eMneBBba/9J
Uq0aKXO05cS2YL1c2IYms89hIvstHmoLKjkzfKkAVayPzihUoSyjOhwSy6slvt2mmA5+4+Gtk9Nk
JKBV3koaK8nCVT4J3hHO8w4rmydMh8eWhVqAH398MSIVAxeENaor+pSArFW0BCiqU8aRW/cFFjxL
Ly3lO8rwlmfS9nRLkpAZZOO1w9gvywrzaGGTPpByisZM+EaJucVm4xkJSkozGgTdMq/sqnl+MBTq
5M4euTDmpGCDRrK7GOfZIHeZejc80M6S5zfuhAImIjX+Adsn1pfT4LDJ6ddiiEmtQod5wwOxGdos
2Nt6QCyeWIUNwumRDKcGK8gbb7opRWdVk/sUZnmYIes/QQx1870A+3v55tBm7Yu7P6GXKyHsgIDz
gmgABAnNUo5LiXmXhnorOqHv9kY8yZuIiJA6IgYlJ5+Tfu4xqUA5B2anJL2HA8VIp/4u7/eBPmQy
fNqO90OVHFKLfV3DpdHsAeqkcK7JoLXJ9FNnXa8IsgGHD7DlhUaKetcDD0KfLSAVQvvPb+CKXRxC
gGWakSLog/0ihNNNrVqBtxjg7Etr38fDTrjIkfIvBMEAawzN9DDnn+IwC2NxU4bQazo5v3zEnNIJ
BzqX6NBWweqD3WyJQNLMfnqk3d8hZv1PLG+y5ufCYL87LuUUHye41cGiVUBRrcFxK2wXcTpGILEV
k4qQwkQOUYyNzlCIZkU10vZbgXz606ZEe/962jIvCuBmO1q/UyRrDRpRKQ4yioU6Hn/YrKLN/PD1
ITCNfLCaxV8hKix0+wk3zDDdEXhXpRWXiuuvGGtoNnygVsLlmmNy2iFaYVkcXefEW14/+uTEGGQx
mZecSrF1I0NKm7yRRQgsSRNFxg+kZW55V7kSIqNCdShrRgI+vZZz+IaFbqtBzVHcitCFmB74Yi5N
KeX93ZaIZrZ801gWWH6cerMekdIMd9hlLXmj2azm/6DFjIiScnQ7S6Soz48caL2daAxjCHeaYS53
P92FTkM6AJ1hzFIL3yPVYfT7PwwB1lpQd+nHO+VgrzuHanpv7Sav5jvkUQOXjalJs3ZxyRl03Kta
RoecrVlorHA8gTxsEHj6tYRBvGjFIOQBgg2QDfnnaVijEsczwxhDHhtmM1le2qM51IEjyrHH3wIH
6Z14xhP7ZisLwxnPKBp3YAAm9O0CO/3xP/X5TtN88B5uC2cwE7Drg2LNsdh9VyXN1DhVdhUpKJDb
8t+GvpvrXTwEAUGqboulyvVcV9UzL+GD5E08IIGXDn7EA33wcvre7A7WouCutlcWcOOpqV6XEMz5
kDTJFEGvXtNjwxJxkTUkUv5pSoMG1ezjAWDi/Ls/JaNa90ySRk2JDS4Lxf9trqyS82zCnB1NNTwy
0pXC9OBbv7pgP8/fqhmMxtclccv/+PeJANhzIwGyd0DoiYIdYaFK7qVEYboaKPP+kpXCIvIbuUzx
MvU6vJmQXP+GvbFX/KVScMOs+3XYjBd22dg2R9LEzio7D/hfy9PiWL2yP0sDcVru0vHuJ0a/iKKA
L2g6hCbVLpB/ZvWTlolJn/26eZtFzP1XqdgFrqloyTXqDaK+wZsrr3999LkNoLOXhi2EAjBSkvhB
OLznVSsLurVhNjxUr7ZTlZglo6seT4T1szb1i5ZzwY0Lv/25xEf81SSm53G4SpvHJXtINYhYZb4c
ALqSDb3eo2Kyi/WikuAOJHLlUkI9UJC5mpAxV1BpXR2l8BJqOU7MBspb4PwwL0itOsjFYIyVaHuZ
zz8BKnyrLJpBaG2KAO45XgFIg3Qb52cf0+gAqT8H9p18sszJ9IDUz+3F4oJVcw1ilGy7cpTFce/V
axAedISx1Iu1MRJcJPqEsmaA9LNfYlEW/hUBYdthJmmgHm0wtgovXPzKVS8DZDsifazqS+I0wAEw
AZvLWIR5ZBBY60/Ae9eCXWiFZS6Bsp/RcQ2gtwjePmNMQc4xzGGox3bi4HJbfdh8k8gehAcUzFXU
iAYnt7stsMeNOriLLgQi2dgXcc3ZIiN2VCkVOiwoHCLr9YAu6JAvvp1hVvnf03UC0h6RH+FA7wr5
dHFJDiMTUHARDwIa8LuBdON1U+NsoZIraJXiCFA/3KIgdNZ+0XRTQHwzKy1FnB2VhC+ztPfr0cI/
ZTUc1MP8y39bTcKv5PoARl1p19X1yNsyVNVr09KQxHnQQEN4EYdxkLqg8e21zt7ptxiJ4d45fZ7G
daKO/fSWfGYemuFwybf22Xa370smbby2iO+xMD0VCIEqQYmbDmw05GJrIjpE+QreBo1/2nylZLZC
qQq9PZtmozkoLtC15Z17StIa0skkyKNbUYb4ATbYddJtYbD1FyWGXzfK1GXaorkllF769Q6cjBB6
IInDw9j/RxGgB9j7rmp63k8Xsv946ix35rYtrMv3nyBlYnBsef0Iw/kmoBcSPJSw2ScTLpmbio5/
ij+wX8vBDduq1MCunpSw1oa0ycy5P3oMcnxjDoy8f8TSRE5XOBmZ+S7NoM3+nnIOARYIWKxzDsgu
fipCThHDM9LMSXFW4yVAQgcFwilITCFe11gilwURjnS8TDTlMQUvt3esJTmsB9cK5dFAob93Wjte
ugqLO1ygoTl7Txhlh/nNedDJaP+ccEuNhDMIbPHDw3Cm2G8ry8gaJAfToY6WhmxvaI+qcY36PgNZ
tpC7o++RXzRJ1xCqLitwmKHY1S93rqiNdmehoH+2EssrVCIKsUcIlt6+u81EXztmR7Ou18ksN6zZ
hOjmBm1Oc6m672qnIgR+qiWjFU+T7fpUak+3oXNeSxVbsjmOHKa9CJVeFgy/yTc8Y8n7ZdRuhN6M
JdNH8Op0Zouf1n5WlrSfQKhEJ5HgQ/pxvrhgOBzZfYA8q6gcgx3EuCWgRrDN0m1PlGNhu63JBzFx
xqY8i5nFzHZlbah1Jchbf2RNMQ5xfhrIQ92dTw1HlEZ+rqksk/nw1sLVKpp1IpMHZ9Zv1DDblEdu
pRVBmdWegdSBtf9iwn325VJGogsJHxprmgWo6jXs8mk6kj3yoDYL0dsQkOfhdyZXbftUa0/LSQAl
YiXdF/53wBImppuxdjyutktRX0ktIg3fXx718zt3NNyi2zU6/0LVIPkTI2XWTMWzGdYUnCaAIDDu
VL2lyTn9evUxwtOa+wEiYtZ6I9pgyJXM1t860+0xYpxSXpHyreEDRDzHpqEZ5vUYdG9dlQkmzhCv
kp4e2mM9R08k5X1IGpyPhkyTFPg6cR66ukIlQW3kmBqH0nba4TqIfB0C0eig4w+uYSWFP48g3O/M
bdIRRijO68dFpNal2r0Oa5S/AYF+cS9H+9WheoEzCKAARiiM8xtfMY5196Ek9tAhO2Khs2IZQ9YQ
Ob0UbIbBTnxY80+lc82KWz1Rp2rTGQLXRe4ngh4dDCFgtwEevAaK0kZ5s35uWdrEbmZ1zMKmI9Hc
v/nIpoLIv/3TWkg+Cxe6/6c+UVWyy5oQlPtkJZjr3zfWzzDt5aMlcYRxR5v9BZiGT1R8/5XrPDHm
DXbZDvhpdA0sBort3UIY9sF4HMALKukeHn1FGOY2Hkih1SwyQNyekvY3ZPQGBjj3rCasMLnkxNPY
eaYy3PMsbO8jyihnU9Sxwn9C0SJ6WSCwJJ3BWkm+5kwWRihT9zn7p+7gJBXZHmjMqnxw+l04mxbo
nC9ZzuYOLla2Rd+bof80vYf8fhJYoKhx0mXEqnCIWeFTTBZKvc5KQM7TJCptkp+CVfEUNMi/1ul2
E5f8VsqspXS9Ffg/JwODUgueWjjZQPcgB/1E5M1sFdQOwp+gegDWzhjkE77boDz+J9SwhXAlmGx+
5/vF/86W58Big2+OB5tz8orRPKb938lhEiZpOOvQQZSh1Xhfw05d28AJzxQ/hQZLqTLxst5jfb4A
+0baXVbM2SBIhO8z3phI1JHeOKcVkqOl9hwQ9JlyBgaq62lMkojokYJH6pl5IB/JijPlo8z03RwQ
pUpOJpOf8cfrBSVyJSzIv4rcoWU7ihgUTG0c23fxuHJYdSE14oP7Hu1ncOPnhgMP5tPfIfrMM5Hr
XhaiM4wtlSFoBtb7CX91f77iluh9vq4b9203wkQexs71Xvk0gd9bgefiwkh8SpbehcTmDjUGI9jA
yo96oBnm+xSLm66fnU6BIwWqCFnU7mFAP9HOZ0717wLS3u8KFAVZGl5VWgTnJfxM4cZi+KcVazmh
ajR19feTBzxe01SUUND5iLxBgA3kTiFLpedf7/NwftCWjtZpoV7vsQBPoh8NQN7zqRl8jdDLbY6E
tnNYPzsr7K42lac+u01CcivObX9dILIgj0UcXocVIh0bWRQYmHysUMBSLZBLyR/jxEZMA1y0JAc4
HHIKRsHWLn6cKIn9d7UgLDc6v2msY+88nEmxD1PJR5qxgv0mMhgse7hDtslrJ1faXXscwxzCP79Y
3Rs8+r4ZNkvgLFP0NtayK/ynAYnPlvSekGtZOQUKcTySgfzsqnh6wmjbE9rC6Ul7JnjXvXSA2sAj
YNzK/obuuPCg7WEZ9Fn8JP4itNx35451lwh27Hh7da8K7L5Gp4u2cGZDtEISRLX0EDUkPLogrESO
p4yy5ubFn6/KetbGsOmh8oVybU/I19JTNBxam8J+SJTa1cNr2TytIuNELUdWD4ORezVOsU3PMDIV
O3Ak5wWy3pQA6ew3zolvYbo+sh6AxGmbvef4g4GhYiV3dGr3H1lLcWlCI5obqFuPIUuRwKGOABvc
83z/hVm67UIl31mA2NDCX26WHXeZM0k8K+n3UCwvZZ9GpafnjlZOLCzzAn0v5E200/+2rmYcVNsM
wHrEbPv7KntPJrYcxgTqe/Q8eV52JcDtg1cAvCk/a2ESf8vRSU8HrlaEyViNZXEgF0KYT9eX9Bdv
zD9RQGfp+ItQa6hV65i+cB/GYDhlz47HW4pdDGieotUgztvdto/XVoLQn5dCQFXqXjnDVzQtM4MQ
MubRq2IohlczTaNG1ZIQ9WJcavFWfMl2LAnpPDNgCiSO0mjcOeMGWYy0wVy+uLOCzOOP+gfKVmjk
Ypn5SxIJbtEHwOkMKmQwiOO4lX46jUwC5CZPjFGIbo/SR/oLbcPjmJjQJnaZ20GM+zQMUwdoSxVQ
lKHUirMo8uDv+UshnZkd8zsY3FzNv4WNTDgssWMrInSItfTehLDNOqAvFMTrJmM+xdknoMNGTE8G
9fsg8vmUTqXhmYeIcLdMBTAN/fWz7Y8bq9L1iYq7X4zpR4R3F77qilQpQipp18lK/iSj4dTS9Esl
dYgTeHuv5c+jGbzFOQCSTVI5g4MtFknCYQWbC8Zx8Hj4B9mSbja8W2kJaINTQ2JH16BlARlsgFei
j5yo9BRamTh6RwN7lBBuPsAR3w+FWOC7vrtL564jboRp1gXEJ/NLEBn98lPNZHWBKwMCBanT0oTp
8WRfDCO2Sluxo+BEu1tv+gvOixvQyDtr8hxrO1ettmSfoRVIqPY/q0jIB8pyEXrwyLNQtpOJxKvF
B8PFIJj3xRuuS4EUXNhGVMSUhRYf/esIFb/mTJIKplvhSdqqJPSkpJOWS1p/UUa4tqdEisF0mxmx
GUYx/abCrFFm3iABE6Y77ase0KNyr30R7oPjq3Xqm16FEKAX1XhQKxAaDanUeBvTglXl/oWkmt6e
sZheVvYtPMKarIrRO/wmULg+a59wwbipDC+rkxsSpOzzwFQaFFm7rNN/fzt8B4f9xmyEkNgRgR/8
55w4Qjk2NEz/m94ywj7BYMeU20H03dsNq+DHsoGAP/oTdOhlpfD4VWtN2Yr1t/JZOOJ5nkh+0ts+
W53vCDYBFVC5n3XrHWazdjshX80xp0YxvNPzmKTSdW1ksoeXITrm4RPRdUpGLCC3HTyatLDhVZAm
7IZpkN1M3jcVR3BGmtvFbXdpwkoYiJ+/G9hK5Hw08Pvp4UPlX/Wxwkssc+TRgSyOhgiRp8imZJzb
9YpRspEZAAxP1cvOBYlfPp1YjvpfWD/qiPsBO49qeBUfNG4s5lyQloaKyI6wDmCpM2avAYKXA57b
Wm52w0nQbj0Lq8iKJdcfo57ZBQxAM9Z94mikkA76Ckw9cAWDWn4N+8mgGZz9+OE4qACjZtrBxx/L
ByQrEb4Q35Rrj2cdRdNoBfpXJ98N0Hbeoi9h2J+q0G6gSU/Qe/scTqo+Wej4Ptzv8SBRmE80FHJU
Cvlbto7xtE9yX3Su7DuFy1jbHJy8hreC5DkrkSCGF68VAT52GaiehbfWbt9egtmrhnY3BYQj/YxB
9NqCOKv1Nw0ogJMSHH6md/a2Q9p7ay8RXvXqmk+sEsflFOCubo2DhQ8n42LQL/y9ktDDZbb2vlI6
WUIpO96Cw1PozCC+bfi6CVLPuDUI8F40v8NPN8yJV5wy52Sn5MhfM8a3wM7t/xNqDSQJgyD76jJq
fAWhRjVH/jFGseeuWzilQhv/R1kELeNhcdA76K0l+Ao5XckDZU7VcAZRjLp47KEXHmkYhaQZmSE8
xHlKxPdQyoXX3BAsilnm5QbzVrZ/NbD2D+YeJWvimhxEgPixGiG/hLa3Sx5lCMkNOgt/KXlDm78e
tpORBfIAQ8nuplCyW1QeS5hECbcU2lyFLI5pOnU1pTVOMp/P/004yF9l9ZQULFTUEgHlsLGvCzgZ
3O/XcudbZAV1bRYknk7PzkJtp4xsH9kQG8yeY6gfiWSXyAAhYrJDufMjit5Y6kVtlGdQLRit5PGv
/KT4m2WKpPRvKjWgzC189fc3Trktd7gI6QGJUVEMdYqXeTr/0lJoDoI8hiFp9xzxV21qIBG+jNZI
v6D9oj0mBzNu0byfFk3AbRcwV20K+2n2BsqiWllOBy/egymTQgOUnvZ9wo/VrJx60EbPdijU26a1
ODtX0hjjkCu4lUGaNB2szczviQ5RLmV/GxWMMZ3Dp8joj0bgpVmriMjyJVLFKuwewtCELiZUwz1b
qYVCUrqc7q/PjWuFDmGNx7EUnKK2MsJ7WUa9mOx1/X4Tu3iFdbvZfTrnlZBt/DtTL8Iuzyje/YUM
hXNOGfYj4Y6Sk1/qAwAMnz6aOTVNWMl2/TB7yYJ5e/mKvX6pGeczKx9xBsXaXS/lQiGHwuAd8oKw
G+XafkAAU0wejlSrv1CozbiMwdzKXCBcQkr77vWpac071/NpFBcJgIp7so/N7k0FTcNjwnR8IpYj
GQiVFATsCbo++OI2SDc8YG/sZQhlRW0cSJcSrWKYZSiNFDojJr+beklU03yX5pbx7z9r0NCpqIoP
ZzRkOr3vK2BSA0ugOegYWHZis3pPKgzf6Do4zu2MUo1Jr5GZcU+4LjKRmCF08DNKPHlK2VNXtGNT
0V2WevT2mdnUZN5+KYhBzAJnMWbFpGzwODx8vtBw5+vwLN+VsufFMQx+oeECBZD6JQUGQXLl6QlP
abAw440re0TrYy7vWUx/GyrJncFtjAA5SEZfG13/KCyIMV8hQtOMIZ1Ditc1HmlF84asnWmg6UbN
149hggTgwlU+GbvCdJTFtAZfdYbNnE2wDQQ6xD2ES6AbjV17hIwXDjF2HwS2LvsxW9sUZOBxQsql
DUL0nnqjkZyPdy2ogqsFpPkb4a5KFKXHX871GOZ7RJIOTJ97GaZ/OAZpp5H5EZhjnC7smPA/jvxn
QPfVqAefPEjdJpH2+k9g0XHLlJQ40GfMSj3wG/eI5sxrIS4D/piKqEiTNATIbLLjOxvNQa98kG7Y
kHnAw+UqEn7aZbwZTh365lAMm0cJlbPL15QhQxKOT16Vn7ax9PlXjLTmM+JHLFV6wNNFBQ51RKfB
SkzCdNKlFCVJuoqBN7EkOzvvCzzV86D5movtEH54DgQldgRTSPNtQglHIgKjIVDrNJXM6DKVgKuC
ex8+sdXI6Ty6qFelxGDT1U7vU8ftzAL4SyzIYR40P0+XGO0XeHALjRI9DtDckKldDS5MuRGi9yOd
ql7XiC37PxRgw4b0QJUVXPeQbKd7XgbFXVCdaA5jjPvTsgikQDLwadEUcw0HVdoz/2Uc5n1HFbxW
9JCU4dPqmH8OVjweMg0eWEmJ0CyTGxqav8DViWqihMi9pqPqqfpT/Ep/u65uzdukDyGBt+iqw4Ht
LirEQO9pWl8I5KazOC7yB/+JrcNL48C5S0UyxiFs4CN04LT5u4idieuetJVRI5vAoyrDy6SXzhvV
MUD/QrdpL6r9HMlCgv9n9X32Qz5BBFE4/Lrc1ihqhcsJLoC+sR2Ks3zq9MaHXdoeW7et2GpSvr2v
3jGGeCkvwthAo4DrZNsuKeNdTXYrmDv2+Ut2SHp4Dc3ZWdfsZkhn/4dO8BLq1aRtvzT4ToHDXEWp
K+YXLa6Rz7ygkpL+k+18WiyAdFSYHELrev+jUk7R++iB7frjGs2lDcOEa1Jgrzy3pOrkmyJp6a2d
gm/caRECNMK4VSSaBuX4TeGcKrj5lM/HOYlLGNcCXdk+MMADXjH/X1QuVWBFDkpKr79KVUo/BYJA
lB+JRcTAfXyA0VnuHrx5+FPkkEy2EXvOuJdnIe/5mukL2umWj8O6n/K1O1wN+eEtI22yT6bdvdSD
WvBb0h+cp3G9bs5TAcFb4d0Bj+HrFI+ZXCPwrmkUmpOQ53+PnuUp5oFQfSL5I6CqeUdZ5CtcSHnn
shjYQA8rXX7LI5b8esh/E9cNKLWFcV2mFHt3Yd3WVn3Yc3D3cMp6JY2pkHSFm4pg4u13PzDgnEQn
pq+QzpmgPJt1o00BBUkUKiM6HqpGnNy7Ag44llUcgt0UKwEplRFHqHn4cH/pQ0rC3kEHT07OTsTA
btoEyniBYxQfR6PimMqIdi2rRi1HHT6eTsdhCaFra3uKlKN+0wgATbUvQ7r9/ePndrtDu1YXgsqV
zNkrmART5/7iS4Z3agHb6DtycmZXpWMWjXg4E6zZIMa6qszwu0ndpE3mPgXzQKP5dXhcrBhQ2AEV
GspUtn4FPgQbmhlfXQp1UngIFnsZuGXd5vEb2vzjKWsH3lxO9w6cz3lRr/HAR/AD6Oa7548ZNke0
b0WN3SNx5pCtSpP7CSVKJliGX04Q2JrRfsfoJxV4xdV/lrBKZjh3YwZNXKytMrbbuUEqM3FgaXDr
9yWlXQg1Owt9yrJxMiHEJauSZ8+TRCubkpwABN9yZcgRsNFoKWmnQUeugJgPQuMPbHy2SFOTG5ng
r5GbEgYI7QKGdIWPOJ79hpGUtC7nyRpbDeCQQaE8d/6tQKaytLqZWaAuViicZLI1q9EqfKQ0tiyD
hDLEZseOyieSNOugy1qSP2HV6KvwDU12uswajHn5149LCpfEha0uthyGqj5JmGhmwsSmb8VLH3yw
VwqTC0xt5EyWr/U1MyPLSKG8rN7l4T0ksScRLP397/W1e08UobbjvkAdIR3kWrEi7cM7xvqzsSI1
N17jaoVvLWv61bTgelM+XY4e+fpcU8TeFN07lS/3b9SVyMJPX5J7K59m3T/3ydtwmC/rLD0icKif
IKh8OMaFPkC8nNxB2EzlRJ/1cKLgoO5NzSyJ7b5qU+/kDob5wfnOmunDVSeeNxweGfStlixwhqXz
eofX/bQDxlno4HjsvTbvXFSjZkKvXDe1YM8jfg3GEkrF9IElRtcZ2lap1XZ2GMISmJW/KNrLWe+U
ftAaD6Kyy9mK6hluhq6VshLA0QlRO/liuJoLuBxE4VRCz1+ZZkhA4kKm/DWtYhbRTTDKlvVPu+iE
vXr4C/7fbAzymvG1gRQZ8JFcP+sFnGDT4yjPAA6uXeaijJNKhSGdRGFvoEasrOJ0EW3gSCRM3Idu
vjd+pERrqaG5gD1Mat73ZSTVjj76ZNqvp0btepa/kcam045djIVOZYexCFeNBy1iRbcLF4IUfl9A
YcMGiczRwTOh4GrYxD4ebufCrCayoaSWs3mc+hB1oOpihQNiahP1aSCpBdXR3AGW8JmFurZ6lzyu
N7eSduhRNBe8eXELOVpN8GsR1jvm4G6LnLXSZuK5zAo8LBy7gdcI511Th7jYYPwuXZ3ken2mGTQy
f5MXnUuGhnV8OVOm5PJY1iQoyOlMgBLksDnyzSoxprYrEeR2n0ypEzdw/AHlyKeM81+QXVrdVd58
p689hPdIuCdYVaxiYfhu1itourKBwzk+GE2sFZuyu/JDIsGkdA0UIqDV6nM1hWIO5UvybrYYbIzL
cbzSKd7tsOdLKWi5A2nGGXwTvRQoipd3Lux53O5NWWeQ1kK7cWJEQPC8VCFFZn7qOJFvWC+so0aP
CJO2h+8Y2QJjsBZ3Wgc3HCKHQGH037kgSb98JPYiX4C3J0pXt2SjXtQNWHCxRHb5OGb+vitpIAU/
aZm1NEyXXIxalODMpSPewZ/INCdhFOozxwMlIp2N6phCu1FA7P80HryTAIuo666QgNf3mfXXesvc
It0OR+/+5xoPG+NgzY7dK9EKGf96eyE7TWS1k6JXR1XgHIiB/C1UWscfJcr3oJOrC+YH77w+VuPW
erCaq0VXFD0FUTGWPAgC8jfYWdjuqcb2u93pekmxD4w948LNCxJPTdODddj+HUsixsB+37ecCifB
mFrsqVBO0ixVXsfPjcnAFwoQAA37NwsnuVtpOZ8MvT0ODV1MYSJMH9UOXZlMGiTD/WnVjdJ0ydIY
azrOM4/wlWBBOtwvB6y96eaORID4KnhcpSvjL3TWA+vID7QKVWKUku/xRYUaXesxWnHcElRdZmSW
RsbjMOS+TskUvWr4vH/o2aMGKr7mgjzvWLeqR9qNgJOHf0zBjbjcJcjYVUKxET6HNvGOX0HlHuRv
Q9P4y4OTArpYztV9cmMca7BIa/I1jGtwLuNW6G5iaX1VSMn53tTsyB9qs5zVUsSvrEux2RJ4mmar
ReJveJbM743xqrt2MFI0jGMyhJIG8vUf3B/Q4sN5xeoSo20WunfsLTgSYtOGZPDuHESUVWFp141B
aIuKYwla7F6ckBBZTaQ+Ppi966RSjAAuVvfzE7JkWiL12CLjDpkIapTmeEAu204vQKRPlAsnapXR
AyrEFh1SS5+WoJTw4w1RjGNYCmQZ+Gct61Pc3ZjwlniFRbgIZRAwr13lLIXCVs7B2FDkXoAt8EOt
R5ZocGfj1RcvFzZ5xFNSC1MAPs6O4O4hdMJGRelpEBXwpkdO+zUfoIbuy8x4jLHsLhp9LLtXzpqs
ETsjav7OTj16Uz6/+OUKazpDlgInZ+xgAYtAx0It8+RPJn9pzjstlqN16HAQnTOdoDDQ01KB7mjo
/0RS5QhiFYXBpnSLGEblVgNruUAWJAg3lQSj63/sA7aSrF9itFLb2OOIb5j4AYB+XaRNvr8S+Eig
MqWJ6uzjU3Xg971E+naeyqPjA9RJg+x+8EneWwZlgdLEiMQvr61xdj2g5FGDf3aH9eyDdcG7nBjI
OyK2g7TEi7PcFMf7EMKyXX9eQho9YeHw/uUmEB5NAvMue8yACVnfNfm2zWEk3LaxUozMRjgNcZPN
X0EH8TLKKcXWPxrf02QV7Fzt9ebNC8en/+om5EpyQ2HssSJ5Q7zew3rprXoYQLJ2/eqIbR76y7c2
2GVR81/Jgc40XkCs0QTdb7jQYBW0H6qgZx9x8QHKkNo81PatFZP+bQQZQBYpJSo1p30MpyAzj9bC
STCfwLJ/64P+z1vaZ6L7jzI8gL8h2L1rJMrq84IWaUtizGczVD09FrwMX4vv/V78kCeZBppaAzbW
zrssPeMDIEbUW9CX0CevML9EjBQUG/5/1keUV2eFRRGWEukwf/NDUIFePtAfC7vOADTWlVjAVf2h
ZtYdiCIRLfc5M4x7H7BugT7E5tP/1n6tYHaQXPok9dmDphO+x1t7MkQ8lgQgnZbySRLZ4LwvNVK4
Su9FrS3s2enHy4A75oLtqQX8tI8kSLF1pvzvmo3eQUwXZ86gL3k3YB95ftzQTA6shXqpn8GIjfj6
jajh8G5854x2EqIO20Wdi59xTUP1B0OU+CilUzzBuOLvL1OQqbq1UiuMj800UyYLvDXI4i4/KIRb
M5d59ZP5h7xzuIhNWU7pRI18Xx8Sn3+QlhiHvClSUVRtDndRulwWeUxotiekxm/LBle1evCBMOLS
2APl1tjVQiSbd/2K/jYgTNPvkKiLFdfuQjPkyCYnhBSOw6buFYjp/e4TKr4eax/3MOlH3iCObOVX
Uz519hBLHlSFXQfOwynQRS5Bg0r3DRIG4UBZFsi3zleBacmp7hOC4ZGmxJWEfkeJe+2v16u11DBE
5hnxacDUMfKwpFYkRK3IPlz2+qyNHZdqvRN4qLysp0QALB4LfQQRnZ/2Yb64p/nlEKbGbCo+4Fwr
lHjHF031pH9RcQi7k0Xg7YMgnXE11ORVhqKoLOh8PxJv6i748kSg+aXWUbz5eu+xA0hPFSZD80Hu
D6vlN0hVXNyrvfLfDhFqDMwq4gSk/dHq8yeRaqj3Obi+zfPZj/0ZaHLnptZ18jUkUm5IvnvYg4Az
TIDiyxk7DiAGDpbwOI6NpXC3YUiU0aBIFti6CZHZSkHAT4fFZWbqYGxNe0LgcdLj0nT6fG6J+1a7
s4gQ6aKa4D6+HpiZdRiC7KKqqbnExByh1dLJJPtNOUSydrOifJu0ugPXU/khGVnTH8G/Zj6EtCNt
T6k/N9mehT9tqi8Tr2pnAuMTfA/X7nDHU39YAgGYbP5Qvtm7qYH6/jNGoBGygnZQA5SpRrEAERw5
OGSK2hscuCGBnmLt4/1Z1OYxDd4CCwONUkQv94EgVY0uAzLrnC1zR/vFAt4TQcVJs7lg7153HQ9O
F2CGgHnfGSMDZtC5ftI7dx+qyQ7gE9an0ai+myxi4fjd91Fyeb2qyMgQTYAMxYiprbquPnwV2OI9
rL26mXq+eg2G2fe7aJZLO+0izuzoa62QPCtXCLwuMNNukSloyeDZbVi+Bxnxb1IgwmiXSf3+ktJr
BK+uGose8WWlvHI/K1Mlx6zO3TThJyIOjmRrNAmWD51Wmk6lnihRU/vjdhWIXieB31Wrw/peFXHu
6PBxLPSpJOi/FzvSN5NGL2GjHXlyg8Xwd8kjANjhsu8kaCWkwb9By+NYU21KFL53midBQ+6LJzgr
Cp8sT6mD7Zs8WguvWFPooE2YGhba7OTXtTp5QqrGMGfYEgc270ue4Yeqa7Wiarmrr7EnTMmS3Gnw
/W4kIllyI5Fen7kIH0RHJY2JtEdLBpFJ1qVXq8G+dS9H8tX+ZGkBJR/CIIiyWjfICHxPNCAv0gal
3myvrum9nbSRLgIeG+dWHefGSNAjzpfgUHLy0/GPxUq9S+8cDuPhClpcqj5JP+5u9goAkyYp050V
Kj5gvlNzS+v9I/z92g8oy+aKM3QkuK1UoCltg5e44a0S6Ky6j/bOFAf6di3QAxSyguD1dBsibxjm
9As9o9pl7xgNQaVrevi1nEhKBmOwT2ayTAs8tsM/kZTKlHkuZvYQC/KjP3q+aFGvrxqZHhB6VTvC
REj7Z+G+LneiV0bs2TW3pCfimn6lUA12eFNhYh+EuSXao9CPXWpq9+swKQIZgEc/RfTSWZSW04UH
0fZFJVdz5G6DSH0j17UEjb51op4T91upm+wFVKaLNE59dS77ZxxfdJ27jE5QhCOjawBQzQ+bGT+M
5UusL8x8VDe1H7ATcpgwfQ9Lt5qwMmBgjpkbsJZ6ML4BvP/aIX++prOfRymFRucGYmhbJTBN9z4F
6DJF3hghGPX1W9rF/knmrkYow8r/LTrjEuV0fZyckD4TNC/+T9O6+kVkqyU6B7++rcT4ud13JWK5
gTKrM87sx5IcXbWbuHeiAIG1bqPRNtX58M9PEpB9Bs2S5e3FAkg2Fd3/NlrXTwLAOO1LVoopuXk5
WriN7eWyNW81uoScE+ykbtcd5qXeFo6FVAlDOxFNiRYUwM0oPBzo1d2TKbCRauR+vqfGMzzPIPjy
WSVwOf8Jiz5yliA0PabdsbLdpx8NTAFZWTUGkSr23/Qm2sq0wbJnvi3lFQp6CoA4dd2wmHNp3uh5
up3KcQNEQj0DE29QbTO0JW6qCRHa0/TTBn7inJ8CLrPu2spk2Ucl4jidobE2QMoZpGLw8PpeLtEs
xJMPNg+DwsAfDdaIVrujsh2oKnGruZmQkiH0py1Y1UM+lFOvXavApeju/CZyCwBxG99UPmrEaxgs
9kHw9y4Tz/hN9bvbUahpavAyh8di/3IKFQp+QomR/hFJV6rrSlUqHHqzCNihll0d9vC0bpd1LLsw
RCV2gNrTUyu8NvFaCURhFpleRzO9El5x/Btm9vz5An7+R5cuxxmCVnD2WFMhkAXIWQF+0LuHYPdQ
RG4fycUUdqlsCQNoHpotLjUeAhThczjsHzy3bx2mEoiE6/T5OdSScgRNQEMUfGTBq9X+gJ7V/QmR
3QuwyF1N8MwGAdIHJmh3QwHKFbjmj+w5TN1mo+dW44TqKCD7vAq9kdT+SM27qQaIH/LblZyT/Bvh
FeDMiz10ItT6sg0iBnvTqVWeKwsREoeOkIv0yflKGSB75ifNl31xNS01uS2iAmGCB4Q3m+FLT0eE
VwXzR3FXgs98Y6Jccf2yBZ+DWR4xv4UL6J6JwsXt58IuZCGFucIuZVUJCHntIcY3S6osxIau5Gyc
ZexFdTzbEDmIKiGihrFqkHbuKcMiVZJljUWVuGA1yMOuyS7M3qJMC/0uyR/2uQLRZ8mYmg2YYryg
eGxXi++iuhxpHh0ea4X7TS7EBYYwVX9BYHTrYpNyPPxtNc7JGU04uPxoFG9dGgfPyPBq/0uj4gBJ
UQ+OAnghJ22CuR5263zbzY6mWydrLtBExfXxuegezvbxcoAD4Qh9LIXfj2ijyeMvcjzFC+tTAXio
LgKCZ16IJ1SO032RLTlV5U8Ero1C3BjGFB/vcnCuexrV8pMauKfC/AZUwpuRQzcsNfV6+l6jeMk7
KuKqGC89q74V+xrktBGvw39XBvgNvoGwnyF5cISF8aU0476PXv/Wa2ZsJ3c6+p58wBOnRorMLvUB
0bEdJoDeKomX5Fj6JeIom842gIzlARyZgWr1YW4RPUUhMaLhxTzT14roOkkN/ljTGhxesg1VjS9y
6aokofjqVR1x7ZaT+HhdKFJEUhGb4/N8GZIn+vbVqQX6UvTaG1p6Qah5yYp04vLUdBg7utT2hBzn
HSw24A41vDqbKH/RNh5FwGhXP0G8yHXJFeOrq/4QpU4RW+38jIh/xt3ArZ4iMk5k/4AFKYKw4o4g
925Y9qIBup6QbfBWdSoGYzSxEdaBYG4E8qhSDqrx+JBtWXu5umi+6pVDztnwmx6fcPFULUIETHFG
sJkhFfHk2wtep7QYQe5dojMvaMRBo4Qhk6otGIBMeHZWHxa/8gfbenb4AiIxgI6j9I+l79wv57VW
LbJc5mosZNR1w6hchrxa8l3eK/tlV5TVhW3XW486iWS+OpIetkGedQnz2dC5mtpnnwfg+x5HWXgY
k0oBnPU3KWItFQ237U/d0MI9NFfWAIRSMIS4XdPEYfmvgJ4tBoPlYKWmU6WmVbqgWYcTQd0jU4ZF
p/CcmcNbRQwjbqntP5DrXAwNaTTpGdsCpRPp81KQNEFhdpkox4wVDrg12wbdSkZ5rW1KyyaxVQC9
UtV5GpEEjRvIPNAqm64MRfyyKogdwddBe3tCwxnqnW4FvMKvS2Lv1OrtMUgM05ayh1h9C1+o+/cM
fqKAmG2Sc7UuJCC3sjaPF4eKVBfg+D9k5OImHnrLOcxRWFIz3ha4wfh8cN+W3WYcAIER7qQeUbPx
vJvroFBXE9jxfGftb8lqNPjwj9MW4hX5SjqGa0SHZ8xIGDlOfhz0++y2gUvEF+hNrPz1mdH9A8Wd
M7b9Pi4zPTTHrjdhWgcEPf7re0ADLPVzsFGOaKqDSdVwEx8WeZJsTdTOcE6tCzcD27wIaHcSgppQ
khtGOIMA5iAab0aIBq6n182N0CoPp51GgQRkg3P30McsEiKLE5AazLcS1fhO+lKR+7wqVLuk9sp/
K8ed+IEHflu2UG0gsWTjDUiVjhn+caIKhZQd+62xw3oQ0QrPAv5cpfO6sCKfznsxZtQjpOyRWXkL
netso5pmvwbopMuVHe2R0AW+TKoDqfNUD9Kzc9alsU5FQQGILkUOBNNPugnHZcSZ5on1iuhHjXd1
3WjfrXw+OOIF1KJiOt5fW2MqvrG5nkYwAWzgBeBYA5h+qIqpGmQjxS1aXYCvT+mSI1OoapRue+jq
SVQh1Gdsb2SEjJnAqp3jyX78Ub5w10hZx2iMGRtiACxqny75+t0M+nQt86TP9NyBj5aOL+PMpY+q
kk5J39x7wc9cXTU03tInki95sTZ/wLIpnaMIa6X995j5ayK5pKkDi8n6yt2S45GKYZ3YoOuBIf2X
/hD4bRW9qNP15L21n6didVZ9fyz3tnNUU+5I3GSKI6sg7lOv+f6xNeL7kfX5gzMILDU5Fe3YYyFe
JNqnl2ZBv6J/u0zegy4I/XRQ77zhnsm2DWbJy2e2JyIs5TIHXNzeO52Ks3RtvmKe/0e615enDqv/
7y3oqfXPa5RhHAlvEeHgLLQQ9rHbeHkrQi9E1xZTBBLEHpOr/gjuN+Ew9riQMb2g27nqgyc//DhV
PwhRD3XUcjqYe6TT4NGJcsXASoUmzCvJwe1FEW+0acBVzC/JJPSZRxS+nuzhyeEs+wpRuk/YDl8S
GAU38ph7P8nE6oHETGk+AGPa+gAIj9+wfnY4eAAQxni20etb4AWuOY80DU0MYrbxtiXV8QFhlXkO
9/Gdg4lZA1Kh5Pe1uUkxL1oP96GZWuXr2azyMFtq7cMm3UVxZ8U8ofCN9M59DUol7BBxo4Hz57oh
J88EnBrF88KD4lC7kN+rNMMOBHA97mYxCuqk4ax/yu68m1iIemRP225ROnL7BaHCcqqBO5shjs6t
vlQIueiFV0gQy5UiedW6AhbCxHdnxtoeKNKI96/9V2V0D1z3QkZknVdsXuxx5gDvUqe0PZmFM4nq
uqOu1V8NVQg7THm4DdCu2ifPrkmx/2s+wIcaIHBuQuKZijZcOY0v2LqH8qCt4u+WjaeZU4hN9I2p
iHR2jfCw+/iscul26P8cT6x0a2tX+jqtLW5qVyfWTSVvUOAq69zAEq3FeelU9Ce2H5lRpwCyTOxp
Rm2lLH8ZZsOhtNcWqnF9wMxuA2FL3k80EkT8TNausbLGCER9Ux9Mm5DQ87bu2jfzgo0tGX6Rt9XR
dKOVqLXx9Aea4MLQW9rntDuObhBXc+gUgdXZj50S2yHBh5h542wqCHLxy2Kt1QtxPvY+5WZgp3Rb
DTvMAWQZD1r4ZF+3MfE/5YAwDMM6PEhahZ1Nt4V/yTA4SDEgCqOUeyC03H1Jvdr8tYdd/7gh8hPl
vu3zw0UQyHoc337pDXRVd8nAwqYs0WQ8St/orZj36F5zksD4I0NU6CttET76LJlcXcOWu6j2ndJn
Z6zinXk+oEn+V4BEXwMz81gqAX33Iu/b78ASuE4ZpBfGHYDV2WdJSKu7ke4oXyKf2/L+2fu8LWLb
F6iZUAuEQlDBHO8Fhto6qIh/UZTHsYzUWvWXEX3XYIFrHdpxr/t+jeYBL7MYP7CGl94kJWVp8CHS
LAs+fNH0lWrDjsIbTu2swqMLZfRBqEpSM25bzNel1K3Czgct7vJLXFNWXkLOtCNzTygxpTTdRJVs
xOVO/9cdkOuP8mtoLc+pkgBj8eYUgbkP2hmmTza5GlJzcEPWHVHZL4Wy5aKWync1SI2suYEjkVnA
bv4EvrF6SXCto6U5Fgz42jRz+IiQpzKztJat0yRz82jyxYmhBQ+g4DE1NsbdidWJjsPYRzxAVT4c
4zZpSYl4mwJjbbZqqAajMYh3bTabNj3qWVuoxeQCXBSOUYMBEBgyJ3vx1lFaFzxyJ9yfO49NJu7B
JqprbLoaiF82fqMLtcJxXAF2OtuZcsHXfESITbA9PN8IddWIoG7+nLXvzSLeYjdmJ+iwTJfospS6
eV5nXCCOkI/5LwFyCeq65iYc/kZLkZN4vMLS6vQFEFH9wjxchy3yszWuO6l2EhAYR/cdCHIjYZc5
7eWxb3POWNG8t6uR/M1yViv6UA2qYKu5px0nKAk8jq652mqyrPkc0hy+emwUZrjfGLUtKVdZxerk
nF1hAQEMN7KyqGg0JvPaaueWpECGFjcU/7UgYSpAK3kkBV4TnIEkctcDxCc3y6ANF9MSttsJj/zN
G0X7S3CC5vqa3lACi+YKvTlZaO9iFL46CDgv7UPPfJt7Sj8kqsSYVICmFFTYKYQ7FfVvyxKdkkGY
Dz7JZ61XlIssMSbm7y5AIfXPyHNOERFwdttqT1XXmhMs/t289H6elnoovawgj+jNzzyJRvDg8NyX
8wM3kdDTgTFGHEDqm8EMBplY5kEvhpCXY+3TTKyULu6GUFINDFET9NwauLLcSJ83CQ47FqMIK2e0
m88Twoxdq5AEN14tbRJDCCt/sa44FSqlXkXTmyRTUo2UAXpCndn8sgIKFnS0msl/lXr4wDWls/ms
MR0SbrEMVj2DhN2LEQXNQ0ANy9sbRkahNupAxU5fj4yUwCkM1ZEHvIR2ce2IxkjIhLM7egLu3aJQ
e8i/KEeW/Fe0zhsoakCTNfrZZ/xn+8QEjqbg7D4xmfPl33tZi+35WaxLqX6qbpjo4L2qqli9H+Zp
cqeHOsoNvJ/TRy5LbAVCizlEweXHK5xzB3dNwotPMjXFtLFI+Z95tm9EPNMazfdGq13Ly/bMmjOg
ruazGl7BmbDzPY/IwDiulNEYLvhaIpV49NGdxWRNx4jVhCbqv02pMDghTZKuErsM8aNOPAP1P6ED
cjhrTkK52liI/FgYXAOqbaCXBPd01oSOKlMTiguXUqsUGq9YDVM5vvVT1m3vl/ADQxNVdyOF42W1
a0dl8GI7VJjEEaHRpK3wv1WNDNfz3hWSvqDA1foi2rieUsf9MfDDSp8742VX2dpiNHCHZfwGbIKj
Hz41aiLxKt//DLfJRZzTttr420FkoX7rAt2Sknk82cYuBNgb1wAehtK9BWegLjrOM5t9+WipPT26
HxgzCzYsS6n+hyUwdUXPsZIxqRovY7Pk5096NzbNq5t5jM0dqBk4168+uiNvODRjKM9W+Z6ycMlO
eJ0RiMt+ks2y5X8zHSfYjuXyNoAwXxLtwIWHiLT8QplwH73sZjlNFQ/YJneSqWPE2/0ZBt0WaycS
PJSY3boQWPGkYdQoAscsd36Qvtt8n3xF+ga1g0RLdbPgGd9ZJyW/hKoOBybcnEWwIgk2qT7lRSca
cHo8KwOYr7s1e+iL/rZCFO9EDXIfhxYS34Dnm+lrx54ZdSDthzQRNE9EyoH/i0CyaX2U2g7eJwaP
h6X/IUZNt1DLjcDsMSNRILZCOk2HT/dMbug4IFKW9dEwDbJZJb+dZopyL3IpSE9N15nafENk1YH/
XFRUvKe5i8Fqlq9IzHspXZAe0C4CWjtNfcme3H7EuNryvgU2IvjD3GXQrypzgaBhpYG706OnCxcE
N9SHmMwQPrlV9zCQfoCWXtOd83O5lL/U8aEG4icIFcw5tUyNNuhB7Iv4ZVYm5/96KusqZ2T+/9qx
j/WuwfKBwf5X/jq0e2ikjk3jiECgWPyzWR1AMo0ML9Z2GmSNivrHWdXyFdzVPHI36/oIta3s2PbR
sxIaDH6khsYj/zQCYlMM2Ybrr7YEKkh0xVC+NNaCUm46fdHPTYPCXAjR6MQQGT9GKzDrCfbld4qP
GVZKoYhmgYo1UZvXbQRlq/WunxgH+qU0d6fsaMFNSloqB2a8dWWe7vUr7a5QZ9we3OWKbRIsSpAG
Semroiz47Xbo5Hy5PjriVWdEsKbAtY8iA9mIwB3yvuXRaW+yla7HsnjB+2E2yqDL3pua0PS26X5u
DlRYRXOpwPx4VMR6Y7seLc9SW8SwId468fkoQt6l4CzxuEh+lCjaEclb+KiVRXTNpHMyRFS8OTjo
EQ/rEUd2n4O68olzMLvCxNZt6v8yDj8ZF6y3DH1cb9xHbmsyOsuXPxNCCvTvQXgXysCYqUw1bhMY
fnWTx3hXbO9qFvaQtl73RBqzfDBMCud7/SB3S0OnQcBqZvZJUAWWjvJeTEvfe7CvToQjqIkQgJ7v
OfMF/Pajlu+FF33SRWVMjA3UomWH4XFEL9Cgiib+bGUqQY7ZUtUpO+vRp+4IOYMul1RprbMXz9UM
09JKWc3NwYG3cIN+Q5bu4wsRTwhuodyISrHXEjB4pFQkqHRg3TslynQcBuUsXQI8KUZymApi+qdF
RvlyVhxYMzXigZSlXT+t9DhPYHtXP2HeZ0FL0Dgyjn4UBiO8kCX6COUAFxNU1d1kgj/6fHEFjiwM
e9Rs4SXIYxBojVvGYKEnwBh7KcHq8p7ChwiSTjqMIpzyHveTy4lNysOB7udsKG1dwkzr+jFOQ7hN
Egdk1tlbELdzyjDHyYeWAjtAQ4/EfK1ilwPQexT6n2/MSTaeCJDAGJ94MFWdZnuSgFXrrp/v9dLb
v9nCOT9Ij16dcfsn/0kKkVICJaLRzmT5hEN4KweLMmWHkzJbYJmLRodXgt81OEVCaG/qmoDD5q/T
DJSJnvIVMyFrSnYDtzbzOfEWRtkyniZgEBRewOGNlqXFCX8E0lke7FbuzzSOCDUHSjXvRBdOYAP5
5R4PcM0afyVdnXhMPEpoglxGXB3ggXZj7gFGKCz8JvzNHZyXMjVzBsbDEosXBlbMkvwo/NaCIj/z
5KItNpyR3gI8zmSmRBCz7oV7OqX5G1GXLXojspV3EYHUBPE8+uA33RIXOU1VnXanyPbn8Q43xaNO
Fmx9kMvWIR+4ZSb7zvysCLG6FFpzy8Trc2jQ+S62a6dD9V2wJGFZSj9An5OtNnlXW6y4SOJ3ti/M
FgHuNfK/JFyLPythf6dDcKa1np2vN8/riia1C/oFFD2ol3ip+3Y8NijxmXG7KqTQTtc95lmbkVMf
WzOBcxh5I+RswrF4NbI/p6wm4BJL4fyJDJW6IyRyefWWOx2JGrJ4Y9APK7OuX2EFLcV6s/M7WoXz
q4JutYKCnPso8CT2nbFCbkdhC6VyYW8HOZWxJq7DEc2vRW5jqik7B77eP0dCblo31S+A7yLO2imt
081bry09PTZY7Tl2JlL17o+FZnsfpdX9ddA1y4FfiiIWOzahT2o5BovkpHmXA+2YMMBWzvvS/S8y
nj1rrFayHtYFrR5Gr3mKiMCrMpcm4hLBz9nblpeHijpqL2PuYY11yOfJ53+z4RFNGVoXbqU2oMz7
lIVzw/YWxCWqFlDzX2ZCpTmt+EXwRTK3n/2YWANxV9FIcTiGR9s5/nwFFDqkM9z8YSRm6tXXyyQh
PoamHgdnSkc21IvE+v8E9d7hw8YL8hoGMdNq4VBvEIQCYKjkeVEsqhBhHf8fNdWa79yGZdXc1LpL
540Q68KwFKBSjW+dCK65hfBc4blmrHySNhc2AGRJmwAf5ALUY8yIex8As6wVPYXbmXPyDOsmig2l
jSZcu5/aEt7aPm45EUP4LQdjvgbwxYkJDpv/SilEQtjYtPDCR3lrZJnQtKvGsZ6qQTgeulMWTsT1
xXloc/K5Q73NAbHbN0aHpk/tHfK3j+XgcCE5/DVa1nP/i36Mdszw+7T0JQF/K3GXBzi4r0+luaNe
jpsDsls5TYz7vN/z35kuEiL6B3G4DQBUcjMWPQGzpAeMha2K0Axnc1PQtspjcmFpzkyQbEG87efR
1LRGrOx+Jqq8lwdWH8KdAeZOM98t088xZpYtKU6fnadW4rarnFFEp4nL5E+PFq9JuUQafUgvrD0u
xXcD0TmxMpLTvKDPO4tXLovYTWbTMDdy96rXxYOmbJsSDqXGsLKZbabKfZ4A4gh7SSQ9gy+NQcoL
9Nt15KwK5X24d4S7nywy2cAIZC0yWq1QL6UoTJgDWtcwJdV89PqXn4AFTg1khjKQOhg03sXCk8Fv
SzolFl8daMcVvX8ED4N1udu29lC3VvgMvkVJDQD0vzRi5sQp+2j/uRvawvJBcFlOfLVbcNtopB+6
zPxKesN0vmhBUvjN2RyTX39C1ZWGaz3t/tt6RkmImVv/m6oCqDPMER+HePshDmwZ5yodbJvdSFky
PBnlkaPqFTgATZUsF3cu4Ist53S8qPLznLK5fIW0U3cG75IsE2N/yWnsJhKGW9jLJhnuCstY6waB
5LOJ7aW9MI8k6Zm0H/PuTC/vpB+qqoWcql/c3y7tImwzp6LI/JBBH6yYFxe4871rKny5jKZ/Opk3
YmFNMrenJFdhl3827Kwe0cTXjye8VHZpsDHHd6/2c3GN2PxPNp3cwsR45W0kzDqgdsduKGcDhjm9
WcuA0t9dKLY+b/b0/RbtAqB8o1VTPXNSgNuI0rsbaLF+Od25gD3rZ8UZx3PqSW5pkfAMrDdap7lG
z9OjZiYhbZaO/PZec6KpIvgi7b8gaSV6B/y49X2V99eMA6+YYaO26B18abt5gscZ/CycS6Qgp/Xk
zZZyVA9mvuJpBQk81TThM0NeJI0KmMqHh7GjXyXXsq+Mi798Jk36A/DvsDBxmr5qioeMvP1HiIBU
MmmJjx1aZxGmO2GGZu9rp7ThkTWy8xBnpv6Rm/UL6gwSzSW7nK+IxjO5QizDDxxZ30SYgqRA5OMT
sO76+ehAipHLhzGbGdWbeLDNNp3yATZ1pfb4DAvvWzweYPwIv/4RX+2JQLnPHAnr+QLVbIZdo8ze
uzB20Bn+QjVURGBM+ELqx/gONXhZHiqdzt+/Et7raaBfjexXl+4TwxdUquBJ2ixYqSAEhIc6DSXQ
BGj4pN5MXgXRi14lDxc57k4qsM95XA6QOO9Gq8u4tv5XlHtZPbuTToTAtjxYCO3osgGt05B+9euR
PBSuoapzuDvyTIevolZlcAVV5r4w8b0dhDbEKRJySbPL3FE0TnVIRPyq+H40HMtURvtq/BLfxw+I
FPF2C1x8OhVJC18vWyQ3C8sHx9pKH2wU0eYp75CLTeqqdiQMw0VOJmIhfVe962lD63m49DbkUMfr
izSJ/7lERkkBflM6IAX3OX7FEgZ6G4PpibiQv/vhFxvRLPpOC0Fq9b8kfgXch3JCNjInZCEHF3r3
n9NZmwbGzNdV/TeX5giP6JiHgfWxB0yohmfVJesMDMd5CYhABmC0F4IDUWgkwRilsBAFmjhZVRDc
3ZSR+Q4lpYlKgIuu6z97Xf/oLrU3wTt9xuV7g62bQYWEh1f0Xx8JgY9PvH6wjrrgKXIrCxw8xjzt
82EAQeHGtuT/3cZBUBOAMx4Wv1s7pB6D7tGLVUwN0ITliXbjEz8rWdgcPAyaLPYESoCqHbmLUXTh
EQb4i4QOimrsn7VuX0ZEyRQZDqq2R2sFV/A1UrDA8d++u/5oCAqCHY+PskdCaHKvhuxnFXTnsMs6
W3Yomhb3+UtYAsDTJ2tqfey6Em2hpESmpWoXSmyzEZt2uRkLHaPIU8ckzSFhsZX7F8Idh7P58A44
jz4YEUvCIVbweh9L6wbb9+LxVp2dRUxAbiSFBqONa4/OZLIwE22mYUJt16Jd7TgJZlh/+kZosmhc
Vu9ntg5VCXMWAka7/3kxIUmjH1V4zbPOCVlfHTqiA9Sk4VlAXVyB/pXhH9lXIgZk/iio7i6oJWv2
QyYMUpsM128zVPMvJdobq0W1eIAzBhwR6e/4Cv3Xd+frSJLwr8uA5Y0vYBhAXhBPBRAiBO7DergH
VfPvF/uuHkTBXez2D/L7bnskkB/abSPTULLPHb3Qwn4OS49UirEEcyvYfplwc8kA9yLd3oHoT4s7
uW5SrDdH2kV83mwfhmw2jaixeat30r3Qn6QyqaIyh2XDV6KJoZXZGv4mqttBKXr5zlgSmDcyRD+1
ate5H8TIZNheJZDSlBZ1IdEgBm9KdRV9RDKZELj7jrNCF4TWheSw/Wtm/8PCWDQ0GnRhXCUiGuUx
odcoQ/kmd43wZ/uRuvd8r/jnx+E3o0LfXhmbndKsQS8nykvxCBYltU0LcAJ+R1kGvI6YqNYVjorL
MKBbSyGsin4w6wpWHWMzDh7S6U1xkMPQv2uzdWoJGc9KunKKw46XbgDY0Xx35Gb/3UHTdO0D4Udj
jEEnlb5pbeO/9x79NrBKyowhSYTKW2ZVahkJrlgaOIW7vvUgem/mgmtkmibHukyXdjunVtvhVFdd
IWEeyTriL47jaHitPEa0HckGG0g+I0zGa4N1e+XmfOm6VcXGWVTyNvzRbqcFgVEQ5EmVuCg5vnzn
+hqJutoejeNQkEBQsnkyRgmNMHAmuVWKaNct1NKvVrMszQ2UKjivXLe5JaZlBpU/qhmI3Y9dsa0F
FmtpxTY1eo89607uRQ/2RhamNIlIPzLwEn9AqIOui9+J4ZXJZtI08rLevSz0N+zStL7Z/rgDOlMR
mdEwjsWx7zlBfZK8CR8rJiTY9tw9Kb6hyh+1wzmW19UpZEM5OkvzNb1Jh0Kqf6uuT4JwWswbzEuD
1LLWrMKyZbgHot0Uwx/MKIZGKs4pfhDpJTddAX4CYuhxokKNZSeSGpaZ5sMeyG458TION0pW4EnK
mQbIzJoBwQ7yZ8vnlWH0+TWnkaPgTLF+3QClngS5/+fDy9rhxraNt4By9zHYgb/FHLZ6GVVEHT0j
JcwSCZUwNlglNMGGD7Kq17qWRAvyrWNotoaIVwt5UB0Uu3ezDiJ0/fdCamJk5Q5DV5uOcpBx+i6x
NNb5y+8xQhughzuCzeP/nEYXT5MCckaff/Zodm2KgXQ96cX9QnLbOGh02qx5ZkWeZ7Ilh3regE1g
JgkxnGpsHru2AmBIWRFJ01W5gZ7USSxRV28bcWeVWTT/+sLPFKzgJWhXkpacTQKiHy3z2tXOQoiM
nNIoYQpY1du5pe9M8qEY7pAkVovj/vjC2xm4//9OGh2bwNPrubOa6KvvCg0U8TbwJ5NgybcPKp/j
U19kfy2oC6BUYHqeCBkdbdCvv4oxg8cFmc/ndYB/bZ0SWvlk86CEcwX7beNrkFk+wr59ZP6cFbaP
XvBvh7FJ9ObWtq/m5jF5evzUL0sCLUi35NRSYcJDxyPQCTb5OOtgT2CBH2rnzzC/BEfO1hSPWIrv
nguo92eROXgs0qBcelqGosklU5/21EToxwU+x/PhF77gxy1GIxsEqVGRbU/lMagBi1dhpt+c5KcM
475wSFwagyGMprN4UcvxoPQxxneRWjhELHmPI1NsCKDta6cYObNaWgo4/dNxfNMxaHiUFEYNsj9v
zLjvXEVEpZ9vrBdStxAwEG76FhLkzAV/geX5mYOJe7Xmoj5s2LtDohlgTTNrilX0ekhwZixhdfHJ
U4au5j62clPPWKN/3r9bPIVWmp0620qDTPPNaVsgpKZMoZ/rBTZAH/byngKsArbyzPivvR26eOUS
y3tlxKCAK04LzDruUvTpJ2kLbl3jLXZIeNF6AO6RKW9O+fyNiVsad1Eaco7JqLSXqXUNW26vI7UO
muBp3UmZclVDKDmxrAzzCXDiA0GHVmy8GvexnNuchjC4xLmyAmicAbrsk+Kd5c8I35Ufm1eKtypR
Vqs2vTTf6V4S15GRVnxuklRUMPjKtDyyz0BL1eEdQYGZjZJlImdNX/BJ8F+b+72zJqRm6hbmtWB/
r71WPmqbIOGUu1h4sxPeR9utnr/Q5waFDjj8VB6GTvPZeaDLZpoAZ15oZVaxKzjPxSIXTiYoCQFj
6Oz3CxInzrGx1byEeNugD56X/Wn1anetJs81Rjj7XSOJies2Xa1J+Giu7iplSBkY8BrISErVFXbE
TBGH/2Msx7rYG2HDe9/4XWZJEdDzyRwhNpBif9TCFrSiamx+SmL9LgDKQIA6DwWrSxVZ8Y6uFVMx
1xg/akhDa7E1mhj0eOVMvFZLOKIEeRs1e9vaPOQaLVaxtib5KjgZFxYEaJVpXp/qeTsy2xpPBcwh
pkS2q2RyPp5FwzF7en7QcoaLUI8lRrud3WOqSfVbJ4QVnXi17hoM2zqRROP8KBij91vK16TOcHs3
EdkEOqvltjVmAAeTvVovOx9SIDp9PlKTaCppV6WaDGe+/dAGtqSWPRnQBUVgIagod4fIzDgzy8rT
6Zmph/zPT4tv7no7Rd/Es4HoQDotqWP1gEadK/KogvIHmkO82aV6+ulBeheGnNyosJzInOVcxsWS
PKFLeVx3eB+XOR+hcCWlve2AsZyL9P1hraGX8Xo1if80WyySE2Bpw/X3ZPrJ0a5DAoIoqzPWMVp7
pMdaBsxdvvOgCUpAPTd3P5Rr0CQHyA58sJBEmm2NqLRWTmUVATJzVGOwavQPr4NQA+rMajg+kRIo
/HBrGHyikFXvfqbPvakfFPH7RYWT0PnGSVZvguQcP3aZu1OXwHHyVZO8A2iawCWvdve1+xDrouKI
9EpK1CW6N9bdeH4BUhqFySVur2EhoSJOjqxPQe4sSx+owKC6+oUUCfOxbbypE+2kWfUAh0dXHCWx
iUwTgFQJoLKm4ePwpSsjC3NATwQNNcaq9LacnuGWHjKjTmiakDOppMdM2TOyE2KPBwE099UDq++/
VMWiM1VqCNA1s7fadiY3EksnOvQeWOcecrLrockCRnEenCADMnnTbUoDSZIx3eSqtT+Tx46HmIa9
GwYB1fLdAdrx8vCraZgr0KxTSntag92iMsCDyRwNkz3fsbP+V/Ey2czXkR5rK+47Hyy3CGfzspvT
WrNny5/09/JweB7Y7DTot7UAHiKxRwno4XyQYeveLJJu45M/9KZaCnhmnqDRcBH1XrdpBs3Curya
uK9pGxvdh1K+k2cJuuO3bFas3j1t/LFbcKGfjmKSc4NWBv7QGnBaTFluLJFearRRT/7RcTdt47kc
cf8McNhzuWP7qZj9vKbkOx0f520s+E5HZ3yHo0Oy5bC6Z5k0jEjUu+vpLoRqzg9TSpAMrjF2jy6n
mZQ+CSjmbRz7vWdx4A0HztUyJMx5d50eYDZPAFb5TY5hMCrEk3yzvBPcnSRGZmdzR2VnQXX+dtmb
+VyGcZWKMm+tsUzFEh7DuEDdhF0p3ESuglYgf0/PUSR5aRijIlifVDXie/DLspdTcyA0jlWeL+M5
6ZWkPh5uzU7y+g7SD/L6eIXPZZKmKYWDyrd02r+wPaxEX2Ynyd9vnUPk74FI+3WADbHPW1imK+1T
md3bhlBUEz6Hl9x8StL7iKOsjJItC+BqmQVm6M3r3DLv/f/g5B2Ck2L4u4slnV6NVFwnJzGAvuNT
AnINjmJgdbwn7WNr9V9Qbzd3cOc/Mqnw8b4FZ7UJySMxQEFS7KNlALQ2LsKytJ4mJV8+49i0P4K8
Gy8obX13zZtFbqJnCX8CwRRCOuq1GLXACPwrGslx+n4wTmYkohAi9ig9ktQGCGJJZ/X6dzgkL8xT
EP7gLbZ5cPO5KcPkP9V/yrNNi8upJuaZbmrWn+Ikt3FwIliFr5eOJfTs47E6mSE5hn/+FfovKbAn
sIZFltwFtIWERBx+MJ+2vHhmEaRkVJXX4/86m9d1bIwA0F3TNtaJQ4n2opdjx7eOyo1znc56q2wV
tTbM8cvwCuh9DcgCGonpRV3X4C3VARfELFI68lFa8Kn2KKoI3k9au7adSQhMGWizMhe3fD5+MWv2
cMC8CAxCdWNkjfkx5xp+lwR6spFiPrijS2D2PUYA2iqtuWzL0kKfCCtMex2wiz7SL1LlY1VFMdqy
1EqJU1ELPH1ka1778I/0HBSWXfIkirUdv+DHaNwhCmnwNYuzPiLtDeJpjr6DkC9Wybs6ZCnS2eNu
B3ZjatxBEJkFh/TNRTwyPCSfIbLNBzSbLPqWLwwP7iT6hCronWN/9THCNEQbiYCAjnh1FlERiklc
3OXjbP8OtRgDVdpLpcJjyXNGBJnV4VC2qNS9V+o6IVbwPidHaCgdhZpKkzeGj8N0CVwFrgHE9Xtr
xlFeVkd6MIEkQC1UiO2y7CjuyQetOAP5D254/RDbWKLf7Z28bBZLTihwlmgQwq0FN+F0CAijMlqB
+RyEfOuEccoIPTgX8VyhSf54GaP0MoAF/8W/MGAkx/pr7GUbzxI8O+hpwSTgR8YS56tT7Gd0O4dJ
BcAa5B2BUs7UI3ljLFmPhVryiNwt2hL7c5L592dv4CB2XaCw2ZxeISo08SmW6bGCL6VMPVI9hSWL
iWlTkSEtah2R2d9HJUvcfxHTu3yZOlD/rvLKGqty8NkH1gYyRsXwQIzBPOxwSeNK31Dm0JevcEtx
0bl8wBmYlY7ZAV2zrcYO3k392bv6sZxEw07ZoQunjheWXZ73fxYiKWPEME9QYI6sss7bukpLvEjO
wZnVgN+QEKJ0m+h+Z+vRn5LuvBc0fQcGzr/N8Av4T5L98bz7sM+dXb0T7w3aAow+7S/VXkbkTYob
WnezfjFdcK63tdYzhjc9UtCLzLd8jbNkqhgfElYTHhQG9bWxA3uImFUfqaDLH8SDI70dalIxmedY
uxHQ2u838lnWX50p9i0FjT4Q1xKB5CJI50MMnRCrferBOUJyr2B8gtg/yxpkuHwNXR1W3GA9bcTq
GRwi7MxC/WVoV/kibtG+aC1xS+72NV4YTJ2ccHuxyceYibIvodanxF15Zc44bV0Z5h3qNdTj4ljd
19gXzqVshdZ/Em6zJ6QFYP+mpy7pbFWRhmuVbZ4YdWNkYA+Tx7U0YEfeTo4lWNZYeJeiO2QXhfiF
mu9MavKGmDiheppewEj9UdtOifTbZNE25oT732NNsgK8mSvOhs3q/CvRb8+SDCC5XCH1fmBpt31m
VTl0bp8S5gOMsJ3E72J4cFr+xfFIWozSdbl62tq8utUgmBDFz9lUCM8sQFYunk+QjAQWow78HFA7
YGA/acLUr9sw06UFxkbWuBsQVs3k+yK6ivsLi4qGMvol3ep1DNhpYCxqjCSRg1qDddkFOzKNN3wP
rgDyh7XhaLJIKK6buH8+euiuVTY0vy5FFWcUOMdEGDfFxciZ4crgMmCuHyfHLfXQqbvnXvlhGWKT
TZ7veB3OaEgbdHakxT9zjRoqfgIydLZDrj7qWH28G21krY53YoVDAt26IdMUj2T5W5bnqVSkbx5z
uKOj2MHav16RNK+lCYwPUlIC/gy4765wC4meDANE/lHQWdNFHbCKHNfRE/O9HGI1saooSgTDlrpR
M82W2hjYyLWn5UbVURhfNs94CcgtlSJiv2YLZyypN0merun+CfsP+H9ImruMbwJWcjEoERWMdGxN
DRJ9Y1wwmm/2sF7sf+yylRaq/pZHboVwajjC7lrlWzccUP5+e6UhDQzi5nT++vmk65cwZLvm0jhX
xwXdT/2W+UFyB88SEsT9Dwkecq+lm606OqkiZnAsSs8arUSKUT+qzzdA4sKUVCf4fmGKHp9p+/5z
XyxvBE1nN72FBmW1V3Ny5QnIYPp3v8uZuY0yE9XJaamUiG2hMo5MYG6QR9xdvcrpAsLCLjRL0f05
wKdBz91Df5dFu2B4SjkBqHsrglaSzXjyZwuvtfPtD1a6rfMiVYBN6fCmOsq3MdZjwWax3UKF/SFQ
P/aFqpfG7MD9WaZAtavc8s+MpejxKS9BjxB71sJUxsEhCNhLNCOPKazKd7ohoFEUpx7oESJj8XtK
eKJfj3SHc5xLZTUvhbIKe9jJJ38KaWdw4t+VmVV6M1iV1zqIOjVWHyhrBCbuLFQQ6+V92YB9JHZF
SkAHAi2Rsir29uQQvqvqca7cYp2Yd87OuhM8gS+R28MdAB45nyzXbV8OlLo36jziJyKsPmcswVc5
3ikb2AtRUGWuJ1iZZ2h3RIgPwTncnA74UroVwUP9FLW07HiISubpIiXUwQxREDE7Uz9bN2TG6c5B
PekqJtZBJsRyXDdfZkw58fo2fe5UsnBxXfuPtgmZgYkfUWHXMNXDYuG0JLMGRfbcPbEEEs31GkRD
gnXvP7gfoJ8hKIU0itqvNIzPX3lT7ufZ0UBplZErbOuPsDv257UvXo8Ag8bFjNzI5cd+zqBKo0Wb
Lif+fTCYQDeRCoC9WQL4KyDN0tggNc6yD0A8FfcrdwB9OG3a1gFZNHF5LBvNulpzzf36VwuPxhkb
X9vn3Isjb0LmtVW5FPETkCVnVKG4AAh/0WbLgJZ2zGKzc9+IOFbhs7l2OjTJWURffK91m+HOlH3k
wGTGMnibLwmdqBEcVyPenvSMwIn1Tg0o9g7CYr5aLaJKDQ3/p0iWAnqlsBSg2Nco/JacXklbFgZN
m8e24En6ABuCCcG0iQl+KPCYyvKCXXonmf83OyXR7O0ESg1hl2ZeRP1P35YcK/PJyP+kG5W8smZ2
3SBK9Vw/uvK5g+aN5SJthZKPAVOD19VhKviT4c//v+u1rrnU8HEAO0Kdq+ra/y0a2kYw1RFDviLv
8QFV9j82tq6hhX4oTRk0MFCydXKJ97UFir9fIu7/ha4t9wPnYxHzyLbWry4l2Kn0FMwbz3id/v2N
u4po3jLLrDMufZ2aoKKTQ8n4Wp1KADMf+w3k20o1VxQrwsAZCbbLNRh3tgXDhnUVqeEvcXo96GJL
CTcSoYo4xWkVWvoNax2Sw9YTZdQbx0+kpbqvmUCIlp2jMnqn2MSCHlAmnKf6udyqmVK5BfgnHg22
l8f8unAHL2fz0LqA2VXUjD+Gjs2kVjWpEbU5CVrTOlbVlOnPbfixqbh05pyO3q97RQDEi/EMgb7A
IO24pd4lCQY/g7pMJO6oU1V1m6HkQ4dJt6VxWa1pj0liOcI8E5duNaQiqNdmWM0pHObRM2sbOtRu
CDLATQ/lqoQGHkhvYu8vSXF+R4CTsPyMCy2cliDoiP/qV3FK2Aqdf3MLbyZ5erRWz0OvpfB8biO9
Pokc6nijBeiQ/3O3HVtyCpFY74RMV5O2eSvcKkWkM7xzwQYLJcveKdV7wor9X5GVmoYteT8iY0nC
Zvygtk28daI42tMoEZb+f3+Bz5WQQn5Yn6whYwap5DL5ceE+ws5H6e3/oIvq4ikRLezoQgd7nPxC
nebguvAzBUgVbDQ9CGAyvVxU2eUKLYfznP6agp3EhFmDF7ToOz1ygckxmD3pxUNwi+f+sUwfkDzi
x/jRcT+2ed8OVWBZtF4mYq9vsbwXo7YImmWGqXSB1BXvAsQH56hESaq3lxsStmRPWn5hNHxaI4DK
PpBOq8bYBc3OpnAL4XZZG60dxQN/VriMjNEJjS9ymlL3AasR31PLfrkcumz1V/FeOqABu/4jNno5
6sW/S7C3ieMr6sRC8NMMrwJK4oxTPkw8+blhbWacMKgUDsx2ITKkrW3SPrkyUZww+dCGcyBHeylA
DEpxo1SE8DYtF0WJZXiF3CFIb6/fhox3GAa0ULVZLTeP5GtLobAkg15wRYP2ABNGZ9DMKV0Yg/Is
CAGtGuoBK1APxcAmhVk9LXT2YGrsISykcSv9Mpr3JrHaQ1Ka1wvKKDKgAy4eSfWwrM5bJy/0PEFu
x3uJfG5FpgxbbevhO9eItdDof8Ztx7Gtl8a73WEObaOZs7alLzQy91VA3DgTYCv9g6GPm3wGR7uU
1HjppfGgEpsG1Xqij33eX+vKimEA3FSoeLn67LiN7u+sa2+rR7YtJ3QkDSYTM4u3FwobDKyys815
4zjdhneV2x3A0oPB3iWilP9+FhrWEAlMBr+mLue4qTQG0nYfjlwO2xLZmWlZgesrndfR5/nywQT8
lQo5pD0lTWsmsNf9gdrAO4y5/u8EotdcbtTcb4+iHxnLI5BGrRS+L/3pUJNqL6M/B3Mwz9tWGQBW
ShxIdxedJQlS7CSO7lGqsXtlmfc0IAO/1OectVF8+AGAj0wVpCwOe3izLa/1rTVJXUfd7wlFhYk9
U++KlRLD0K7TGOu26vKUIDzVC6WjxnUJ6zhDPSMGjLVm4tmFZRO90YZvTt+jtQn86qHdtnZYVIro
HCAWdrcKxSiJM0Bdo2Ij8rSYzyO3W5RwqfuGqR0kK5NODxZLjIB55tRCyZbHkXc3eIf5Sz4HGy7j
RyaEA+1FemsiT9c8uouVWU3X8j9fYQ6kbN5Fuy6t4PfCj/TQUYsygMxw5SAuiGADMUzlXvLrtoV5
PUFmDswa1RGfOsIx4Jt6aEV7T/oHqZeotmbd2aCOGsOT0d1oMRKssavrYc1Yjn6cJn5fU6SNBN4y
PUJ3DJ9QIqLwKZhtw1zJF9wQSovvn798PvqJr7kpapjBSOZy1MXMyDqSJVYvvKlw9ZTZm3yi0OA0
iTVZkiy8FUZAZkVLgE6rrfzSLHkiIyb2jt5gYca1fI9sim4hVs1E4PSnx0zTeW3TkiOs63fv6Nre
cRWTcVTcH76b8MUoYzjfiaPBZIHJKs33rc3V6Q2d57IWPXS5Uc4N6Ohchjdg+59sLhfDzCsqHfv2
J4GpOpgX+XE7dMQpxtnVsei0xgNJ2nSo1hLrMb5AwlxIa1E65DV3lMrvtHmPL1mP6FG6C5uv1+CA
uYNMT826bMwVwGVxskER+XsFMfl1yjs89xw92WaHJrIWj089ZqPuzP4NvyqLPT13N8QEQGxow0h+
bYYCWnQ42kLtHWDsf+oS+hrYKkqwrw99It7vYHUr5ywq+DsV0hb+7hxaLPJl4BwLf+h3+l8fvqte
u8Z7wSP2eXXpRpa7jTt0o6jS6qDJZdFVg8ADunL/S6gIH1cZJ/3HRDePBToXpAJscYATdkummphE
bJy7/aImYoBYTF8gPnooHgWpM0jxue55KVH7SMeQpfVfYyuajmR2Zo/IFRFuYUsnaiuXvUtJ1kzC
oqyDlIxRT9NifuLeEuo29sS4GaqR6i/R4YCp8Bt+ydbcb+BSss7mpMksHBnBxp2mU5O42CUIoP9b
E11U9ei/X5cpuZoEhVtO3V5oGVMjzx6Vle4e5Z8d3gdeXNHesp5C2AXi9nvumj+mP0uRYrRXVOdJ
OMT2FmI=
`protect end_protected

