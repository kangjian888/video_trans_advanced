

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DKaw2YF5X/sI0l9aLdTgbK/M5GUdtEMTnIFmxvSMohXCNpaRunL9ipaA59Dc71YrenIGtec5QT4M
zCoGKmFbyA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QRHRuF+/6jbJdc98CuDuU1RSPkw4Mrd2rWInSv90clZq9I1OTAA5/xdv3Hk99Vg2prXDV3YjNqoB
pcpnTJxql+YZ6VAzN0qCk+oUeO1cCu3qiinofcBjVXCdgYxomUKUeE7FJeYz3Js2G/kJGoeHFW9U
+zAl6jadwyF9Jbvv+i4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Lb7wQIOJLuT7MorOQ8eHbXO7nLYJ4w6DRb/CRc0KXgD29tV/pKu8nH2e+iVICJbGwJJtQ3k8P1j/
LscOU8Hk23tTbvsi/KP4jYIAhUNpSlUfm6H0KJ2yht05tm7/nGOSq+YwUD5ni46LH6TZmw9wRjLo
RAHSpBohLboc3y/hVTXta9kQmKPnqAmdZWZqkVyyS5o93+63/fdqbFaxxtwx1mXeZDQ2+2zbTCKf
tbrO065IQsNhLqpQ6GmWS0y4Yk762FiY/PW8xLoCZ1V1Fh8ocFk7LKyATUlQjo3T4vsNks0JLfh6
k4wW0gpjLf86zBHim396ye0D0jCoECOhPpGtaQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZXacKhqAwgw8zLrWO0Oej9oQ1uNqsfSW24Ju9AdSqiO9hJgeX3QSs/Auka01BXmxZF02hREfAK/G
6uXtwOuytUDW3C0vu69znjuzfKa65iqAvitXfuV2wV2SBDUohxstI576S9cHfGPfoJ7tVzjIg2t8
+fXxMYGWVW/hL5Dt3LeBc+ul5BEG9/vwugVmMP2uMG9nGEtDEQeLb7bWAsdsP6jyz5L4K49swiWc
6TrDCW/53r7o1y18s7qcumMrH+8e09lZWlV7gV/qSGCmNFjNoXkvbq7X5+RT29nF6kaEY/1Y1wcM
sqDv/0rI3Yh5PZatD+o2YnHnz7Es16C87EBZrw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pkb010SLYsAhKXcWm+QlAA9Be33Kx3pWG3KQ8c4OXZxiNI+ziOzdNGDZkUALVJhYeeODAczIsICK
xPobg5BZJdmnFjXMkYzJiVNc7H8OtQ+xwCOlZfGQy0nG30bs3aCt+0ciZZz0ed8EJ3QfOUNUrA8S
ACDctQvzk535zqal7JGqVOcbax0rksASegZXl9TYHMAWSFXsQNDtHG7HCq8QaEGySiiJnEz1Zygi
CXmAaOXrSZ/75eRU/jV0Zmfl2uX9M3RD4WyT2L0mtTPVI1Jo5riNKDciMqi09G5yCgGBizlVK0Le
ynsKW0Fvo5j+TrmGuES2+DcsvwzxQUmrQ9n9YA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
saU9xQVocYCNVhmm+/jaIKt7f7lGDiBCwD7GUeN8jk+fV3dDx7VH8BXnwqh3bO2UtgQTq4TYazR5
PsEJU9lk5Y+2uIztywixaUOcY0t6PGvi6DZ5S1UapcNaqz1GzVDJNMdFrGWeodfXgyVpIeng6Jtk
EKceFNW0p1SgbLjlCjU=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pbTosJ4LwLIDFDsIbDQWyryoCwFpua23V6z9HaJa95eQ/VgCaYwQRc0pJmp/UgRFI8GxRIcCfLjR
nDQiDTQUzYsgXuFi39wSqyum1ybk+zJc/c0tfa3zo7fAh7WEKBR6EfegxJoOfQ6umn8yMUOq35ku
5cQGVgAH0mV2j7kgcszzSTcMNu1shLKlPJejpCdXAsAct77F4/JiYgr35R62Nw5TiOPHxLGWKlD0
S4rOzGqDzYI4jb5eYbnrBMtpHWXse9ybFZPj47SvpsioKcFIHeUE7GrNOvNDQPdNPahScNll6gSb
fa6tuXH+3Q3DQNGg7RW23POGEp2w+WE6Kef4qQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74224)
`protect data_block
S64RFxt6+8N/TcP1BwQMLXZiyl6ySs1prnY80ZDs+JZjn/pUttXCGOrfIszPuS7SJ02VOwUFnSvH
/fTXvL3JNjaNV9R6keej9xU6gBtCShLRbOiupHkbzhRjliTgluwwrT98okCLr8TA4T/CzQ4Hrfss
t/o+jwsRIPLq/J3MkRkY04dQIzXFaNvRXepayfCIDz6CpYQvzDJlbjqWGnHl4GfUDK4562qvbIj2
e7idt+ktDg0GFhtdHWS/rQf6baurEnp1ZSBHs8NZU6QvTK43lcxngxbvVHViXFmmuJvGsUJJsLYB
gzq8SxSDBzwk9HiCO1s7TI0zBJS9YtvtD9gjWHHFmsepXty07V2T49GHGzFogd/mbmLPOvv8QAqF
cgFIaoo/XI/coBrQvQibmk9BMEMCLT1xILJcL2KMMBb0y0DROZboUTfz0JN8yTki9M4qDwPIzqJR
VuLogw2CPkPtKlXxSeNwDSsJ1RJbIctdL7l7bfWxfkpehNwmezKr/Yyk69goIog7+32pL6nmEOZc
nU5faFd5ka0No5jBkD80WDHCtrAs8fne3kU4dxul1CJ/YcgQEc7rU46hwjn4T42Y4+h9sZqAXo4k
bl8ev1fnbGn3TZVp2NtcWDyoZYpVRraiQEF0qBlE9iT+lIqDvnV4LbsY9Lvoyy7toD4NoQRMXTTB
jM7yRl6Frg1ZQS3xOS6wHB+BNrgaSbsOuCEhLV5ezFRbDWfjwzKzqS2j+AFrbSDqHpC7wa0XmjO+
fUYPHdn5jQC/yOVVQW0JBEVnE2WOVZNwzfNb2cPVP37ii9hJ8sFdKzZ5JBaqXjF982VwAWItJY7R
cNQrRamLCXOVM7qyFuBPTlNgWdrseuSATMngSW45Pa7GoCmNMCp18WAYDWGuxW06anID1+SYDXt1
Tism/am9RR5WAHLJx1ONJMMbb32T3cd9oKuCcdu0+4i4Thyo9vwJLfxZnCik5mwTf+sq2Di18gbD
+0Ht5eg40ciqfoZXLTcwrxPK9OObgJIh6tkQE7CRZFCJTGz3knfEKbQSzJMGA8JKT12qiKGlqF4D
+gPk0g9ye5OyLPvKInOFORMXqaiwPfp3xhrHLhMraBMMEPMi1rGDkXGGtt69mrEAnmnm+DzV5Spj
crrqbjWfNqqYwHosNY+/PAywrEc3q5kBTf7ojUAczArpfjZj3CxOz05NCzl549WV5/tjMlih6A4Z
PkClS28owP/HaepfkcIhUZ5xJ9wL5rI/FNqvdvi92brakcgwkG5zFUBpZkVXVpfksHnauHyYs1bI
1nXdTzXTOT01zJ988UpZb5sDZAvJdVsSz4WNjGaJo92PY1Tvz37UF39+39SrCWBJg71ytndmajej
oIauX0ch5Hp+YMCyaAMBYb6mjWVvQW5iJP7KaQsp9NGTGoU6RmKyawhdnDQylV41o7gVi++U4dP7
y5sywCDv6z890lH7qBJ9W2A3iZCEK0gJZEW/7UkZDK9yWY8oTQJFM4k6zDEsGoEM7JxMHK2uLi3U
+dwXhxx1nYOP14jqHix6RwerxnIamBhmkU6sQQiDNHUxVfKzfIWFyPhVXNs1fOx1/RKf0PxqBXzQ
1kufzPtwU06MQ+gvhhfvORgxOYegjT01pITE9+GvuW3wUA+VNSbnyqU4Qi/NViAU5Y32vRVvpj8u
1CmEzdROdOnEI4t11d1voQE3qeYJ8bZCsGf6YC3Snja0qzx3sumARmvqnDrxMWCs495a0Ba5UWlM
3ELDKwJHGWs0O7QUM4D0MaL5mHE1J5fkgdaDDJ8E6soc6WLRRgpeSpqVhXO89w9daZRIWzqKnbEW
ay9a0XPu+busC3TEc7VHek88+FUVSnkZfkoFMO1vsa64T4UpIwOu2Rn1fNKE/gyV6tq0WICpRFXl
V0Pc7xnWv76/VoRpQP7Iold/Qo/HUtrljgJLUc47jkILM8dBnvhcod4hErehiSdPWgcusA4kmQ48
7VX6WeTUwyPHIYGdPJxIaK7lx+8Y6mF7A/7+dY1QaauSENPo7G1C6wyvlzVk0diq8yFH1Ne2qTbX
MBdfJ0o6Ou6oqeMYQAlGHrGzvvlj6W46Ggmr+TzvPs/1D2i6CGTgF+SrxgsFhEZ1sC3ZBQcHba8N
ZCKc6vqUHn2w7pFm//iwffj6h8w+ImgH4DthnaMEd1u9srNt7NM2tLHSHIoVxkC7PFZu6ZW7L3K1
pDIcKVaHHTlUx/LF7gBsipGqhV0o2uq2huAS9tTQdTHWYCl5hn+4bNFDPga5Uw+wArBQlWjErvmm
hJknsyd60qQziGrd2o26/zgV2YDWlfC63MYCQs4MTLHLjxvl7cXPLqliCFbbbie0etTbcPcL3Tmo
1vHMQjUYhysVdKrcKTNM5FBVO9wVKx97pfnF9LcvD9+FycMaAtpgy0FSdHjAA1+wpH6uHDywNdWT
zDobqq4FRrOLm6PUl6PGP+fdxzKb9l99owvLfuqhP7ECN5B2h5X1ejVWLyN/DPRpJgzNjQEwS/+h
blgG6KCY6tuRZX/TZOQP+1QiC999NXJKMB64suFV3kDhS6qdt3v0OX6D9ehwNPB7PtDgSDZcHCMd
//PHkbCIVIQhSXM3txfWdTznW+Q3QtCGqjXxQzBdiDTfRocHDuePM4wNF0fB0v7kkqdH05GKvMxX
ib1MrK4PdNYGNysiOOj7s6bWrMtefoMNOXEfQXlY9I3LDJ8sF0/qwNRb6aipKBirg9kpPXT+MO3e
uRczshLvPZiIBjhCMUsaiFrjlQw9axFAGBsXf9hrqWtRWdqcHlkAD8cUx05PCqz2SBsVMA2uaYEZ
NSlwNh//z8W1eRDfi0w/KsorooRSPSmeitNE/2PuiC4lfOo6xouXDKJl1OyDOZ7XrJ7lPCjOSTDv
WEH84yXkIacJkGC+bJGpeEYlhJjCds1pZ8V2D+6tXlIXYP+Uo212WLXONDSmI+q4S0hBVHh031T6
Q6+Zb8axVNlefMAsfqhtPyV04z1cuKSBcIeZmgqhYtBWr+8pdv0LtmibH5Svo0EsYt+IRHFL8O0G
M++AHsa6iZ1TgK2gRPHoajlyuI2x9KWWMvUmOpVWJeTMIsDv4AiM2rMvfs+mMd//qsroFtWnol/H
5RNFPU2w/DL+SAvqam6vUOzDlOwJNsxHU4jxSdvr1uCO5geH1N3oiuz/WAZhRB4mRsQj0URNyfka
jIO/dNyZa4UL9zX5gMd7dYplFvUs6H/a9tJrC5RoKn8siqZTt/TUaHYvqUcMTZl3iR/eBbAyXH2L
WUWYBU7OLVWPScf9K+jOi20g1eT3E3AythS1F2D3IIruznvhTlAsZkmp3v9weTkssbdu9/KT8zpc
cJEmNnegHExYdV1XXW0Zcfv3U9NmkK36CNQfiaemYfEt4Qgim7Qswin+sOdl3PzP6NoRQXBIOLTd
yxfkMZ+qaiEv/M8FnJr7EX7cJyvdI5+T+0B5dCPu44ZHug7At8PL5YfqTYJtx2Hf3RRIYGWvvEv5
Er77ZhFFVDrcWJ2Uv/Zl2ip2G2YqvFW71j9w4LslEjgu26qvfjOQ06BsyJT+IsNVz+1ntIHDPpo6
0dzPpSzeSK85ILRW5N2rpK0crNwfogt9Ma+rEFdudycOixAZBEB1sly2CHRl7OGumcPc5ndQSJn1
WEag0Sz2orKp3Z0aNh5WhqxcC8peugdbHQguQHfAWdVDVcqsYNv/h64BpeTwhF/5ESmrdXcU7C7y
vkaOyj8kOSb7gI8komAId3iffUHm6Wyoe2RkR9gyi9LR1iYoVXzNncr+ia3I1rNxfNCtlO435hgj
mhXWePfdSi20Ib9WsP9Fcx8qhS6Zzg3c7ohtjAC3HYFka5cqyUd6ZqBFN2jyMy/miXrlVu6+UdKN
WthKjA60gOk1lFR9vdMQ5nzS/UCfVFkHjNICXTqLJKkTFvKhxiIAMNru3TD/41q3Uw4dt2YHULxL
KlLZeQJHGskL0kmy7ggKEFGxtX/0UabjmgtSHgNCaFCCfzOswrHIbtTkCUCvMI9cIcm1+0dwcyTW
r6C12q3j6chJmLVfJm0CphlKWBdx+2sUlrGQDoeYTTJw6NgLrEp6Ug5AxAAmX2m8gsWMbM1DJqWv
gJA+i3AaHtBmcLKMiY0Z1r6aXO5y4MJipKc14a7MBKw8toQxOUbAucR+FGSuROCmqBHuysi7RsiJ
u1SqFkLBsJDDV18UzgQa06hIcm9lku6bAmJNzZUDBfO3B9qk/SNjDWZ3cnE2HAcSA35kC88eLomd
UuWbMuWwUjOhaCYafSt1HlNcDbFrrJN9YxyZNONvezR8IYO3XZ3IuU+KotSmFYGwYuHBS4/xh+xn
NuUx0m1uPqmwCM6Lo3qU/aWg2vdmYNKLbeARLBJQID/WBVpQvMdeV9Tg03iOSQvVDuli2Aq8VlKK
HxmQzbLXOunj0iPMO7EbyXAcOOw+aNmZSDQEzJ537CUzlT1TtkcDeZ9Nir314j591JPP/s21DKTw
wcghWYGAuTrwJYYx99gZS+IW1EGVq1tFUbelnQio6jQAD3Sk108nh49SiOtQK7Hi8y9GBy5HdkaQ
RwdUnraXXGhW4lkK0vectIvB/LRXp+cgh7USBhDflut3PezLfp/4mk8VsogA0zsSEoaol+lUxgCr
ckFrzrANzEHVbCmBaR9iztfU7KRclB13Ap82ph/9qODpa3Z8eN4SCMGXUcUeqsUdg9ebO1vWC+bI
SxL5n6dY9hrRpZn9Dz0BO5ZrpGIPyZHsnnJN9h6Z6Q3AtQwHnAWHi11N7rx6StPHJz4cogeXn9bd
rQysz6/gKIxljVLhIyu1+rLtKtofc/Oj/r3IrGaebuIO12bpY6gAcYGztxayqJL//jvSbHl7+vwC
+qJWqr0S3RoYb0wWuEY7Z4+I4w+7n6IhN/KQKO8cBN85zFpc1uE499T8sVm8hc55oyWDVB+P9i5F
UGSQJN1S/Uf5gSPobMPpTljkv12ZBNth5fWE0eG19cxhNQZF2VUQK2e6SvlaYfkdYc0LoNz+pVOd
r19eIOtEIcgVYz8wDlK2UQ7l4HqPmisKEvNQnIQLw02q9eClwlOApv4Daqs7Gz2aE1gkFvTwA/pV
fDdI6OmUP5NyRyK8AKqnjD5NPTC35tlaLEoPsOZvV8nVMZNZcs0Ej9YNrwA0KisB0UA5p8W/IWlp
BgEK9xemfyjS1bj0H5YlRm7p4VteprYbuF0ryTmbvDsVFwW+0Q4C6DkxNsGpryqfReXL/1J0wA6d
JQz9dcZOpYFPIb7LmOSLZ/UsCYCYahRP7Ta8UiBPg4epgEHbRnH7/ynD9n/B9DeukJhEZHcvUUTZ
n/CnT/eouc0Pz6l8sXXO4cdSvwo8dGOFp1YBO3rIFURbGJgUOgpCeHDQ5avoj2y2Tk+fzPz3c4/Z
Ln0quyXhjvj3rYtN6q9mKySrrZIyn1+wZrFzJOIU1lSvwhet8KCvWmefotEZx8dot85WGMVzRBVQ
3I65MqRJSqHoMX2P8q+Jf3BwPtawO6iuD74LRyKutZhoeZxK6IHBkpZ3Cf2a0L9fyRBENZVS8i2E
6jiTFh9pPn/Ngt9TmX+SQeGBPOHYi7YjOylaiUTw5P6EjtGC9Hmp6XMN6AzXNC/aN5U4n3ZMZG0y
30kFKaXP+8dNMYIxc82zNnkphKRGTvWt6nqc+zJf1q1pO+QjfgAwJIUziaSQgrtr60KslhMju/ZX
HibLtxptXS3p+8b/rySvxJ0E7UIGO3biUWlBx+rS7pSRH86Llk9JaGw2wVl7vvy83Ikjuclfp1By
3WkikSBySssfGoG5JKA6gbzLz1KJLBUPG06Yg2hgdlOqCdVnU0LhymI9W1TgYckTO5EQ4ZmM4ZYb
H8sEIkiJfV4QDwPqp6VcV+yedgySOa6U1y7Lz1Bb8oGkFEH3WsUgHR+uayC21sB8bX/UokX45aTq
nu09GPxjKKYyh7wInVIFMDUbxT7/vRdgQS3gKHlCwMl17CknXKiKEJ/Fs+UENPYqEpXqlrIX1JZR
bYQY7JtgvnfYs1e/69VlMdQmu8BN2M0mcqXaRBt9AXl3jUyOV9o5YUgv7YdiX/c9McbywEfXIWXb
qcsEAlsY/uYmASVmHI04LsxiKnXqmhKCNkDsyLdLGXwKp8+Z2XkaPmJ6qmx4hrvxoLYqXW7sS6jS
Bf2vDJWRNFmox9WclzLOavEjnOAdUeXJ4e9+dV9jOwjb41jXuEkgITakKSD7gX5AQL6wv+7Bqq0l
zwmCxJlk4hUHsS0Fee43IrD843V99Q36T4eKiwl7ngzman7v6T8rI10O1VfheXgHkFxlXaYm9FVn
lp2eY2yyUmyWcgzxAsNDM9J+zUOjkRnceCsusK40LHeyOPchh4/zNZKwjR8uMUT7pJIf0agigwcj
Bn2w3cB8N8MRAikDUt/kT3XBhnbIJK4WaOHXAu773Ko+aHv09JHCVbimSlLlmoF/mu9WztvTXCOS
2hWoeKDI/Zf5YfXa4qyz/lnLx8Wahe2h9KJyqLfl6KgbrBjEfUplr3LnJLCK5rKJTKiiMDuQL2x/
XDrF/Gk1kt7bx60J8FMLcLxNi/TDD1qb+OXyevquuiYA7HUEqJe/jD4YuMQyhjwp/5KvjmIpJMz1
WCNgvQKeTxd4CzFpy7i1wPfZ2grkWtafB1f6ldeBpmJUWQCF1/4v+zK81vH6lpSzuYGhEKR6M7/h
goEVWmnXyjoo0tKMujEe2y+0bIuHH47hr63uOW+AnDkOdOTYqADoszTMTZqk+00cXgaxswGSgq9a
LExobOugIRFqXnYPoFzFy/DcQEP8tTeuKOwKrsXuSK2YSD0trZKsZVchb3GBDfJkiu8jz9shgc8l
qQG1SEEdUZwXSoE/F6MXRxNMzXvPfJ4fkOPjTJezU/lKQhg2+w6El1Dk1FhMdMYj0R8G8eeWlBe4
qRe1Q2fCKZA/+yK5rWMfFBZNwnmRssROp1qyPvBor4UoRDLd5Lu8uwVgTGlrH0dgmZESDygWCQbi
e7HeGw2tk5gaw+/86drnC1Q7L4qbJxYNCDE4rttpSDlIQZNHZuOeY67oglPzHtJYtcHmgQZrS37f
3b2WpO9Vea5rT8QL2g+hcJPcFO9sQLDlgShK+fD8CpoHmfD2OpaQi5KFOzoERqlp2PQjsdnpG1+E
ItKvxvANUY0T8mCu4Xwv1xDrJ4r8ZWnP1gJdz4uCgRt8doZ8nmAv2B0umonUNxYGkCtsJpE4xmNV
nS8Pmiw9IMcrZtfpYQEotEOQdyuKJdCXHYxIseOtjmDExBp/8alCoOwd5XDBqiTvjPbQ9xDcycmv
gi6n+MDnYERJCD4LnqLI2qCVUWYyb37UTJhxpHt99FOaTdIwOrYjtt+O2aNmO5G6bBSB2ZFCLKUV
VRI41ek6r6JQgbVu4AaHBlBudLpj1xa3rS/B68BRT31wI2kIa84hed752E//HYLMq+oFQbWR6DG3
wbJi3fQep328rRXRpaEFSrqTGusa+oNl1i8grqUAXVJVprsWwWECiwCVbzHWOnOn5VcjMzNVCvlO
Zacrng9A1QJZ0RsS6jox908b+pWOxj9nXLIXah7mfw/vI2dKUsHGmdQQ3vFgKzCdtVeUQ1bkP06m
PUhO0nu1OnicjDMwfFL1nHRvczkVFt1T+HZ777XJBVMLXLgGfMwN+N7lDam6gqeJcObgP/osXl9F
osNbOlYXYlFivuKbzqMR0U/Ad8ZGXpEGeJrUPCQnUmpuPh1CxwEgbbkqEFleVvqEWIIr4qxuF9w5
uJhH2OLSzUeDijX6e+2ZwjppuUpovp5yXmoiDDoKkaeYUgdSxnDOELNOZPIlcxjYsHjxZOQ6e9xz
13cG2ZHtn5coUOe6UBTXZt9NupR1+J/08d7wYY5zsubAHWZ906CVgzkPIZvYKethfmYCH9P20niZ
wqfTsx5lF+w7K3NyUgOA9UoMbUIlmKjPzIaFW4o9FzkkyAS/XEBrQFnG+s3vMAPNlpU3RiBy5r9w
yrJlJI4B4ocNrnvlAzMgOdDLGTynYoaWZ19Mu1G2eMhuVVGvWI0QqTcPOQdhGtXYINtxGivJC0Kt
8UUqVRbaJjb8YKrW5r0Vp0UPK6sJlLtC+nKD53PuoEFHy4nDZuN5Vm3aDRA7WLgfFi+U/y2tx6T/
Z1tyENePBQxTSA5g+hkCnuT84rUS+yTRKAK2vAu3ZESoRyCrCykcvTteoMack494Xqm0e6odKrPb
DGZZb5UK1jXGNoSpkQuMX6DDxEJVGxa3NItLsbtJZACLVml+oVaKqzwFUBg3wYu0QNza7J5UZUtD
x3rVeILr2oTQEGZlCxYZt/10eYizdlhkf3Cft4Ha2O16IdVnTyFkOujRCOGZR04hs8xc9399LSzS
nGYcrLRaWdXVI1MorSELtgo4IItmJvBMSC1z6tUxHYDsWBGp1SfdalY+ngbGsl9dk8+S8gJ/IaBt
+5CKsAu/UKq5rXJGg5DkFKfEVPWc1FOl9lQNWDH/C/8MLJgKvtKX+pnRk6drlVDyYTukPmsBmaBB
qN5LCI2ob9VoX23jgHk8/XuT7VtU3hC4aitwTpX4lHEUnsNMvXy4tO3VlLmErA4bZVsUCIU9bBqP
xkf0/V5GhUui32+bTGuaQPIJrSITZh6+ue2KVJqC74b9V+RfwHIBvEvnEMJ+aEity06Y6CKPLxYh
Kzk62PkB5Y4YGAGVqHFKlisV+GNkBF8Uj/8o0AjC9u0X4rYvGTgiMd/X006QAJZpmU1NWd+BtKik
y09bcTXMZKPpb8Sc6zgzHTfdBi4Za6B0TFj88EFdvb+IuxBl+xHbXb+djiMQX25QjzvBBfUxKLNT
YQJCjP/ZXbjjbFcmrty3kt6IFoEKKTAfAkonGsuuVScY3dIV3HR2iSnHTCztx/liCkqLTdle/PmK
Q3RfvLloUF/gr2QF94TqMWKaeFD9cwhgU06b9/IchF2vYRNCmJEoW3zEvgN4C1mGARX2hrNVXzZ3
UVtdzFEJLXLwp6d60a0Crt/fgGD9C2KhyPJiIAaizx+wXPcCm/0xw00zFadP4xoPp5q7LJ5/XNRA
TyEn6mA17X2uTwXOGi74FVK18QGhPcop9MW9iJY4w+GtBtLVm2G7y31fdznOx+S7/TIp8In/B/PO
mtJ0WUMmDa5rEXc/Z3Rxk4RdLp8CvUQwhM+Tmi50vklt2eVPMSHZa6eG1EE3trmXjdP2uzSdk+gQ
uNp+R9Q6iKC/OJOczbVhDkQUisxu3Ev2re4sqCKS44ujYbO2JYcf1edgpsf0u5ge2d1iX5hAe3hL
kx9E089xevvS2e/vX338gSRsOVr+Qv1+09+VivGgEu5qr4eoAn7k2bCp3/DjN4RiAWBnOaQFSj5o
34vjM1MPlmUU3Q0Fltd7HUCZI8sMb0nAc/NYCFxSSSdhY2rWHlayxTM4gX6I1tTyk9JiCUyiTNgQ
Lv4FW2ZalY3TUmwkSzeOwpXJLk2eiz8x32Y8aNkbLWmVmHPfhed3LBF4UzzOIXPVIIPU1GCbcZb0
JSLatttnpwwS4h2Ua4xyTYW+/fnVkvBretzHCxHIQkLdQpwYcy+p3Vjaazep2F+rerXaSMWX9dun
9LqulUeQieUcNXUJUZBOX0/OsciHyxiAbDGzPclv2mD9mWBCNyhLLZKZ/sK+/gUgF/uKTAhUAN4R
5NNhd3lAbr7yBo++jDkutWfAkvmz4TpArDcgK16K2NzGt+uJ5p4zjcN8pGs7eqwsOkneMnM5FhDH
31TqA+YDiivhV+JF5E6xAVR7l0Qxd5hH5H4ruqWfiD9ysIYGzmHp3pL8gJlIQTwIpAnos5YNZ7UG
fLJfI3Fg7pEc6nWF5uK3DPNDNjrj9MpzhaFQ0qbbbEHaEwlktCuz3fwMvJIvrcWgrpm90z3v6Gpt
jkC1H0EwgoZUK/hb8BajJS2th5dtkdwU09B4npM1m73M3iAVYww85Yv3dltMlEuzpPiM2XpyEow/
Va+FlvLNPCDpHiJF4IftFX1XI9JS/pHQ5EzRqkSDkVrV58PYILzoCBs17W0GPb1oZ94I+jtVP6lj
a9t28MjM7/QG52KXKqKbwpHeyn1KtCzg6omyy3Q4lcEeM7+kAI8fXs9Spdh7JAG+kqt/MIxHRm8b
qjvvm4EyG/pTn2ZRgalGZNId/krHWTKzPC+XIlQ6uriDT4x2Qp4gspQlcqXumh72MzM6ZALNRGyv
ImA+qeFJ1IGniV9JmsX/lQ7GfwmpyW7xn+FkVZss2iky/5UJHAMgshdM3k1V0dr2l99vaOhoCBew
fXFYoPCYZ9VdA6jS2FKbfspUaKJ5GwYvit3EkB1/j/9YdIAvUNXWtz+S8L8SiP9d30o+Wa4KYh53
vSfMtocfBXNj+ZzBM9HHaJrwLWykP4Ve1gZUue1cnDKqR07hDtB6jvdVQmOdvMhEFgt6l7PrFfQm
6tl47d6HlqXZZOfRz+fgtQMguUiowS5r07OBdJf/ufC9CSkaZAF2CAFmS6pWtJ5AiaK42BGM0bsC
rRWt5RlYRTHyDGK3eMD7LnDDg8iLFCNqi5TrUp/kdBu8Qot2VgJa5utLWXXr6vyz8pgh+K6EalMZ
3gzoO1Dg8pbBhHH0sxvT+ZGwiP2txcO7y65TB4HfVoX41izj1xh4E2cw0Ydrq9GrSoVmJCiTkPWQ
Ig1/YyCT2zApXPWjs43B+kiU05xhKxIXMktgqV7dsNjByML/5Px3L3ItmcGKfvBfo8R62Mn0AKfS
XsD4yHLTdrXB3DSbE6NDnJg645KwLxoL8BMnMdJ2M+MfMr/pZCSfq17O9ZmZkVxI/5lkD7qnoFut
WonbCFLfWTG0NlhTx4GbdwSkI/HMbbNnq6cTqpqZgllNcj7l7L78TwNrfoqJomSHcW5LjqehVFlg
LY7ldwNi4ZuANAi2dUo5vNYTfP0go+E+2B0V9B4S6yALmaruTHFAVfw1rtF/eyQtve7TUUoF33Nv
iqsg51k2EgI33uXXgzT9DdYBpk9dmpuDg18A05sIlmVgfwslu/Us+gWlZm/2mmI+qKLV8Nkumh+p
pzxhmITX2IUsUVa/fZ5ZBkeetHB8MbTWVihHbbEffmrYaQ78sJRF3QKDqxhmYaZIWn9xpRgjKjDH
F1zSjNj7Y0OmFUDbjxHlCkEhE0JXrCU6xHhpUYzOriOsrSH68HdPerwe6noEbJZ2PDYcWPWwaCEq
bl1bf44taWskB0p5wLnk/WsqyFVnRsHPQhvGU7phKsKKYJHKVOIqw6Jz2lnajGYTkPorbYHFo6Qu
0B4gmFf4h2GuhQW6Tv0vJXtXR2PKubaLylwcxTqZEGn9YBvRqdXjWmtlmldWemGfk9WuFKteHECc
bQGYVPHFTsZTvtK4CRisCXo2ssPz0g5OZvwaun0fuWDNEztiYkJIAE8tS6FsCaITKN7IKm5ndzI7
jPuMlpfSv8whkP4AU7Vvljk0o8dr8rtq2slo45HNNs53c3LFIzeyRMYRKs8n8qWiAqJ4BOaJc9AC
Vc9uDU+IoA1Py3R4x5u4MznAZIQLi200KG73fqRiTS0ETjdYEXEfyAuRzzkAIA1ymUHDHVWXphze
vxLf7pgGEaWyFJAB+7BaIzU5Ua0a9fqjzqNqs3kCyVf6rg4u1lvHoXke0sGRS4KT7h3/+sMsKa3p
gYPQKjL82fZhjFCQwoUh1bPfH0aCSznAb8+K0kZYH/sJsMz0nu4m8ZOc73XvaP7LTibPAeou1UU/
Nu6rFn7ShC2Ibo+CBBnJdvWcZTLYRHpWerYCvjB3OIdKEbql6oMqXxbJsf/H51S+XaQA1/wIdpwR
xLbYi0cp64FZl49gkZ8wvsEgSW90d9ErMmSSChNKPSYSEva5+2NPYk0TIOwBbSYEWD2STPFiuUoj
66Ts99XXt/+LSR8aF0AgHtW+Pf2EgAFd7LaeO7cI+SGb8eIDV9BE0lpOq4Nw9NkyiDEH73dAmo4O
o34AtxNDW20nu2YqB5rXOWIE0TJHw6FSjNoJd3sNe4B5ujlxhI4aG/g1An2LLGglY3CfNcX1Hasa
sWyRGxzYYUBQ8yyWjhlK+ttfvUpVqux5LPY9R7XOprPgd7k/yRDFENlTx2QECQNtInpihHo1wnVV
NzE8ZBemJHDO6KwyHDrtbFNagT7k/svtve4uJyQDpV5J8qo8CW6vbgL+4qMOIrgLpS7pExj1nyCw
nwYSfwZmD5tGNclwAt4TCAwPAMBS65R2zrP8Wi9IvTkgOnCJi5glbRW+ufj1IRko1ru+UpFPOk8w
oinWHqpKLZzlBXRtqVG4+3LX8jpCW8Sx3yzJ51hl6nkV9ImSwxfoAwQYnI7zMiEpReQv1urlpwD1
j9uIqRXOnNqgLVX2pKpioAwnekiM/oszz31ZPtfmxORNRfOze3D+2y2Dkrs3jfo+Sx4HLlXpY4Lz
EKvPc+VW9hj/ib9NJhQSQSse8UgXogEHsT+Bkp/evx04uQ8SRKVR18D0fCyZJgzru1TIQ0Xzgj/i
wLzVN8yAfq+G9zNTtwP28n44JOpaof2tF5btNVfBEsjdclK/YqxygfOAEvZ32cYDWGyRZF4x9G1G
CgINCMilntWUBGNkO95BTk9uHseMZF2o2dV63X60awWUsXuRWOGU9HRbmrjGH1ND7kgMD3xn4RlV
Xz+Xa0SwJH0iAkIAsvpcfq0A8II+79bLgCAcjI9c5wTVhjliWA8+EbojT4TB2z4pzRo6j3C+6Wba
rmlpMTQkXWp7jBTEXBBuR1cxt/XD6okXsh/WJYW4wKb63QhgcG60KUtGf0pGP/TmeK7IT6LQvsAA
0ONg9QUlIPPQLRaKBQov8ZQbZto/rDMaOQaIIwRev1Jxzjr518mJLJqGAXlt3FOseQ0smW+93Z/S
/eSWYthTG70hh8yVrjML5mLJyKMFCgIcVy5I+hiP94kmKQu5GwkVDwBDUpM8ld45BR1fW7B7L0ua
3AqWcWoN81C8nF3xDCNCsusLEZI0PI9usMc7/PcheD04AXYqWfUH8J2r92qBZesxZzjPFmjnSYck
lakM2pKU/cgU6cgU+kA/NtkCV1lUeyCszsfEeG+6PTuAU/Q0ASWADClDQ7pNLpGu0OiCQWXCMYat
3ViokahNO7gMtQ2oj/+QUerBpDjtPjRviO2m6UXWsYHC8HLGgoo9JaLpC0EvP9BIA1hH0MCCCeQD
LfpCV1Wju4cFJmkcrmMgny1kaRYvG880SMbh+dWUClzNMQiDc/m9x6n9PZLuaK7BINwIJXEEwvCU
okmz6s/EBeNW/TfPCMT3ZYRZJmA7eC/wTasG+fBoWy+7Ri2mWcTMoxp6qkrMbwnbQ3pDxpExbir/
24JJHqW2G3sf/yAFPeoqz/RJRqPA43MwYE6H7kRxLGhTmhNLSdF3MniaqUuyFUoUKp9ISbpI4eYk
6mytxYoH+kqWD7j6c/bpUpLVeyPxohbfow+t8B2dY7Uhi5kZVyDNVnkx8ductTnYFDceTk39dMBS
IomGXDGQxJ93c7bW/CaIHNkDVjX1OGEBXlThYfzfzBwBP/8PgCoOzh00AULuZqxOJkOjcLLZx6nb
jPSdABF4EORU3DwwCcsbKd/zj+6D7OMA6+mRtM8XWCPreH22WiupFXz7kDoPwL2wlrl5wX5g/K+0
ay7OTILEoFiWYV3oLvb+/WITJnT0Dqntt6oqzSeGqf4/RUD4rAMlnB9FgevHSVZfwEAILmRi+pUF
mX7rwW/tQzpAVYa0KpNs5/71iYRvH/iQupemttLU6myQx9FukLPg4ATxg1OBtUuMqCqpuxfcs/zF
MQYNhf06QyXKLD4zq4bxc1GZCW0kX/N55YWec7Q/h5qil+o8jE08FtFbrQMBA/PNGSoi9mFi7/iC
UbmBTPukaLKu3VYnpIbU+RTwbeWfwsQObLmXvSwttn5dy8Bg50G9+SfTtzHs9igcdQTCUKKDoVzV
xphpkD5NtK0vMdVga8ieXefsWG92XOKHsh/di81F0E0BPD985FTgyszxXaNeSMnvSTilj+Afu/hL
UyCTVg6PjFtVzoTs7JZ85L4GSN/zCs+gEOr8wyZjtZpWwSiyw/V4hBHaPjENOn6UZPFHkEyXMTNp
ZFTPjJk82wwvTtePP/uybWOLyJbdBx00G8qp7tE9pgT/PHv2CB2s5WLquZAu4pOw7++CqAvSpYyw
vkGju+jFdCghX5hq53Y0rJzhb8wGOwqhswPJG9VJnZYTy/mThz8nYqLwiVtLuR7OxN710fNuTpfh
gfUHM9DQtlykGnqxr/CSAnj8sw5dH7+OHPnQ+Yku8ZMgdPdNIOb4lvr6jbSvvVnV43wVHpa09T/W
4fZQ9MR5tq1mOj3F2N9q+7mz+N+FrK+ev39duSRmNaNwwjx7t9pg3Xf9gcV6zucdb3/BrXeXI4dZ
0Tpq+cN5Pib54ENOvfKn1qQVtSBM08KXDhGJvXz3gyHV0YIz7EnGh1kpJp3DI2RLNozpRK45EAx0
flUF8h3dccpCY0EnW6ZxPMhNIwZrzpO5XjoIe5lgI2ManyBJfgp1dRu+wFL0mlVwwcEWa7SlfDmM
ogt0QiK9YXa79Z6HO84HXM+ajtg+DOVGqYmzefR9zTk+aGmWxeX39xEUs02E+un5Kxap+h4H08p5
bqsoWSup8KzOjNzvQzVhDiX8TTfPvkqxWVigtvs5GRe/z+peCI0T9N53b78tJtFdYyPjjQMPspyi
dk9Q1Ctn20n5aVq2vPp5rEG377CKsv78fnMbzGYUQ70BXDYvvtbGmnctDbk5vCgaFGSV6q/vPmsG
uZzWsCpyIr1G90OT7j3kzMQrZL/YQIgperHsnsCNLHw8oswGrNlj55YqI/ohj3xi3LXlCnwL5rE1
FVrPMv2boquCcD3zjrFkSItjFtcy5jbkceQ5xJbVKjHVSXKwCIk8VVei1z2hJFJEgm4vnyJQTLw+
2AYLWpaRBzuVYCl6u9tt5IhDCA1UIuA9afw3m602h32qqACOD5/pzFE6Biv8RFpm91UCwqvME9XU
RXGmfMdP0lEHm/Ri2ZyTGLGIePw5JL/f+H+ynkw7vIDQb8TuHG51rXOWPw9ChP0EDTKp6vkTc3tr
95ZgDTllkfuKg5elhr4V9gs60i8jeAaQV4aRJqsEkNsmmM5FcPzmG4+Yctfzxol5bx24wXEvdUeK
ElpuimPuPKH7/SkAAtTrvur9s4hzvHRL3SP7Dd0Vxlzarquj7dLDRBZmujXSFkwGxZxX/4Lh7U+0
Fp7+E1Ot6I5t552iQOd/4T0DihHKO+8Xc+WCNOJCl8a9xYqcDg4SEzRictdTltCW/33WvzFm6Te7
lfMVeQzAPN3O8iVPmk/7PORWfKwqm3tN5BsZt244TvOUbJsSdp+yJCttoVCSktzgVeqauqqxjn68
5tTTKozjb20hraQ/xoh1fIo4pdIZ6K1P2EKN8U9Lzlv+SOGF3Pr88y7C8gNixDMB7OFZK5cWPXr1
00JtlGohGBxGQDp1KSRXjSg+MbTlZMBdzfsYMKu/5BAhvS8XXF6CDFcg3r7Asb/MgOg7oKgoBlOv
Y34tgkt2eR2bwH+Hl781hJQ0Q+VUheSHH1TA4zUAyW5v9GNeA+gGCAZXWHRQR+CHl7c2UDbgECeq
0PyTYRjTDCTCEfHl+UwTK1mP31XEnaOG78Tb0S49bg04f1EY9tc4LDdIqseLcubvh8kdzQdiy/3E
sSumBmUSI5OFvzXEQJyon4nj/SpTKlryecTXxBqex4dd6JaDNQs10xCEIGoHqsaODzowo0sEdrs4
V7jdgAXwPzFVFEXQyGL9a1C7qmlJRkOvs9cGSoNpGTOOAXc2WHT3VypRS4FjVJt6idzjMjh4hm5r
9O9B8zIe/EXC8XByXvGk4Ha+s/D4C46YVRkZVEIwzbYSB8ncC0xtyt9lZUO/csrDScGULckicuzH
LJsWz8NYdyxY6LFqTJEy2i9f2QpvtFAnpN3qZWMSzxZzQOXX1jFrq/1NfylulftweenYPyzEp4A2
AY2c/A86Iw5ozJ1NaCMQ+95cDnsgJTzIQjdq6xo9sklohvdr7jUg2mrXzNBK5PaPyC3Y3PtrJ0zo
t6VJxrTDUlICTok182Ve31NSgc15yuKwyVBwafzpAzGG59A8rt++G6CsPfyluMaQV9FpssDnSOvV
vLkKsG7sbXbY9KX291cGzLBTnBULkoiOOtUVtA0G3Z9S7O1SSTSEcvyKHmIrDocl+BfThJl1Q0sa
1KO4cc0if7Igh/JdJgyVs9VPJk/+lbN0T5UazqYOUfPJLbqgdvB2TEgY6NQW5TRZOANK1ZquBjkq
TlSQaDmiOYA4R6qcmNNkJitBbNFP42aWAl6Y9zjm2L8JThkw2IaAGQYpMW2XLnXVfvjotmF8qRuL
Gg/LjnvDFZYmt+MrSTFVUL2Q4/VtRdpoOVOYVlwYcQu9uHK+GkpeFn+242yi9pqeX7VAY1kFV41Y
1t9mZRjDwKxyPUkYoGpYM7YBpXS7X0m4Ak0IgAPwpkR05CizrtDYPIYKVgOYddSWuoOo8Xf8d+PE
Btow3rmYE+fLpNl7sapneEL2G9jTihWX9N0N4D46TiHQ+2fq7u5vpqd/+/BhV6OeWGpgipN5M5r6
EOxsnZ5x5dXWifLVyVZ4etYSzec9bMoYRUrZYn1Zs0ObTv7XtdPB9J+N6b82VjoeGDuUcZ/kiIxX
rAWzDFFCqCtCNdkMFZTQo9nmYRDQQZuSBhnqqYe+JSHkAZUIwhpbsD/5rsmXCd6KE5ejAp5uYgNk
GpIC1iAdjAKKnwEj1HynLb5VyO4p3WZ3Y6R93fyEO1xSIfPwKBb5tTmPneOrF8i6vkhkEG7k/M44
udLFY98gZZ+8QwXJf82D3jaDPOxTobRlnk5PV+36RhUL++2t3xRE+tk6n1ywOUtJGrzjhVkmAz8E
hpoOGR+U5hPZ+3uny+33h4PNIMlRl72sNgl0nKhu+Um7N+/D3KuUY3JCo/zVwb4/xOAHe2v3uRcT
M7DfOCjUdw938Jhqjk/JI2B4gVqad5xz9UqSwXHgsHZZ9DFWKVpIpuYE+odOtCOuRtN4b9/Xxj1X
0NpcHzCSXzhFxZITS68kPE+xovhoATGvAq0pc239tzyf0ixRGdGIK4vwaqOItS1q8EZbVuweCsEH
XgDiFbomPBQj7nvbA6LFzaaGV5U8ry3bOJznpAnYMbRHejddxnX4heH82QxwPUxveqgplcx5YgjC
4kujeJqAb53sYE15sDzpghtKmI5CssCxfoG+esWN6w0qQfjUd82cn3mB1d+w0avjdJ7zZlJqXHly
qmC/aSJ4yyGXyEb1K+UybU0KzbXalGitGmkUR4P+4IbMv/2NPZJ4xuE7ZPplLfEgDkAnzArnwfYe
7WmAo9GKOgo7Z+vuLGGhABZYEf9vQ/QHCKbhq8AcTBCbzsCaP4ypTpEDZGPUt2gH7kBaPS6CrwaG
8ttXFJFmc+UkLQHfbeD5bfDQ5fqD4E9tDM8b8NHYmitISmIMMfLhMB5DpSuhUPQ1l/bxvleT8LUi
XbsugKFjc3Z9nUDq2nJ4UbT/rKDaWeSXHkc4doNSs5pTLUTOQ14IdlPLgXpeRuW/8KbZaYKCBVVa
vulUr8t1jzkpVB3J++dbNiedUgciKL3UCDMcx91MmEU6JJ0uSKMSx4Ky1LWgf9sRxPJvU67UN+SH
XTAd7oN8tvIYaTFwCzseJjcKapmoCoETAh/cg+mmm+RauwVdRv6RW33Lh07xgd0S+bBEfOiQyuU2
O4+WWmQAmMcvyXSUBYSKdy8+KDbzkVxPRylqmlhv7rDDumqgiA3SW+gtjSgBkZTEB9SAnMLC5eaa
T+0IrZdAJEKM9WlRjEfDVw0JMOPAr0XQTrJfH4dFZEbZZDMTRmTd6tWCqooAxvZ8f1KYjq/Zby07
LDmjGiVJfKvdiWDjfUj0qteko/NwcmcZOwaiFK3ofSpISxTpTRnDvBLmwZEQpK/zBYzfgfk19ekE
v3FfCTYUc5HIEQWWc0naJUuHp3gmtIjUaY04mOBkZs5u42OvFKQo8/NHIlkKe5j30guJazTmOQO9
w9024IcUB6qaFrZoycS6z7ci+YYgsJggeMLf6eBGd+yYbQhHY4SUvNg/bw9mzFJ3eudr4ICbyz6F
T+/Yd27m9K+zBRsM8QEkPI0jVJORYgiSAEGGL9qYznx0LQK1cE4/9RYe78WxAk7Osg2XqnpdMh0Y
paI2OCVAGICBWgO4qjG9GJ36PZI3rMl/CNgI1HhJLEtodMsxJKnkf9dkdzOxKe0MrKuv3DNX53Pi
s+40NVJdbN8VwY/MJyeV6b908/hLgh5aTSFDpjSF4SQroWkZDKPKkEppAjVH+zpfkPOZIEi44qdH
Sr35ILN5goRKQQDtjpTLIS/Ej+lyh0HyJESdrhb00R4i+LW56ucU3Strdxvogpk6uTCYkBgtS+Xt
pN8qGrsgC0mwTs7EsIF1qntxxVey1/7qzGckgPsfguH12SYUvWTRDMXsS2IdqUYV/DrqldoIXHAb
LXqB+3pq8yQB076bfjSoqz51EN/ZTYa8uq9HEuRglpRgP4Cz3/AQQkGPu/Qei2yMPB86YBDxVJPj
MoBEF1DampQxemLSSqVDkVyWx+2Njd9oEbl9gsTclkMuOog0eQw1uGz4YuOOXjAR9dwkSe6JjO90
kenw6RCOhwD/pXjJbLaSfFevQcSyvnz2TRStrHv64Y0WGHuqXBWdWzdGMvDEi7mLyXrEDc9Y3595
FXyjTUZWCeKnZzwA8rfFYMJNnK6az47PPQWkHxrAOKrtjT+NLGlE+e5FgUpo0qYkD7CglzUfPzlk
dDF385cULm1bSiRjdkHiDtuE6U+4Fwu7IZZuRp2W5H1wZ4NB/et1dwKW0yFr2r84Hba0j6Sp2s58
XN5iHdMAUp3PBqu5iYwBS2WJx0bgwnh7OyLMPSy2HUBEw1qE+tDoWXDFtLJ4mTJAWUGAAsYuJejq
ivyqv6wIdIp+rG6DiceNstAITMpp/VoZjRqEcOT6rjAObvFT5oXk7r+57WBJ7a8WxWmP4zyVnDpc
Ul27oGkrSau3PHq2BjI5D1ZtQGStVW1z6z4KpFrp5uJUC34rIKiFVhX0Jpan21MVkZsmXDNFqDoW
XNUJRyeLfPU9DKDM1olm+UsTO1WX+3lbZbFYJuoR6S8scy0zbpT2MnokhavJyVw1aK2lBcUvcrF4
02NlbBcVCbau3hUnRMSXKlhpoOWE/WGfGLgNlIwYBgG41agou86VcwdheeOEgq2+K53OSijZQSp+
iyvlW7TB7ujvbflRN9Z38TTLbY7WPBugZGjFd2hFO4Y6EPnA3Vc2RH4c7bz4O/s+Dx0HQkuQzLUs
i8pLGvIVcGkcB+CGwqlvoCtvBPBu8HBxvZFTPzKciHBvPyFP0ZQBbAjcyPjoJmQWPYjISYkn1g3C
H7JySjcTMPKZprOJC8hF7YuQL00HuqjA60eDjQONOH/XnmV2ooA39i9Fn3PtnEp26ShTA2QwDxkr
R9u9uKWBXbsKOCvWb47nDv/5YXoQrPjneHHsF8+6G6iVwUNFEIlfoOC0JgiGihiLSt75S1p/tMnj
ZKNlpQSTnkRU4mqV1CoP4/ZT4V5hG+L5IimgMAC2wzYipmK/65TaB5rQ/dVKOm1vw1geNxTKS+l4
JnfElz4aEIo4JhZ7mr2rBTOYPtNiCdPjbxd1csKYnK5yf1VKCi7dUS/LTRJFBVUHwRcm1HpqYDid
bzDyCajqf5h9s/3FtlZ86a6RzxQ2SQgFOYbM41rnKr3Hdt5C0hfqauTRqVqS6ExIOmLriT4m4Utg
bnd0llddtxfHXFUmFjJ7aYWrLFrLnztPI40oKEdIqO4V3S+W+G5lw/FaWzHkMB4gUGo8OycxcRgC
N7dqid56eHV3FYTnigaG8VtCYRutI2w7pAtlwtwRQSpzA0y1Cgr4ADHEuR/Q8BImEpgcqlmjdeEf
Ncz7jepMbTuVi5bfXtGI9A2XDKfK+7KE1K3QQYokhjns/xs0sRf8kfkudF5Pih4NeIK1cUrsVtr9
+suNiMSgBWudSKNNHhU7N+Jwl9PbrkcQWrC2SgA/uIs5LHRXR5Cr55uAe3rEBcQxyFnW2XwwMKQ8
xtb1G0hVyyLpd074Gy/RCssldKCCVNLBFZH/IecXHKDa5ebmcE13tJw1B56PQlLhXTBukgfH3rjO
mZa066g7gaM4/YKQcIzlNt+O77WozTnsbmU7ydoTwNsQ6sgyVRYr5Xn+BIsf7aOE7pPDa9UWNQRO
dnpHZmiz5EtGlTGsNJlF62GD1NqVy2AiKBsJASXoJJQuu4K5/XVT3O7n+cOttOn8n+XH3j0xQtIf
w1lV84OX/6iUL4vkpWbCgy6n9E06xPw2GD8O0GG53VxA0ofONkjQTnet+NydS0p/T6e0Y+zcQm7V
uwTjwpkx9Iry2cvoTcDkXkJHJMXMx83lOwHQx6ZHl7HFvKAyMvRSI9onYOP/ygA7uFyz78ffHLzU
q55RINO+/vI7Ylidxkn2bJGbHCmobwnXDdDgRvAoS4FM53cMjTL8IHcRPul+cohg6QXMKOEd+9Rw
zS/TTNLgBp3jJp0o+SzPrrw/TW6+/Hw0yEuZ9Ef7T5ZEqjsuMVLnJNf0HnFRfcc58SpYZ17zYFOl
J6+ewTXWCKcjtBZGCkEPA+J+p0b04oMD5/ouUS+fg5SlE7AVVI/yu9qyAoMzdEwJ9Oa7n5p1H9MY
E64ED3h7twmEgi3SSw1/52Vpo87ImTtM0SMhee5+jd97w17WJOtrpGjj+75W4Nf7+oE1O95jDfB+
5txewdDz31Yj9JFpKERcuced1vDEyyfHLbI9qS2AJ/IuhzUDL+LH4lHujKGVTnnIWItyEviIBNLZ
Q7tk9ynqHfGQ+Pd1bsoTWvXs1wr4p3HtYlVkV14vM6/08CR0XQZtfTjwFSfDN6JJz58/pose81Su
a6ORVq8Ns4NIvF8JjMoaCDNZuARZGA+dCnypMgswpG8TJBNhBakYFbfHVdMQCEXDTgesBxEZozwf
9pBlVmVHnblH1AuNPvlpCMC+pccG9+BmHzsalHNO8a1UJ5KOXufE5cyt+sHw5cuVmucC3Zt9Y4HU
hVBe4tEg2ayVvbPDxW+nHmWNu0IAqprt6unkGJEnA5ZKbvr9veHcZakFg3kvrbId+p/exWDWUDye
qDT8ifn07UBkFzJwvEp7gnXcbNLXa2/CgLdxVIWeo8H4t3dKkOztoiw206xSE+OjCHBvUq1o9HlX
qTYOui2m1UkmRs7dG0YgYrQy9JA+S/qQlMSecaM3qzAyWBXRV/3oixeWSAClsh9+ViXpOZqgglL5
HLogumuvqsS6GDyzGxF8PAg9xgv7b4el/4/7LSSzbdqyUP8TBvZd0ND3WdwMh73WahhDRV9NrX1l
mGeCCTILOpL+NhMaqIA6Z2IIyaWoIzBGoCSffV6RDoPRRliQAy28JBwODDeNX66nEK/GHCz19UGd
yzA3lCe5lzqNwmb92eRwOaWHUmbwXMlPOTYEqheOp+13L8tAqo8uwvpwictHRoG0Mrej4Pbs4bHZ
hLbOCh6RXX1O8WB8G+NaldMsJPdT5ZP0W2Af9UPpQAwuMhQ7rySNkyXjPMgINg93hIdj/bcOJPVd
FNpupyBOoSPIC8XRcu6J+DQbqanm82U/fydzErO9oqXIZzGp7h20rNv+hmOMatQ0M2dEG6GXiEss
f4dCQS5Ti5FAyNpq7gpGCmXxDsDCBF8pQcf1AXZxF3PsX37VCZ3lS7CufrOyntw+5BSrX0EPTPdV
jnmpap6fDIjh4BxUffRSxehLDD97wxALxlY+iwyHPTJwyxrVA4gqee4LTc1UvwmJIzebfbOFZdyZ
REEp5/PczNriLYzGgQ4ET2RPC1RVOQarZCyaRKenduyzDLtdvncqJxGdhczMQxhts9Vd9MOvteMS
t/EBmqnaIslHu3ah8TeMlPyiL/Yw43nxSIPPBfeitQ6EHeDIpxKnyO7AYOm4uf+9PjDzL4zeUHlT
yawE6q/hpOw3UE1sLSd3zteaWz90/IVJfrYo/ncH5fnoZ/ZOcnSQNbctWNQoaNWj+MVUrYDdQMao
m7yJ88GeL7Au4ZNq/fpqdorFudNXFYK4pRbzxtNetkV2jx5Vg6j+RA5uPYbnDjadwihaR0JjkVX8
IQOglLsU6L4xdOv7v2Z0SRONvP00HMEheDyytDI/77JAqieO8MPBMR8EkpX9NRUy6OU2iDjyX60y
g62P8GkcxUMqKkkXB046E4Qxus9Yg6fb0eZ/CW/8WvkK2h9H/rK/1QigatY6GRE4oZtT1BI0sdqD
rH64npw56OOLdKl73JnSaljXkVQdoAi6pnYnWvJLXKxh/RqhsbbwdBwK9A1pQb27YeEIiQ+trL6G
VptQrEhGVgmzdakZTgAIG8FNTNJtaDZdyJvE9GoB/NwO/l9wCzfNqW6s2tkuyChf1sFGpkyIjiJ0
35bZsbR9mzHEP371LHP6mEpajxpRhzLiZWdGQ/u0SyM84RVHVb/RQtp8bYpZm03V2bO2q7/VtjXW
8P7pCgIaAdRp2ev5AlsBpqRDNZjrpT+o5twwQz2t8GNcKUG8GdSq4hEC5H9Pn3Q+EcIhbgMnQola
+g+IOkY+aJg6wn0Zzv1ea5d3SCtk0Xz6eMx/LsielIGGTncOaztPDNYqcvB6whXUagqmAL2Lujfp
ZO0wzMB33ikdxFI/5ET6qBfhCTa6fbxqrSYl7455wLmw+fPYFVgjQ069WiXQQJuTln7RMVZgNwW+
ZlPKI1PjSziQWmKbqzsmdoT+9P3f2lgDdY8b43pJ35Ju1czgsFnDPyxINjQvIu2ClAmJsuWzXdXp
tJVMQ3DFR1CKEE2LhQf6TWnGnmVeMHJarkqnORyxoDOiiEtWGqgHDXYAMLomWVhFd7e2TqYe6qAk
tHfEQtuTgHmFUTX0n0tbIGiL/a/Nb09KoGUvm2vg2DpFkj0djdYl0FYJjpGW2ftCtAjeRsQa5+VY
OsQHdiCrPrfsRV1niVKhA8coPE7f3RaAa8OtuguNHauFUf1Lk6yHeM5bek0gj4pTuMW1eO3FSayO
TUErN40RFWM1kG21ksM+Oj3f2AjsDo9mhuQixQNAjdiXqdWzjkmeIsTNf8K/gnvezlHTCvCO5S9j
Uq2QWKWlNA17HDKdrsiVzQVFezudMpIfqzNwh9VGXotFGUGVKDqaU20KCIXRvlz56mN/tcUPNVSs
zTk07A2WZQkefXFmn+9426MGgpYmPNSQ+HOJfrOyX4UB0ox6zN1Wfr/pBUblf4sntwRdZdCm6jk2
kDFNuK4gLQqc5LhJw2Za04SuacDdT/R9Z9RJ2kByehKFxdnuNEcfTDnqlPVETkdifIlRVUN7Pse4
Zd7VxPBgOaz4v/h5W1KKwKRi9B5083xhmIDY0Yv3hRjl5ntp154FrL01PIvKiSFoDzNOWtdpZFHK
1/aBF59C4wLWIO1O7pLzn/zaQl7rStrTXWuX5t3obUq0yqA8eENrhGST+j1eDWApBimdGEb6Mq9q
69wnYihHYO4/0Kd4ZXr0QaIfMg8pH0LBPw3oyonop8swP2rhjtjB5Jbqv56GSE3qPffW1DRmsurc
aTCW0g3OHK0esqRyqpWYBbDSv/xQFWoLy2HjT5T/Y/lL3pf9Mkf5YE2hmhq1sRWtvIPg3ShFV4He
1wxZedUnCVo1O+VSnUjZOJV2tIKHihdedXwbKzblqg6CqvwonbQ6OU16ubGE75S5igRv+pI77sKp
1Vw5R5jUn3tI+3Oj4/j7ozz+NVHWdT5PTznLhOUywl0hJ0xy5g/2TpDTgv6Y8ctIK/H97Z7akZRq
Xq+VkiR+ZkycNJaV27cUQ3wMH8u3CYYfcAzxExwYDPDRnNBEPgyODzC9iE4gdv9qFabBOjZKZUWH
RfD7ryaWDvjM+u9zTDCWijFlTMzT/oPYrxsp7yUEtlgDUwJuJ07T+DMEQU6q9DcSVW4mp2BfY4iM
I+cIqzrZQU3jbEXyY12fWERdyjobIgZ5QYfpTZaDFGkAUR/J/GjEQYiCCCJcOu7Vh2kQO219mkI9
JVgUYZvNpH/XQVpx+L4gIAjAkECjHZunx3/pBhpi+MYz8tj2UimYxzz4BUs9360mDZer+56pRtEV
TSNWgbE/9JnUyoVbe+fiblz1YJef+AD+hrGYrISwzqVFgidQ5cKJ+QFBjpsFo13b33RfqHHzojfa
Pegw4eQbP7qGAjGtKN3LtS4SkHzLJEPPKKoRYsJkO+TwaJuqbunoIj2ENMf49WbNAcjfrQa+EMSQ
XLj0ZyB5JjZsdcWbw3sxs+3PLdxMF8h/nzbh+qQvjyVLGq4lVgpjg+qFa6UwinfLVtKiXoI764Xc
ikqvq6VCxzekQ9TvyhSnuGlwzq6f1dKvppumLD48ba88hSabNnWX/mnrehg2BOFQH7ry/w1Ll7qm
XpR9z7EKzfcsRWQH83PQl9TfUAKZOLksJlyxFEt0wW4yc6ChckWz2Dt1M6o0BnNJX4FjNwKf9f0J
zWLvHEFfqz/AjTRqczjgEMs45UuIoyS8aQcEHgWxwwHdnqdQSyVdt1kxjz/0AIxsLkkcE8v8TFct
+9sGYl08PIE6Vr1QQdqb+Oui97AyISvFzQVh1VoGisaydSFqoGO3f9kMDDbzpl1QEuuyJ9QoYyoC
l5eioT8pth8Xij2sg7QVfjKxcqskma8euCR98/SdD4W76BaWiAuhyQHr6JZ+6wkkzm3gXmCnaHaf
B9jWRFmapNhg4w2fcVE97Qw8cnW5yJ2g1PlfMBpfZgnwWpIsXPJq7DGVhh0vmpDK7vn5Fc1C46E9
YGx5HdSsBZtdkRf+UZxjtRDGO2lsuyhun1iDTnYmdgDSpPAQKWaMmmI855+sXyYm91VatxABeFA8
lNvOXVyHieVaFgP/Y+c0TqDAroGp7TA9xEBXdRmFTnRqM6eDLewfRy8VRldgEyLNxTkqw7jI3v9d
7iVIY9+eM8onFmT3IqNlMdFxj6efoiiA3+GlwOEeWuU75Uk3EJtPcKLPfNVZ5k2YkHKTe9KUO3B3
WntUwvvCvK+Ww/nxhOormPRStD+uCHxXtElqY72tKmjvrZm7LNYQs2msy1eOBDsztGgWcQR7uGkZ
EE1qyeiaqxA/oChegVjwJZZPsUUrCIavKIcZTyQTvs0u/7PZmU3WxHugKQzNUOB5LvAOhkMOMFi5
vyixPykZsZhIHfFQBNtSUiw0efF+5zHEWKkyUNA/Vlt4bUg1DbFXJDx0yAhqCEWbpfNWKkFuEGI9
N0e654b7Bhfh8VG0vZUd37/pBsDKtIu1phzjzGEYvUZyQxII4B6IxoHiuzt174ypJH4EAJL/q8Lw
tLz4WA9Z3Oat3VuoEqZdhtgmXlnWelHuQ9sTV1jv3qkgTvQxj5fCdwFcOgCtFG47hdw7Pl/2L86R
tIbBGncTxx1r6xzFPeOjgHN1zqGTXH6+4KP3pE6rkTFQcbfosiMymNYkEjgsOqjIitAHqvf4nD+K
w7AxZ80CCKDtuuj05N1ET106IzWPeY3NWtcKq7SN33d8DpiOfoiWBvTOx6PD5ng4Ga9si+fiqwG/
x9GEQKe9nJ3CSs9BrPCK4J8SUYNfdFQSf/6EGe1keDbiah7fSSgHtL0Oigr1BP+9HKYGJrfGDa0Q
q9tM2noPvePZS5RByw6wQIFyEEyzq1kgXQx2Ch7foMHtZn/IDj6bIMbA/jpHKvcgPJ9nST53X+k8
phX05B6Z69XG4GEPBe1yQBleXN0W/bK0qQINMqijcYcGV1ANbBGUg/+4xG5f53FSnM/GTM1J3Xtt
KR215fAJCfuccGa6zLZ368sY0NdDNkAgSd+/NSeJJrcPucGB/hrdRhz/8VmsBRypmVXMo8FpnRpO
Dhtc6mrcxfrdIuUnuqRU2POeSksqc3I93bNG8aBbCYkTnaJddf/81EYiMgDOoYTq3Ow6R2yEKYWO
CI9/1Jn0NKidPCx1DHywbrpkh0tNYvWyP2PmwLyZjhrM3wNhTjseyLl5tgRplBMjoP0bOOzdrscd
SQv7bO/dYGpWPpUeaEOYp/0WazrgyAQabNh7/q+Mrjv5CgDJ0tIxsVbaDbP6ggLsZnOolQ6PVddQ
e1HngQsJKaFXwQXCUg9ArR00KxDQRvaGqpgL7misKfkDhyOs49x482kv2/1hCr8YGMtDxeLSwFA4
OFRik3eU+sIOuRzUmtOGAT0i1E5xBmPTBcqxEOy71JU1dW6EA8MUZm625qDrwuoAwbNi1Tr9FbP+
dTa0TxfE7lbUJFYTJpvzpkN2Z+A1amhsEs98GDiqEjcMiq6tu0iwabiOz5VdWoJHnw/M15Xtp7+i
mIPahfMB+wahif5Lnj1psnYXB9ZIShioA5nNesyiTlpWAigZA/EE9N/an04Pd2iMqIO8IUSVBG5g
Y+SBirJCCLDtbjmvFc0vkeREruj5/ZQIA1b56ibj2IdEBpniD3bUAuMUaGeoMbUsDz6K5oYfmKFf
jpnEZQoXzc4FVKZbUUqsAnScOI/8aHDTpoezxQv0hiQmVo59N/hQYmLn0ZSWhDPoI9nyS9JyTwsv
ytkM1S6Ttvl3NTs/nCrafk77+VItOc4kjTTz5oR9IGPYG/oGGAs+visjwp5h+0wEsI3ALrF13TXY
V/t4ZuzR11F5GvtwjO4xGfnzELVwAJi1sy90BYyNSCivKgyX5CCRgUx1YiPkwjvpLMNWcwutY1jq
UyZnfdzrg1jYAmIZFZPknb+xeOkhLKsmQ6KjFFiGAuVfQKEGLriDVzCSkvEldqFVG0rv2B39S9eK
74Kei0ulinIOOk0hzvaA4pL0ANZkMz+GVykh3iRua74WTpy6VM5YB6I5ZdC/xKP4YixE2aw3mswo
ql6RsaNXub8hxQUekosKnWYbunjJeYyb68SxlKMKebsDIY06CcsLsaBy/OFlu/OU+KRZy5NdDuFP
eOcVEytRtG7nrIdRYjOtWt9Ad44KjIHBxBX28nojE1Z4+rLb3bRhsS7YtFUJ+IuMa5LAd0Eh9s4W
Ix352ghxx6l7iNWuBQVRFH+uEWQXf8b50kQpNU93eNyN/ynbxdB24RS+sSk968DlRV4iS0b+fViw
0Xp81VfT8bIVX3QpuNGV2cS4LNLMmgTDvIxzmR3t8jb2xV+qU4PbOL0dVt1AhBVc+P4IBIOHMP2u
cpBTacnTXcuby2XcbUJBnnZXZVhgSzc7ZrMsgHtm3nXG80MzCNp0WeGLSQxJLIryCnrBjpA9lByX
ccQ3kcc4u95qx1E0idmUgOujLXe28mJibhhdWPjadV+vkKJPcagdr6Nix4GBqbUiLL6+yqqKIdFU
JSgr4KWNGF/ubwNcDwwQ/1fSmclupd+co7GCHD5qN1ypt98/YQvJ4yHpg7WOxaMvXE2up+tfhJHY
vF62uLaNkuaLAFO88b/JR94ldWR4j3Ski7U7xAePUn0x9474oD5dw5dvUY2ffRQG7UQEupj1MyGw
lZtXcHFojw7hzx8l6BExCQGw7rbffZbwye1mZs/G94FoflwtmOgkXA4uKDL2C1ucroy5/uXMyLsK
yeluTuivuqJvAhpGCTAK8dcpVK2uSWnSYZ9BnGDbJVHWHzPSoPf3SD/s68hwsHER0rQGJ/IZakXQ
wMUsi1s9eusj2jbThfgAGYyWc0JG5u6SZ6r+W1bbCVhWewaemLDl1B6Q2C+0A8LLOSYjUt7EEaAq
MV2qUtjUQhGaysKI58+q93wtripe4f++06sTcmWD6b3blsOXVZ+0PKqBHh4g/vgJYthH0KKuL/Dv
YwowDo/xrfYnxndEmku5DjdQOSnC5YykNmD2bGHTXeZ7YOSwTe+cYX9vAPqt+dqzPZXMkMVwTovW
4N0b+XOJPgW25afPW5zoT6ModJOI+iLTkMAzROrFd3CsKrHaH3xIp/1WQHDMC6abh56qFze2MZR7
JmYNK9hDkTKJd6xbEN7vYgMngF8nrp2EHEKkZ7BzWDXPjZCzHE2HtzhzjqLSZtk2McEncOBOiNto
U6yYFJEVMpHgbi0F9vQ79FG9LuXS61IuxtQ+2IexBgFc14nsXnhkhGEd5o780UFLyMSihgeJghdV
rYCtjtkrtaAoYE2/VsTTt5hJoAgqk0Jqk//Cj/cNhv5RUilULI/HQRhba4w20lGd+S4MnJwhIGMN
DY/jA1/FcoLuZzlFxgX0RqQ81jYbk+G1LGDtD5TTrYBr/E0RMn6ou9bRx0SffU/DSQ+jTdjkM6FC
5Vc42eda3Kp0BJKcRDaNfcUcDKXicokPR1kWOKW2ELECqsfxkk1W2wfY8VLPdWUOOXUv4Z7nU6fZ
TYliiWiNLlte4rcMjsQrkSWL0vK8pkFE01KVDSsURZjcskphwWB7OOZNmIgGkwO2Pzv84Gfvy2SP
bXZ//wtM2uvMcVmATURv5E1u94BsIuflj3jLKyjE7V3DA8jw+9gjIz/y1vf9lnM7wNqDrgp2/IkS
fGxLFPAU/k9IAV+kn18NKl19La+7Mj9c3KC4Ttjb2rlvgoUPwLrdr4FQub6lcciCHIVHm6hYa+FB
yDaGNpRJPxpJbGxdKCGmy8mKGJsx26oHHgFXU7OEqZoAom2SPH84orw6yysvJzrHaefrQIGK6S2J
U5byS+yJpDUhS2NujlyzMpNyeOr0EmxRRIBcEE8czCKKlPFxmzJQnLYATy4csIHQsgTYgYaVsTdL
WTXJneoGJFDrdfMpsdDgfRii92G7hg3r37DSEIOrS0Fdmi7BBsvsqCQyip6dVIS0I6/fuduVS70W
pX1j3/9ZYgoDceVlNXK2PBk+fQdsfvTm/UUoJk/XoJrMWTlJRlvfM30Q5KgXx18eqLAdX4CNe5y0
Egm57ClKEWtl3LG6/as7trbtlOjr8YOkw39+RL+cdOyX/AxfGBjUht1M7d4zT27CgY9EW8qAhhGP
gCHNU/Yl7azsHGj3m6vRchVgPuySspk6Z6l8AL61f94uiTauZv+1bOV557aQSQXu3uUsywrUYpNG
nQqszCW5HxYZU3ypSYRYYlBNFGDIbGWLBnrCnbS0HMvyXyOQ0ZpZ2rFXbOTW68U9W8ic1+k793Nm
HsGWvUDdqHVwXzvtSsfTASpE5u0nT3VHEQ5EKPIw6lpV8lDP01GwZhKUEWe2pPV7d1M7qrz25b5h
7Z+i8NOEZBH7LE0AsL/AqebGFPDg1bIzw0/4DEuhuaG99GRb8SWds5OKh5nhne8YXOeKAGgx0hdT
/Egr1O9QL1Zxd9Jlyrl+zEZ8ZkEp11i8b243e3BrUFS+lIAHhZywOM4gXK6Fa8ObPIvquTx4UC+2
rK51u83xqFsg+17t5dHE/k+Sd5jWdEtfituxVa3CLkyGe8nsElvX+OGOF0zhBRPKthretsHSYGDL
KvYnteIEcHbKUg7nbAUKOmMjeBIz7Kf/g6Eo1LV6a9VpatlBlzmUW93UGeVfHEJv/QliPduz9WLF
jUAidu75Ij5n3sUJEa/A9VNFUxbWWG9DUMtl4IoQzLbm7Vov1IyaYMMRDyXwTXFOKYeLRoNkX6Kn
su0+7tYngIscTezxXWz61DwVAm+gq3E0Ju9k9F3zwJpJczHcrRiJBVereVK6MBDQreaOqph84Bsa
DoN38PPgRSjvaqx0fGedBBTcVEu27afpZDMQHf0J9dwnl1BXXI8dDWvS6UzRn2pNB6XOrUGxtqEf
U9sVUnIzx8qhFXtNndxPmtDjQ9T6w7bYFcE2/etCip761WFiDBjIBGVCFlT/HORaxHWp/LdHnn6N
ufSCe1VzHWyO1Pz+NaDD0Chec2q9a7S7Kt+UDim3u3S1zjnhJxLaEpmKloyUrUKiM+k2M9nnkm3z
4ulMzAKLOLTy2cCT+zgJHVr7EKu4jfHstPNEBSliD1r2da7Vzz7OwtZ6FDUfy2LVMyjdv4x7OZ28
VjBQZoznSs0c7Ttbd0UeuisJUGE98BPaRCDuD06ZcjA0qe1hiZtQiWkvH43tGoB2iSeJLgIF88nu
Gz+Xh7bQVJa0JbgM4+odCLaIu1iaIviWHyl8NNKAXLrzCMg3mta6tWvR1WDOey4NcZca1BahduHr
dB4BfI4NFW533Y5tLzDU5Grv3K6cohv+WwOSXWppMbccMaXdZ9OBpVKx6fY+84m9Gd9KpfmsS8Xx
zQa5sAm5Ey0HsJnhyLaldRkh0SRrrqAq2N0U5KV31Eg0sgI7l/Q4ynApUZV4ujtewA6WJxZ81Bmm
IjLklsIK6607c1mq5Br5W2B3GSKbp0wrElj0izd90hGG4ZY4s8WKUnxtg8cAjB5yiwiVtRuqE/WO
qeDUPMGYl5SRB99oCjuFduvrKRbAl1uxI14H3nX9r/mzVXtyIpC4tuGmSkwvcsbWIv1YSIGtJi77
xgWeSwKhiEHQAjfC1hHekLBytSyZpbnmRT/dO4k31Wx98Zv56DX78yo7Mqyd176km07VVYf7llAZ
bdizVfcrhHqzyMuNUmLon7XATDwfaoCQIeHyGa/fzIC0xKM2MAEqPbIqynZbdYvAosyGPkvw35Xg
mDSUvqdDOumnif9HUvRufBWrQE2Ub8zizwnXHzow6qBz4piNWawCoBhWXLWDs3r2McwndaqSBGFZ
iAlcSmP/h3zQlQcAcdEpkqDoETu341UbY3qM3rIzXZx5vrAGk5IPsLj8CBcObctoKZLqe0diLZmK
dAuSCSeizoiI+5Ao6I2t9CLAHrHAHl9JM5Ufd1LnNk/DY9TkOuX+9i4Did6Ky5vp/u7QD3yHW8VE
H/8KIBs2KOTYSEb2ZZhY8PkuefwjdG8D00gSrtq3vnm3MlohUdCCte+mzeM4B4KxT3hBiw4vk0el
T71oqy4xmgB9pmj7y9C4QC5ys0LXwaBj8NJC1PEy+6YE+WU7anRXeo3xaH4oh3AmqN3brpx05dRK
qhnyS+jfj0VnISPm0NZwIi5ndBGBoVwr83sNQn3E67mUQm9akj5ukqRSJxXzDac3gJpIsZ1rLdcH
aMSs/Ik6GBg/S95LdytLrs27eKCCKDSnNa71jD9BSOMMSlaW6+RREqIzUVQzzeks0FqJA3SeQ0K0
PVkzX/d2H6X2OCPyzgP9oxfQ8bCI7q17vkp31ExVpZgHi+el5/Ua5BsUFB4eJl1Y2NHdSd/QsYfL
Xaek3Wfki3A1pdCCStPZUB2tlNFT9PsZox9BlTwfs6ADRo8Jx/tOO3JVsHFQ2Kf2vP1l6Oy0qK6W
e87mOG0JC1UAdIuoWy0ixPjfLfClYua9rZGp6XsBjj52TtqDG6prkkZDx5JnrfNXs5hFwwz1ZNF4
pnwl3DMDsJ/ndEPzJ8mISyTHujTaWeeuuVfUCVDy8gF8fLP+1TL5q92sv6m1Eo6GjZcMt5CMltE9
TgWjQ8A9zlXPyYd64xvOXfoAjb848EIGGnbeau+1fwwfZX+L1mGpivfaaX6Re1A6O6x0ubnNKj2z
BZedNyLqPx90FDBAI/sW8Rsw7URp8VaAlCLmHgtBCxa1l3DQc062bjgyRyV7Vd0z2SWDO25/Hcq3
pttGy1gzNoLJjCt1pe0/zllpPIzz2mqvuAYJEYu51EDcrIU30Z7scVSwamdZiEvfOTY8ZmwwCgcx
BfhiJ0WIQl+avgkBmdfkDihclg9ZjVXUNAZVrUp8U3+L4b7dOeovK+zKxiEON+eRijEFcr4AFcGe
U2PBvsG4Cut0Wqed8lnQfOnmBRXuQLe1CZfJ3PUPX4wpfPOhZFpTv7nEXtni7FPGG8dWJCGAOrJJ
W5l32N3Y0dc7ufT23OvVpn+PeigYj/jIGM2bAG2z8XjA0v7slVbo6DT9QJBOpwEu4BSOt1ed6EdD
uujZM0IBlONlQhg3z2Kkx2uZNhodecLWeWWcZnOJRjTBR6Qh9u1H+9uzK3AOLNvVbBXpamxUVlma
GQ2Ta5Pui756Nynj467hdLYLAjxUOCHIUKFHRlZPFMkHdrC/dB3v9H9pN0d8lFCBH5tNF8Dk8hQE
E/NR6JtchIRAbhI2A8ZI3iMLCkbfnBAyIUuKI3qQOgcXJbeLgzfrtJ+7srPEzBw6qwnAsYQgBq7j
0BpMQabmanwMyZFy7FwkXAds942aEnkrBP70EL27UgcIR7TYPTXqUgIQaoXx9ysvJEJYySVATpYL
fbYRO786zN+qAZM9nQnWAYQsmxTm4ohjD+zVykNie2cza6K1ZmoCI8p2qVrWdZsybq0SIJwsuTpu
aJm95I/jXUZGGn09SyIBbt6K3BJKLpKMDuJ5+QR7CP2XsCgOHmxSmSV6cHXObvKKh2lw0/jsRwuc
jMQ2YGS2tQ9mm2X56AS37T8Pq0CAwIUi8Oy+z4DG6KyaxExk2qM17gOrn4sqn3Ain5Zy5xx8udjJ
6bVbbQeWyrOmxkxlTRqzuwaJ8RZrL0ygpFiwaN+aGaQ69OE2CPsMg8igYSLg96IKj3gX98eWLxE+
TWW48+rwno8wuRhoAJ/77H5j3ZgkiYBYCvo75tsPnN/w9YMoGGLfJmtj/CM5fboFXdZRvpXiFcOI
/C7Enoq8PO081YETai6PvhcnFlLK2MZsxDsIjaBkjSCOYddLktaAZtpY2DW/p6HKuf4Sz1fmdW3H
OQY/+4z7SxK6SWsoOa21aeysW8CjLqSbsizkVEc5RXHCDfXZ5MFc01zs+ZiaATGCatCfV4A/ux/4
Ui1b+J0YDOyGpVsS+YBsaFS89djcti66hfR21wdg8fz09iqLQtsHD3k3JI7z5Rpm+uJ2qWiEZDbI
IxQ5Ln16HmhG7HyCf6Q4+u3bBACothfIlT2grCFwd3tn0p3enl/RfKtIrqsyHnhqkn2lOMqVokS6
ktCMaXlt691Udl/jKSej/pyg6mv3yT2YPVCEcqaUwUfXAat8rqCaWxRk7EPc5OTnA8UP1uI3AIL+
czRbgW/NIVObIvsY8xuuW8b1Rd5QQ6hv1QtwrZiEMfJUtac8NwfbC/MG+TfAmwTKjedO3Zw8vjoJ
t5/fudWCtEJzzsXKzarVYB6Yr26aCTK0PWr3CHBo8IQyI/GIy1ySECPOK9e3slKkcg8LQ9ULM3IA
9tP11KFgSCSSUzYYPboOJpAZm0bwC4s/bSLAOHOWoxAwoHC7KOINU1H0dmygtxudWVjGUYJjMWRd
N7axz/zXdGyVytoWNSlS/8P2xHQsL4NYaBoX7XwmlO3O4BhVj7Gwim9ccGfrO/okYpOT8gwAdr18
U2r1EdujsPw0ZEjNpwFM5W4lASNbeEA9WSCXbXPtKN2/uAW3L1CTFjn7Xel44QQOzn3SjkAtp7gH
0HcX8c8rNzzDlhjHXbAumpkdKj1hAuz2iRQlALgdH6kDNZElVaJTRF0GFFGqXa5U7J9FMTAo/TCl
gNbl1UygSdfV68CWb5ATIqRJcTaFiJIK+TNajQjTjjeifwG7ao/ucWyRZ+THmBKOd2+eld8E1rZP
ynziBrXrxCDDtVfpJdEjZLI+juh3raIvoWqZ93xgKMNJJNP/IDdEU6VKMOMs2iXZlWmwyuNCz/5O
1mrf8fiok959NBZGLQ2cyZTpXPT6qcDuQdjXNtitzBxKozzb2rR2emfco563nJnhnCYitdm4ND9Q
W+eAP1Q4AUP0a4OpWOpasulxZzUSJhnr/bcOslpXIkgm9v06oxzvwUdtbMuZuG7Knfy+lZyfwu5R
qz7IEWfT5wY9TTLtMfyar2OB6Y12ok5V1M9cw0MMkPDGZnS1yDjgNLoTrlM+CHLQZ0NPnYM5V6T/
z0igicpesjBmk+N85/IW2QTzcgSRprUvABxu2vO5UW5i6OE1feSsNzhhkljfGZNqfbiphWPI9C5d
VVmKF52B+oTu9eDMV9dl4VmX8Hc2wPQtxJaIh6bgHCyckpe7fSHZjOqj9DNaw84sitgr0HJYoJsb
z0gwQXdnS39m0TrP0U80siQzpIgFnTLO2gLFZY4t8SUnzk4GJd2Awa37cszyF5gHwBAvyoG8JaCX
JyCQngbxMmfWOibclM2usBy+ULPVAaNOXn8pWoboJswxMIPY+6AqSrx01imSQcuX8F3guCp67bAr
BEz2ibtOhiYYJ0DPtwcqLcfS2xkhCZOTClMveKkYxCs+9mqqgAaS/0C3ApWv8b6JG2c0nb3TP6p4
q84UKi/PeaMaHX3ShZeCPeoEilojSg8dgzXukiVMHofwJ6+sV2TkL14DBOIBXUQ1zPZTu8I5iweM
YmCxER/O0xIO6oTlrUQTjWgwFuXCq0DrUXQfofaIqdNPIJi+X6IsPcA5iYBTC+/3BlDP0F1G/yis
sLe6Y9asr41ngK3/IUQq5TGKaI0myuDV4jaDQDyPEX/FJWiyb4966miA4a0tQjhUqQ4rULwUuqob
tRw2UVK33951tsP1kec3m06mEUrACFnhJqsEwZJs2s7khZRAuGegxbIBSvE09GTod4XL0+NJoUHu
xqa64CIW7qUTKoea4RFjkHyPBj3WJhQjOD0rQWQ+UGQcTYgEKUZA5cGFmJpifvOCulRrLwzrrzfO
2mLXQ3sCTk97JoHNISRICCdWyJGx16Zsi6xTbTtVDKPHU4iIRF051aKxUGieakgggvxuO2xeTvWU
G3RNhlmPaQW77IAzO3SMt3B6hH1jtRBLhEqifoq4/UjvbsduiUs+zeH56/3mlkle6Oct8IBGkEdw
SDeTYysfmzICfotu+MHxifUYmrlCMjDgDGO6s+4Sn+bSdDiB1efhb5vHPEkEDIJsI06KLNasEPLI
4ckt4mvKewCfwPLDliel6Wul8AhKB4/TXKgdtbM76EYzVQmf69C590vExU9eEVG1vSn67Oax/MXa
GN6lNnitseM2ehV/4eHI9tT9omI2xihBYV/JrK3YRu/VrAEPBs/2qkk01WJGMQ1weMuFgnOe2mDG
mnoKtlZ8cKCsfrJatIH2J7OhHRrJSCC1Fi/AOlZ5XJQr6iTPAt3pgYLsMstlgG+hmjL9EnwTWoU8
1d8maMlVfXrK1eUn0AK1iORsYPHcU0sX+8xuLKAKmB5w4ZxoaLeup/jT2HF+97zp1rfLA0a2mjE0
iPGpxGwGcW6Vp+ma9Me+Ske5AHn4ChUEJxclzAyaZBUdOhKOK35YjhuMTehe2X+9rjeXILuQ0Q3T
EkUlAoWmrKaUQYxwq2pnxrosd+FqqYq6aoTkv/DWI0/a8Oy5e2mW5s1igEENtq+hQvg9Ngeu40kF
HeV9yU5DAKd6BuLW23KUQ4HnoWWS1Ez5T5xBiNVwM/FnTzI00Q8VqwdTDxrJMLdha+OBSmBF6R20
gYry4hSmBPCiGirUb3447BOk0XUf7/Ox317FFOBCZnhkJP61Thq+AMk1IDbX716vWGY1pMLWH2a1
gEimTlb8nnvDLx4Ly/5AqqshnPNGXDCqJflBJEGoa2Hp2KCdwh46jzDL7JkOZl5hrA0ZmyONu40z
23JK45UFRQxIF+iv+cbQr8gZiI0gtcqWFC/YFMC4slGSx66WbDIL1LIA2rRq5rrObgXXlGpyLezM
ZYWW5N7sBTuGO1UzVpTLpmzK0pEkP6IU0//woNszPvg/DYmSNEQHUztJM3miv6uqtn5MFVtgODfc
PEbGeeInRYv9QcbUu7/ip7fwdRYX4EIDrn4vPU+7yMzVtfUmKhioVsstFtn4WGLdwLovpFQFnm9e
t6YXMtP8xjZDrzWCG/g+ZgQ42CkVa5LX1h6AXxQYpY6h5UbtLu0mEE8u98ltrFvPtC9wVkmZBSHf
nlP+JXyGG+LUdGMJsqF7wnKLa2hogJ0ZJjGODE8a1PBUYu8NDMzedBzi8WoaHl6jIJUNrFUC5quC
QUZnlHH3DGPFhAlJKFpFxSmZhY1d9Q6hAC9JiAxSaRTWFi0gEEto8mm1B2YJGF5+b75qm+8sHfGY
4k9wE2Xh9jHNcme9TNOitZZVmQ9VOW7eDuQf1MVWxYvcD8XGTmXcgrFZHVUUKYGvrjp0WRpduBvU
Omv5ocSlv1ytbJ9KO9hDRNzMEMbF2juT3edHFmZaJFloAXAdIIntOCMxhQBWXd/nOW+/dNt8McII
K4efjnxzZmqyJcHumVCZzzHOvj/AeTBBWT4aJx2QE1Azel9YetWcsSd8sLOrUNWridMC2L0JKgEC
h6NTz+mzja7EZF11yjQ5Uve54ig0m0v/QtvWcZVE/+W8pi6ICpUvVTg7hWL2hwns/xvIglfrWO9/
+jwr4/NvOP1qcPyWnbfQVqXtqQO4g1+YsztNEsW3aZvgWUZxy1xtXU4t0yAFih7Q2AMmylMog4G1
e4NFJFaH+94X5luCFqz8iWX75+Fp0PI4m/wOvoHxGsKi5b0R5aKsS3sTvDxzS1AEC6mtHnrJwtfz
6nVzwZSWvayQqD90oCUk3t+vM5isGBhMYvHTTEqKdABopSPg7Q8dv4JkVvDbBWQRGKF/f2mD+MNr
GJo7HlIjR5HI4e/Vojv9KRFvqf75MeW3LCwtOSMlQ1rmffkoWCtXZjv1YCWjwMDYGdRPCZBNkVht
jWlPt7fQmPXE8JHFBXFS14Bdrm3ZTv671C9gnf98ItkaHnrk/UwKOD/TMF4GCS8MN1M/RBepR7M7
sT0tr7dvcN0s2lKDt8Lj6LI0omNg48fm5TnVGTbWZpwwKUmx1dEiUhHXCC9YU3Eu6H1z3oHYE/U9
NeQeTClCQXdTC9IgvXdxRbDXqqvjNBISK1cjAWIxa5Q5nqqiVOhZtSD37uYjkKTiFH6NHPGwyxZe
XqEg28gRCGYF0DZyBItw7dVx2zH1s3VTPrWiHyjTMKNhxGma4iUllMBO7r/FlkCDoSUGpEDhmnBX
c453Bfs5MV8R43WNX15tCdtocOqGQL+K5GAruo4epL8ZSfM8fPvhGyuel479aWpdTNrPZPJwMTvj
5bwzXfJ7xI3DoqRsntsCQq3BLQJjFh3n+JGf6w24+hvT057u16nFvBZx/AavEfHwDvG6HHp0V+ZJ
HMxdo2hZVg0RQgN6T5tp3mLE+/rNtJXtL1lM5GUWPLACvZsugjJ8Kl4tT5kVnatSphr3MKFBKU7m
p0tXgFy/2YRJOooH7OWHWMADLX/ETX2lOqBnT/VoFdFz6OOWF2RwSMyInTbasELohTCFEIat7FTt
vUpea8bmxG26i8Q0exJOm/upF9yAeXT9GsocayCwXLnc/z4kK1nrw+bV7BeBevpopL9y8vEl44u0
FpZRutL3SQgQSlB3zKMhUQfN99aWa5hgKmkruMv3C5otr8J36SjcoO/J6DaKWe+NguS82JKpI63B
SrWaNOFn4x30oRuXbl+Cg4H7BJ2AA9x73mPMdAueTeXXC1rVlAllix+uU40exxq/qFEZSTi+uEN1
INU+YEOZ0tuFnKLWCsIMCFZyOVMkFb8oMJylnuF5FUKFQdxn1c3PUhwG/O+bzFHTUzY22D3qBrf2
dy0lnbnG4l5DGwP7MHpnvcSClNWeQp6NMiJTbOawdL2ryLm/wCHaNkaBnGxG/UAmQfqNEKBHlJ1L
aUBjVeggz3wYAFDppEdxg9Cle+y4i3u5BYZUf4ZYmWLiCFRP/R051SBOyD2/Idm9a7L5OMZEepRs
AstvFfhTAH4kQNu82qSA3D14vsft53slRcxSvOS6TMzbEx3hMqTShpolSLw6inS9SR4mChTqdhoo
K3uLLPQdjS7TUEIpeLRXUNJ9E2aW7Bq/U+l8M8PYPUttEPp/it/2yU9J9h/mKfkvrfzOh9ZUIOgO
XCtXVZu/MmVkJEAR0XySTnMpjl0zT68/RBHG/9qDHM3QDQXJA4wXcYM0tF6CYqsFg7NsDnh3ebxT
y2+usGZ31J0Ik//7erLDNtUYdRwmUPL9U/hY9bEXf4Oa4hLNO+seWD6YsW8C1ATAbbBYhy4D/b3S
LJiCpZjPnMOP/XETZf6UEdx6lsdjY92RUzMcuHyxi0Dzc/TqE1oD23PPm+iaZgYuY7nQ7fjDQ1cg
sgIiKhrfWnbzWSiScEgdYHRtvCulF10DqzhzwiQZLbQcH9W7pqJ2AKFpPHtkuWl3EqIYI4y8XNAn
xMuBWbnFclbMM2QHLOgyIRcqZ813+Z+U0zOCHslIkpv+YJRNwjcYPPMQ72TUQlpaZxeSpJUGSOdI
V6IGYsfJMq8Y7J1jx/kuGTdkBPJmrlO9LCOocbccGk9JoLWHZCbahhXAkTvVlXzXhgG7DaQGxG9X
vghfYFFFPBfEARPnE80xBdrE7v+TqTiQWCuTiKRj1VFkG5wayV8BtQEfChT7lQJXo3nUCZCv0isU
5gOUhO0mwBxb4HEX7uYkqJCuZ3q1U0YdWEZKxpIJXXi0e0dpOeyzcTbA/5SDuPfhe800EhbhsN5t
Jibh6atENZTpZP88+o7h/bOtnuNJN6U3PdF450CJM2EVkttNaZ5D7YZZAyJBm3/vyKMuvUz4Ko4z
Wz0J4czINfE+/QcjJ6t3biXwcg5w293HfkQCvVFC3x8OTOIOs2bi0oL13NC8hXjO4vsPKHZnnrcz
SZ3rJd1N7FwUfEidzABBoU1rsXZgIXB43uft87T0XyKZKSs6quKRUyZUyK8m/vrf9QwmOB3wMYxq
3nBZQq/EZIKquRsis9GI2sAaudnQOr8t046vUUzUVETs5O1wLf46coQtHmFQXK+RjXWjI3I4+5rh
w0TXiKdBCczuE/kgP62eesIhmKzTKj11n8VBsbuPSKSPiNSbz2j+tYUGbMhxob4as5fPrujgNVPx
8+w5kuvMvaQ+A7uehzLEei/fDL9Sxj+oLCT60pbvGmj7qJ1u0DQX6C3IlfIXk5z+9TP1hQz0+Hor
DxYuwUHvTeuHlR1W7wIAFjqDS0xEkugxkeHfvxEFMBgc4eSWtF7ViOkGwFqGK7AqTDEwYqqNHVuv
KYmUrH3t1DfxY9PtEfgJtC1PFRymC0qIaIAwvLFzkjBP/G+RFvQOeKk9dElL3/wVjSOpzyiOgoQ7
HjbmoYFLN90j8UT3oPghjmVpP1oSRbgSnlc/vqC3vww+CJydtYvrDtetTIw3flHcaW0PoobrYOeW
6AUBoZU64qjbuf26RjM4s0RqUblwspUlFcLpjLnTtaAJ9uFBhGX5EgraiOs6L9nnHl8cWcuCuAy/
9Nv59caF+c7IgJk+6P0uqnIxyHEVhLCf6wLCydkSxYnjo0T7Y9+lRnOZS0sP2QO94ug1Yj8PXct6
kt94n5JzGTqGgckC5z/zunEdxYuRgwTzUSrHxr9LZldQhSzX0hgnHhmgDXWllNZZLOkbcd6N2w5d
a1jGrDvxcbZyPEuC4hY9xv11Tf23/Ry6+uSqG/EVIqiPLFGz2jzRqE75Xm6/Ix5EohnRfTah65JO
NriB4c777joW/sU0sUEV1Q3YemKj/0uhAb51CcUZJYg3pk1ERJX1V+V8ksU4qCmNv4+Hv6pJw02l
MFY7Mo67fcrsrdgc9iRZRmlaiAaiA2FyY/w4JOlGaagLJh4RH1Z3VmXdMtJC/Ix6tmILDMkDjOtN
fQlI6OCg8MRjsq4l1nKLYzAbRTVJMToxsNVblMwy+xjhJ1d7ZtyEC/lGa6qBj/gvDOo7MiT0z3Rx
pWXRkWJT7PdmQlrYQVwRyDcVN9icNxGkYs4h0ycPPIzygnAQlN643+Pqbu9AqTuPntpWRjc7EIGk
iIOzJWcLlhOOqTAZd6B1zfJb1DU7YnWlSNVtVN+SlSM/aMziP/QgoGbm0wbIDJdguNJCUhvWYGe/
M3Fq3WRVGu6PUctmZKQj0IbDze9ojmtrXTPL5Yk+9vDi2ZskEDQqTKj61S6i07vZRlq6a734t0z9
hFi/EWjZK7wTy8O04ayyYDcW2IyzkmlkmQMOK2lix2COl+4axIc/1Hum36R8Q6p7bC+CK4wl351u
gbKkk+wVKlj/wQXBQpLnMilTcYON865IHiOOcVrkVLTC2Tn0mmyQbjPJwE18deoZCg2vuAgXTykv
mBWWJouuKbjmRMTbTae+ULAVuCU3eyzmnhDzllc3JgoIhjKL/13K5B89NPurq8kkIPejxQV95nQP
sd1k4DF5WOkBBF4Nep4QmZjPlG1rjjoVxNJxJJZQnSWaNcScpg+4hsV2adzQN65vckAg7C24uhSo
P82HZ4yy7BD/OtK+FrutvqMZ9yJ+eFo56EROfK1vCqufuwafynPEveXi2afPo1A3yuPpirSFQBXR
zX9LWt7BG38TV6luEMuqzOJn1lB8snaX9gqikkwNGX7J3IotlJ/I5MQ212xqJBzrtuo24aelvqAp
WQ3oZpZemj57y3zTdeGOt9DLAfrjbHsQKsPmNQDATUY8T5Bca0TKmPpdPqLQtZeueAwr0EI8OeEy
24CHLX7bgHLZs07EheTEDTLEEW/x0WZ+NgmTEdrUAeIJPMXooqypn2bWfhHTmkktPpaMvJfyk53+
pn4WJGSTfZ00Yc62fhDOMaDOSaXcKGPexlxQn83xXOuMS44AEbGWKj+uVxTtDD9PjaEC15M9dMgb
v0ipHe+oRZMXR/1hIcpbpwtPYC9UCWblxjycXG+Sq+sLUngFR5MnIOxt8a0vL9z12KqzyZYJikMX
MHywMu6ABgAHXYdD1FMIGwFmPxvuZr2mLM++I+GfyRaOq7V6uVOOkumlyUQLBDH8CNOjekTpDMPg
Ka2Bk8VGywsoUtIU+USIq09EaE2WODOm/1JWrB10w1oFlFINf1VzWmKMXijcBG7Gn4utMTwSyEvF
ZIgaiTTm/11H9flKxo8jj19QZxdsQGnn7rezVefK9NWNaxXhuqCKkE4YlYqjjtqSme/4z28ksd0X
Ie0eOkLnk8ggVAk4oTMVO8/Pa06e891C1QlsvLqHM57H/KRBnBvqph5YHUbuB8h//pdc7qR8FvIm
9n3E2T+X0ihFB6knfAI6cKU3VZ6N/t2EbdulMhluBbWRoiboJoddKZ069nMrk+JOr1+Hc95LlQvd
IhtIZJ++SczSU+1cUlyz3utNZz+qLT6WmQSNlHQVCfAo3kvv3ki6qs+/i2UMJFdj9ynLR7abSo9l
z16LUIUeFmh3xKkfXTpuxP+y8uUxi4LU6DWvHu+dr13PPgzoWIEUYd1BPWMMwocyyyS64BrwHDu6
4fR8mJ7bJyudKlJG8Mq8yIOiqKbdu4nWQAadZey+NEHMYB3TWuFWUDz9awXD3AeJFyUxcxmzAG2u
joGscTXHf4cF1g5vuwFaNfLIriUt+gTj/e31UU5LmIUSTZSfZh+FGhX0uMrPfm06ZDM8PQwQIthd
8uA3aoJjjRVJv/224KFPHTO4x7CgSaGEPeBZw4hXxRHlOgiFldCJ8H9Tu8CatV3LnqRDTQpa7G3l
a5HZaYx02kkN5F2s36Os2E/gmo2wEXaXItl0pPSFwwdFRnKFJCFFkDdJSuwAFtE105uHINCvu7XN
m6mHXUuWoCQNLNiyBwyusV66Yanjtw4LPWoRA/Vmjhox0s9J/mjDNboXQrb8Cmvgdlq4qErwXost
uLvh/KAFobdW8OuLCiMW+x7k1RV/dagZLdTbCGu71RRR673GBFZ7AfAqyzvHdA5ikUJBlBW061M+
jC0Z8HSEZkCsNUWzQaeduELcPJiG9EFzInqqzu11C4sE0neLkZjXCp0eQcCm5XlUKDGvuyaojm6Q
bAqkPqsIusFiE7R0vzlkUkJU547o2VwQ19NVu1WFSeY0yu9+esamTwS2sllENTGg2QX8pmcLgZjR
rBnsBNAn5eYihigb61uW+zR5+6Lf0hf5Y1I3XU7epiMw86mK4mcxina025WEwtRXvqabvl0G27LV
PNSRaPfKnPv4MjhyFscbeABrbVQiSwKB6+xOiSSbRgmM2zJOTXh8Zzw+LtkkQwJ2Jv46npeptam8
dE5kXug+YzlVMj6wozqz0Ho6bDczwjV+5q0y6IKC5ojq23JKt21zlftoPuBfGyz0OGjOidBTlwXS
ssibx4UvQMtLCfINE4sfyeXqoQtJfnZJVIRA2MiaZ+nafq+I9zc1kLbJMPSYdicezv+sWCYgey5z
LDC0Y2B2OkfFCL/D4z/hQUGPM1hTDp0k8jG4aJesnDuPnF2piCzwKMSP3pDniNlkG+lwLoAUFA08
r09tRA8xd0u/tcEoqGBmn//oz7UWJ/dfpxIDdxtvKEvj2YfQDEXWhMR695GzjHIOzphG0z0vrZfE
5M8r69F/B3GGnWeJTItQSoYskfrPDQpCwBfHnTnbIU1+EekHgwJ5Fs4uOV3A8zYGGX92lAR1hxiV
zEcN3GkOM9wDWxu5CFc/m4xScYuLGzDQIU1B2OqW1zfLsR5ARz77OPUyqgZLfxIezMidgiAA1jFe
qSadTfNOQJSGP3mIW0XMiSzeNk8KaYDOK0QVJl4km2AQmDikJ0FLPS3UNbivBP7m6KtqPjpwKUuM
/fdqEj+Mg19V/uae6nmGzFoAemO4yuw0JKdZSDX8OcY1UEdO09T3liHX95yIM6UGt5+QFOut3phI
bv0mStUmBEAixUYGCzZq2uv79B8HubY0Ul0qFfknI/88Z1ZxcmN67ROx1tOZtI8Nip+hgWAHkXVX
Io7UEbyRk75yxUE2KNELKO7zAFKt2mZ/mRf1p/el4A31U0VP1bajJtTrr8Na7t8mQjTs1c4Jh4yW
QBIDrE+O4/Vw56oiw33aw1suL3dp+RCjK/awNkdw4sEmvz7DKvHTo/aDm8/lEz6U/pcJ+68olDJm
5tTzhP59G+eSRQAhn9r74rubcwHIU6Ursf9chuUf+Kx8gR7PfKfDG0p3ODa/qNJGovz7yWIu2ssO
W2pZatDlmaZNUORi47eVkxOG+7QbkqUjpp/zW9Zr6HSj7FaVftu6cNk8yNS5PhbJtzEHV7UKOXVH
KZefI6QDis77GfoQGThOd0+MMHVFgWR+oSlT6hGSKrAqbHCywBVYCSdd++8b6T+MF8SiR/SEP5v1
PcezrIAb181AtdtllpTAd65EjAU+r1bPw+th4lU4DgCkUL9p7ZO63ZQg7CjDTRdUtzCosJbnMKFP
xwUCYUB3A6hbLovNMEOMPRdi3okXVQ502GhpOLnsm3S+8DxZZfVqvCL/5n2lQv5wlp1WCE6z3Kff
yL/41+yFirED2ClEI9ZRwr+ShTzIKgCiUJqGkw9m4JcbjCiUDyS77AWq7BAJCqLFu9BW911T/Tie
RHnWSVEFoDrzqi9DKLWzq8mQK2lOuyShH3ybN7C2ZbyHIK/TTh/1EjGPreRxnpClNHmu8texzOhc
NmXGl9pZevjHTXQ0q1TJrEmzuQnBM91d088TI2rCpVQDusv7qsamksJl0RPfg14vy4ES2Nptr3X7
65C6eaKzEup/UgMfy7K8x372YDz4aWlF3/STv5IxLcP//y1c+1JVH/UzALYrlNVtxv40ONqpu9lR
Fv2RimxKkLduyAzdp8S2+q0zl+woT0P9Y+QC5hPCOXoPL11qswo5EtYbYUV6ny94YrrTJtlq8gYZ
I3QJ0PsGCVUDQtDcd44EGVGl/Lzu6zzgBkm08DITnTEFri/Ke50dptHeJwhKlS/pw5MkHBO9ayvd
0MHsEY75qYdbYDp9ruFZoxhK2IN5Cc8ZTubjM4DXx8HoiRKkGKrE7prIFtSnkY79RdPcwzWKmdLb
n65DR+vAoo4aV9jZxRl8fmwJukWjISEtJ/n6P02py85+vcXi6dtOVFJZ7iy9bYeQmhLZTQOEGpRu
SHSpTjLxA3dOdHLy6bsicXgDUPYp10ENCm6Zws6UNo+/1QAn5W+nRmIoZgPiBUCLKhdwSgkxwPpO
aU6ELl8fnofW5sk4PEeb6ZRWUH+PXjlJVwoB6M392j60M0ACgJvcOJIiHFY8ag2gqKN7Ftp3D7KO
aFuY/xF7qTceDo0R2JwJCIk8t4DSvURPkL1R2oXziBCUgFZN67RJFxxzKFgAvsv+hdjfWu15FqiV
2BGENmTMYfeivnTYkaYNYsI+MBQ6XCz2jKNXXSIcYQjWP5VUzi23ndc9JcKV10RITsfciH9GfZcG
+8tXNuGUfEkbfpMKdX6yiHadsTK11DIf4dIDnVdaOYz1q6eLqyotWhrr8fViRoWWr4bhdschPqt2
IFaldtpjIQlu/U2sjLoVmGHhFIUBhzJIY3S/K5cuJMM/BUXmrcGFF9BkKNdObKTPxEGrPkdP9lD/
U7xCS83U4oKRQToLoKQWk/VTsHriclPl0eDl2vldfEKRP0VeuvuwSTJNL2zJEgr/Ks9/0GRqtK04
Zs8kDH/4Ia4H2oS9m4v0JNghDKSI73UrgrqSC4gKZIp4QHzWJ1Uh6aWRuYxrPv0WqboJUf9X8QX9
YpwNX6fVeX2YMjSgZrZ8hpzX88HNaxI7AGmvMqPi64WbFPVHJojBmBo2vsZhtbJkj5Uxa8XcmGSP
E+4rpGxR402VdX9C84Ah83mqmL0x7zSxvpxlWYyT6n/txY3q3j/HEoX/iguVF4fcyFLe3TXSnn9d
yNR4SQXyZJSuDTlToTet9sLCas07Hc9QHtQ/cqUNRnnMAIo9e5jkPhgE/x6gnbuqGjeYi2qGStTE
uch880cXym3MAhhE2YnJNWbs0k+wQvS54nL1SLuaxwk4EoNcQOaw3T7ttDrs0mBoegyqB5z/t4cE
LS4eHgGYd2r2BNGBgHr7q9s7dhrZZEAhqXIutApxbS9wpwAvdRDGTUVzaULCtz5+552Rod6+eGwJ
BciLLsfwdKuXBcGBr28RIhmhVIoeSpBycMRpr1ARms+xKCLT1RXTyqa3pMi8t0I6y7+H9pPJOuln
Iga3n59S5p61ki3dz6GnNP0Ak57+keGVL+1iVNYoFuTLvO27/cTT6qkaVabiTHNB44pCuMk1jiSp
/nmBMb32LC26DUtPGBb4frc/lGGLdje5kYtlWjM8yKOrllYq014W3C2BOecYaTLfhUMsQtWXTFkP
tbg+UEi+8FAYVFk4EXt06alQV7UFbUz1kRwtwM+U2piQtg8WBNcLYbU0kiEi8FgYnsNfIU7SlOmg
LJvcIfVNPx0PSws/habTErqnvRv4pYLYfqpOhgWQdgNJHI9CTTYyEpffUpym8T/kTvV5uPCWMbkt
mbGyBLMgTmMpvV37MXsuk+Jc3G3DnxOvE1mKJbb812YSz2q9bNi3/PEZFI3GzsNz2dR/3A78zof0
xdptjgvedJQpDvywL0O7GxMPGlAoc+DxGwrtWQPG51+zdkNRl5r7HRo94zOE/N6GgGBsHkoatUIA
qKmZEK068HkMMQeMnoMFEOYw0cm3Thgu5T8rO4beNJ504NaFaH30ygPP3EfgOk54EkbwVhYU1AKZ
CbL3oyesctRwGEOF2Fs8yjSzvCO2wwXHdGqDKEmgVn0XiDc+DnEBUxDGjcPmuzUgYAbx11Li+KTC
kJ/mzelQXi37sRDccxkqlUR3n1rwGWgva4S9wMssBaRaP9SpTxNVxVpw2LpAw32kKabwfPIj6QvN
SL8JaSu34VGti2yslM/lsOJzS89p67YOBbJXQzU42q4xiwpbkyjjSGc0OR/iHaCl5HUBZTbQS4H1
afZksuv/IacfQ4hsi4PyHTrt0Qj0Mz2QTgjFjNcm8ztruQX+K9FJ0BRTnj1uXCxIM9eqcwNNdo9M
kZQf46ZIjngEb5gZv3hyI9xM5yLTYDRBVJC8tzQZ+2x5rVkDME0+Zku6gCABHxFv0kYiBP8Lvvll
TtFMsrQ4YhbKJ9oTC0QcNofG9X0RziMWs6Av5sq31oE+W+bfWQDXktgXfjFG4hB4gfZILfpNUyoZ
IPOTqz6QSPtLV+U6SZtDZn46N2X0GKrcT9MfYK5yaUzWcbiHs+GhSQPehQHpQydaGACD27GHmfwi
wXCzcI6rCfF48lVlIE7u8ndqelyrH+swGTbG8lidTcvIrUyyg1U+AMV1qoi4BrTPkd/vyV+JNIGL
9fPYZqlpGSrzkxMRD7mN8kmJQX1gj8m404o3OBxHc2z2HmVoolblKA+MTRHgkojX5SOq9BGmDWxJ
DAXZT46CPi+0PrNLuGWYkxhjk1ImE+9Hkwj5UGREht/6/+JQdTN1QpnCM/vcVZrVJf35CDqHKb9g
JKtyMTOV6YLRt7dsoOjGix2L/V0ebTs0J7cL02CE4U2Czb9EeWnTObFK/Eybx6D+1wvKy+80o/IU
YZYnUELSDSKjiQ5iB7TXwKZMesu7Q7QEYcq1NdF2nJOEoBHBjGMMQkjp0vL0r4h8LZICLJQGrCMi
q6r3InHvks+kqT11HNXYxMS4F9ecGGBIEB24HvsQiQ2TCXE6RRlPs4jnAtEdMCQlDs27V7h+fbvD
KIvpgAKBFp7uGxge0X/WyfNNBCqUTN+bfVGghzF8yhMdoXg4SyoYQ5j/U+6Z8jEVFKxu1HKiIQLE
7xzA0l1LlT0QBkqWATfZ1g3mkv+4jeKC3m+VNOlJIfTqjAsNE2PWlS7ow4wJyuPk2g9se2SDX8h2
5A0nRQ8GWv+B2LoaVu2z9aSAdVGXgUo/bH9Uwxxm3qElHAAZKUXxay9uA1Xqio+BH6MLfkkj0PZR
bGOl+x0yk9hOu93tL3NU3yfzTfFojt5wnzjw7KRdGFrfLZt2US6HYRlwiQ7CHcBt5qfFo4AN8l6U
UCKorrd18xRmqnA3sXYB0IIsrdXWwiQedodb593fsrjwNEKoE89qfDK8rDlbrgmaouBVJp0Ze196
/3Of1xtasWOO+TdZKhJWKSScgfXp7/NJSYW3Ca/e0qAvtH84wA5Rhf8Yfj1FggBDuZglML6MU3zW
c+XVT5LrI78BOvj3f13SO+oC9um7Cw6f8Hityx2v1/06ynBetCW2sAJkeauIbXuZkXKtFGt2o2si
pIxBkUEd/Q5iLl3aK52qfD57dgfAkECxQrZmDSkavY3MSCsd49X98C+TTiDUelRhbPRL6miscp+k
sSv8Hy7oYDNCJClTx+CuGxSe6qxnP/MTbmlZZQ3+vgiM4m44jkNGRcn16f3Nkxc8NAAMlEFEyzdr
o2fP7oyYiYUOhFYBHkzen+Gt2pR7C1XCqrqWUNyvLdI0r1NBNUynsnTF5wJhSnltoI3AIQmQT9Jk
P7Uetjm/ubFD+9hzr7ceMnEYK7yXl79uk2/c3L6mo0SKQSqWRzzuOPlyEYiZdbi2cj7rwKAfBGOR
50cVquR4wZF1beolGvyuESOh7AhUE0l0J1sLYTqagbX1tPg3f0ooQwmHSW9WfZmAcflujDjKDDkl
5pp4+EEiaxqcpQnQpBCYGaSoIl90J+fs+QklXY8rUPy1RqAfzPSv6CEL2/ei2hh1v3PGx3j0dGrD
9D1920ck9615Trr/wgfcFiJAijQ+1opLod0p+mT9cqPbu9k4hY3Mf5R5glKy5jBBZrdVfUy8r0Qy
oip7tTAP81xcdcCgJQn6OfTkWMp2pmn8qaZjm88ocDgPtb+U2z/TRRKxHGXQPXslYSGKdOLyCbWX
9sNamEwXdzf5P2qyIlxo+QNmvlL6Tnckf13sI26VZPGDTGVnhRkXw0p0/uqvy9ptsacaYMVv0goa
O0dO/ADTUjMJNW2L9BHhkhwF2YUR9SCSG0qnohPZviWutBSkqRQkm4E5rHObajvvsdN/FJ8ysiGi
ccsjbtuB4xRsY3RFr7BwPeSs7ceFMeBgRSp6sPD2jOBjyzOfaICFRDXQCI0vpBCC+ZdgohV7nWIc
nR80ZyNDVF+yaMcy2ADFo2WZg9K/f+hdQmOIveNy8iO7s2VZzMda45vbePfpcEEpbYWal2Gs75Nn
cActKkQ43LpNK7AWq15bIhm01SDhWUgYYYbCO3QKNDFtfCBkBlXm49USb2P+FFxJqk0Yrgc1ljIN
bbiK5nIyhgLuCeaXSIHxvZujPTvgMFB9hbSi8hqw0kaMX1xigjHkD/zSKm9cy97pbvxLOqphTozE
rQ26Puh4Qzqlf9GKKYPhBP2rbRLRBTAiVMLvgflrLiUUbULndPodjYf/SgxelKNV/wbQzZ1oQfXx
JRHYrGHcZr4/2x3rSAsC0Pc6FsilnHgTv4HwlSTIwbJvNbbSvoauGDxM/LxFp85UH8sFvTJPHVSc
gk8nBOsNKr8Pz8x34/5Sj2oMynwTgtl4Xyhe8wsQ0eM4ZUW0AI0x6YzGPEJw/gOsxPHSg9MtDTe3
3ASZiQECuMn6lzW/IRaZfLThn+WQQHOTS/RurGTlM/6DCPFuEYpAAQB84PepCFvWtOrZH0qu38fv
vz5chZpABPltk1LbZ3o/C9g6N40Mq1oZ1gtxrWkYe3XFi1GeXPoQtqP6EXrMhuqmEuUpA0WKSGCb
wy1zx0OdHgClrLjAFXhS9yfNKEEfm1V94jTosqeCYAXeSq5LtBx9iL0LFyNfebvpoNt0cEQeT38b
LvSjF2+2jTbHJGW9uWPcw0nhz5CXut2wLGlX3BWUFTSw//carSozKt5h+Q6j6HC8D4Ego+9yYu7a
cDRGXjmaYi3rNIYEQoAev4o3xa7oRzB/27zFs5v947oJFuNX9J9ilwz0ULa5idWr6qeCNkQ+W2zq
N652fktwiu0tBMMirZ5eUC+oXrSGR47tRvINswqpGvCn+lDTdc3kzO3VeG5yXaqQcAAG6a//ITLh
+OlAL/Wf6Es5t397iKNCyDsVMpj+qTclJF8DCM3aeRVGxwVuHcs5u0blVR4/Thf7watXqvZkOi7X
dv9V+aSn2i/ZPojjptDwbPjMTA0ssXtE3i/HHUByoSycPBqGdFIgPUs3qzW69C0QOCQvbH/O51J3
MJgO78NVBlf0Nu2pgKEAy2+Q7ryQck1b799ZUBbmWBUAYV7s5M3C8jWXmZ0ZaZVB0sDxBZMY21ij
o+qrDx2JqQeIHVn7a7GS1FFesxzHwjAdQkV/O7+fiO2parea7cOdBHBD4JHaWColh1qk0vP/IzYY
5CGAc6CPxZl7/GQEb2CM5kwgL0MlEwrdkSZEXZ2fQlcO/VjfeRfBreHC2eAGUI/N+2E3olVeS3G+
hkh6uRznpa/FjVkH3qrM3rlcwFsuaaEajbrlTo4l6Gq6QX/SNxzMemPNScttji1RHoM8QO3DSX+l
uTrzaK+uM836X/M2PZJVXVAlpWM04879mMNn4ZWXY9B8BXeh9nSq+cKyl1bgZO8q0UoFHWvbyLxM
AcY734/ak8OsHIwUdiIR9UrzvfTILQ6TnryEa4awKnC5pUtMZhpY05PBTNXveH3jpvYT1j5OEO/8
10EukRbMd6Ck1d9hNwuapzB9x2xb+9onGmXDktFjKMWlGWX3kJaHfLgFizD7Q+783F4LcR1SrlR0
e2NVwgBurRpWVWVBgJ1T+PQbM5ZGF1tMTeBZRdK9m3GVYofwQUfvkY4RYHHko4mB29IUuf+TL/7D
3pl17C+0j//EfR9eHK3Fx4WE6W1Aw/87is+/xovxWdVQkUY17w2npW6XHocFW8Q61QTxGHgJUvKx
keQPMp18Gb7f3KRhjBNC+NTjBsKe7iGyynh2qdxL0L3LgsDts1fWS6VjvUbVd2ldq3hmf/OYvDWx
PCxRRe3JOWUyPFmm5g4ZAO5wvqvVQ2AnPtkMKKTCdPWcJYwNZUNXZvtJKHdrKe28wVmIwFzAlR2X
udVsddWYv0oo9rM4tjrp6nuw3OSQyBqWA6VkO5GmM1lvjZxov8sEmg1b/mXA9TXTdrh86sSeh17R
3cAltA67CaCtrajbVxQO+EOiugBlCgay4pG38B8jzYaOEXLfanCfNHIqc1JlJBhnpeMc04hcdpW7
YqZySlvNE1ie1+RZ7PUKwG6GnNfQKGP/IFLO6cl+EgPSAm/wUaczWSZ0GLov40nPk8lDwOipA+2g
zJ6xBfpF4E/XzwZKGL0vDwpBzxi4lNcA1onsHfP115xz25J+NUL494Hoi3ss1oaQUuEpaGVgmCFF
qZwNW8mzbfKdkrhzo9tRokGNRtTziKa/Pn/ISTpoB8Ahp4CgOKlQpeMRgoHWIXUpphQ0/Idkh0iz
3rOkDSRvI7vHzkvCQjgEHNqtBteXxfXIBRVfVkf4hTruqyCHg8GRAHkWHbLxNk+GE5+iP4+AD0sw
GJ3n5NWKLg6GWdxQLm80dwq86WvOCwFDuTWpnSBvzJi8xh01sxk9pCA5ifyDalecR9YfTmVydn+8
yGZMBDjaPJ9vHo8HJGVd21Jsft8VjJkHzvh0w/QIMncg1U9eJuPreV/y5KfKwHD22elcKO6Yls8r
hm3K/2gHe58JYMD7dk+CTQd2/24XzhDr41cGyKq4LDHPRZDWiCsHaL6ljj8CiXyYi+k47Blmbyt/
77gYz7jppJRM3RTveczKCITNCNNdki4SQn4/ROf3tZFTw1qRzLZD5Cnmn6t3hZ9kpIgT2XPVLt6/
y5st9FJ0GDBxSBC3lsar3d2UCxajPFpjBOBXWW9U+hCn+2gqs+r2vBgEffPl5/QzT1dm9vUrzD1D
rT75OdvV0MekHFcYQLq8z+RiiDznI3+/bnxYocImdI0SN8AOYG6QbA4swsswqrJ+IA9DpjsWH06u
hiIq7H1i/1CLwMcNbID+mHICZXcnFe4hSDe5mIuIwC3/MU9mo15M5Wybr4iFi8aYko1wbe0iD4Hg
KhPNk8nJJcv62SlYP8AYmuAvNSN3jbyNA6byayob632n5n9NXaXDLECwjWqpEeJQMOTMB/qkRFcu
Hfl4yPgApnWAE5DkJIj4zAO/azKaTvL/DuhbGhQIqxVWYTAG5lDC6zY6q2G5icElMbAaF3N2M+7h
ztVTIsDRnVwexGXQg76QzTIAurFgWCmTZknBP224YerjmRQjeYL/OWsGLWkumKeFBZswbA+ybtET
xKBxYFmfhg/p/W7ojG0yTnb/StxHZxFYfE6nkJd3VPSfX9vF7bsTUTcvnzjweuuhWFQm4FEPMW6t
icMLr0l3xr1NDUr5ikXO9dRD9d6VABxlmcXT2jZWDdAipj1J+rvH9xodHflROpBuA1OYSux6Trnm
ft0z0O5bkd4bUAjzaFpZYqXPoczXdr8tajcSznVG0Fmn9JCKZYUftP1vpQFXr4iwkhrlSmQFb/fX
8B4VlnNSUEKhX1SrpVhcWo97z4OXItMGdqb9H7+PMSnS5ScPUj/qh1Mqks2kk9oSMNuBf0/gZomE
adhZfR+OS5iJ/L5vy2dCPzPjlnqs9Zp24pAd0faixck7R6AcT1YBxjjIH1or8ObkhwLtG+yCQ0us
Cp9my/0OmhfZI/YkA3tCmldyXsveRxqZT3Y3aSuWEMzFp6QpFehfuNiW5JQNemmmPR0e3tV/FbWz
cN7GwoX6fDTo/6yEq6pNZ7O6eMPVbu4vE4ILMZm60ldHvb35LGBCv/wTs2H3ZsGeRonO2u6z/VjR
x4KcA43Gjz1lG4S8Pkc1KO4PELO/ozJKijNhHYSt1o1SmZjctVN8zcjiyBZxOiP/wNB4hthpjUs2
6yGi4xSTb1GKtLveebSbxORFg1e5uE9UB7AgLpJaaFSrVZuwrSv4nZp7kpMkFGuppdRw71L57zD6
j3MPhlV25p/Q4cg1VZt+F6ML1fWaeRnB35bc3AxixTz5qmzQlVr9KceYJV9Jw7zvUhk9r1be4FuM
veilxur+im58d1x7PEhklhhw/WipkrSU5jCv4ACwI5eRKoWygq1vMI605d6WcOmturjc+CzvFo2S
QJbIwO1ugPC+jFqA+iWvu6ec5PcNfWjPugSi6fvlu66frteEHZstoS3T7xR8JK/yhC9FSLZVjRyy
3ICN15Uer0N1k1tMs6NKqgWIZVd/seIPGXyqRJnVqsmQUY8+KHbrlQkRPFM3dNFFLSCmbR+2hWFs
zaQ5sl8g27M19pgsCDnHYycxxd18hgXdH8tRrRFoDeUC2DlVmKuwNEA+zL7zX3jLdKZRilp7j7O8
vaHPU1Nc8PoC7f2AnTDOSQUisWSYDDsP0xoFWM9HIwmVOTGsYfjZszg6OjcpCxICk7yN3GLCrkL3
KxfWmwmRaybaWGUCrVsIa1QdKCXmsMi4S+LEpc8fso+pYW9tOGQKaIQ8UzHutbrqHOhTwoXZKrHx
deaRmqty5mJssWiB1WH/tR8f4Zurhts5yYLmr5ahLKEo09/NTvVD86UZUcEHtEHnzqlpmBoHXuAm
O0bSIe6LWm/+7g8tV5MEF4EjeYkPHs8FmQqkBMQyeRChy5EytujpOoN+Hv61TUu4lPJnnWp7x6qi
nhLB/5CbiZt2xbQyHK8edf5Mv4nXUzR+bivMOQA0uJ74F7xmMqA6IiPf69OukSGWfLxJK4LhSFSa
EylgBZhC5HQGkRB0OfP8IVq/7Sf5TpEOCwt0h5D6oPYh0Okl/2Nuq9DQn32tDZ4bOELy8WLF/VVE
wQfwkgH9Nrf5c2RxwOoVd+cEvFzt5mwCB3JvA80sQzC9Q7kc0oVXxXuM9Oz/g5HzYhK/jlPf0Nso
ShInqtRMShvQyTExfAZ/0VmHo8H+txM83qc7NYhdSKUG9xiylyuDZOc+rDSscEZ2u5tpW9g3GIW8
yDwldLfiTBHBsSDi/N/eLG4kiSczoCzucxHnoU2Dt9p1Q1lYowZ/Thkicv29FiL6jhB2TYiQFtFf
N4nBF5XToZN3zvxuRxyrwubhIlJwPVk5cCgu0DbB0O31ef7tFDS1AMOBuxHabVtLeQSAjnTqX8Kj
iD5DjRgwgLrbO3UOW25WSm0yYoWrZSLkz92EyvL2Z8KxhuLwFf2hW8YKRjxfIoec3zljnlDvxNyo
DPiagb/u3KZiB2XxcdMhAqix4ROlZTYo1snzKBHgCRq1sAPUacW8KPhtKZ0YDansyRsq/cz+m6eY
Aoeul55ykQHPs2UWB2b2ATqS/JabmhtfUM3PHgRWO2nsajvtx+IbUUSnebz7b54McmD/cjiCbORy
DINi+nqv35MhSwIdTdl3UHk6y2fx2Y61VNcewcjABumFeU9c1JO129wZNpHaxDMinfJp/ahnjleF
CbFIahMsjzd5Q1SMnziBrVj6XDL9/Q79lacE9vBGNJAPMTxtBMGrxCYbdOJB4MHexthowrHHYAyi
ZGprW4ULEATKQXnf0IwajYYgeI0zVEsfX0yeGu4sZr9LswUi2hF3aqYEhz2jvlsekqSmtIVJnER8
GA7Glr/jlgcMA+EuuuMSIRl03KBzCKziXKaIK2llkWxUvu8xYmHSmDF4GbZAIdyFAPvKyejoJVRl
cRYVwUaVHn3Zd7a8nsOcR0fWzvy1E8jEJT7QpM+E/xBJ/bcBa4hGB5CgxOriPvaJyn17YcVgKyUq
7ja11/qYTH/naDu49ec75Z6o6JZ0RQm4p9Zx8UxU64/ljgd71YwmWArgmvcvxfculgiIj4hzSqCc
Ho7CQoPknBQTnOsnnn/LBZqPTcahLEB2/gckHRhkKF0muimoevWBVlxIs+iRBBN3BQEC/cp/alzb
shv7SnnzRZzbDfqsTgqhuafTARj8ftxXjRKnETG0BFwKEk9sYfkuqCQEgxnsNVlp6FIWN6MfM3uW
rVfDRRw/Ako5hAUt1+FHmD3A83VXs3yDw3lQh0Xo14KiSxYjaKm6NAG+uHEEAk/fbY2NPsMB3bTv
oOvbzDkL1dvG2l5uFku1UlHkJg+4pxfnw6zu51dD8P+Ma1gjjNe/ruEPhAkZ0wQKbWwM9J0kAGDR
+GdTcATPhB3BCGj8I2gNW2caZEBo9HfI7xOP8Ih1imCk5eLeCWvUGjtjPdPkrAPizxBYkCMHevXF
p0puZlfCQ+sIHc11QmUd2CBzTmcQ+MyM1pQvI3gYJrdWY/VBLRVruwvXQ0d3Y9kwu36vqPUnXiOj
kpu7Q6g9toHAuOhOiq+M8NVTZnkjjAAx70m9AGT0B5Tl+v7n3t78WgIOvbdit+O9WWOX0/xXWviS
rwCDOm4j75zBbL5F30RXRNHUxfiv3X0ZtCm+qNWIUkio2p+4FGud6Ob6LdQ0mdd2YabbiPK8pN8R
4l6Ei2kHjd5nNeI9PnYrn41q2TMnQLR1LX+uZ0sYOetv1sLYI5FR14nibSMxOBBVAaDqceXe9soJ
lxA2g3WhOtBhMA/zBLWT2Sx7t7zNTHiGapJkPIZSTp/yh1krjv2zGfa29IExuBjp2/Ly3pdOalP9
trePfAeunKCLDzgPVHXd0ZdQgcyIRBgMDAYcKDauK1yMQrI6WDhoNea3tO4yvyFouidRej2HSL31
WOu6HM29S7logYXZumksqsxIbDPTAmqCOMcXwp9butj7ikx8yOWOCJBr9hZMYnowjIzXOenfE4JP
mOLmmg0QTqC4OWFAhBoK48vTlZ5O1IQLnCVlu0ffiNRhcodVhuGXJvQgC39XBs8iNob0KcGp/WWb
bfrhY3otz3qlYm8GnEQMzeJqpvcpuyWPZrSt1IjDKqZ2Cv6vwHH25OC8D6fgkgfz4eAwQQVyWwiJ
d2qMnQyxuF2AtALIneKjq28bNjdWnWz7AWBCt4S1jgASPyR0ezQNtOnLWh2hzUFPT+wLXaVTpdpZ
3lz1kIkxG4NubtEJ3YboQpY5o9lS6rDMLq3bEGW0fgpL+onL6BcGVP/bP4Rgs8V5K1hIkMQcVXML
QtCC+3muPiK7OBd7aG65wS92BUyiBSSJMIUsON0NlG12UDY8pIQEF0LN3YhdkQxCOOsosjRqLZn5
CLEPp+PDnWw0VERdK/7FZ8XefFRl2P9lcaz/5f68vYiapGHm9pNXlcDW/W5Yv6ZwFD2kVTTPkNMt
AObp8MhiVnF+lAK0CDhWjv75NqnnseA6cnRetdkc6VLUD3ZTNDf0D2J7Oc7CwG7hvUL/mkDlO9ov
hgmOSCFhGymPKGNeWKG0ubs7A4m/JEF1cLlcLEourh9Z9zf0OUuYQbQsAW+dh7xToOnJyAhc2Fqm
VdqxsQH9XtdfKWr5zGvmHP7psxMaeacoUM1631EAOKlIUJLUYWmQsqxEj3/8JHLMg2U/2TT6PrbO
lw4UOiiXpMIcVQruNW3XTgZLRxQmlOi8D8jYCeP0Lp7hlsj2/CKb2S1rOhCiWYmF0D/cd+hZ494Z
sHewBF7sOfonrL//e8OQogr6kiC4ow/M2UMGD3sHSME+EOdRevENQPKXmYJdpk1uoUTMBD3ajVW2
CaZ27pkzwypJAfIlsqEq7Jn/hW5GvqBHSGy4drAZddSaXpdgb3QZMFkKZB3ROSfK70/KSFPAWw8b
Ybb0r/QUYch7PUk0BY/ypS22yzwiI/6RwjmW1ROkll8p5jRpGerYmEb/D06jBJq5X0s/73InMw5T
153urQt7HMRltYT6kvOn5uI7atbjvrn95NHzzSC9y/0kXsDMc8Otrhr8QC62mOtuE7FHG3v3y06i
+AbNcQSyb0KzPx+o6duNrlDhousggWziTw8Lgd5expC91ZOEaWnSn07XkGukWLEpDEu15Xxwyy3g
mLDUCB2CWVttsnJXL3ztdN/dhz5cR/I2TgYiQGpQN2D39VEFsMhaSwCLLYDnFc38oRLieum7zd8a
oTcltJjdl0iGLDP9aYFijehXllV53rqqnstgAdB4okPtnRKr5ytVwImkVEySoKiY3caCXEzHtz9+
UTS5L3rl6VOzjfQOPxi/oR+l37VI84Zs6IxIz70Ah9kFTFToujrCcVMJktFhdS7ngIqJvwQPEAPX
31Bb09CC/seinA9ovQfw7j6nRScdd9ytVJPzdLffAIiAPNBJLL58KX6lycaLS2YI1t7icgSne4Hg
NVUlf3tdSeZFuMZ08R2HdqSvOaR8+gZJ5uW0GKxb2HkQUcaEi+kDcsqi+maFWFXg3qouH2NSv0Ra
88GBhAhkNTgzoe9HBFsfXFeW9urhCfoMH+qdao1WQos+WrrdrtFWmjrTGhgncN3G5s3r2aiTMeKw
J5MK0fTAqU7i0xfMvzNbP8TEEmOFOHNafZjpE9mxsG3x1wv2s1vf03sv1y5uyTMDYmpF0hnSu94T
GgkDZEoHuXU0sZnTaVgWB2k+dslbsdqOR5yuZ0XNAhg/bQzii3EsVX1NSAHgwbmRAPlfQ2z02bXC
A70lQRR0Qk5ZzFzW/P4NUdfnv5qTlc/+M95XG+nbfpfF+bd5YkZNW1PGmG+reJemsgLzesaY5lD2
EZvfHtxtsRni1KVEebsvSTDrz3qtkKQKTg0avajDX+wpTMgFScD22bWmATA3pdVwgL6HlvYqcg6Q
yCNk0Oz/vgPENMdXDnIb+ATN6HLR8DWl+8ViS7fSIlGcAnI68V7gODoxLu2tjpwpbGFVNtDpFQLZ
yZRivXeed9AFMF1F/RNIQ3XGprk7OSdbz3oiqxtVmHnQxT8JGr6aFGUw3Qf6C8yZHbNcJ0sT/o7n
SpFgLwNUnUBbF8Swh2+53LOCAnlfjzkM3HjPSUR0NoQN2cz+wHQgVCKq2nsGoJMObt484op/0/5C
dXivXxU48uG7BdOC06ksYFO1JE/z2ruYnxjAtqb5TG7F60zeRHwtfPT2070nL7ioXHHzVjkocpwa
ESde8UuC56cUJh4ZKroEYiHA+ifb07la/EMHZ0k7hnSefKQ992ucJ15rk8ismrPpvS/6QJMEBpJN
uS3qvan3D4quEX67tf157scCJmaAWMsggOA4WbIu6ZzIsaYH+WG+SWzB34AM6SlhtbiI8FUSOMOP
HT61IzlY0+SRj6wEmWXnRsPcv7byBrVE2n4/uUYxU4buhIVyOf8LjOPGo846DiNW+pNoELf2/HcC
z7SDVZIisLzRnGRAkynxWAjL/ZnDdxipu+y76GyTFvfLdFYSLARIrC19RyZz3kcAYzg0qzC9is+s
T7Z+7SA9ZxR9Ij6uuEY5oXU9/mAGg9b+i0hWdL1qZKRv12bWyz4U/6ygjGD+90r9oahmnSlx6pTP
LnEIEKXohmM78TALVHhSmLjmOziR/JgfRJhPO2jdOCx5Ucv0oH4Nf2IzYOn/Bk5J1nIfphi7Q4+p
WNX4EoU/3ldiQnQNr9H4OpJPZsnQPROZqp/gaOE8c32NIZ9XQDFWt3/kii16pNW6/fEsF2aBXisF
e9LWW74zw+YD+MJMQWNRqBAo/5CpUDzq9iJ767Hx6uAGinxTAMXAnthknUZiRiMZLI7BQeLTsqAv
EZLx/ZJ+7F4wmjY6RpbGBE+OobfPHvCPhA7FVBruHc+xch+MamNw1H4FLaBiBxIr1cV84H4Fanky
yAHaO7OGdlo/mndojyn9hYS9F53t48mezso447jALhUvvQqAwjE3rvCkDuVJ60JWr/uf+S8HmrI8
mMCEKrIU5sDRles2IJD9w34dwmXfCyHLpOVXIfyVY8QmvESBHkC+VeRomNugiz9hAS2xqAfQaHQd
bpPQDbDnF4o0xZO4v9RlblnmDnQiistBVhbuxCPnwujTdIgEgeJYmWSBNVP+e9zFQjJgLbTu6026
Irgdw5ER6ADkkB9Uj/qV1ComIoAXUeAuiujoZvyJTh5qKZB4OXD8b6Pts/5AU1l6BCHfPD3FYJHW
x/+TJxRD8Pv9zgmmFrd5cZQOmJ/LVRSH0fbmJ5dKheNlVOQyTTHU+yxByq/iRW5bQofv9eV3a/EW
0v0AgpENmZj3jPwICNJGgXLyYYCo0U6zC901IbCd1siWAqC3KnGsEUaraAvoszjYw6wDsKQffGF3
mr1om7UFpGW2q3tItGzZaFb+pOKCIJbL7oo09zwSSQMxBezWchw5sx0i4XBWPMjOA0zmusbvEbJ0
mQ+7sSp3QcRMWlROZRgYHUtO/mbysXBbt2v88pKJiVKSd4mw775w27dtwcRfqI900B49zL1o5V1b
XEWxdeHTVxShcu9OmMDP47J9beUAkKdAy9Bhezp8S0ezMtBksxH5LUMwZqJEAIWo6nOSi3OPZ45n
DItotnENVrjtE4heGDEDuAB8IVAp/CjDqrE0pL4lBWVzR9Vmfekx1RiCybq7mgosNun5eCW6a9UD
WBcXy0GLGtIy7umkGtqRmNsBN9nPMnSjDFIqlETDBJJGu62m13RRJ82kArfRZb9B9imTSCLYic8p
ip2GMt/GmK/7Rn8XYwkcmNpH0ej5D7WvOIgu8qigpT/0cE14OZjq7TzHX1oBFSBipgWAR/eMn+Lq
mjdzmIkIJkpQy3qp+rjWEI+VJzeX+7ZPGFy4/z/bBImokTe08TxL9fPlPD5JZlTQJI2MLw1DICVs
rMMXiT2MCbZYF8Iq3epyVQkaloWRs1ZVXXjRWlWJuqnLyXr87/oVxjNx0KfDaX3NicacF9u9aVaa
GcrBhY2/1gexQdxZE8bihELP7fJnxQWOPFLG/qUzwsu2h18pfwlnDVH6gtOGakSI6GXeFyAg+TDE
XOtRa8o/Wtb1quLzktya22vqjYfX8x0hHfTkItlctMRgd4aVGVEm/LSqd8sUD7AYp1DBVVIzlWqR
BMq45DuqiuvhV6Op1da1IC3LfIR08yF+A/GyT2juRXgDXOtpeq3a47EYRIdWrR7Sv4u913bW1K8J
Oy1pTqCuuqmP80T5Tm+HQdJv4VBt2EZcYfzskOmJ48BM0CmGTM6DuFn/5Ac3hhQ44mc5cQLre2lK
1h0qC66HIpedL8zDq4pY+MU5pVf3Ya+LPwR2+9yUci3TEs3Q1cXqBBqRHKQnmRFEtenFcr5Zu1X0
oSLzFAyKsxlSrdwR7WWkp67RasdQf/QHCVo3VtBEe/HU74XAWV0uzvZrI2OVEHgUgMoG7LdV0TI3
Fn+2RP6cZaGXOE25dq3DNx1wNbKcW5CewhxkepsUupoeoHeC5Qms/BNlpdbRcyR6zbnRdM/tYGRV
7RKoWe8GKK4v9NCNm1THG6GwbQvP7n8vaaIUILWYSjXhhWSkgy2MKP0Yz+NwOH0znhofO8j5CO9E
cjReS+7e5gHwvreI9u2BrS7AQvTXyAmhWVbEMDIsQOxv3wtDuT7kXThVFhgvIm0joHsB7pSypJ0o
zCt09/y5lCx38vCUuSHhghQqd0S6y0+Gy13zbsJ/840OMiUucMjDr27S/VmK6t3dCoeVYW9cOnlC
8E7t8ryhXEBtW8fduDJR5KmyJcfDPbEtETTTi5Fw1PmRhJZr6LIAifNlkm+5qzsF7cNKjNfh+wc3
1wMnaKtwfPT5rrwqjyDbCEnmhx2HiWao+x2Q34wQJDwtF/67GjBNfGDxW6fOI8bMBr/rAdx0plFG
F5rWSJJymHoH4Yd4mHbo3nD5PuajtpbYLtWU0/Dkf4VOIxBgsrbHuYqtfFr4bhf7nx8AN2dA8CeI
S4Et/tpsDEkB7H6QvPmi1Tp989h76JlClCi7lkvL/S9fSuPuRyIPOUoMSBJYPIqNKyTmlCIr1PWY
AMIuXYrYzcGNyQ/14PBPFdDjUooTBZDY9ywW8r0l0wewJWZPYSyxNh2wbnjf4dTreK40It/QV2Jb
r/8LYW+d6ktb5NeABmmKuFoURMXvTHrWpZA8BZt54w+O/gwbb6pKEwetBAEIk+mnw2PlL+OyH6PP
mIKZ1pcmUN4doj4BaqvGKQnp31L1AXRfbCLM0HGZaO7e/zLs6AefMMRYB6cMX4H08gKBE6b5QS9S
8DMd1iLwcdbhcMP1aIN+Ubyw+OY6z18/g/+8/xZg307Ftmkbx9AqIoycG5ckyRRidgVLQuPxxkSO
Vq2B0oQhvbYIf5EGQA4QtCc2s+zpAG2tQJ+HQqZKCQw+DOCON83AeK9s8mGxEOZpV5XBdqnJPW10
X+r+87FLyZPQy13wZLWfKEaAIYtrpkWFcgMdwLZ/OyK32cRa+SsytiqOahR4hn4eg20pP5ZqS5S8
wnc+DIiw1unW4MB9T1BF7zXE1SFSFXqXcCAeCmEsFS+nna9uoeG1iRZVB2QZ5WOOfw4AVjaUschH
/BcRJ4JbU3vuctjYkBoAqrRDG2dz0ON6NEE6059OvOYmaXljgwbaJImyo2mCkMBSO9r829LZEt7f
3rM7pLN3eD0kRCjXu/eF/nfrmytpUDhFKapxrl1YDP0G565sElP7Z9LFI5C8di4eAuv8e0E5ATAo
jVDXnDftQMQzZaCJWgshJCcq+H6Wj+Zj2/1XHMfIEvc8rfN5C/mzxJlp81YCJPgbvrVqjQh38fn2
+a4qQBYDok0fp/0yU2HM5qCuVOcoLuO6qSLpWORTZPfGZl8Y3KD6cdXAS5TRSACViA+bL1dK8+2I
Jrq9xlsNZpSrjC1yq/8bw40Ak2fmiUOndUpWNfPjK/2tiO/2rjUmE8LVHyZrIy32Cs9xbkg5c6mR
mati8UKyLN2wvJ5YYyWPLEfjiXBMpvEI/2bDyTWkdzgeuvmH+W6Its1YTCo1yWEtNmzM1jZUT8rg
uPEdw/CvLqHkTbisMsX1HR8MMk+nY81Qro1q/jr45cdFvrhnt+85YTOdn82gumjSqtgp+J+6coXA
KO7nwpxGhH+dIAnt60yPGC4LzfQ25MnRpustPvxeagaGZIZV9GC3q4pNjAPoGxH6oCeC/0oW3O1+
G8rYOvD0nRBCnQhyskshgk/vOY+3XusKaOBbPyIfVE/Wa/ZB15rycMGU89ia1EctqyJWFjAXPEAm
VOES/4NoRFBB8cN/HfLYFGJR31+ag8jn8bdIGvOhmeelZcTlzOMwFdNxQohaRrHBo5kAtwkJz/Pw
usGRqdtIMm+m7zdyH1NfApzONetUzyMEPSips+uY48x5R+BRquj3N7P7iBbKLcvF0ZtnnBq1S0sg
5WEi63NS0/N2i9yoxmD2frAM4THClaQ0DffzW8S5r/7YXr2gnTAsOVtwCvmrbD/G7AOoEsren+pC
j3lU/Co980V4xCLtn9sjqnbTgok9gjiTjT2s6tZB5KYBv6fbiw4fNvxeVOGwAq4zpbueLxWeS9pj
7mE55se9XGbn5ArTHnDQEVLnHMkCTbu3ixN2WOvuOrr1HIa23PpHckFLhiMPhdahnPnJMDSQmlet
Y5ZmG7GdfC7Nyljth5OuTuuRLkEUfGLm+YIamlm2bwjr2peGMNl3iIZ3vOaNvMeiFrw4yQaaipe9
c8GixFuHa32QPIUNw8fUKw/BlaiWbE7/Rpv14/OkP10VqAbytW5naC7ZOXrgFlT2fQ6/X0VjZc+6
Yz756wiB8o1fgOCGylEEVeL2xyBN2OhakOFqD4yn9IRo4ofnx0KL8ScHEWLjCQuDURqZEgFJ2vCw
r2g6wSDgNac6dcSibi2/zZVcA+s8UvAIbQSeUxNzRvdWWSYGEKSTEMGhkvAzKT4bhQq00XW/R0OA
I7IrTEeUFToPezkg7UBfKQnKdS0e0kK85mA1uSBQNg1zp+RS417KRLJJ8YcMlHKHJnWqpMFS3tu9
NH7eaKTDDBgk/dU2P1CvylNgg1J1Ay9AfqKfZxid86qQZErqTC+xHmaCFwedWDpy+tzTBTu1B9BF
T3ZJzHTelrDtW1ZyIkFi31dBDUYys7ejuU6YhBdOCRS3kB+ckuVthpuMnw4rqz3U8OGRE4EBTOb/
cmCR5txmbZmS4Mz08XJpQSLEymhNI5kl9tu8oMxqp2RWIa9B5LbF3q6Q7tyhD/jvQp8KWgC8oLZK
AlgtDwNmLmTENTHRBs6W6UdeBb5FGJGPzX+oOgcvGu0xitTKb2d7nGaMrjuMVXNaUqOiVlkQ/fh0
TrzKPXxqbFDVbtVuJqJgyIpC1ILVGLv0PLKtyOlyd2ymuVi5wgJ2HYBivObvh9vVh2YEPHa84m/M
9SVIalkiIgNdf306npDGfwW+RV7t018+UF7dWznx1pT3LNeMaL2AojENNYjHKdLE8ZcXOJLrFXlS
iFtv9vi3/IM28r8Zho/Q/BH5EcfOqbZOxDdUQClhRKKJpRrbi/gCBs+tpkt92/eavrmNRlGT7MlH
7jj3MUMZyl1iO3SsnkvAbT3BjY8iocVwnAk6d8lb4GT73/cZdbDwK+NHglnonLBRctdb/WGQlQWm
ciTrVELE8J5VFh64yYHWDdcxcaUkoqwY2o8HVWF9amENqAJ8uHkS2vMzy+eGILG1lR2KW6h4dZeb
JLjllNX7d8o9oHTgVSeO8HoHphD+AfrI5+9LmOnBXux0nl36wbFNEtmNcNcK3fDyTJ1f3HkSK89q
iOvRgJoIJ/y/ZL7xf8gmkSIabF+gtpDm2ZyBkpbrABVZazqyBCNOxiAZyxuOjLFcGwlfJawiUqDc
ubv0ucIDn/pXWNeU7Gb5V7fCwAbpsXkP9JdHaVSTugYtjJUA4Pclke2sWjdFnsEpAr+7KHYRuqtn
Ndk3ZwCVg5PQIW6lVek4aDf8EkogNFg5JdcJuy1HvcTdIunLKkV+4xPLyjgTDy5+9NaS28fSl99/
mbQiTJt9V6tuCVKnwsOsc3+oLH5lqoQDI578Spjv1lELrzn69FXFxKKwVsieiZBGkQjWXAglhE9I
lN+fRuBpJyOsUpr0wHclheDnJv/Yq315R+JG1evcYmVhLMxwouItyAn/vHs+8G/0pQ9BYQ7xkLdm
JkheWemyPCprzDp7icSFZa5rGj5W39ETaL2/0NKhzmiU+qz2rVEKctJr27BCfqmBRVd4BFYnLfQo
gsXZlqewM6iduIrQd1yiyjbhO1FtHCmc2+CpWh40cGb9EOM2/8PIyYbNM0yPAAIPekN9w4B4bVxY
w3Ex/IV+HwZ338RJZcmQNgL1c7giXcvCmNhIoTJm//NEwJAnKaF8hEsg8d6Ymdjvasn4hxSylrk/
y0JQjOmEdlHoKRlfbV8CUIYy3Jx6Gw6pN1NSzwvQGulF1Qu/nyw/DzJxACqjTuWhpu976Tv2lVOp
MwxM/filrI/7xiaDmU5LpjoBBYVbMqskAaSGz4k6AjeDED20DSGUX7EDAEQ+XBwAvlRgEiPXRDcR
j96A1/V3m2z3KvJECOsVKe/aTyuomT/8Y/QjkTYY7xI+agDphV6PZ4aKKDG/8ZIlrMrCyry8Ubnt
RGsovXJutfE+z16nt6uq052+YFq4OmDEwmKeh9dF7O0+6Rd94/atPW6rfvXyyE/qBSgF5VSgfdxc
3S4ybmIoRdSE2o/QdgMHfL42ul+akfUntcANPg40fF2uoac0sfVIYkMH82FFKLOIBVlP4veHQYLX
0ppIb4o6LENH4xQ2Iwz6+T7UkEmYk14PxrA0jsttTBU9r1UZhkSnpJHe4JR5mRQX150QPb9fq0Jg
h8u0V+X4ymh6u1r54e4Xbjnhv3iIx2HY0H3TBXEeyw3g4AlQNkbDq2IslLT/A8dgaJII1/DYsbHl
TGtm0wY+KDqug7HTmZ3zTIXGzjb0W3hOBa4UCvwh3cjRNOoOhEjM8RuSSDG6XdlCmLoi2/FPigIG
0YlPzGXWQ9q88tVoZDjSeHVmGG0+xU0kpcJMrszHNggOZdGNPrYrmYuoYOGJgnnqaMgmen8WeSTh
7DzYcqdSsnciu1pcA4hTIm94TCHqxyQEnmO7uewxs3HXIA/Ky3kNGYPP4l6yLbFgAuzy71mLMmjV
cjpHUhwk7Iw4CKsuCNFe5fy5DaZhF7eZG8qIsQ6TdTVgJsd6TiEsXenXO9To+Xf7Ei8jgtRwbgzX
BaAEaWvleQpbpMmhlv96GMaVQziHYun8D34f7trxCi12xJxhW9tF9rzBodZGpvxJfD+gUYbBRMsS
aqQhU59ETlUHOpwVXEmfVtVmUeepV72+0VAJ2AZxke3Z/4FjkdbfaWVi2oQGNEAjoa7hU0PaP1Uo
NWyJvLIpradkcVT872ru2c5NbRg9dbEydQ2B18ROCqVKprQbWd8mWB+d+fIQqhnB9HSS1IhGR4lo
Mv3VfET/1IZsGk4wNgG/3w0yFXBqy19w9kXTA8RApkAstLC5hANJJKOD/A0AzDUG1sw3P0umMKbo
0oz/60ScgyfZB+NonDecoGSqnGMvbtOGkWMSZQ9G/XawPn85z8LAqwb1vQxHTEx4orf+ajxcTYxD
6XmaO7oX56JTtB3z+CygtqALlh5Uc+HSyeXXK12/nsfMolvY7/t3aL+2YpAm0k7UfgmFzgorxoLH
ntytjM4x/tVPraaeNgbqMq39mOacQaMh1IlVNRq3LSoSfoF/thanCFvu+MoaXTyx4Mc+1lmwLze/
WpZDv/0b/v9GAoJHZDafFrHWwADwhO/TIgcmuQkheu8/+nvUGjU+nKQ6pnbbkKHMYONTmnWatkFA
0FCNaPVerx7f76xZfFHAoL01XnNTuUkipuBJgvWyBiZdMucUYoRBCk4G56oq5ODJU4e3n5zGD1f7
bQBMtL+Vh7JCNzEJmvFP1X/UFChvonod0L7sDoo1VK69JO4/ENfioVeTneg1gAn4BCntNW0vbsn8
FG5oWkjgjp1ERgcV4hCO9mISIc9N5/xrRQQnnC4/NAZuGXymTSAlZUfKQJGwqD40Ke7AVU70HjuH
c8TUDA7aQqsWCLsVkkggRJwgxBYTZ29bYaL56T1slltgg0BVpRypqnaU5cRwAdzLDHtCdXFCOKUu
fFCHVhxy1daPo0bVBgkDDjGEZDFmMiw9UQJb4HMiFVeTT9b+BHKpMrSgApstaR8x8Iu52j0ckNRs
GakXZ8e4xPgI6p1uzlQfHyBOhkEopzYWknfjRUYIuopahksl16jYPPIBwSac7ehot48LZ0kBed97
Cxb+s4gkiqC3Zyec+QyPyVeTRcTEu+a0WFXXSuUIzKnuUFQo5eSsqDSj9gU1QsXr/JjfqJxtciTr
bX/S75aX9pVzdd2Q2X1dJ9CYDCLNqrAbOzbaocvSLqQtKmnMqdRfLED8oM/jRJTakqOPpvLuAgvK
5mxizoGO6UXldowCQ5FcNcXTQDwfucj05n3ggOP9NoGj6t+ZLi6kvx37RnJu2GEVESdKL8R9+N5l
UdICWDMnbR8YHX64z0so+9Gq8LVJSY4RT7URsW+E7mwFoXqzsfBxhB2cXNlXvN/7dmCUpKE6O0hw
cVxFPn7wli+F25l7XWY7YS4OnF8phYysJQx15SJ9qV5fuNFtv9PwnzsNShEAtGb4dwmtD2c+Nl1v
pwq7iQZdm4oAMXvsBmivDjXXH4DxDOSRv0pZcSEW8sm6qm6SAzu1lBj2vbnCgyUUyNkTEVcdHxZS
Y5Ks2DdbnvHFufrKxibCTGGEruW38WxivzRN/j3hj+SLkQd9vQGVbyT+P6KMSz/n0jYRvmA19UE7
rvvf6sqxXZ335jUdyp8BEM5AsZ6EdUF0ZqjCYdRMrHZLTj3P+Dhyn0snlgZF0eShi36Z8XRSqxLV
xAZRoyabD9TIOshuSrJVFDNPAPugqG4WWJXuUUFgzwbyHGlA/cPCaU1SunaUZLKcEEtHf3drvtyJ
NjMGAYZR+WsJSJ6Tt3zvVEk6GEzQ2fg1f+sdvRJ0G4yI25KQkNYg0Zb5FOZgZAf+oh+Bh1BcGGQf
lQCaDJerFA02VFjPOCbnnfdMy6QHUhqble4+e5HP/JMlkFbVOx/tMXMYOm3+GSy1NUm1UyVfwpIw
q4yAkusJqBJORb57p7+kS65tsUttF0VZ39gU9LKiDmpGobq3WP/Sf9ZoHajVKGK6y5I6aZmfvMZt
gTUpiMRBAi5PuWjjJb3dFahjCE1WsO0KkYXLFbyhRy+WbK1wRJtcbhoPzjWKo94wiCHjkqk/c+lF
QWBREv/NabZFtrDIw8wJS2Z0LIn3vxJ7JT7tMsyeSSVFAYqRvwleP6dTWDtiKlDW0GPMNMXHye12
gfN8A+m41AX/zQoITpHEhwYi+bI4yj5Qtu8AiMjrcYxxOaKoXUk+XY5ho8SnUAEzb/OZrHN7QBiQ
zmz4gDSaf/jZckyS83A5hrmnehHgFzmH6wQM/ffY32KQUdoWEdSQTlvgMHA1I7jybaNk7kfKXYFe
51LpgACuUpKqwg7qePOU5zs3IJO51nIykWVJ/w/mTg2nbiVjWX7B+n3F0OtWDMC4k/LDAF/wP15m
VP5K6w+Yp/pzXWaFo2cDh9nqpckWE7+a3HmQPn2beq7k2E5GS8OJ1cCr84We7cAl1os6FElizqBs
JivDK8PJOZiW6TzXPCiNyvmFRqsB4BT4P7bicQCNBnJnm9EITO+xtL59V8HPcK7QzVHIUDj1fLXk
KVgC66dAMkp06YSHq8C/AnsLFpVXfXqYxRB0QPkTrdq3zb+9Yu7zkFc7CGKcI08igiT6QTtobZn6
jFepISAvizb0HmsRhgh0gvaovHrv2ipXDkpfvK5ShLym7+buJMlmQW0ErM9lyxmMxMIJU6ni785m
VJUmjs4lkezbG0J4EiXByymtBugK7qek1V9oaw+zVB/ZWIElMPk2xYQgVeQNfseXLzWXaN5hyiOS
2HKNuP8pw3A9WGGulP4cBnaHdgLGd01jyxTEJjeyvmbC/Hn0uMX8S+HNljUNCh0X3YpE73aP8gpt
LyKzrXmYZ5zNTbhtDObyOCt/GMIriNkYzv8j6L1AX30YhtJDdV50GubG5zWhHeBmVGC76zTmk4Hk
dczfe4xj5fXWHkA/qZi1vcXH04XOIHkyaQ12MC6c/Pud/n7IAD3BPrGs1H5bbbDShXmFcBMQhxi1
/GbXfoIyNqDhyEJRljNh9B4Qr3asgYKAjJAqgMZEyV1CAgSHXxmQGxpDSiJNvJfJq5fMB65ESe3e
tqX+tdLPL3h1frm4t7cIa3aghRU5T8GaJu487TzY9wNUt//ZKB/f/Ts290JOJ5F4OEt1sT0f94mH
6kJUBj21WsGAIcqyCeANkRlUy3ebZMo9LYAduJVotZAZbRW6zXShHfuUD1sXJxPOPK+vJ7M6xqPS
jGaD0TC50ugSh1xcIgwe/qsyWcB0uwEH+STA8v2Wbsl5HE/cFVn4HLiF2oryCWLrwgDAbvDIuOU2
kvIGadIU9gP3z5w1qsRCUFIU7tyu8iMDVuE+12JFnuEdQZiyWSQLLfjeooJrgeCNE5l7UtrEG15C
+vDAgPefRlkCNSeQnH+c4fVxuF7ry/7Y5zzAGP98tXpWxoBiUHK6HUykh0A4WTVjTuX77gtfXyK8
lkPdD8ilNu/1Zeh39B04fXDWEGQUQVGpnvzgxy7Sz6bwqy6FlyScq1eA51BD1PXSEekzYoVDLigZ
hDftYuEdXcT9fYmqPA+fwoggUoCXd7Shh1j4zFu76mzwM4lnQ5NAH0+QoNWxrW4R5HltgbWuRaaf
0IdxQz7ldlHdMMpOuiHx079RDkoUxANDOUqh0N/WzCoBfLou4GU7waYEFrcRzWzufOK/FaLoxMJx
bU634Ff+VmjRBsA+wYxBlV1DGIWlHIt4vzQ6m+yZqJTDJR9jFvcfDiKXYO+ocY+EtqEchF1hzBCq
o6Pcw7xUc7O6VaNm3fzR4fUgk9CuOyLF2q8j0ftSEVc7EpaoR0/3yKQK0KgOpXid1zpUI1OwhiCb
hj1Q/2skj0lvwKij5/m6Za4lysivp7nwGa4yW66RwSbV0LAToFvTG/HmEnBxV+2LwLc8VRHwT4it
cblZDU4/O/muCaCC7ilyYDqkmoBZKAGnPxuObonMMZg/MgMYxXUmLt7xAhu4U//phmKI8CE0UaCy
98FyGNclU4W55P5Bh6SLWJbzk4DcFWAlc/kkwinv7OHLhbGfcwId3iYpaRZI0ivPoDzqWtnRfT+y
qffdXBtNjxtgFU0Hg56XJbpP3ur91KR1m2PH+Q7WSLz/zH4tLVlKCR48qs60xX9pptcCtA/lDUUB
CFmd1fW5GVO3Ko18V1mBKHDIEdqdReb4BLb5EP//PXXu4+VtRyAE/TDhoaNlDy50bix5K4F+WXen
hUbffQz5junUkNG6IUVXQDlvlOMVbQUF4Vht5V6eugm5GdkAcv0A5sURJrkLiIkZAj5RSRrG8voC
yEKRYWojeikz8zGAObyQN3x37yMVmzBcD2eNoDaZ+8V3UGm754rLtoe/Fne4bHJif+3oXLYp4zfj
k47cLEHO8pxSCK2iC/g0kVEfzSJDa7CiRaUXbNWtLlHIN/rpEADU2OcPm1xaGcpXaSN1sqwKc6tl
XVtSR1zhWyI0jtKNB4TWoUkWC2T0t30ISHNTzCt92Rka9v4ZjGBOQglVRhslY440dUaXdJ9217cR
WwJ36XAgfIZbqkLZ21IB6G5CxFoyOH3EqP5pR6hL9yqLbFmZQG8htxriyuFndcUCYu1cArq45ZCS
9P3umKhi5lsAeq5El+MhE9HCWWlJ84Jsl1sK8P28ZDshqyghK0MdPjIWa4wdgYXZ9I/wCTbGUc8q
zrCHzmiDHj0JfsEUgV6Q8iOi/pp4suhKYUjDKcEEw6vZ2KM8MwKscLnuo6+T0jlT9FpSKkxMdxKk
5Hi5qExihow36EHzj+ichOHie75UEyQbkvX62jufaVR36LeoJTIDIfKgWi+HHyaGsGADxVn7USfu
2AKSnPq1z0LzntpEbNIQN7qVQb4SXF9a4J1DnScMQQ724SCXzomgYIB8FKhPVzD0S33XffWq1oJV
akLBKGOsNm0IrJVvjlvsDZQHWr1ajEsqG0gf0RNn5sHOJEBhAXCowo7DDIDKQwKkt9REOvkT+XAy
qC/A8SkuQKNySCVId2JTjoDegInbYQ0+WxG9zCCEOXBk6NM3btH6ue46+cOLjC3bdndV5vINMNH4
rMlObSHctcJeRgPZ/4VVB4xL8vP04ajWOatoYqVrHl7xn742rhZMaX5X1D9zf+AjcwaZg51nNVlo
heFVrMEm59aj+y3XzAo76xCFrRPLlT8jRpSt+UJPtySxybw5kDhBG3lNPIvPDKMDi5UvZIMsWu5u
7gVWOuBwIO60nrHSLEYIA7PknlB1Iql3ZrKHON0VPxQ3DXJXCXFlF2SnV/0Cdtfx00D7fywpNFrX
ssgmHtouH0CWlIhUm36WKtC3XYTtIT8t02KeM10LOsPFV9eWoDZTg6lAmAwdrU28AfoINflc89ef
xiNTp3GKDEzdc9e02OSLNC6C1zmSYWSDUjmg9FS3dasOCyHOjWUZ3+N42KR5bESRpMHOJgz91uUA
PRWIKuRpJgcmuitxFleEOODCgXANbG/lAmdp16zJ9ooua4DmJtG27MEA+M1RXvaRJZC1tiibCqVt
J/92IMQxZK4SGRkJ9x+J/hrKq/il7jylosHE5M32qWnhsyEuSZQcSAnQbL7dgNFnv3Fa6xsl4jXA
JAUGUD1L5pQfVkh9zyaE20sWAH7yb3lnsNWEGFEir4PMQ32FKEiDkJbVWX8S4/OUSvOu+z8bk8Dc
b8pW0DbDvKM5KzthsbvBdOgSqCT/QN6RcGY8uaH1aVtg5eAW+C3pNRfhp+44Wr/Wy4X6vue7Nu1U
QLCfYbswksHpYk2KNl4bRe5ZnWBwgujeTQZULPFINM0sHTSMpgjJXx3/EHJ8mlZ7tH7XMg3TO/H/
p5+phN/RY/NVy7Uke+jbEt/gEFzSW/b6fowQ5ipxw2cO8oWOlx+F/VMoXL53HsJGT6s48KKknYCb
pXI37pefSRNGujHnntJOKoYU/7n4qEJKrr7HR5su99afmd38UrBPqSbVOZE06Azmv/7MclmuBYAY
GvP3XlR3KmiLJoosXzplXyKJKjldBseXjAdB2BIMiEbfno3dS7vmGhXoJVmMqR8o3QC8LCDsRgQ5
MY2A9mWrzvuUyLlkuNPzGfK18vDyNK0eqMpWo3iezJwmpSEZKuiwH8lIROuZluBfUGJ0S6RkKOwO
oHnLfQCfvccZL1ZF2ABdM+TxQFndkRyHP7vC1oj0ozaRCsA5tt7Z2uGYJci7/ASsI0s1pFH6OsLn
8TS+d8gTKLeEPitbsKeHYdEkhJ1/z1Yt4Nd2Ru4e9nmkgYyb1rwd/JGx9xI+AAS2XUKcdwPJon4h
uz0FAyq1aypig8oRJiBUEGJ3By+XEMGBWXDtjDC4AstROT/i/80jWHuWLtPNYCv0hfs7ZkL1ScuF
ehR3N/NdPEXtrzpLv4Vpp7m5FMpp4v7TJ6CzC6fDp8gFQn+owghoeUGLA08eOTqkP3YirqpIjuvB
mnkHqLphlyMXgmUHK87L8jKTte6jwR0p2DdeEd7YXJhxvdswzie6HUheTSnCt0NnjBirQRxGasx4
2uB2bCKS0OIg2KOYfyLJTnIlnNSyZ09LT4X05b27cJ3eFhEEBSK+oI+94Vqpd4ELnpRsKRbnQjPh
yp22cN9hZ/peVwGESgCTSKS0LvrcEEqgl1OmjB76/xJMtiardk6mxa+v2VLENhFjVw1xYtRnBQZe
LErPVidCNnEt+403Go7OXf+v6z1hMeEuvdp9zgaRfUmLWO1nsBF/Yw0/iDy+9UTCwJyztKdcwUR+
psBwNDUhS6vpwWLgZAaJOSpkTk9brGkDKzeJK9C23HZihjx3cUwhtNXrnnw790t8AqnPfw53oESn
/jyCi4vyCvxemDu9YKJB518htNAAwC/u3fWT5vbVW3eUHss/+E4S+Zj23gn2JOoHuOe+2b4wAFGj
jMau/Aupn6GSycO7zRQI53gCCnUVBGpSOELUl+Wb0qqwL7KR0I2rFz/YAa2J1nSJ4QA5P2ZzCc7K
kj4ZPgtSOZo+sKPtU47rKBoJf3+AP5TGBrkCfrR6cW6pFKONlwaMlubQsq2Gli1j2g3V9pJNVEhE
eskIsng8sVt8maIfcWelniBTP3wu5N242uPkv3qT5LBuMqYjoasr+s0tpFw1GHotCnvUTudvKQRe
YybJMqsLiYPVgRVPFf10IWA6ZrgqK3RRcqPr3DxyMDqSVrPN7gAseCi/NZX+zL79DGiUjugyxgbO
ReX3/oHroqItgDh1wBIGlnikdWxbM1ZCX+ppekenRLq+5nGxfhZcs61EnZsRj3X5uMdCGtwkNlXi
NnCakZqrLqo0tbYx0FtxxM6j0eL+SY3cbVcuQAR9fTvW50l2tjfZq2tcXiETXTBLxifYdnlUh02H
j8jB/JYMvn0Knbat28KJpoolh/e9fZJG7WTjDI8lrk0zq7FUg8AcPEXinQ5QViLbPPNaj3yn/kiK
TQLzdoZc5aSANtgmlmMq18kIGxwIEq9fnLqaIchHPcqSAvIgbsJUXmt5OS4FXNeYIyXmUrKCmguK
m8FhfWQr0WMSCjYZGf4qBuCI2Xd6PDiEc8NhjirX3EY7HOWepYrqgfIK/IvyKufaMbZuU9LiTB+K
nyaUPYzRyrniS2PvMD2VJAP/zHsTqN8Pim1s5tjcTo92D6zgytkF+ILHmhjhwwXjpOGkmz9jPxBU
NqJzhL2OpRBFboXvUb+mlvi1JFRmbxWIP/svK9DCYDYnkhyubzQkGo7Y318dm9wZSMKcVeuj0YTI
QxAKQ+xxKp5YwTwNvZtiQygXYiAlXLbjThvxqyuC1LekC4s5DNeeOjH48gWuAFRMpGKdIBrIDaRb
jGUQT9LXEGlCfZy0VAttUIftsk5JScAs3h2Bn7/Z/CROxuoxHCMI7aWx6+g9ssgL+ZMUFdu1KMFV
1XRI6mcJYM8Xaj7+Frn1dpIe5J7nf9iZJ47zzbsLWMZ1ii0Kh43SsZ057Or+g6mqTCuUHpvpdxWT
iD0ME+kHrGHIUTdSxBKWpI9Xh/DuOpv0UqvH0krOJvE9e0vDuw1U6PGp5BDJW3T5YGyCkOQUfyrG
zIAhFXstGVRxb7HyJiZ5S/1eqXD1XFqC6e/YkTOXT764hpr3hwF9Azn+MnY3vGWmkJmslcm13l7K
MgT5ZQOdODA+xPYCJnupX8NQGNPyV31p5nYdw6YP8FstY2aQs4DUctAeHiItKj2QM7oxQ3Z30WVW
dZwlW01lXXA1CsyAaF1qRY8DTxBskl8QqhklIFUfxaLoF8CPMUevJ70SelVo7QULNc6gBvfeddZJ
IWXFUiMjryBwGrFc0O8z/x/gvWE37RDJN7SSbm0i+KpLGIvPluLSTwrHpf3e7qd6w+C/x9NvP4P2
jO0pY27CaxUUOwt615HkPZSFghUgIJMIKhLq8iMJdbKBORlRnJInmhDDzp0nJTLnvl9h+gSu6fnw
JWmMBeON2Y7+uQURMuHzPqOmJzhXbMwOipC2lXy94gRIxIFaK4p92GaTYmxM8mqVg4rmELowlknZ
euM4rfl/Q128HN5SZag0Zz9SQG+6fQZRbydHZP6DbiqwyC4VOIxcEwa2MG/PYr2gfRjg8pKoqVKI
H5D+TlbsKuKt2YBTMnjmD6eR2QNPJlTYhDvLy0ZTvpR38yihXcNJ3eTxxPWm/HzDZRQEhg2YIdPg
45+Nf5oMPoPbcwgcj2Q3gz5NmeZR9NcNJwx6CDEehT3J2DFSuIoXjqGtvXsnJ1fqdjZ2nt22pEtY
/G4v4EIicm4bNo0t+0FLApB/ycH9PQclDnvF9DmWHJMaP7XvPaOtAnwfJ4p9zDfiblSTvy4H4KEA
nWBlGyHIyRSszrZeQveDVXaac+QA68rgdIt71AHlmkIKGDqKAn8AljYPE7Bc1Kd+E+dmVygT1vuW
ba8sfJZCrZeRiqWURFDT10M9Jtk6o/U1KAsOjj6kTjEW5wHZhoIHPQfO3Bg6zS3HltFc/gQO0mec
dG2sVKbUBDS3LGnJt1ju8dXUrpVFxcOPSxHWlpP+/P1VzhXDpIVAlaGyFGh3CL6MAMT9dRR21345
9F6g69vhzhIgb9UCrkvpRLUkSLz53M9cI0CrQrnucwwjU2a3FbqpQpL11dk2wwQU0uJot/GNDTe7
/cJLphYBHQpWSlMKILKJZvzgMBxws668kgZZFYibpU0xXExb2sDXH6psdLt/q8IrZFgEjOhAXxvB
MxYCH/QY4fMABlNu9KuQ+x4QWaWhM6j/rxIpXCbcb8gLYjTMIbSQjPuJDEf8bRyP7x8pCzsWh6Il
4GeXh7Km1xNrUPW67McI/9mFqSRQ4jEeyjICZdxbewz0ylUdXR1FMpDIGaEGYGjGMN8SkkApMiSd
OhnfTXxCZ5ewvXi5tr0nO8W7JE2iZNeTmW0VmUl47Htwult1cBZPFeawlaOByknkiRddc/aIdsN/
mMayUmWqMRxaIw+zVcTX62qrMYxxXzpZokQCoomS6XrgjJT+h2LoJBjPYFyRtwPsX2iHXxX0Mk4y
IcHI3zUuqOvUIfRTP2lOMPTzPs2kif2s8a3zDe878u7s5snlOComnBWB6Cf7ONs6zfRw3MjFX2lD
0v2vMaHU6B8wzhAA2ipgbYPaPB8sVNkdVxtvMNgVT6Bj12tB0nmOBqpnp0BIzC3qea75z2aeoYJK
u2gLSlcT0b8AnFbGolu8WGlqKNKF8l7CUT8idl+c8unyQnDrA8gwuASQkhZBSLlvBaQpTTD4hzSR
LQTmY5y6pfRxjWTE8U3fnJT9kGTxdf+0Cgld39tT9mVPMp09Wq3R0ZyG11tBrT/sXpehMgLsh0m5
znpPBv+loLaZR14yREMbpAK5sgKm6ooRyfeiBe/jzXfFaRw7K4X31RO/8LjRdsZ2UBK2U0zSL2eT
f+fTDDXV/L1jtEAnzvS6HRlc7pLDzgVfUuqlgCTZc6w8fvMfq6llC2ojKfSntcBZDZGCOfDSV7EF
rAh3IZD1/oeXHI48fYXzBXW81J5tLKcDpzCih+URCYzOj6Kflkni/42wB62g+yBSGksE/uWNIQ/P
UDDTrCBM3rpQsEK5Em2WkB+/MPQj3OXSWBUZSIvj2h234bBLGb/+FDKl5f1O/Cqi8nDAoIH0o3TR
ei+L6EvE/hCCfuPAoht+jCZHy7zLUbod1t2XaYcKS7CXgSc1TXfxGHLpgy86Kv/0RkdKvGAvuNnn
yvNEP3bBG3nlR0JeEYU8YwYxLLc/TRKUCRHnDDZB2xTTSjNh1hZpTnT868mCoOTjfW44cB0Gl1cM
SXapswAkUktGyoyQH7tx5+WlOUi2DFWSqHRD2FStqhFzRDoi6PIwhT5sqzSk6dS51ww8i4S5S33Z
+tBvITHmGzV7cUQjxl5nWzyT+rUiwYOi6bx6fDRoKLIxYP2jO0FjyWa1dNxlN1yE+0uYZELdLhPB
gO0PD4E9yD58lQjQM+bI8o/E8b+KyjPLyCYsLXqQoJLm1y9+8ZqEV1MeAxVe7dmBdd2+0PJQ9Y/r
beBR23vyIsKS4lv/jKaSqCIBc6L6zSvB+UKLzfZ4ALJO8qVlX4kU2G24wB/LJ3PMIebUh3lAQXhp
0VwhT+B7XHGEes1AafTycmLOYlY0Aqj73nU3p87sg87srlObHhEQb7ppPdozo7f+2WP46y4HYwEA
inY0tMjdETEvl5CVZkPGqUBp1i7o8MItcrZHSR55gx0bWWlMcokzfJsk4U0hy8SUmMabk0Jn/x4j
nQH3Yvia1co1xOxiCcACBXyr0+kYb5hirrT5q8gFwMiAMTrTvxNNknFCGVg3bdZNjBZ/KPqsLdse
jXh3wqm7G3TbtLbwDEAM+jm9dgMFYD9BsvvskwSNFw7V9psPEhAjqmY5on+zeslHaLy+/L3bPYNa
6eNQhUSbDoq4WLqVstNtWNdCcxI+oDDN3c6UWEoZGbScy4MgJyUaceR1x+deUs5SQky0osyFebIX
VVvh6hQq9wPAd/dNmqVxSjXDQrIxFeENX3OQwjzfmDsrJ9HKsaor19zHXnorre+rShgWw0CKVVG6
PZSHSFgqVnrkstSLnceWPvbtjfX+iF6UwxRaR09rJkNJ+LggUpMKzQyl/8xnixG94XieIjOHyqdj
bt4yMreEK9ykOH2TB73ostOE1kiUqPIbd5RAdx7uqszAnLKJ/dabUhGMsq4QSpgiHkL4eO7y37oq
xwYUyPnImH7rAX9K40WPa8EchoKv6E2samVSvaodH+GPwjJg9QiK+DEnl3eiNoVMIIM0ZRhKbmBr
XFXwmfs6xJ3XErOfLo+E5iJ0NIiu5t8DPGphoX8jsUCU8UPZvrSz+qT1fsqODjUEmGRVy4EgaSFF
AyxQiC0IyP2iUDWT98Knv4U8mP5IVGHsnIwwpfv3x6yhsEkhMQYXeXtzh+YDXZTZGVK/SxURtM0Q
J4a3+BnpdkTKUHow/OoH8/zDbnu6S0D50N35e8l057y42zTv3JcJ+LtO99cMw6RH587oqwkUeUNj
mUjtHtcgTPuHzd9lgq1LLpn1It6E2f19HqIOaJtn4AAp0hzE6MS8Y7wx4BfOADLP/X0ajzzUD7z5
my4h/KDJJMlikpAnel0pzp0QYRwU9vwsk0WrAe5TnCOE++YHnwCq4eZrNFpZBq/Um4IrO7hvo5rQ
KmMCyPGWXnh9e7egfskAyKTXNZaUvWlxGQpDsKayBrlBRjkO1FXTsQAH/gvDX6fDu3LS+5nczD9D
TzIeylteTHrO8d7oYp60js6lsdnAAsmAqQtkzIVex4gjp59avnhUFqCwnqDTEmU66yxRrnpgXjLQ
mPey0IwDLPEPLinsFoGuaDtqNbF/J4B1UyRZm/VwKlGiREQFEPZvwKNdSJgu0i0CBMFsXKd6msxR
ufQA/0P6/EBqW+GvbVwjnPqgt/TLMbOse0fgKKGxJHAMV2o4wvOoTy2u6X9/Y0Rd0BxN+1EigY0H
5mmCn6m3SwnrgHOawi2sh8ZMgvzAdgukAhtFSbT2XWyifVj/ayI+ECYgM2v3M236IAsAHxOolSZa
qcx8o7pD0LwYyd6lyE+nk0h/DEyBbvMCKxP3H2DE5a8SMLOlfa+y3xhHf736XUrWe2e3L/XLAzox
TEP2NwoZBOVkFQEZJ4gMSAcI9W0AevyIcWB129kBaWOvHgAxfgL5zBMre6DIBCFkuK3DuNrLxm6R
PpbOsV2V7fTHtKIhsp+xMvr0yTurCT33B+xUCfnsjlAZWPUNdE1lsGsVht4uJyeQcfN9RBhfZFik
gzPOC4Qv/Vm3meYSSS52yhC+HJZqMXzC9RDdxa4UJBidiFg9Lb807Kem8/Qhibp0J053LquJutY+
erkZNhoYM5lCvmAW/Z0h3L7f1ZBYPHAwKdgpoKnL7bjVcKhLaB2zaOSpUgw7FXKgx+CO6Icmhngi
msWb/WuiDXyexoJPNhuRLzA8ENBV6LF3p38sKyhJe1EoM5ahdvFOvwZhgwihS9T1gmQ6fZPO0xAn
XnnXLMy1lRpt4huLFgWsuxTPDss2cx0pAwUqBYbmXlko6mQa8s9PVSNHCB2FectIehtDmgCNDWOi
kDplfQmeEky/gDE5vVseQOQfFAsPvfhej67F8fgZxm2kDvkk588fzdGe6LcsgiwGg/9T9+S2mqsv
rIMVIWEkUxJjWt4ula9dTTX0pn/9bRl7gHlVdpUz3F0MEsC4pn/lHelU3WI7iQbyVnYqZiJe7AlC
mlIq7emr2oLvpPGw/tcYqik4je70xtxwvtAW0YckCeWksPsPcIhWUEkvu5SZvMOMohRt0YUb3Xtv
XU6CQMnQf1qLmYEY7u5PlGr3Ugpl6BoQP2uvnoKAMLzJivG9PhR0DIjDjyeVOKEtaM/OK8M0iR1U
LlpKklXH7WFM6xi4kewvD+Cai2Ri8CxBmNEfqUCbtPk5We6/N/9O6HhSKDbxhg5W+lrQfPCsoEdv
DjAYRH33Z5xvqi+jMyfobEP8wnUcN9wuVhil7o3DVC5xLl2FXuwBbxsiih/AwHgnPi8CK9ffu7ld
y4Aw++Q9AEBVq7L+ZQjIRDD+88ufWQ93VIuxiNds0fPo0kLJMxXndD5JLt1QjgBYBrIJm9VJmH/5
YQGD1eoIDjsEwuMLh58lXee7azDneQPhTKsfy1btpNvKqhs4SgEocLrv/U+L0yYWJIwyakiMmN73
VvvfMhR6eFNUM7GnX8V6dzKuh+uQQd51YXy2kUE3reiG7NBkNeSmstuHGP+9zYhY4EIS7EWTadrt
E7zc4If5mTrLPAjgikgcGpqcufDs+aeb5pFX38Xl5P5W6h9sFzb7OAOManhPbYK9IcWjKK8vrBMH
wXIqENRxoG92N+BDvf9GA1aEH5tp0DZbnWlQvFDQDORtDuaNjf2CIV3aEJ9IwXvIebLBFzDcH/et
EeervuaOWqH8SKeTA/fmlOKyeNEbbCXu/ew7Skb+XOvxSH3RARmcBnDxv2eJilStGp6yPUHoLylf
clSQtLyBN/G+ea21AM35rZ2R9+G2OX/0Mp2g99It9wZqHU1hXBitHpGuKqwrN/aOWO7t22mZ1VEi
AgBHwMpnz+tlPfsPwRCUWibRmHdeFzShnHUoKATNwLWVfoZD+OuKtDrFDeBG9Oz2OForUSmzdpjw
fLLpCIeJfNleZY2gnYTYWLml94I2W/Cg0Er2u5TZSRMLLXCm+ABkDAUVPSIY+yrHQQ6BDrrBm24b
wl/oSim338dTxZ5n5dtTBJHvHo6Xn40HnCopmGJjtZXPjrBSU88HhA4j/n3DXEM1h/tGNb1lxhSS
KP+kPrgpMDZuwCSaAlhUx9Er0cceBeUlwGBtW9iInrrmc4fsaPaUMz0rQzg8XhIv979WYDNU5bhv
ntQ5ytAUU0byDFS2brFaqpetjOLo9kvIiThzvOBBGtgiRao9UDVM5+QUjfMLjB7kiu5mPuX7Yoxe
LaK9NcOmyZt9OrtNKtexeAhoFwA6MpgWFyodISn6P8vINHZ2U+FmdW6TdlSZayxxshb8RpjKduZy
jo1pIBcMBNZ16xWu9QtLQ93Zfo1TOcSNXzJNp2HpHf9SCcmBee93eCAfno0TLofSr844463xLi9o
1tFdeqPI1zEy+EUe84pMZqT9y6zlWt/fkWy1Z8J2+GUWVZCbse+sBW0Sg1/LSb8twoG79Oo7t7pi
cQEulZMaHczpstnhSRryu/1xrPRHncOnOpOSrCgl0mL3UFBumYiGidhqbCgNuttMO6EnAqpHrgSX
jytOxg9rP/klYLB9ntuqW8olQGvoYLyct3BmGS1xse/G3/B8kFbT5lvEVeVJIQnn/8alFkHW/Tre
tcf4SwP2FatwZrd1LNJKlpw7ApkZciGW2XaAeA/6Yhy2FXf9pf47qGk6ed8/vUlpmJCpKNZBLXQL
N+SMnsSmi/cPP3UjQBzButSWRv+FU+Vd382ut1K8jaLVT4hV1z4zCX3jiTIIKPI1p01rLwEPSM0z
gGJvNlcWGZYqNPaIJjDWgG+I6CDCBcmznxeZhP1UxwPTiYq+J0k4Beyonwv8NSnElnBAmEMMexIE
5lzSZP/8w7tW4OAxd2IQO9wvPQUjlZwblRSS07VnsVvIuDovpJdDDdULEPb9Q4YznlgOPfqqq+4/
4wZdEl2LdKW+J0i0AbBsDygRd/AvLFmNXZArSPAR/DGsqWwfcSzTTBeVwW5rTI68Mdm5ufbHC8uC
0RW2xdO8D1Agl4uE+UxTSDufvvsYipNmRZlCEys1bT6WSbRwdLqn294OmsMz/5FbFxY65e6+pTTH
HK0Ch6XrEe+TDfdWG/2NJw31YmREnHR3tm2uNZ3KxNryypleTYuHZyyh/HbN32wFk6QYyh4OWei9
pODMtWsVaBIENGFUgdqB+a2ZEIIUHfA5Q63o0F1vVOcgr83rdlgrbHvT+/ZIGBWVr4wN40asRBXV
VJRvP8oZ06fHXajvvf+0d7QET5b2hSX8PU+hFKMxWCYtjUU2JOjDOp4UnFUJWwzga1V8vGifqcFE
8Kvg/vjj1bB5OrV1bJmgwGxkjywvGYmNrVhJbFLcuW5JljUh3gVDUZpeeghcAVfRMd7Zv0yeGfcn
zqyJuhfnw6dRoj7cGVkOqNggwmpM7BVie7DgZLxJSiRB6+XQavCsJ8z6l1R8lno10bsO9lMFMbfk
seclD6fMIUs+rvS95jnJNg1MEJtt6z44Tms8j2sqOBKCpp7LMEuk2EJ7raUPJTB5bZktDsCXeZak
UfdxL3wdfxfu0Vb+YEzqg0QHXPTmlfH7YHocYwi1rK0iTbqI5IvPvW9HxeYQoCG6ETMHd9iUZ/a+
7sq5Kx+Gj7iE2AftTdWwJ8Rv+FOk2lSGyRuCvPtXXQ3E4PNRQg6eRWv+E269tqIn3OPlPM3Nx87i
FBQLYitx+nRISu1mXlbwq6WPciV9AIzIXLCKzE1jWd2nP7AgJuZJoQlJqJww6NkgbSkKE6TcbSkv
jwFh9WLuraTnXA6o9rBOW738ddEKC5xfyobvjPa5qpeichrVRJvTdNjXKQSTAOF2PcxHJN68tyhH
2ZAXdnvO4eiSk7kWf7+VeSKalRD/AlVjd3QuhOmuab0hdB7p2xfkl44hi0MtVSgBQ2LvXQJkI1uE
5tZAyPzDst719E87+blR/Fp8/rNKSwRoCnxxgkZqf4jFGdKB7gIfbk9xG3tOmWGw/ADtnZ/Be27o
/IZ8uFRkCG8HxYeqtsn3ubAKuliFhVA+X8fzlhgG//7csdB3Giy8UO5x9+JEDADyjJBXCIt6eDan
19RfXReCrQUKb74K8vmGpruXQ9QR7bAUNQOtcZY4JbtPLgK/qH7Vb06uHulmzvH4oU4desJBSSvA
9OZO7qvzjj9TXQvDLaDlniCLOSNwZES6mx4dEF8giFLquB2lAosOTEj65JTC/hYgf6hU4pRIeRvs
y1KbT2jgkLVSmn6WtXoW32l8pFsJ8eitKOv8SYlOVdUr9F9QZMYh2eqqOmUD4bnjDxmsvy2C4d0R
VNK7eA+cEFaqCII0/W5+nVUTwtCvth64oOMQlw2ZnQhpTStdIPmDH5/zm9pZcDyNQREQ+FDWh8PR
prEQ6ZHps5bIl7SpiQNNSljkcHAFSeFjwVcfhkF9zv19l4pTO+3A5ARp4Lh/g2JyV6jwrFp8+5wz
ukslaIbSv6sUlwaKEFsVdbDmYpVOJ0JcO7PlAWGQ/vtPPMwoiz8nCSaMaDHoQkvifHkXJksLL4+t
zVIFhtQkf+v+E7JpS4oo0DftLBXwvYHR9WTzKguECcVLBIHkkjjQ6A08H05fJjrJIvoTKq2nGmTh
P8SQJ8DSvxxA6qBdvEI+dzjxhV+/Jk7J/qtmDyt6UHP+z92ljHN330KVXiHqoMfxtiwJs/OZW4f6
EoIwNxyvfdTif693MHDR97t5Ns3WdUcSk9rLX27kQpyLNqHqKVM34f6VKrevuaC0U65tS2I8MuJs
rTE63D6Yi081ILZ+ZoojWpot2DnWOKNXadpb7rMjgg33oS/TeO9ohGZi2XCOw67itegScFv82Jpe
ookSrKbY1toOKme9ge1/TE0fX7IoTQ7ld1/gfoiPA5HnK8JViZpm+Z4LND/2P3FIH5qmfj1YsyoN
+QoavZdjO+E/NlopjlRJ1SRf75tc0D5im0OJ8mJFggpZPMCV9tLwDYN4MqSipwIroap7zblZp/pQ
9akj+hvTp2FuM782x8cvmOCDWTr8Rdf0L704W65zP+S4VYiwjO8IMBlSBaegKnwtgkNSwiEWxWuZ
svAfsAKp5Bn+PA7WUfjWBp3jtW4Dpk2i+u8Ivg3vg696NP+JnDnj7NdMXpHfMUniRrhCgLGnT/Q8
wc5n7XTynuJB+Kt3ui7Rvx4M8nx4t5ITF4KPOLfzmZkjfDObhzi/KF4+aL7ly9zqdK7mNcZQT2lf
QZfEiW4mvj9bz1jWLp+kUrtBwuDUfH1TJQ/zntnTsdHFnnFUapn2eb9fzf1XeDUuoXdLyvSApGww
LshQYeWfbVuBzBJ/TVk2UHVfzyH3a1oSNJ0VkzHYlczJnDV+fJQZM4FUK3d0Glg9DvZx5DjmP0i4
waFW7cYBARwxsWEaPVnUwq0xMWFSGB1M07TBTViUXEPCmqP5AFGJIIO8b/mpOSPBkQoXpr+UUmd3
9cwemlzMpvQs1TSlQ0qjXqi+CfBJNspLF77+BseOBT37JBOYtp2mgNLYKZEZCoqRJl06ek9uAj8E
UH2NGAOFHtcH8SxYfwWRwyn3rJUL8tBnjA3W5NdLswxe3GcRTNMxsS1wHYoFB/5JAEu7alZ6YeAt
apoe3WajJJ+nbg0Few8Z44iWnonGNB54N2QpKBuDE+NU5TyIzJtnE6JxS+kK3D6epjAf3Gpzd1W/
jBAdEEJprBUDNgn0zbqHibtfGoWH2ARAVU6NR0HTSHte6bP49rKtHdKcK6FipmLqB51lbWtTI7dt
eJx+d+wsLhTEiuzXUP/3cHr7y4qWMDotP0f/EeahIBWbaUcTbbDD08ldqeSDMc2llKmIenUc65cM
6HECMqyRkcYhhwtOy/0eQAvXUWv4rSnQr/phsw2RnimqgUY6gXlbPXIcA3kn9DOwaH0ylp50+78k
n7vkFHHiN7PvmSKCZg1NNDwTM09CgPFpAWEFEr+lOIrbSgLlDugun7DptbPCb+CaEdRyMVbIkxek
jBNABczbZLJ+YFnTWZtLV1R06oLaXPmSGu7Mq0M5k7Ef7EWtAKwArF7Ckx2UBzQgrXB9Jq+ITDhP
9gQT2WZc7c04j3rpDIzfWF+D/ALcPG+21tKa/fqAe/ejAC1WtwwjiTVT7P4LS67HCs+w9MHafOfl
Ncep65gpCdyoR6bVx32zLPp9U5/vhv2/fg8RVupLPlE/yTnAI/UeR0lqvUHh3ZD3JjswgGIF8qVo
mvqwjaDV2WchLao784cqViXCOObp0hOk8CUeF78KDT2hRDKLkS2AZDBwNVKeZs+mZthHTnAwn/Nt
H8WdpH5+W7mX3+61Qnogpn436ajJiaWTmIOyKoTe/e/oZNFXfw29/Ks/qN03bi7CEA8rsdqoAobB
OXR2HVQsYw09YISt4k3W+extxFJuINseupE5n+Fc8GQB5Ioyud/lffKUokhoQeClzY9W8wfoVIlt
n95HralwojzJ6TbDukiswHf1Rfvc21vuqjjH0fSPjrZf1p3nHubmvg/eN7SpG654REiUFBXzecoN
g4EGbCvoOcEqnwZRunNDmn0ml7t1yZUrBJPggxgEphNHusZcKCu0wb3tigXdNWbcwtXKpKU5JdQw
6kKLnIC/pn9aF1427jMVvm0D/SaSy9OzL/iuV5Qgf/3wRT5xtBhZS8/trfI4sDCgWzUakN+udQ1M
ll39hooKmnPwW16wu6/4qr/KsblC2mLsjMsWPOp4RN7Jd+WiESJXmRwnVcXDkfY3LldTfmk2/eHa
oZvYWCa7NIFRJXgzCzj4++bJ5GU4txYYPhmuH8fJiMVyo5ovTt0WHRGBmi5OqmoVcbMEhzTqXBr1
6FvTXe7SFwhoEnTMyYg1bdWvHMZyVOmbmEdVvwMJ7uXa0DJvwKScYstNFihQiP8mqTVR2VHC+Nj2
T0Sy2b99EVZcyyjCB7an/Rp2TC9B+MCuztd0kCSTKgrdyH6nKxaJmfcMpbAKuxrMsCu/LPusg+yl
HHYgSgFdaAdh/loi9p9/fm2DJQuL9g/5wnEx49xenKh1qNp3HYw5GxPR9ts0t59GnnczkMVQqdVi
9m353/g37UmZhbBXswVYTECcsgkwx1BEWJqaDqBTSncl9BLcfGEmhkQcYuNVuhMJNX+oM1HodbhS
44Sp15zU54t8RgrGb3alvQGcON1vZR7uI0oJoM612j6hM0wTEcvfPP+S/hhMGaCmBqdLpOKG2SFZ
nfWaZn0yyTLPIxj570A8uft9OLTfl6oPCfi4LJ8qOcE9IYxbfraM2LFS0l5s85S7JhK4IvIuIm7G
+W3ClK1Y/4bHAiOMqQm+131NmxjCCFqVvSzMTHWTn3RzfvhbnkYbOyuGv/W3t/9OXFyWh++Wj+v4
px6kMmzT/6glC/9kl+4x9N6fyLeBPU1ytovW/kRfkeLNqLYShAQdl1wCN9oHFqF5Ro6wWiry0RAd
ke6dE3PcefSZCFSNuo4ZyC3RFo23ZE8UfkxNJNz7ZAc1sLMS/nTiHuOiWFxvsX8APsKOQn1Jh8ul
VOzmpvkiI/vbZfZo8sIWE3EMq2BEFCNFG8Q9un4qGRkDtxaLnFNIBddvNj6lBKzrPDW9QSvnKIEd
k3kDL9Nm9NCjN1oxg9T5B7Xmi71RnX2qV9tv/FOt+6sU3KiUGg1KQPbqXL6nd28OYVwjiQ+4ftGC
IiCZIuTfu7vcy8xWWgloGELHaFqoB1ypPUxwUo4NP7qCpwOI9UH2Ncue2CQyMdVBk4YWGyBalST5
fAabd/rHW2ITRs5ix9qcs6LzsRtn3I6usLzUPMdaJwIggMC7oQnYf7HHsotWmeR5rBC0tPaD2HAB
HUJwdtwfpYyJkAv7QtFlj5F0ZdgLmSeMw8Diquxp5mxx3RAiYKGGCCZX0WH5s+67eWeaIP3YYJcE
+JXxAc3of7QGGkGJLuxt5v+GGoQ4jk35CQTA84UZJHFLxbe7JPYe1oDrQpU3jkZa2kM6ZTGFjFID
qcfKj8VGJXuTWnP4NLvE7hkB7vf791mnIZTs3gqPYUxWB6uz8cQ0xlrZdEfxI15uyqwdwzPzU2gA
wGNJYUd05S5wKIOki1LBq2Z5Putw7gFI7tzBkDf1FrNdxcZt32yfyJndk/DBGJ9bJNz0yTJ+kg/e
2Uk5kx6mozL2D4pBLRDvqwoAVLycyuvjxXwEtkp9zDVyZueO/kLkrfvNcDiy80x6EqFLjhzcI4HA
KPxtWYj6e0aXLNgAxT9mfEZrp0RoOn5iqg6QldMoISv5Gly+zbBE1v+HLtfqT0u4PLbPb7QW0OEf
GvIMc56dxELXNZTyxs7KTVfOikATO5evO2UhznprFQ/SA9QrRku16NiUV0DHmE8pnhMW6l6ZmLFX
F4xym5sDyiU4SaiEwfTWoFvxN2JhrOPsCGYK6sXpBFNSKTSAn1AYzXLP3MHXEjIMUzHLjLwsCdyh
Ul8W70XfrQ5v/A3FoIwz4Y1jrnt7b3YOczAMtC+WhePi18tyaI4FEIIh8DzU1BEAUlAF1n0NF3eA
wHpXzFLVY7hG4H35mnnTTrwPLNBG1DytjEp0L0w/l2iRqKKu+/YA6ug2JG4mF4+pfrSRO/F8EPd1
muppFqPz092dhjXZFUBze6F/NSp5xmK9lmIlXZCIYqljC/Rvbuoxm4RunSq+Hx03WJq5gMwy8PBZ
mTnbwxBViV7mTvHrMTtYImBpSWuZLYyLHR4bwQaDNVCd6NJ5ogkKMUtZX8bfvGspQtOm9lMdWy6n
P3j9+Z7WxLNLvmIbQ79gOgK1faNXQVLt5X6972iEXVAJuEHHJiwQGmPkSc8TDJccKJALoUxQnJ1v
8eXtb/v2OkAX34zSm1g+uFFssoXrlnBawgFO/rNFiHocZqDicajvH4km/ESvhPXk5MXxmJXQ9DDR
D9LXl0NRqi3Vd2h+CJvCgQnIjb5jbxvCzZxqW4FBONe7XH0wo8BlCJnnByyK0ueefW8xv+Elf47E
2VUGa3y3kjuWiELA++zdqd7j/KJDgqSVG/UTnJxrDN9gPkoVqa2qQsWXtZAsrYRlzpkoGPj1UtnF
YE0Yctpri7Sb48TP12NhG9SroS3S/6kSyBu7rncHOfS9LnXIAzuS2+PZE/3woo1ilzOTrcE48oKD
qzE2Zh3QhPIQM2XVETp/AOokYHDSUIWZJbNGR6nMmc0BpcjCEPHqBOp2dXLjVsxWRRjWbRMwU0Xg
fgwf10oMF8TWSbJRX2Ed0af3Q/23UvwzW9oCBmpXhBFp7Cl9CvtDV7dj5FXADfSQ6xNPBbquyVuk
GTd0FLfFBow3jDujvt7dilviAB4AJGKmsqExHMGOU6e4qUOe2Fb/9J6Klo0l5GZoPhnYTdoofmMi
fVX3lYDYWypDLEELAOoXXsRGrBmE2WdNIXqamMFLpm36OwNSN5zicHk2GlJZ99zhMKCEbRhKooso
ZRuAEbepAjtX4iqKtimm/bEq1h2+FQK7rc4HmyLMtvoY2vUAWQVuqKdtBX53QgWRCEpdmp/2dMRd
zUicx5hpNQlmwj/OT05jbqEemKGB8IyF3WjlT6df62wngx1BoEnPQu0DIPw9HNO0J/YJIe5Gg4MT
oD+KJfixMugCEnLaqy0dQjratjrDS4d2r/LEcSBTB6lHVayvZ4h87GtVuJlkR34ksTkTTtIoGtsJ
KqGE2Xl5BARObfLHG47vZ/GB/6MxU4aDKYjML523C9X/9jR2+jc/+p4KJ/ui+R0T7Wvglfjun3KB
HMZfXRbUcpxfhBHqhBgyi4SAiX97xEBWbomwqFTc1nNy2vQ01puR1GlcMFub+q1ysiGczPNFXn8C
CqJYMFZPWC6hD4yb+A8AwxvpbK79DivXA8ALSPD10iqsvL+jmlPuzZeMcZBdeJEdQXq7BZPbVe//
VAA0Qpz+zFU8Sk+NCtVooCrgahF0TB5IBM+99Dw4whRjoiyz1Zr4dg9y1shVkeG5TH7BA3I9COb1
0PC8OkUWRHyALiO4HZoKBYvC0k158yASoyi+XxQyLf2pWMuR4KXEuMtZ0cm6TjoAtYYx2ByQkeQh
BYJiWx+DVBIOZv6GfugH7o7AYisnJ1E+Tup1+QPkhAA3VC9pVYb4qJOFV3iYwXF04A+kG1HDVT0h
fSd9MlFasq1Ys7AHOi6Ut8+kYo4FSL5r6OBFDlZAVwLDEWH8AK5xgkkvaysY10EEnKgVMOWVCzVl
Gpw4FsRGJLJhybWP7rw7iXis6xIk+aYqO9MN9B9QhMKIWdbspGD6OjT4UMXXY0kbRLDEvdVW0Nnr
Y8X/crjexaJiCSFxq0T6NdpQNOpJ1whb84KrRoXRRqZF9wZdHyZr+HDOXHEGfPpY9B7ULPhPJweQ
Xmh9gldRYrS/h+aNyAYIvtBH45NkMEmprJ+X96tDkhRZC+SIBktrotzowQQF0k+/4kpmqxkB96LH
fpNRkCb4ZhTeOXBNg+LI6gMam8EPeaCvNfLhW6mcAwRQhtZY0E1V8m3maEDJIlI+W4YAtgNPtdvX
ENICjOWHruET2LWl9pbJyJfWCuop+JSAyM7LY7dA6oH9/mqgVQdrIq/ydcQosVkJoUNJqF6cAymh
g75O5YVMH2jZrSc/Zu+sTNujB+yhxEcxOcrDWCsBgzgVUbxIgUlP0BV+x4xt4xtSENRUeyeITmrk
4oWa4RU/NpuyLNG7VPjIeeF2f9TeNP4QkDu7lBbe+Uwn8SO5LC05gOZa4Pn7cmoKdZaHMRS0oOSr
k1YIiX3ni0+6RqG3xt87VMro0CduvNC1h4eMKy5WathFXelLjSPHaWn1l1V3IR0fytFZPDyEHCg1
aT8mWYHjYkdHRtfm5tKsyJvQ+Pk+cMoqWZ8twIGGPf/CBbOexVd2FaDXksNsevf/FZ3/wfg9jWEP
wZeea3kdg6j2Vj0L0tyPSQkNZIsugy9Rd6OTgILbNxnxF+dfsx0XcoJ6JEDlXGz4jlT0xLBoio7h
Ju+udxzcS/4/bbJWTkKXCgZY/3ZL4hCeFLj1TN36ttqp3Wp8PM7nupM3Xs2SKhCW1RzXktOkP2uv
45x+NNv+XXFtkDz2lLC6O9Gy+Jw5Bexb6q6+Kp8rCpUxmVfwYANKG+Ze+sAPbGfCclemoG767I1J
QjQmkNhvQJZUa9+9Io7V6xiF36eCyUMRZPCWGTnFg8VhYqsfFs1uDMVUHtw8uozhdjjW3gy+USFI
/g/m4P3AAYek/oGuhKsjKLWXGaIweVnRCK/tdru0irt3ZtB2MbY+zV6zjyhvvMLGMKJ+0lwRzPx/
9IzqJ+ZiOtM7L47zWI59sGS2iIB6RZrcxxz5dWTKSwEk0LlqrPh9R0N+hzXgIyf7woBHhHQVE9sY
OWdStHQF8seINxK5+5mpaPklgbpBKQRwMkMjprtYjMZVYjbc34E5rGrft4QsRmQxC3ZTp9Zpf8wT
v5fQtd8wkTdwzoXCvQpatXC9ZQA5ahT9Lauom8cmUV+xT5RjOAqZn3yRXtUZpm+D5y851U4z1L0+
Szh4XQyjUxISvMoFYJ9OUMR0pOhDpWftfJGqgaCxf4Zz/kiZwNxZGnLTbiN1riYjl6Q5nkNAYXJM
Ff4j0bNQqN2NeevwXBLJ7QsYT8NxqImsbCwtQkYaar4autIWH/EdOGxo7JBT1CbKDskBodm0icJp
j/suInu1G4idrXicVd+cyR9k4PAFc9957S/sAlWs4I7OvaqrqUEFB801wlU5TqLYegEBgig0th6G
Bh4IGeRm/WrA/et1uAq5eQq3Ocv+2O/p+mCU57/pJiJ28Av1YUFHv/9MRoP4oY+ZvukO4DP3uEy9
2b7j8AeU9/6M533DY1cm/a5ryFDBLoZZ0TBdN3ZiubVAh/tHSo5vuyUj+30AegjY8yzI+1yk9BpE
iWbwq/UHvt5FATkiczzR+P2PWIe+UXRcPzetBZMjMRHdiclscLrA9ddfWlB8nq7XDXNrmQbL3AI1
t4lDaKSyOv3mcAvH+am8vGHVNLVEWFbUyfkjhl0ZSsek3r/3SPYDReSSUrN2iIsVyVFTfE+t7oue
HAFmRo+eInGdsVYefgaAIygWtC9ZQuig2T9UKhUYq9OOv7UpKPh+CGs6rZlpIb0OPXIy2qI1wM6t
PhJS/akogHPphWfAlCMBvakx5kVAb2zFsDVKZdK6oEQci8HRYlAY6YOMn5+ZmmNkhfAFpAevlhlg
89/0KVU7ScONUb2j7atwPa9XNjK+mx4rV/5KPkGVHk6r0tBeeV5FH3I0ym5kLOY3BKfM0Th1nOuW
Kscdd6GOtlKEvjErj3n8C3rmdAbaeOXwGM4Y8erjNVHfDO15bdcyx9AlZ3VbqCKW+Gq3sX7OvpM5
x7A9pWhPUJ+Fj/jyfzNqKHD1TN5fZYUc+8cAR74wAojNBjxsS/FV/d95Yg7PCYmqkGCfxF2ZXB6l
DJ5bnaffYuC8/M2MA8+8Eurn0gbkbBFcT9QW1BoWhDZHK5bv6UkSmq0g1qcefkuXpgh5x3eoHjpZ
BvAskSw9IqzTUhrvdbie+Fly3APQZH4PuFjAtYlHilK2QC59xUm7Akb4g1X33/2fTDIxOKhKBQWK
/ATBD4bN/wSe20dAyAdjQOYfeo5q5N2RKf5iOvz85WWg/hiE2tGgP3Wc0FeFEQ730H+Xg/c2My69
XI+gDdHhlvZCI9YLKWwnnXJUzetsBKgJL9TIMz00nwANmIC6Bl1tnUNuPW/nJTy8/qgaXvYErUXA
aTepWRmUd8aYpC4Mb1tdfTIFmTMi2Wa9wD9erwOz1zSOAABI2Ipkg1D6xjmysivl5EVivHI4XNy/
FosDEuNG8inFA+kEsJSyOBrngJGFp0WVjDnnZOyCX6cq9i5KZdUNftlw51Aa+roCpqlStXutOhoI
hONxO/mKC3SBgZsXgMCbH6T9IZNK/YODhaV3I7rPOQnyBquaUdHmvMduRk9YOdpnBBev8PqYcIK9
AC+X9pyw2rXyYaF5HwNpLiYM4yF0Q8L80rY7zIAgG4oKbIGt2kIZWgEmH4UQvXlt6wYizcI+5t2O
d1ek7r4WAm337QjaaA20JbKPM3iJP6IxhtWgln31dZymnesKhPjrc29JtExeIyDoAfST2/DWWwXH
du8WzzoqON7VbwBR8TWbi4XZkFRjOEtHORnjQFD6mTrVV9yNHh2vIA3OSDvyXyqPMkRA47qK5kEG
OgcOGosS4OUGxBQrBf4bL8bPrrkIT+s7WCLbQNGBF18AlzduiJuxkMaqRYIffEN8dyldbCX8CEPR
UuI8Sx3TWaSss8UlRJ24owaSZNuUwmz67+b8kAFsdwvWAuYUId2FcGQilYSwX+Fnq9G6AbI4XFHO
44TE7itKJmKdMBU6UtrRpvLpLbhIDcvXmFccotWnr8eLBEheTG6dnavPgZGxvGWG8FBmXa2dJhRZ
yIXLGZ5JFvTTxMaCVjG/v7uJRxC9mYCsi1wOlx/qFDreVjeuullPYx6DsOPlFrDnSYR6+O0H0rJF
iobjNGh5wLMUB2v0Z3QuhzPqEKqcCh6m8KlLUXIjnfLrnOp8rdko0zugsyrL0lf0rlOo9OFze4IR
Qlvn/MTsT2Hh8u7yOBBQoifbibX4CCWJfiMqw/+qera8PKvUZHdkkKVHlqatZlTVCBoDd4UAlhMS
LAL7i2erkKDcCaUyprQC2HE4FMThV/TjtL1iKDq0mTX2lYYifsmk0tVnEhfEPJU/VfV92Qq0qj/x
PfpZTfY/AyrZJtc+TxKG5klsYMcv3wIdeVgH242vuU4ll4oYyxy/M1TWoPR4oQAzTrbD2t5F9F27
r474wDH2v+Y9/iaQ5FFybxuOFok9qTP109Tq0JFPd9Qegr2qFjpMnKlY+BfIMoxL72HX3B6lvnSf
LHNg05cM57tBoF4iU1Kl/e6u9RXTSvjqNJbwyWmyDZ7ApjB02VTldbzy0cC/9O+ZaTLr0Gpg3Mt5
nl0Z8n8B/itnwWEMmV8OwXkPdxyRQ7AdYJzopArdnvo9f1cBPP5EWkvkN6to9Kl78XgcoxnvM9Z5
YERj60JQdYRHTMXfR6acfG+bxPR94IanroagKec0QePJgfZjzbTr2+37+egGuWs7JyF4cvZF3uxw
5E+nTel8n2O8dwIrbIdRslXrr/YegK/GdPwFCKib/ORV74EPUD+VmJDhtQiFv3mAPQdYpDrW5P1K
DRm1ZMMTwJBq84ijwyXN/fEnlp979OREf05Y2/Qg0PRdvBkId/7WueYfLCWD23pNgnS3H6cQIh5o
88bzvpLPMUJHumkOQQA7l3f4oF0ug4h0XuhpvUAtx+dBqbW1w1yyEN1kDSVTKHUFF4024lgo5TVW
MD9LLiCkLSnIeX6oDseDar5Vilr4C+5Og4qtujAr9Cj7+Xkyetbs3ORQUI5caxLhKCTittXVyDhH
7AbaV08EB4oRtthHTyZ+ZYMky2hJhtdnPC1cQktdLpHJ97RDL5CCjDs5zYj8sbIe1i54/wJg7IWP
2PnnEesSAJexpb2emAZ/RtMN3ayntXyHcZZpP3EYKsDekzJ6abNJHOgyMQoM5Enueu9h6uD81qW4
POqDgxN98FH/E0qwOMqpI/XfUeflEMSbcnwS1u7cUUi0RO2i/vXNbnrigk7cSvttF6t7JjzC2+1l
BcXhT6+inZv5STMJ9HkoytVDJNr2RRzE0MHnJShB5ptslGkJ0+imtyRIIYzocrSdFh+DyP4mp8dx
KMx63b8ScdXF487pAa0+gpW5yoqstfP564ISgD7phNRViOsBDAqhQReYhMNmRN3fpvFzwSFvoVmg
i7BbWxSj43i4cz04Fv1cpBFse7MhVCTYXYPO7oVOJSRC4naUUDbvwvOWc9XaMH6G/AUHGus5k25Z
/DetmJEZAjlL011sXv8vV+j0Nl1k+oDqAFiMvtCUrT+ZWKpVIKbqhWDxEvAA1ILhq7haDOuuUg7V
UigQSLIrBcSDLt84BRA0KzONfe+0+jdtX50OzICEaCKC9vvDBde/JcCnm03v0f5MoeteLjlEvVLu
vNBc43sa0YSxEFlCQDATZ5m6tjqnEbtd4rGt2Gp7SDBvQqjo2FKpoIKgDJ/6brAupJIzNJ4EBxLJ
meJQrGGBUhWC0DSn+PaqqfpA4rec3M/KrF+uRYv//mZlLLnZA+kGsWNFpimcsyh1jjqNXK/jTnRn
/JwTcsHgrRlNop7jlcTftA8RlK2iPeOoZ7PDI21vLb8E7NYGt9dUuTMPF/N8axvZWDF6P4B74/0I
wYsT8YkqVCigmCBg5DLtjM3C5O70/uFl8VFXBIxsiueaoTQjYDOzgjLMTx/Ig32pLNCzLEPtTb41
SJfz8morp3EY/H56H4xoXv7RzsbxVaBip+hAu03QuKdO6Bk8RxYOKnV2G27fLzRgV0VZyZhdraFh
nFUJJuY2DXajZhncQGbfWg8ZNHT0nw3LkTD0UCiOHoeYV+WXWAYQSdz/E5y69XRo1GpjjPILmwey
vr6QduXHsqu8yvKqaXBNhWKemspflWfp4vrpBgB2voDtD9FYfX59tpshKASKE+81N+hM7k8gNtGq
vliUWvr3u06Em/NZ0oNeIWRexmlWYdEEKZ6AjArlHtUbHI6GycqSimNTHmI6a0Vifvf7U5BBFKvD
KNoGn7POBzfRhz91Zsm1tWJz4S9UZgjKSOLJqvSy4hIEaXgIP0/hssHCavN7Um2/mzxzJioI+UDa
ymntYTJBUx6ty91s3+TyvpY+7AG4neD4+YXhRaSdfNM3hdxydWACTvUBxRp8fJ/Guazc6UMOFMnN
csObvgQ9cuN5I4vTVU7li8+3gNKVeYXgQNZuGIA3IlFuN0C/FNkrD/jRRlRFDMx56JX0jP4zTxq3
Kilie51wbTeQQdIN2iIRw0dIreR24CHuyNHS/xZpLkvubHNpxj3MmJacyvqvQUzPF6eqyq1XaTho
r/yIqvSeu1GyUNrxwPmHxBeK4YVHH9N3ojwmIpHdVJeFhxXR6hVjRHd3L44lRO+UgCf4yrSiaqqc
03qV8SenBKylMjs1aU7Itrrc8oe9EY+Spnzk0WvjBWRRdc6N86yPCxycA9mYvaZSmNK5m4wYIGho
MSaI8yV2oeXIqn709rcSytM/LXXNdAqnpL8WI9U4Rbe9F1tNfjJmc/bnkjvLnkQQ/znYaWExb26f
j63lBN/lL551LyqwuhvU5901pYOuM4beIRUgl847KhTSuYJkPwno11fnLG1LT6y4JAg21onfnHrO
8g8BHaByZ/aTQJpjtF1v7+9zz2fAzDOgSv3/vtMowlXTr+CBx8V9dtJ5Kd9Jp0OKt8UshN7/gCNO
jLHSNhnuYo43Bw1aejX7C4JPc1nGJ9Rn8kZ0n1olx/A2O/546lccYzDYypoam0lyfQtTI18hQd4W
SjY5sA5hxogEbL3zAY2h0ue4/MJGWACj9FNiGlo5I6EIHVyZZlSAb91Y50b0G94ptyY8BxwsZqdS
22yVhcNCN9kG83oB+J1Gh7shhePJ87V4xq88R+ZZz4GK9oo9cibZ9X9gWycSnXdlpHBZMZLJW+Yo
/osmsBrbMxyRi06NSBMLhXKVH328JVSWspmUVq/q00fuk0k9Y5LC7MCI2pRRJZI9w+tvQKkg7L9m
ZFFsP2Zk1AzbQHdKV8vNbiFTH4SvY/2bm2jfQnyUmoILUoCRoap4nE2lOzWVaNR/Qw7hzwP+FGO5
5PHQGEcf+Z+jodFSNW9ty3xJsyCpvgRdlGmScVQ9/NRRFoPRB+IbBclnV5TULMwEHHULcuTeIWsz
e5fLHZGlHHYs93uc7aMo2gxLJYZiUkpzz2hYRbhTKhZpaMW9QVdJTsuJSmJ+/kEQe6RWx1DjawoN
5FpvaEFaTyc3kMn/dfS64xQ211OwXnZGPUMp0Vg14+PBjIJWvFXhrYxKzNgP+tms6hPnoAvNtv3Y
tIlvu0m5cVOYhQpLc+vwdsBQT0lt1h/T3ua7JpM7iz7sbPPf1jzGeskFE6e3jft6meqg52PkGiXu
br9fuT2FNRB3ZEG7zOWukk3LVTBOsr4FBcL4G2DUvvKhtgt7c+UcIQMYliTyQ69ljo0gHPcxijZS
k4KvIOEoyfvT2M0DP4ZfSj5TMIkXDECVZ/7ZUh1Hh30r72RI88oLXOylkxGWwFLGeIPhuS+bpAdA
eH/4ihObKqtARhDG63MFsNCJ/w2KWKK2zAK54COUA5UpV4UgiTXzPCY/ZL9ywdAa/9SvkfZOIfTZ
IITQC0IP6lIpoOqw3i0mXoBgdfnwGdrW6cFmNprPy8kcXfxCg4fG34o2VdLO5WkqzoTec7yPQMwJ
HRpKO02dW2sGMEpgOXsiL+lVGQQsMY5CDV5Fs2I5o/fa5D9P4r3eutEkRTxznCbUfgCeoslQ9K08
0gXlUcVq8tOYuzLp/vwdQgsVPgy7PgqpkJOgAzN3HWWyz4yoZPSz+FRCOpe6XuN2a25lGORAzc4b
dfUFjQA4v+0STSx3jcO+XwEoDrtJoB7fK2XxWUPNqZrMf+5pJ0pPBFCb5nMimDdawgbL71k/VK9p
Zzps4djtvXugQ3fCCka7kZzFY8ngJ4zabyZqt5y3IyxSZ4VB86sMUTnX6H5k/jNsTjp6bf9va1x6
X5M1kp08CZMM7LOQXIyIfheEidDLb3hqhr+aInEz5zkNdSjj8dQtvzMXAtqZ6yO9oBIrmGk0rJfW
MyDshaTZD1oo9+dfLSsTwRMONj9LpPZG1z9jjgaPof7fsCSGSHWAdhcWZ+20avy+aZXkh8tcTNp5
4egDqed/f4O/S1MxfJOgjDB6s1s8G6ZC8MaaE1vuO1Tp02+oFR8BIC8C2WE+DrfYY/WH2Xr794K+
3tkns7GDNyuyTKQwa0wQWdjCF2kU/eOZJzXbpKvySRJ50rIvLmKSmbgxYPQdVYCfQkJWaFmoyL4I
pewwBzKtjY3DDYONXJzNUFnCLqX9e1RhJaiZ4jVlYyhGI8dT54chrInk8bl+W8TMxfNvcHBQ6zxI
yEAlBP+Jnc+is+xr7U6CPlwbZ3I424hJPsgvyYF0rmM4YAIZFO0BSdRCQNRMRu9C/zSuYE+en33v
CLZFpCaHUPn+TzvFW9ic48/X9jijyqHaSxR4eK84r3WK9xUTndsE3vdwYTqBoJP5WlhQFNABOkHN
ns2Ei3mL4p+4f3ranjfk/j3MSMhrYiAWUbeDouk/V7PDvkOsmGlaG2/uSw69eX08HXuw3dkfcrXx
/zy34J5QxSlqMu9VlUjCZwSdDTEMMG1Bavkuj1PAxhosWnM2HRhTPVSe4YSE6wUCAJqJYsiBkgjM
vesurBpSYcVrv7G1VgQO4D7nMmhnlBiZ4+FoHvoRKa+ZxLpo1yRCC3Sjr2t8bYP5p0fQHYaekV9h
n5wAT0oDsUpnApYK5jOteofFd0Npai6hRQ7lTx7AKpVw5ie2u2tvKnytGwuGLy7GXZZKIg9dgEKk
KzTJ/DSW3+bHYlnBW8iq/oCoP/phoegiDflNHmtgPh+EFP8cxROSwJB4Tkt8SRrRvgDxbwzAawS8
euCP4+d4TwjCDjaTrr5O7JJvYxknaRFnevvPo5o+vBVbQZUwWDZtQG7ZTRUkVWV9YDM5+W3LZdY6
hQsAtT9MlxFY363GOOa1cGjovhE0t+hWK2eLys5SZ+LryIZR0kMFYOnezfbXLukwWN53cykwUkO8
nIiDOmOk+lrxGlu1MzE6Ho/kHZGwgnvDPrHTRoTtoDXwHyoo8cihuwiLC6R2hHS6yj15jQjrqmEp
3AZRcqJaFS3oZD7uMe/hlDlm5FQ4z5Jvw1ATzid24ZVs6G97b/yhS53+mKj4Q3bFEboIoaBegqL4
fuB3mb5WxNgjOZbFpWX+ocKFRWD0hrcdmxEIV+sAfQrsTZCXJU2ZWz6zOMI52Na7rfg9DRbzcoIG
zLjsBnLcxRPaZ08w8UzU7KR2/yTA5SAI5KxI5fw3x1JFh0Tf1PRnISOua6K28RHTDoYEkLXCinHR
bF4ImtOsdWSHBsTOwgnwsZP5hGvWIoMwobzTYRo9+6bVjsr+Tp/xcto6txfQL9eJmvc/hhYR0d8B
BFVIU2mZD9JEtVp1zKP37fJWYPminnkyZ4o03gPFdgaTkt6N73dkCUhqjzfOpQCzMw7XigWW57Oq
av1aSpLjBfwyFrd7kwpkttFJSB5Xheyzq8iPskD2/SfVVQNwtSMnpKgZF7HK8OXREKLyveibH7vu
UiPFp+AIoQ0zpHxLBp1hPy2vNuNdo4CaV4hmRhLavPMBrUX1oddwEPyDhMTSXQsshBUl7OcN/EA2
6Lveo5FD6ISmd26LX5vrH9iWS0aXg2zOMsf29J+uylsvGeGsuuURyBHWYMB6ZpfvGJ8UrNo11vVt
5iiR8KdabowNcX1xv/ORDSoN5MobPyoCscWnNm9JVuIlctzCACB6yqRRyY+GAx/DM6lf7bRRQ6mn
k/Pvby1K8CzwnbtShupyxMMwT8FUnb5/JYMT5bsQdQrmAPlhLkQPoJgfbmNHJKdj8r2RYROhLLYt
0QX/noKLoZ4I8qRN3RfS+TMNVCaEvfA6pKALrTtQeskU/BgnRvDMA9Rw8GsUpgQasSg6nlMGXgcp
NGcP/o0WzbxruvkbXhUqaW+eVcYyefRLR4Rc6qdS+f5ANMWgcWevRHBngqYaHCbZLrd8yr2u9NTz
MgQGzx/zWm8NlYiN6IlUdffJ/+CKsmjNffFcn7jHL4iUqGzrv1mo9aKzdX3/0pxoCoERXPw6zZTt
fy0ldPPtFyPqAergK5p5yM84/rhQMRFJKkaaxJyRy6Cc4ADd0eq2t8/Bv6oe3WPUUhXIEqBx9vdC
CnOaL8lzXSGvviLXjU7Mi6JpLECYKMPimRB+KFKIucuCc9yy8wD7S7KscFx8mHNmmRISrZyVFJt1
W+0SqTV0ZHZvFyjOYm+x9sJqtGwr6XPmNhjDg30ykYdFxSzn28tKratJMguukpN4+KhckBnmNo2Y
8WsF4e3Jx/yq/D4KyvqhZVWfSaUsesBR6W4FPtWo79j0oNUD3FZKT9ega3mclEq8cLNvU5jnCF4L
srMec/Oxrc1vhM9U8E2mWza6cf9Il+yciXv4OyEH0W9+6u1V9kiDyZC1eVabjHyd7B5xmQuIkZuU
vWe35PLyNawhC/ijVLYhejW7fhwTVKpVVVZyX6MVxmq2/L9MKej4wzabZdlaWECLt6W67Ax0W14Y
qkOFLrXwFk1+yMmE+IaHfVP6vTK5LLh1oJlDiKRHRoX/Dg1SpoQerZyQi3x0+oQVcu4qVjaanu3G
v8fCz8mhEKsQ0GVfyLBDbH2YbXxnQw/JiQdk6Gu43Sm9SrPsqXyUqpYKHNj1tPWtkCetlyPZUWCu
fGn4kvLI0yRzuB9sx1mIB9JUiuDXBDlfTmCDJKhrL2lvk6p+i8ku9nIWJ7KELM10oS7RkJ9THGhs
Y+V0PRzBoqe1+c64UvfP9DTm5Q5f4H78o2Kp21q+5ktYvJNtgUmeIZBQTNXuaZzCjc05Shnyjs2k
YWgf8oXYFgPyfx8EKXbSV+gnyTImqvFtBd6Q7OSdnp9lJuefHXh42tulFqrP4mFQEkhLqG2ZNRTk
eGjqa9BcRrCaTEBzi12k2VYdC959k24uGW+j1hpSz9G5juJM0q9oltlEqfhr6ZPwWK28cBSET8xh
ZPgZNn5eP891ALJ8Ca+IyCo+hzuWnuDrui030C5mOYg5+tHMN4vJXzvb58H0LPCj2Ij9f5dYbe8X
/Hnthzo7D0rmI8xu4w5Jp8atqE5AiGj3nJmZd/eGHQu4pJ85W22inwTanC3h1EPPO/2ZdxT42xBX
8znC7B1KW0syBKz+PhX+6w72bZ1ywLRnue30CwxJPPl3LQLl4xOXQ2Eo09L3qw/m3i75HzIgiLQO
KLmS6qHbznBhn0SDlMVgwkXkBlMY6LWGldA0bGEOupyNsdB8Dg7kGItudJ/za5Qi42f7E8GU2aXb
t43jov2byaDJyZ2BQInrpao6hoKBQqiMPlsWH89dqsEoDvMz2tHrlZMj96Y4VXedIXD+OKcclkcc
V2bal6iYswYCuXvK59DIjTm3G5lyzvnKlcp2+OI8tJ4K9XwUVHCcnkJTOpkprNhPwxb77IGJkZus
9k28Nj0srMHPLa9h5WXPjIYage5SIkeL4P2tBNGUxFcWcWjOl+2LiKGqHCTb5OvKCYn6T6gc9dqJ
4+uUyf4G7PjIbOFQaHzhl1RhQf7YDkANFDL/nOPUg9ZJtL2ZFAlgeI5wPh8K3xbKCcXtUgjncg22
LpAnKE2y4oTanf5GbGy1rf3WCmULmrPz7wXWgXE4x0QYglLhnfRjg+TsnQtLzZIxEumpMTTVBIU8
PoykL4BGyZ2ssXAs0V5fhJmXCrVxuSkmNE7N9EePUXlDYF0EhI/Aw8Js0bkKsUuiX0wahqny9y/u
fHX7NhyPm0AKmZl3LtOqipwCKQIcsnnfbmJTop46fnuDOiqUspTvj0bRwxr3DQbXINOoyl804Tfv
oUwLOp5qQGHCc3Qy4y1eYGMwnYQqEZyQ7RZoebo6dEiRR6XcR+aTNhLabHIAg8ilDvW+VN1kq9uL
wnmh7OaZuFVUK7uIeaMp0Dk8MHBWKApjQ0uYb0eYXbAXfiNUJYbyJ1nVpcndsUCijqKYVVlOs9aa
emLUq0Jqa1Rwz2buJgK/V/WKm/Y5l9XBpMvWvEeFwb9zElDsxGveswvEfsVUURGuLp8nEmnGY8Lw
whdnk+M3w+UQtCsudSq6JzObNsbgQnWAJGPK0wfDYVQ7JtU3d+joz6MLpp4zARWwAWoEULW3UNfz
mcuOyxk50IUrSD2i7cad8MwLBdfM5ihhYCR+D8vCVukThA5ziPVteX3yb2aI/wNv1l2mMhCPPY9J
6DKtnpVpO62FA3ndYPFl/5uT5lAfPsv5itr0aJ0a+PPzal7dGyJGJLTQuPnf7e/HuQSEbM0jWpkD
EpDg4pUfxLuN8h1aeVoUQTOvLTYg+HIMH4ana3wZhR8PN1k83gEK8KMwT+unEF/FO2BXTilOOp6k
JSe6mqXX5jw3e+ABf2oeakq2SOTor1Sz2Vme3U9u+3ptsuB81t6JRiI4oCSaFnU+I9hTRJKZr8XX
MxthO6AjwYRDAEVI1L+yd0VLKz+wJYmZJmDTRLGcd1DDC2DmPFmmdpRW8CohCd+Eu9RzmXyE6KQ6
oQMf1hQhqZXfBG6jMEMqVzF5tCf78fkVw8ymYxPBg49J8kAVrm19mp+lkXjIp5ruK1mH3yMsapZQ
IZFOMtqbXD9vSKHlEBiDFTPJ7dpApS24+zqtlxFSfGP130ulbxTI3qBkx1gF0n/pXDjkrmlivLmU
S8nUpdhmnJ/EZNxfw6g3RNvWNsdg8yYSdYd6X9z7ZP8oy05z73sar64B8FKxlSbcJ6rXpOrqmToF
P4t1gQBcGfmpG2oe3Zl7mR6bPtxCyTdVdAYdP4VXEpVhvPQbR/V91jO/tFxSqlRCssaV+B8+K9an
tulsk8aQsQoqea1z5SzpQw/9E17WYNhRycYgfzXEfNekKNKCQd/i7Pyx5ylWhlS74pxQJgXY6m9f
4hJKmYKFyfemyRuMfVU+Uf0f+B5CrtVrHSWFsy+h1DyFxZqC0J3SOOUfeKWUXmxtt9mkEiqPWz8K
YSHhmhdaPyZkLBKFJWm7ZBY9jM7j/odbmfTGPdlL9WeKRQkJFo9wINOs4EdT3U5JYu6F3hg8v0pV
MwbYdsFu5NeMWIEKjygRUED0sM8N+TZSTIWzjCtFB12FAVNXTWhF8isSWkc43KIrr6EuWhHljFsu
VUHZCffwVCShDvirNPr6mlPUXT77OiWHfMyrzRJIVA+OK3iYdAp/ELosLedXS6ew1EBfUKqO2dFi
m8mz5CMApxLwrAIgYN8pzKUYU/g6jn3L76/VTaAHhumDOBVEu5IwLCa7/0yFmSle2fSnr++WOTlX
hP+KF1HoqiLyhrz4rcJ2VfoK/EQcrFD6WGT835EwUOtqZ3FnaY28430Wm/jox++FB33ErS4XtBBc
bFdtPVbFD7idCHw+83/A9tcFloUvKwiCgUSbOfdm8swfPKBaUq+46mszl36AhtPGwjQRnmZji9zR
9kc4jw+TISEmkkVqQ6lL4ue5zoGvvSu1mxvKEWIMbpX73Hii7rVCxFZzt7W2TaorcQ89imRSexuE
YQ6+w7Um21BYh6x8BNDSQ+EDIs+z6no9mUgkppsRF73xQB4VBv6Ey41rNpKNkuSLF24F0IgrTDSR
Ay/ubq3piIzphNLR1FotZeV7mvgEPbujrtX8JAetWSjkMQwYmNyp+Qs9PaPg8/6OtmahRcCZlPgs
C4YykOGEMO9jEG0pnrBl53AbqSsSRHw7H7y6o4ZFZSICtmrxBfcDEBlemOdvcJJujDYufat23K9U
5YHFp4gwSWLZedGmtiMu2IKdZzIvvx5spAARAaWnNizApa16dZQGyGdPmwj9ECKwLQ2zp4k6L488
I7I5ouDEoF4DGkEYP2BSEVtAiyf3w5mFGZiXOcbn3nAXfgr1q0laIcUdelT/L8JB0kIFN3sQFWII
qYS1l8LSHcbQiSE4k05B/ThSf1FYtFrDGXTG/EsiVWH3ESf527/gggEVOsdJELlGMrpEEEFDCRfN
6h85mRyBXf9dp70RaBPcdvMYTmhdQB0qhcdbhJIHMJNlxEFsxMC2JJ5TI+MZR6mH+hAWRjWZ0AQ6
YyiMD+lfpc0syF/3cUN1u0+M0SVvVvGVbhwx11m7cJenYxzkLlCMB5uVACAreKCeiKZRpaAzjLvk
KeWuKfKs0GQg5sKKIASYkLSBHtdOunA5bwPbQGnAyeXMGQaANdqmiwNlbly7oQAa8RR+i/TBqq0C
B1Mqi+KQXKG0M+JB2ft7K4j1wywucnwvvdb2J07Huk3bidOIHU5v4alMIlNgB0gW47HmAzEQXuTp
SR7zaFvOr1phJpj14QwasVHZbFC6fJ1e3ohMoLpq+3lUvJ0wDx9pZKVyuEI8oubpEp2Qtg0jTHaz
APhT24NYW9RBWyTHeSKW8fHg4ZDiERwF3oOA4y5LtdzsI9KlX2iVO8N1r+vW1rub/rhdDtDYB7aA
83LGiC8Wv90WpN55U2XEo1+oPk0j0eZvWVGeGfXSBhUX0Jz/SU7hCqCKZ9B3DKi1B86H95OudRTS
3OR5AbrK9ISDgUYHAbvbQRRkpIpmonoL8ILzYwBJpkltJ1scMwAoL7D0OjoRXUN4iUg2c/dHIs1f
xR0HyHznIxXR7w==
`protect end_protected

