

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SFpyA3WDAkH/h6gENMNzEC70V+GWX/AuJRjC9uuhJRzuSJx7LjCfMePfd14YnV5eJpUmzZ71W3kb
9tnOI6KXTg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FappTG7uNGFdZRwaHkH1xaFvi8BC2aKkPLd6PQ4xkTkeceiv05HkyC3+B1zcjatywH/Tgp5My5jL
RzYpXDHCiS+WLEnVqDpcElLtP6A/XLl3ajXqKvZhmMUVZsEI6d4wI3wE8drV6caY5dK99YnGiCxy
c/wD5JKxsx7IEFSu4qs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LRNAkwpKrud10Lp0Eq/NqP5B49JnJU8WkULh5UDIksixm1tOfz3iui+8sx8gHS1R0x2iJMsSndD1
7xzPuxZn4a1eVkZa4n4EghKA1iQCL4jIUagjOF/A226osIvTkxPBVZ56YpbMiMwMMgRLER5z0xet
LPBfedO96PfexivUiLv1asz99hmC5fi5UUap1VwJdrnsIHsC0bEW3N+9FFvOSldno8glOl5txGSe
hOwrv3syYadhoBtySSxq9fjTH5UTCT6nikZqZkVb5yhHF7eaz/U8CnmNnm4+vrB5n+GG7KIVkI6G
7PqaCstXyxVZ0I0FOvUz/cqAZvJcffVN4NdFGA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
u1B6Vk0Eso+5EvY7kmrlz1476LggIIsaO8lHvFGJ+HKHly0lYN/LsIll2vy/lYtCwxTSlrDsJgNk
NtsXioC5DfcQQ4kEDu1f339J7HYisXvM7Lhemt1gBNgHhAmdUioIYx0fpzcnzuhwqs4zH51jdAXH
PU3S8K0B/J5Gty8ttFjVJwRIoxIqhWdYqBDiUuGzr/SoWf0A03jx+7IJtD5tY/voAJ5g3LhC8YQt
AWy8nfe7i7XNQN6Y3WxajBwMrXsrAH821hCM6aadbQ0v9Rva24HNcIHmfKUDspzFekOzU9yGfpW0
fWulISNFKBsu0+/BoJRhSZ+oJMcibfGGrXXNCQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ufS+qjgKdn2oE3oh7EcYzivo13DkHjOXZdvg+7gUZzbjFQGb+M3QU6lNcH0LrOEXll22KbI2ohfG
TzYR0mnCNIzsPfjq3uw6taFIWJM74+oLYtSXEeuY6ANmuCGlqaVPg2smc7PFDAPdH082wsWirRmd
5thR9q4u83J5L0asBhDI9ZTgri+q5MwrlbJ05yQiFPUliJgl6amNWt26C09sTCAwIMPW69iBKeeW
4vt5DSJ6XyglFS9MDI6DvF+Cy8vysZSNzc8P7lm9H64JZqo1p7yTgGY0TjifISAPXC1fHwrwfQXY
BsZz6suWdJqjyzpfb60JVTQ+/k5D70Xj1MXLQA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TI2B3m1FrAeKaU6k30ykyHfDnWZXVLw3GYVFmPwE7PU79Tu2R5dzZ8wRPsdfoPSTye6ipaIAsPtr
CwCMHFOrInoC4tES+00nqn8BAlNtkgIns4JutCAsylfO0tbo1jdQM1s3ZfLRmzO8TErqp7qh34cJ
cDScSpPoqwYzQG0FgIs=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pRy8ixMxliZyP9cGiEmLhkLpE8BPUs0NUJLS9EUfKEgqPIYh3TC0iGkIkNMUl3FvP77e0IxaktFA
/jqS+a9b+rZb/lQQUSJMP1pPdZyeKNO5EYTlJkeq4M/QPt/jHeYrB9fa/fTRWFaLSO4suMctHSMB
vZbG6s1wo4stlPecixWiLDS8vMBqt9xY7MLA6d9rFSok/TUkwwve+vf4FZtQpUFEhypIh+/V1Yj2
bwgtk5lfZpX3tS8eSCYcpYqNluL129jpVqEYjJIDkcuxvvuRJPiKMpRwiViOhJULCVRU7pAOu9+4
kiLxod5VBhsHJGbgGwc1XTZvGawHjedADbu7Tg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 124208)
`protect data_block
GlBrxHplPNqXezNKT5AYF3rhULvbjvKXlrvHAmOnNgAL8KA2PbuI+aoBaQhe5K70zJnWcgA/JU2I
KWskhhT/7HeomAwXnv+OEsitwnQJFXAOw0VmJQj6wk7Y3t41sGaUyqOt2S4G+mMIpymUQZrei+ba
PoJdFaDqSWqRXyUHE0NAqdSWDe5SOHNujGXhnRfRqHyfLkK6hrtaU/CEj129OuvFwOAtd+/VsD15
4qVKdGr3RyugyPRiiCcWFJUgqlmIx38076mJO5W5t4NPACcAsBT10jir8tDgWLeiIL4qnrboyqTO
gVDJzwRrZwVX3o9g2nkUykrrEmv8qoNgmy7VbhF8tsxbonDmpoCLyEVNiK6epWD6KQUerrYHJ3iv
222Q29Cl7SKlSQDqfKEeFRBkRwP7QhCxu5+JCprsyzemI/A0AL2WtK0HJN2sXHHJnNil9oFEu11L
mogZA8wdMB0XJbXsfNnis2bG1tOoUBVujjxyNvHgNI5oIMqQOoeWTyivpCbLUFVAhvSqIHRMqMKE
bNljj4L0RN9m/7nntdIymFNMO5epQztdpbhn8JCA00ai4Y0ygoJZ5ur/qPH3u1OnY3MinT6klJ6o
8JCShNdgPjO35kMat9J6pMZUMb945xdR5a2WRhosqmRrNXWhYHEH9PH/NeuV1bZcKwwhGO8jxQaD
oQqt60yWVp6/etSHsXWdKB+F5lY2euDz6AAjgiwwyO9fRk3r63+nDjcIAeNil5+RI6tRaTd1VYhu
RSPmvPN3XBT9NaJD7PH0r3atLyRxTfM4qI20s9jelYEn2jSpwHPoyJQZk7ogk9QkbAXDAJ/BF4aM
0FcfCfM8jh0XI6ejSzFJAOyqi3oNcPd7Bec8axQRYYw8bGlMWzE2Q5HpFZwke73ePJMn2qz/3Cj7
lRCjw4UCYalprVj7LBf8fJD7vznQUhTF0AOYmgfAjwV2j926+HMaspNxnj7dORUmmf6z3K2mUGrb
GO4heClxofn/1FLECYlaUfo7z23m9jt//kz2obLnoDYVtrLNIllC2Wf5GwKYQNPlsrunNBZppqlR
O5HOdliSAiq+1oriznLXtS9JnLj17TLeWtOS1Ynwati0g6AI7i0mwDifuwHyHXG+IcSEO5QYvy1L
KAS2ICu4xscS/p7HmSTh77q9N3xsYPuHl/EaB5CEPa4W8oAbtBRv0/MEBNAnaJQ1Sj/rqYtPPfGX
edMxK46qRdlutFL95/U842HOrWpP53QB9H6WB4z7psGvuoVZOr4lgFP79b0Pu0LrTENWk+DzHaxZ
4zVs5tZ8L8rtxd+YlEQwMqQOdOLGr5vasf2jdPEwFfDq1NENwZZMTAxYwG+ap+2vioiSJ3U/KvXG
Pa8hGOwSnr4dfIjQ21AkEjXCBT8+BPuzjxpAuVKTWJnHqT0U6WVTGkgELA20Fez1nnLzeQvwm49g
wg32DvjZWdaK3jCukUFhDtmsUU1x+SzXxTlQUgpipvUIdh1NqTIIUJ0UgV7IRDDdNfXcWmSIuKMt
bfvJUVqVGylYAhIVx9/2Qe6IhpAwoyzXJtQWSY2bejrFpl3oRIrshKoFcU199Fx8ngmDR+H5AAIm
MUxdLUpkCopR4joZLkrLcdlt0hs/53OqRqsWSYWhCrZvziFJ4nRHtfK/cqyBs5RujcGzr6xwZcTc
KiqMhaTrzMZu0TMPhZi8ajWCGHkM7FnWMarRCBBWjM1A2xcEcT4oB/Vp+rM3DKqIye768dp5cc9N
02twsw81MAywN8dD2Qdyi0oB9ugrxfOBEXGIdE1DqfJlscod8ITttx5czcvTnNS7ygW0EUqvuX46
Bhp1CMzq7T878yIoT6RXJpv1bJcUF3Lr4CzSNwFrku9v1PkDN/G5vg075UakfgSySGRD4bkvQmBj
Bgp/PwD/7oiwcz/qb8Fqt5CvBcr1CPp+iVcGE128NhJcZmBQFbPvY1cgm7DhSPAqLUoTis4yduh8
EZJtFNr4hYKqEUputQ6CqPBPlaA6zFjZdHJwR5MppmYodaQBKqVKh6WqufOI1V4RJW55vRfbSKqs
RooUZ+P7oTz8HvB4uUCtqDpNi22k6qvJDDu+s0xvRKA/A2tysxZPAyxaMNtqQ8J0m22EE4JEcERo
BpHwwRfX8PDttzIyjv/3QrggTYMSi0ZQ7n7d2h5+EblS6py7gGvbQEESS2SHnCqySIDoMxvYnM5i
ZadbShbrbOFHd5/Y/y63c2rEz7Ya4lgTVzxHeeaaU3i3ZAHPID7EKeYLiHvthlFM/1m4L8tEP5Hc
lO4ocGquVI4dvUZDYzSFr5bv3vYuBuysgw05frfILRpZWVMg6jl3kUoidFFmzElGxR3E+MvhrnWN
q/DY7vzxpuh9QijmaZMjSQPbA8OcYZrQBefdyZIr85gROUrux7M4WdAIlpg0RMi7spBIKhFKe2eI
r58TlIxgQWFZq8YSaVUIa2ceyA4SC3zKDaGWvaIS+5lv4fyinuv1y3PjwEPAfbqo2aDxBX1p51RM
r7Hx4K6xTZSOHiVDoiik5mRMaq7iCsY94t/wi5Qna6tbYWrFvQnBPE1vMLWKVnQAPa/B2ROVpGMZ
cPdzXIbwfwWOTZVgNvF0p7dzA02DluyTEHe5r8hGdSik1n5hgsdEiQbXDXuIzkv0Ire3tRHOcCTK
NsobO2zePqe8LIPbwGT8/3VgjzB5C/dm6y4xkVwNXwln4lcs+1YYzCYexGE2NUDx6Lrv0rFhS8Zt
ZiGRqLPSX3H/HtABWGuNLbV/v14uon1vtGg80y2fRZZn9OKYItOCtEe4Q7V9ryaPhIsCWSDvH03T
bktmxJr/zERoHSONsqdQ1ftQN5VyIntZTEfR/H13wC32H4sEjkR8YnrKgDkUX7nH2ePfuxv1BLIt
fpFA9uNAeSURwGHXD85UW6VRKm635oUbo6YjvAsBQzdBi7B6GFJBTkBjFmPeFid9BV/LlP49WORO
jYYTrM6mCxiP0LIPx0AzA7BekchYMhmaoH2Qq7xOr7tgZUZHMGTF7B6QpY3X2xMChBFqnGygY6oa
ABlcZEp7tNmeP7qnt5XCzeHQMxX/GTK6vE+u9j1y3UChQag5+xUIuzUO16r89bEsO07q+XggiOth
JbdO6X0bJ908dCe8Uq7rEdwXU9VlCcgxPwTzzUoSztupOcOntTnW5/nCyz09annqwZh+e0k1CLbD
EhAEn9QkCOVCENaZqOLAqdRp6qavvNwhbX91E2IGI1xEE54W8VseC/iTfT8u18kBXljEDESvDN5b
C3tbSp3IPAimtmGNFFruoi1D7cfryQYvWcoN2GhjWQKFhG9bT4d1ZZn6E5fM1/lHUaRNMGphPBE1
bGVnsAVssS+WLkc7ZC+NVe+XIc38K6+mpzFDhhVovkWSOX4vRmSfMGGQXKZ25iRSRj9yw/YlUPi2
Begf6x0KvWGHKTrt5FEkZGl1Kke3kVH42o8i7x9i29Y4MjOT1zNn0brenvsejCqBvKuFLjwQoH0F
YmjieUirZlKd/R6zDegGunBgyERmrWestT8nS61bc2Gf/V4M8w/G5+ICgEeQX+MDz++CfTnUgG0y
xUNWQiVWI1fLUd6MzomupFyOsLrmPUkVIsh8oYftNrVdfX8Di5YgG9XgljcjlD0CPI6oQ80YCjwZ
V6VbfaKfqOOMrDTvcDGveCjYW8fTVDpWw4rrXsek3oi5lhPHrvQs8j3uwzUZME5k7Dan3sjQM570
vVzLUHw3NsavgbYvWJidzcn/HY/ePYu/BOYc0c6O9fPR45A9MCvEKQBV4gkJQt2v1rr51WQaRWP/
9vKtAzyK1BPqri3D4fZaEsQh4Isya/Mtt69L0mlxJDPI1PaAXujTs4ckNkxu9r6HpzatTd3h+bWc
8UeBWJ9OkRCz19HFVygPFEdcsAeNZPXO4fHg3pqJOUP/FhNbnQbixITuJlyYMA8/qF0ruUqFJI5h
VQqOP/mKdKYiWZ8urmU4NPoyxBypD5EaY74z5OczYe9fuzBZd1qFA4/Okcu309HeegI0Pwr/bhDB
AIX+BeHnTI1wPjskT+aNYOjKgwiH1SYUNv5n6SN6A9aiDwaJAgUMmFO9bhSjxzVeO+7XHYcL9rnw
EGsMpzrf2mr5WNHYCV+IteFVopJcnklaGT0XG4FPndi1upKwtkK1n5m/2n2QXJVqwBT/n31wUyVk
KCD2/uWSBZ+pEs1pYOHtvpfLTrmRCd4ywEbT96u//c90EYJXVnd4f+Is5v7K8X+gdVAHH00Dons5
hLS1f27KvwgQkzHnuvEqe6VlrfyU3tbB1zOPf/IzUlvNM4LBMCS95xmZemvKhyvh84bb9WM/EmeP
IakWK1hybTEtV9HKc6CYZXVkqhpagUji/M3z4hAUqP5S2Pv2fwP0igXxaYj7QubXZ5p+a/34+DJ7
q/tQm/oPOWg0oy3w16nhUjRzO4DyrYprpdh1NEtMupeQGRSGMe1XA2mBW4yU0zegBhyqk0ZHvEsJ
XYjL3KApJdVf3A93DURO3CvgPA+87WHLy2lTISi3TIs70wLjFHxfG552i8Q3+48mSJNn6z2puyno
e01V+xLp2KNgFjQoUlnytIflkPe2/FxblrH+Zji+opHfZQcw7dI/2ARzVBLOUuhcYo61qW4Y+6l4
DBEBqq+66S5f2b/q7tN0YgmBqGn38nlOKIQ3uaPoYWUf4K41TK6HFzf5kA72L8LklkTBKscwpqRD
PMZpdJw/b2jQZcCRERRXEcCMcyVCmqVa/WBYbAJMMrMfXf+vUj3JYXyvZVjUEHKwtyTU3e4O9rjO
6giakkx/GlDOQCn6SASLU5d0lz5H1t0fML1hrO7PPcmaoKxKz+zFI3gusNYyTC+Uiuk8BipvW8s+
eTSyzvinypXvnCrRVF0Q2Y78RxOm0mHQ6tbSeGKplGVgfPvL6C9KRf2oRCCAvkO12GLWmRUMhC3h
IqVB0eQ+awkxmzLKJTcc5qLqbrMU/pVzLLj4TCxO+QVFj+Rt0lJBSNJ9f2AXuzhnUk6Y/rRLC/I8
pd/3NfbWwsjWpP4D3mSqUlVJ20cG8tjsuINwPFvJkMqt6MkaqJ/iWeHsZvhhAmcEJvMczU09cYHX
FTrvE+6Sq/Be0XYDH9OkeZl5folIxWfYF5dliKzXfX+6+dtKGnJuRqA9ivW1NLi6q23EXq9lZsBG
gLJRCWSe9RXbXVkorPKOwMfSW30v+mbqXdP3BhrjaTNbxxCODNu8lCZvHjL9atfUfNs/A4+3YxuB
V55YaFySixwQmGrEbIZd8lTgIHcLRsUVywq7FCt9xJ3LIQ2UcPfpHxq1x9AsULhVrhjH0a9Jhh+C
GUS2BAAkGdSSk6MUUMAW2ECKleDa5gvcbrh5q5M8Vr/HgLGc5ZT24no4FUJNUYu6jwS7iH2cMh49
3jVJ6SxNs5Zpei8fvIH5rGU+JxNEfygbd7mRya+8FG/YP9ZEeG5wAJZbG983NSZBSmYYegZ0EtaF
WOKCvMxE6fcYDrmbDZtBpPbzjgNjiubQk6ovn+uNw6PIkKV6mqIRLVJEitCKctki+n8WhLT4Y86x
SPGWqSQ3leEThz4+fh/wzB+TxkbZw19ONCPr2Fr3268Xcv9PO25IBX9VgtyL54zzvsT7lk1bsVmB
TDsAyw+8gHLzMc+uzvTM5hnVID1TvvKiG6R2gZBXWhxaHixfUZMdvyIlYaXk6XB/kk9IAV/XeVBh
stkDbj2AqC4Fe2f8PvbP2l+10DKwbahVvs0+lo1efn1MzkSv/Lzaks+KUGdLwvs+lyscp6137o/2
IsTorI7N2SANvhBrysH6W1I7YMAEbSkDZVEu9j9dheCgJVk16AW9w+dGLXO71rkQwzEQvrISktVa
w/T8g6KuM6/kwQQeD2jS8I7mNRboBbCWzh5tczzP/A9gDn4DzeLf2eJAPOCNhcXmRh63Ty/yMbfW
Wyb15pjMqjsRKpSoFZ/6iB4QxtTjTOglHSenBhU/+tC61GxpjdOWFDj0ewGuf2j4mVv/jtNmXhBe
wGBwcz8Tho8B+ZwVFOnAJqLfKgkYsk6exidp8hSZWk0KRkwJc/dfRWJ/FyGGCpvCvj0jXLa13XmY
nDmhz/rGlrj/4T0hqoNl8ywC1vjTS8wgqCqHgfNRc+qNMFZ8z3SsaktIgFWKz3kA0AEmRzvlB2hx
kQ2hBHVdOMQgP3oTS06md75FetEfYf9EaSA1K/oX0CjdEFbTXNGZkl/Tc3Rdhcgtp560lMqdVTGz
sjp7i4rD3hvFUCii8wPhegZMvrwPj02ibhGRIjN/uXuEcfsqeNmpDu9QCjOCNeTSVzDzVeNb7xqX
txadAC+B40MMjjxT9PQOWZzyJnViE4uNTtcrL3XxQ3umijWq/NF1gLrF4NoEBmk89QHvtlhhxg/V
ti2sBt1j9IWljI1fsN4yeCZ9WL2woE/Hi1PHY/WDMS1UBU7IsWaMGvh89C4JorxG9L1v0LcZJt1d
FzqE/bwO0LYCGGHYCWy1DTSTQMdkhoM6MRKuvwFznKr5APJyfHmMhJydaEiDkATmo6/yY2UwB0qp
aUGrQV5n+mJ+7LtKJ/7vRBTtvH3xkGjVAgtLEUOlND22WxFR32ZoE4v1tDj7LzBPrLOiZVLEIMAa
PJN/G0Bh4PS9joUzy1/fJlkUFKwpodif5DiBYojnnEKeQeMHfs/6Y8KwQhFGGOzT/xXo+NiAABF/
yoFsQp2maVLFOdb9iZ2JBVcMA2hyvpAThRFBvxujezrNwoyFUKCRN+W8c6/vE7OeT9hzzhvWswHJ
PsuBoU0iynXd3o16MiHndBog8h/ES6JnZNLQMfO8oXZi2+74CF3PDbBmS/vX03C0GirDBmjilLmz
WtNqSNcOUnV87X1kGoGAtVBd0BiR5bYciZZutT5eJqQRa/xiWzcQ+Td5rZ02X7wyK4aqTxjd/pjE
PezTu8uGCXP1w0Xi8yzk0mVaT5wna/gkK4iM0c+V0vF13qYX1nUuOGJTYggvZrkMIX1kZwqI29eg
Bh/qYkyGwjherL5rLFPwV+3O584RFwBnXOnP0qLLpJgR8GIimpxfOJ7gfF3zaz/pzIkeiciCDNaX
rBsXNBo0dNxkLX2VtWwtgXEXgG0Tj9Z9WSQ2/QkySb62njK6MYTOVTEE6AmFZJBmBpA6MiyciZMJ
VkCMSanGCBbd0/SL63xoREfGfAtmm7Xa99/lI1ghyFT0lbHmmPaXMs/ov1A8qFNGHLQ9sfdNUGoa
ECmY6oeiYxsB9H9WqRKZM3a8MDedim52h6ZZwX6RBPMOOS27zQXgEp9QZ5hzxxueOvNONRK40rna
dAyOZjC0wra6zzgxQe6+OWiWrTCtY+cX/S3iZ+r6uhZQ9hNx6bWQw4qlqQbasQ+rJnrgOg6ahnL3
efuTD3ki8QsM3SHB3OwAJpRVBO46MgHEZOfPr1fMLSpw5eEsss66g3qSewWZLLF8ixXJ9tjvfzlv
goUJuwkD6pvuMJ0UmTxB1NxyHhHgOWm03iThxkEY6wwfudfqrrGUoi62HYMcMP9gVMlzoGCBnXB6
Lb+EnBX9BQrAGaqTVYyzv/G/qv9YQFf55kWq9Jn1Ki+vV0aHncydw7kgXAhlQ6Wngxv1Cnle7qN1
1ZYJW4a+N58oHju1smagKA3xtGKoTO2Cm/OIPZE8eI43/oi1eMPZRrma11q+HZpsg46JpYjTwwoW
EN6CalmXRAdGcaFa5JI1AElfNf39FEiyqapNZgbI/i7lxzMTVd41GqqP7TC6y7T/3t0k/T7OU87W
Hwo+/8PPTcp4H9WOnn4f2Z4QU+hJJJHq4JIfdbpT/zhsvRiusPEKNP23IwkGruNh7dkDw31BK0cQ
ficqW5FoergYikyHjWUwMGgwlBSnekG1LRtfY6IWiVHWj9EjKVPULvlZUrNdE7lPLRgafbZ8z2OY
NWor/mesEnCspvW8GmjPPjxHLwlKnH3GPQ330BZ8V6ZUOh9Ms1//XKScEZziCzG3TQQAFmceF7DO
olrMm3xFPuiDyUXFBzNGeFJDfv1h4r3SvTBvDliXe44ifG+K0h4ok+pARdw04LR7oFSfszTY/Kyt
tFdfodn2pY5NTDPhGPrGlIbB6TVcMrmFcx1VlFs9DEjOcMQO2vfrPUfy14+DitigmeF7FFnWtLM0
rfCNJ+tKv10WBtahuqBykvabLxlV/WYwLrmzFGslvYcWtgy47JxoL0CtrkYfdKv9SGPaNdqBgopj
7InEeDz3OWqcBssuf5GGi+rxlp+GrAiUcjXsOkKH6USFiIcrxxyJHjGQBuWgd10wVhApa6cW8uyk
hpddC6KtEHPLAnhc+vZm9IWTK++ox7xngXGdcjtWw11+vDCkrqS3uSm4j5Hl4+rLgy1WzKqo3wjf
qzv74YqkYTw2WibTqWs86sxxLMRHpwBFnYfj3toC7RwYVsz3Rn64bTBRcT61b7IpvzqhcMEpuRWz
l0Rp3IlGQgzreGriBfcbFiTtJcg+eOZOMpD4Fz8LPa2T/e9jjxQ5Nnd5fWisFgR4hY3rD4o0PgSP
/htCi4hUPxL7JLWuhsL8b6+VZaMEZcv/8+q8doRzWXAfsbUHn8Bap1HBd+oQwmcklSIO450Ylfen
ZU8WnfqaePNFMSK/2J3HavPDsNboaC+2Vuii9eNPLeHj+KSK70yqrqiV0hrQasPif9j86TZ9F62f
hC5LOr4mHCvktL4cAkCF9AQRAvK1cHncleoU781lbZ2v2MBCCuNa1uvnoYQwXFFjh1HWG5tYWsjQ
WdK/c8+knetJRdjbDIUJrR0l78REcZAKtDnFAIV0oLlD813eouSbfE23VXK8VUDR8Ufz6hmxXEYh
uZCzu+jZF0zpKejMa5A33JLEXAXxkABmZFh86Yv9FdMQMLFi+xoSABm7rkLmDO4JWcruE3knn6NF
i2I0R0WyJTq98tX0Gpy+CxZIf4TfjCM57V/JAm9eFeasgrKVcCeTn+bQ65/beRfLR3ebdtNsqMg+
5NfiMzz/kv8H/l3pCUXkelZ8CA3E7n+v7piJfI7umnMQCDa0z3yCqBh7SQ7R16bmZwqTUwIsS4nN
RhxIqoNLaWagfHT2gk606iXXUwrUtAr0d7mh9VTTI0ZEHlnHsgnEHhVbqkX0+BcLsUfSuuBkYPBg
5x1FylFZcWNM+clg+mKKU4Kf2nuKN8nKgMlsMsmwal++VZQdHX1Cfhof9SAjkKg65x8ptJuspyLR
WzR9uiLmLaKw0CDaEjfGdy/oLJpWN1PM8VYl+ohIB7qREeehSnlPrhg2aDG2CbjAFWG9PhWuZbOD
LqEfMs2xBwcj+ZddlIQrYa3cONHDtiJ4gf+hKmll9V/1EgS9Ycv0AtpeRdtNtDs4WKlycmKTAguY
xeJHrbqMKi/a9x0wtVMuZAhmg7FTWgZm5XXwmT3JbjlNtKRr6wxPyUWMt1Trv2OvcFAK3gjrNpzn
Hv8r3I2M3E6XZs+SAm00ZGjvz5UOLTgpIxv4vtq2sIeZlex9BD/cQ/pihV557wjztRaTWJd+kZOs
Sb0731ytbkEvhh5izLPvgjOaSU+sNb/oRUdZDx7LCr1Em//QORWOSBrIG8HNJWcwJ4bWdApo458r
WNsIGFVsJDPKRbOew05ZGc8RWEMr09fpjRa4FGlNUbQQWUlfF8bta2QlFHwfrd74BfguNe43Hpzz
itVImRg3NwTt75AX8IrkFMhSgj1N6QaX/eScF56iAVryM/IJeAKFziKtXRtTWlZ9qLVwaMLNYPOT
AjWYWwml4M4kHwB7Yq/9LJd7Mu++hZ/Vh2nREI5+6TXCUYPtcItt67O2IjnPieL5+qt4lKvv7bX9
4vIf8AUoQqz8YAmCJY4vnKfxLqFq2NgFSyIT1QyJwtUfm1sYkw4gE4PsHOV9JztHQO1OM2V6L0Lz
b7HRK51bB4kuoUlriGcnWvUsGHrF/R0Erl716Dll7BdQl5/9/po/jyn3wYBF5LGCA+Af8AasuGv6
JMC56OlZbSPKA/yCJOk441ieYFZNCk4dZdlg0uFznn6Hbc/YqyPYD/K0c3SjsU1j56pjfz8yv377
LsIVrkAFRurvPznjPmfk3lQEYdNxR3i1pi89EIPSqmGf5hA99Hi7OXmoUZDyQZKMB6jYWQhMiU/+
8QXZPjsZqKf7agmZ78DUH8W5oZNx9ug/cyvPFI80zaT691DddosDRzAXJ7xRlWREbnw8pCdj95/y
6TWK4YynUAioeQHL5LraHqbAba/NQo5jgS6goQMfoADr8NCQtr+dkuJ+zVazD/1zOsmP9kn8Tl8T
P68oLDcaByU3kt3cJ5vgO0E40LTzNS8GaBq5siAVjipjJwOwKQEvctqA1YcJmq+60dBp3OT6Lusc
B5Str8AUSYw0dHULpvJ5uGBHs+bA4+iR1USBp6qx3u6x5+LoRqPXt7VCQxK0XMTnxHg4At1M8Ytl
0V/16kuHghEQu3BtWa7EBtYxFxIa4EItrd5jSZrSctQRTqRAIcKE5FUk2HJvkuSg6065SbAigI9+
Ip1EHEuNmI9Fnym7SIQWibTxJrnq4ZymjUDAmqMZdNYH/8PLmgPasQR6jbWNtbwE0zY1b634XLKJ
+9uGXt41gPbu+qEFP0zsK5cdkkCovO4ArQf6OQ+hM+3r7h7NP9GL7kQaZPC8IiiGkYMtiezeTzVk
DSuNzsM6/1jKNfN0kmrgu1w+ziD6HjB7kseRMZuiZnz56RBw0uBeSXyckKHXR1sGz7XOEbzLzChs
NpsWRqNutW3fL7eWHlDsdmyIi0sU6p34gDiZ3qHPQogKSXcxQyjFy649Ru+g1tWMIRb5KPmVi5yf
1oKRdEYj4q+Yx4CjegJgXnzqCdJ5rDLovDsG7w3yLOiTtpt9IdTPbd8PIzB45ttiR4KcJ+H90Iqi
MTUF1BDdmmhkjllUIDjK996Q3l2Rdj5eZq6R9X0I29Q8RJEqQVwUea1NbwonT42cLgsBvyFIIEkk
nPULoTTdUKOdSAOkBNG1o2byr3EPoYufXP1OLUIXJZWfcYYUpWgvBpo/wrIAJObHPbsCdCcDDHYc
rqKaiA4PYgwuPP7T5brIuioklKze0Rw4ZjacxUGoczfh8BXGCZYkNXMdbEJA9NzJZrzhu3414hcI
Do21/gBKF0LNBaQ6lFAuFNeozW4FU4WdXLn/pMpBhkIbcKL0nNiKQuRGvwcPd6n6BrqcS53yAO0Y
wBXm94v5NKiwU4nGeALTkzTSaaejcpMqVqLf/Cg3RiN7T8xosj0aVAufi1V7o8KZkCi3odm2CMMc
/zl8Ki0y/++Ug/PR+/TyVzkvzOU3htUO3Od/ocTsYhZtFjUn03zwWnScwKHBuM0MIg5jMh7B0aQw
bX8S0AqRn7P0IuvnUo+VM314TbPGeluwcSO0aONGeRil8KMLZ4xBLxK1AZwwQQ6XhuSkPOPmHQz9
7fAIhsz/nU7HoZhokD+MY8cRXH3hib9HJ3kls3toAv1KettVAooMCibiuTyaXxl/PxAYCEBEqK8f
zqpb2K3W3UR7YgZbDQtf0f+hB9PHcJAhzBehQcdHybynxiBshSl8QSdbXGLsXp9dU77Thy8dWdUs
2RFcBqRvM6LLUiFx8S6/3mmvzvZpOOmGKsTFXVeO+MAwJO2K4+0cbP3PcBi65ePR4M0mk4UvtvwB
dDMgiUEVFKnr25cUUnROWW87Ok6CEKcoaBt54bFnjlOanqQu27fCtV29zZDSIRz3DsmsjGt0k1fR
nX0EaqtnYg5b7hvN5HQVyKM3roczLZm1Des84v5/uHaNYoSqJ9SNfGbGrdL03DwlZUgYDM09oJB1
HkPnkOGVhEbw6IdAiOSldiZkkUhY+B8PXFGhBFokegwdDu82jrYoZ8o3MHOy7pvjSQR+2hOAbNHm
bwzKlymMwgk1YQ8j6eXpaN0BOe1xOo1BrnMljI+aKenzrusRA8W+ML/hv+GuTooGwhU51o7PNL3W
TDhnVHzNUpniFHkGyIHU+Z/FkUMmlzRaFggpmGH+KbzezCng8dfcH/h2rafSBflNxx+dXp3Qg9Yo
wJIIBojCMp8YCcB8lSWWwfRMQYbVFz/Bzurz/gFpl3sslYJzbNJH2YngJtclyeiq5rT+tfWWQj52
ApQxa/lIuoqeehVoA7EePoN0U7SJP8lCGixFQFkaP9CUIy1rF3i6JU+vuf6XBXUClhZSuiZLOLeA
NweiOepQZ/3zhOLzdoRQNJTBfxXvkn9w4Z6KaGKcdF3u5v4lIhEutavJ6TdiTz8fdD4d+gJH6PYk
GtmEI3fNpZJEmxluG+nfKCRSl4qhSWGMPqRVzAzKwzs/6seYvZW9g9LZsodWJuq8nSnEDNtnJt+r
0a5e1B3kbRG5IwOZh89N+PBXDbSrHGOwq2sjkNkrvdPBZmtM9KIHBJwOTCFEdv3U9qCNyl0C/dPA
uVQNtAJyb//Rwjmre0nYUcIxvK7sGBoSz2Pwo3ztIzzIKJSe1JF3nTxCIBFcFrCxzb30l1S2wXKQ
u0jHZnf2Ft5fQIgqk/tPIZfNM8CCOoQkOV/y+VsB3mvaAER4tK8yPf529bRPRORAoZZCU3IpIQZ4
rLri8IVgFjXEUHl/TnFQgtuMLkd7nYh4R4ZdDLqvwWL5Xu/vAHylZ8l+mWbl/E67pAzJsDv7QEcn
VcxP5McGttpQtgnghAhltdPiOpyPg5VXSDFWHNRV4xLlSEOs8XxUi4jtCSx+HF/kQW4oZf4PtMbO
b+shpdFzmMP8S/3XDTo3/fCOvhfLLW7japV1G7zUzFHTXLLKkMfjWf3gO8YeeSTZj5bE0qiVHU3b
ezmUfqP/EetuzVHie6KXam+X7DnmCoyH0eSqf/hrsqL0Xlaj6DckXva61YlipK/rKgcUG7sE3E4L
6LzYnI31JqKc8C7AvyUifYD8KIZdBYNpqoQ9OcBBn1vPkuZxmtIJzn0TtijgefULbMhF7qFQvVX4
uSdq6d8TDgfFgDN9epBRdcwMYKABy8+8VfLkSTHOB2d10oQAS8RICwC94kWGXmOAVXMdnKW4h3mf
h1wieG9ggM02oPhXiVZZ/c8QTVa0qxYb9DyM0fTYsmOFgLhm3/n1PuFYWpFxA0sQlV/GzNsWBz9f
WjYPLNvLD1SHrfsqEBzBwVls9LNXuQ+asnbcPW7YOeDxZlMbTO+Q3u5i5Nhxmokz6GAraZvmPXdg
YJ0KAHJlyYN7751KdIEhyu+nBaiaXa6xK3fF5bzNtbNH+Jk6G8NjIi4D6zVAZ4JoWS4BbLLwiKP+
pKlflQJzOOiRf5P1hLJdorHVq/7ABX3nzZcivi5Bcs6zadTE6IZCAFFuTTcQ1gF8qrpoUIFfzATd
JAOfmo8BVHwBvTuInejcCUDmZmmmDrvruVa/1bx8WZ0fpPQYsle2GCfXRIWLeBHXgxovbXAqLMGB
WTvqNpE3NZKq9wM1WVx4O8oQB85AMWGcuu6CmEUWY7iqKXzgz7UapM5G2KtkBZ22MUg1rvX9gNPq
/lAEfSLt95yTrTiGeA2LHsmfd8Ms7AzX7bIosjp99aolCkc+E3kaDeY9pHtgkzajsaKOX8HwimmY
QT5di26nBPPW9vA4sFxbdOEcT14H3yIkSFCwgzXmcSkMdMTt9PkHIdHgfyVWDpUdFSPSh6iAFuwN
gYiW+vh+kyiFlOrLWzAww7JDC4D7chZrkPejGtnOg5aphCFdXnnGzx4GSB7BxF7ug/nGFccurHVV
AH3RANv9jCxhxSxSgsUGTZdt5zFYauZtSoxrTJR966NOVkwuAEePVfkqypJnMMnMwKNp/44L6Wcv
ySCskwsNXSX5KX9mk5AeDQ3kHQBKvkFqCw2JstPWT2HDH3H4wflo1tigBn+DdDjvUNUmcqwXRSpQ
WxKJgMnZrdjJ+dOnaFbqku2s7bYAgPLDK10VGP8Mm5tVmExXoy5VYsRf/PI43l94DQhGMvUmzyPb
eY1WImqyL72vKSP2m03dM42piX7foubd3vMZCdcUKHC5fiZOH6LjZm3UTsrSMl9+mQEiixVXL5Sw
RKAf0BfMg4E19n9ihUCrZCHyK+DJesvLaGpkMG71UafXu3BBz6TJythqg3nFXitRAE2ZUuoBe4RJ
fO/18oM/uyd8gURrcRcmtxtrzIZjMgpwYGtKHLHbGWmNLrQlzbc/NwYmqLJ2P0ULprjheayCZyIp
cU7B+3mdSITlMrtv/3WPICfzefFiwhXyCRE9VDKv+mC9KfkgUc9IVnc1O8IYNUX17k2PJtW4Gi7M
4yqwz1gAdGUFo389fznXvm+/q2ZhGQSw067yO/ARcHJM6ncwuHjcpxiHUZxfrxtRi4ECSIGLYDNl
rJqiv/EWGfBY0tSDCKSnPqommjpirH4wu1cEqt6ezQb1pglO1emM1rJWckbEkvg933DzY6xtzmpK
l+Y6ZykAulSVrz5guK4Bzp+CygEAW/6pqSzj1u7KUpcGuhEU8Sw7TWOQZDVmLVf74FyHLHDpNrmx
N6PSHhEsy7kjSEc3PHCd0WiDHgr26OBanQwUROrQxlFYqGoCrtjq9pAi6yNpDBrEsM4E4VMw6CuY
y9ILzMuMBxIXRfzq3E0BOdEClBUkIcu6gsThIBTYXmEMnyVzK8YIqq2ONnpfbMTLDHDGDkgh/hjn
RJA/b4fbozZ8gC/DtFPtIowhLkaLu2HQsOVqpcC68uMW1YrIpIEWlMJSp+ovN22pT7LRT6hjz6mn
9U37K3BXpzQiyzdIQUNYI5Mx3XaRwWpe6/lEPWe/pcDgwishslbdwQIMhCG+uE3OOZA3tUrPsB9R
pszvCHPjbYGYVde3BB09vqw4foPuX9EuZPrCu0Awn261WjC75hoXUY7WizcqdvIrgECIXrlzBc2D
bCsaWsINIDxgEpLvUJ9GvbTwRh+JrzE/cmGzJo5k6xWhDc3Az48rv7vOvRN7Yg/8WquFBwlJNFPo
wMNqPCiJY5SDZ5nhIp07IJktpVZ2KimtAraO2zPL57iWsnx4Db7Q87F8OX4o8+RVDAdd6W4H2AKZ
LkkPBLL0ilG3hZcN4iyoQKifDljqOBW0B+89WAInovQq9X2tQPBRQSxc5Zq9820KwhSPJdLMMC8x
OG1e5bS4tKVtvmgBEqJHGA2NjPbH1AzZuNlB24fyyQ70JP8WFnlv3mNr1zmA4AIAVtYcF/g7ZQqF
JCzVKr513wtr5H1Yvnel9HGKW8A+OXCSAdp3Aw4rk/4skcHZp3PwjR2VCUXXdd99NVYeZVJceut3
4tl837kYY5IIk3iCV/RpyG4OFOyjwDUonYO65woZHTYxZUi0ZUz4cuBkRVHilG9akDlsaEgtACy2
7VGtt66JY6lfwejYFO/edVCAgaUtEmvLGtGu/akygf4/nqX+aIR9+1bw5bKBHu6eFaaYD7aGq+7J
AnzjQpyMNR/PaPEVfQXCOQVOminC+PxPHJuZ8IDI5p4xqMxG0TrnIT7G9aYHJMpz2QQ9A/XZ5f7e
4aiTsfoKmo2E6ghbZydrpgi/BPdziTutP4Aa9lIOmYRKM3Jl6eKeXr83fzEKMRdf4lc8Gpm4uj5J
KfpjFfJaxyW4csGrWHa0tm9wlYGYrVY/nA7xPpRqb0Gc7sa6x4uNZRhjhyDbAgM61Aivoh/mXpTa
caYfidqA+yrGtRGP1XDZIH7ZjSLZua3DnowCTyaHDplOzFysWRtMnQtPvjlRMvPNW5FFRc75Qv2H
FNzM6/EQ6TOXkt8SCe/Im1w+fKB5dGd8py4tbhXvyq0I9sQxYcoXMsrFIsv/oxySmUsuc1/GRKVm
9EMyEfiEKYbTvwHtJKuVeCu7gAujb5sFdjlVk8KQXXY/PK3kgwmakgp5KfpHTXyqpo4zXygBBvgy
iXQIcdr8hIpv0eO5+NUH83yBKOhateyqSYUCwJUquZdqaOybZlvzcTQvpIFZ4iiwuioUWTagevLZ
zn7kKFo6Ap8LWr+NjKH9xgAGiekw0iFuGr+r7UiCW6O73pKyVTCP/GIxaPJA1g4U/FP6J4fb7uWP
RZFq7/1tlnMSQ0dgCLkEMvQ9xP1FPkdf/BFQi83rLwDs2P4aykLM/zUU35bpUUIWIPc+ZriOgqLz
eq68rVAl66bhyZPUIkAwXTUr4ftUS6ITHYkn4sqDqq1/c/1epkk/SN9xuOXtOcyeUDSLwQov0Q7I
V7HyQcHE2vH1DM1QZvVXTubcb/B0vnN7ghDP1DDbn2lnspJ6seCnAukTpWLzsCluC97nNJfSYVoi
q5PmUUF+DA8IRWT8AInhIWV73LBFF26u0vaUlBZDj5ECAWczmAP63ZrWLQ9/16cZYhcFicqZGhza
CXQmOMeA6EaDsd/5qi8HwwOEkbzTWr9tqvcCkVjPiudcfcvywPWuSFnTVclNMbhHZenvbWyeH4zv
PiDSGKjYQfTsyUJYhfdKYYMuC4uo3NF9ZkV5Ap5AidlEycJppEl9Wo+Q6fm5UUcrPKTJFKj6ho6+
f3ut5DJ/P6rDfB7Tt321oNWXp8XnCfOX80YVhmBrpwl7MZV8oQYkAmYekHzMmG/P1sGrJAj/be8I
SdqrOEjquXBRG9SMd6PPfqtqrqW7ohVvzm55qpa6JPYjmY4/T+06mjTPtd2Z7T/79BwNXsGS/3CN
Qli8sciu0haGKYufLlbECzbQ6CPPxnMap5DR3WHfYbJIwW0xsj17NTXhlKEPKNBlFjYcPtXu0wwm
WwqySlKilNI6zjl6ygpfZ3wJ3yMX80drCF4rczTQIqNH15Jkrj6MrsXCNNgQTrZoXVxHZD5SwPxl
nCNRwvc+Fh+t3ZhTKuet52RSd47QngslopREwTjmXh3cPIqbmceTp6HumtjiU2qWs16LuspC9ERo
1cOHlnXyyVLdwZ/a72S3G7b1b/Gh52vkhqtaw1R2JaALIuXoGM/Tbk/tNZgt3k2mr3a9L1Tn3RGH
nwUggiqjy2L3KpmOBhtT3Cf2o3awqP7+gewC7sJ47q5sX/ih5SvhDWsFZeXDnlaTCuaZqzjjIQmN
PtR5uZQzhGHtmgKFICOP9quO8OPuTr+fjS/eJnqe7zdg0XnAzYcK1f+NRr8FIDUbi1DOxYYHiaOI
GLa3sjhd1ILSygaSSsQsFRr4ff1z4ECbfAMYsgCLd4hwCEDNA/03/s5kwn7cbQn+2JaTUb/avwVl
wIyCA/FsSZKyCNMoYWbRLC5wX0z3ZmEYNjh0+r8YmiLK4D1Um5yuViU/3gE2azBqzqHhTk+pkbw/
UXbduSYoIDSUXmHVLK54zGQS0eOoumzhGXRY+pO4PXy3hRz+o7N7ekjmssK1i6khTixbFyDqUElb
MqTD2sgvxbky12zV6Is1uHZqow//ukzo0En2azNE3J8zkheuEuMgdQsRZ5wGSd5vVWjD+C/0TiTq
KSTh8uUs562L/qX91dua9UnB9sHO1xOnYDOAJImqoXuAI+rJkQw/l5oOVvZGxB+3BvkfHlvKcQGS
T8ImzGmdA8u0/hbmO4GLy/PrxwQX91lpuZjmTGdDW0ykC5miUGrkGodNaEU/Vw89JiS1ccu6LiMS
4M9SlGE8L/y1d2TGai7MPyaeZO5CZTlDDT7uCku1enzQGWFCTPNOD0SG7zlI74lDFhIuzLPXqixP
hdTLkVtjtnsKQm+GaG52QwUZYhjyXxk1uhoOPFwZINoWIiSpHqRSnb7R+LDNsQPQnfjdyFFozML6
qP+IZVw9lUMa5z3iQBFtG8qvl7YxLkw+HC2XZYK+c7kbH4QgSeijWbFRGult54M5v5pi0BSryq7o
IsaeWR5ieKhsSuf3pZx9ruyk0KdWjFsEjVjfYHkEX98xDm8wr5RdjDW8+YFJFoN4QLFqyD/bnH1C
DneOGwiaU5mi/aR8jv8lF8IvBff5QWkHyjNfZtV7xpdcuc2ChHm/ArZeTSubsVYPknHWivA2UDOV
+KltQMscU6S6rc1RS+aWjqj3pVoVztrDNlRBLiCcutDfC7Y2C67VMyqhI+Zoys7R6b4nFQp8befE
vCOIsb82oSDPh/jfJUNDzIDyxJvbVCY/zoljfa4LJkfwRKKIvfxSlBuIAgsW0THumCJKsmp/2zyt
bqlqAKIpSTjj26NVO/AmzughTu6MUMhFxzGaGR0HBmBZyeCh0LC/wFNEk0op6xSelNeTNxtR4+8A
+dO9tJlPHndZC5greay2/a7bx/0pLR2mjVNQbhJak70vv8W9Hsm+3vjxsYtWefUki7U68/hMdB47
XLQDLmEPXSuZhOwRu36tZ9M629SmMAmJwLFpEcpg8ioDn5PBzOKAecOkGy8cgD0NzgGroh25VC+Y
39fQZ4kLV8qH2XM+z661yJDAaZaDemz47HL1RRESilgUeaguAHb4pDsCKLyE2EKXaeJ4S7Pc50gW
/Sdb0SzNMPSS27OdeIMMNij/17iy5W8A0A8MW3WoMk7fTfRsbJpOtrpARLgIRKxmFZ5MCGNXFCLl
5OC6sT26oY4iIJC+Is0axyXr8FrHRobA/fkYMOBTS/3OXqXOOG2eSBQtjcAit+CjBuC9CkXnLJzS
+JQwQz9RW/vPqjdtKIsin3K56rOB4TdqmemnyEm4RKaA/vMf1AcKsO85G2wcZD5Gat/H1XloASj+
TXbMuaHnat7IozQTI9tw0O8w/eg4yBUFfPjXW7J4kVSysPHWzBqjSIpuq4ugybclKkQSEtZIurBn
kOzi7bdGTjzyQrMQFl2iYWJbim4BOqqTt9NAptd8YBO74PPudWZstZz1dodTmfMlsDrIhXQ8Ia/e
EPii/vCh9OcZLAjKuHOb+HeNALZqr3/qwyhTvDbqc3dDjf6NkkLPWq3pGcGxojpSfCWEPFEyW6Mb
QvA2lN9+xfLGLuRhYogbvQp7Tzp7xuf/f3od59WgX4To4emO2ZnsEN+0U6WHAEEOU78h3SktAYUY
aFbg5GazpeJAkitKzE1zO9n2ml44P24Q6dyvDLdbvtj7P54B3L7VhcH3+sWFffnWRnSCWCVbmQz7
32Wk2MUCcrXwWrsox2PWJLT37GYtokBBSdYd6n0qexg5c7x45FREPQ/lz2eOA351cgSlIdfH7TOZ
cK7YYuIsaY8ktEtbMnTxWeKEULpZoW0aIMaeAtYYS6AU6A1abxOvcDpnnsy9h3qbVdQTl6iMfvmJ
+b5NeHEqCONHmGKa1CiIcbPOMzUQQ2/K1MzzPUadLT59jXk8ySmGiu0gVXXGFV04CqBOneQQeb3c
S97HETCeLw1uiSABm3vN8XG0G1YYE+0OZr+9kFD4OziLf0H2euOy/9SG3MGkjwk4YQ9lgxli+vAO
RtN5qOHm3uVizBz/nmO2xRqFWnWeoGRtuxmT5mQDIhzKxp1f6ng8eRXXFGGYHSJmb6ZQuxkh5Ps1
0iTNQoG5IWwZMxhTIXCAcUHxEO6mulRN7XCCcPKD220jayk1VRrTFb29VeXRwmM4EM73tybSnZI5
BhxmF9hF9e2ZBnSZ0NS0Uz+i7TYAHj3t/RluivpbrxCY6QNH9vsQfWFKgsbuaehhmbC8/JPKR92Z
HMlSY5tX/VMb+/yOPg57SVX7pC6qElRPEDSEikoCBpLSNX2S5nA0fUlu4xNTkO+K1lJQRdedDvKj
Uoth4xFzQhoz0gueiMw/aDnx81MsFo8fRBB2PGm8ZiVUtlgFu9ZtmUBiaXFjkw0XQL42Xb9wkNWa
MW4+5GNah8y2bT4ErHu1yd4Ww3i8SKkv9SyhJydXoIGDw/Ssy7A37KJ3FyzjxZRuLhZEKo9tFctf
6TXATFFjRus641zID45DsrfPfPOo2lMKD+j+h2UiTsphQ1Fjud3iM7ZE/VIikXIQ1qy94JcV2LdB
htgR9bAlwRh+1P7H5JAZJP5cWUyvXSnD9Z5Kl6T/xKuNm4OYeLocQU2YZ4Q97nA3+DzCHaTEyBVh
QlL2t07lwRTvTOeu50uzAv2QGhyoKAVAWjbFuSZ3lgghUKRd7n5b3cymMZq9MAL3+3UAx+FC5tEi
6xBHjEIKINcSe7wJCzNPTqiSTevhaPnRjT4ymkYEIIz5zA4HSBo5Ppdpkl5EH7ZzAxs7Tgs9eozv
wlOu+t/opbrLp5p5l6rNi6GOXdG+Vc/scNm1DGr6bSyqoMYV3ZbgzjNVjG1lbBViPOVd5XWmdnOO
KA/dR24TCSRIn+Bs/4tKZzqBnvj7KyZcW/OBdpy7QGhl9FxWxJzKmGyHnlMuW1FFiEV39VAQAJbH
amljFN29rIbnKwbABRuoWbIwzVNzNOfa89YqWEVRjv7HNvAgLmxxkcbB+zXlOw5DH5pnXAtR3nAR
QNcsMrjTAnJMyB402xJTDsAQ4vv+csHp8H/LUbGTx1gqLQsvN6pl4v1TX5yQ0Zi8URmudBdVorj9
Lxhff9HvOtks9PP4w0iRMFLsU0TA83WLUsiea1gTlcmy+Y7hlGWohCy0GVyYeSpUSGvlviWmFBEr
Hwr7KWS1AGXD1fwPv3ErqvYi5tGxganXaQj7iUdqeKgD9M4N0LGUrXFB9EH4WDEj3JQ70pM7D+a9
gd00KJeTQ/nLOpW7LmeM8bDgHgUWBXNis1doRBzA5vOXV+0fUZmilFbUH5kcyBJJ2xcfI/ISBPr6
Wn5EzxjqNSohMixj182WU9QcCGGGdHIT4/uuafM/j0xRYoM2LE7SGfHsC/OUAbySdCzRqGmsL1FN
dG/a7ZTE3X/znIYrDaMLV2CIJpREmCI3/KsNrT5wG5A4Fr5IMfBq4o9M2zI4tXlT7/CHUx3zotni
m0zgCiSG43BoSOFbproy3sxLaR39I0tkn1BU+nKcSdxPuyxKuj7Pt3sO5TkXMYu87KpEQyHi88Pv
9yjzmMinzud2595m+kwkpx2Z8YASZRDCQvsEkVijHD9uDgkuAO2yTEOJWSzvATxJqKL/1P9rcrrU
HZcbulmtzI9XkB6lf6Y7DnY3XNWZOkN98b05g8TQOegqF+jWMSfUvDU4eYPMO0TO4w2Sf9oOoAXx
91OhNb3CQXzH5KAdJu5+oyjcCr1Fi/F2VQ2tD23MSYdWiYCL/rBgs7oO6gphWpavNHyVkog/NH9K
++lTa75yN0ARzM2ez/RtCp1eCwfw1RF9P3ALtLkUiSFHj3BzfoVLGOJW94kNlmSFA5cY7idSMN3O
dOR9ohpLYigiOEQrmz9+/CBS2JHJaKPmCBaJPeWaS2WonOsebjMneP3UyFYD6198QwPhzzSL2DBD
If88Zp6OUacXVIKqQhlqdLuN+yB40acsDGtTeTxg8btcJnHzy549DHbUc424r5BXIVPOvEhTvqRk
QUfVB5SQ+htaSwRCZiDBf9B9ZpZV/rWKNEvy+dWikIUjIYX8PDwa1i0Oh55wyu2zF9h7+8z4TyNt
9CAdV6JL1+a4Tdrf7NBH/i6UeCKHeKHcafLYDm8xa6ETRT1WkffF4b2AiY6vyU2CVvmyAcC2fXdp
r3jabZNTxh8QqU1g9YIYfMD9EVjkP5ynfmV2JIgF7lmwLf2D2bfXkWeD7BmHt+iDr2tnfoN+d2oc
iLFnBaNAIcpryCnqxD3D56vKqq7Apgo+ri2vQVCy25itg0CFIysocTmyo36FuTBMmAzz6vY34WJh
BOxR/DkJuEAWVmVa8FZd1RkPyo30iBDX/yAc+J/cy1s6fp9T8yKWOXEAHlTaMEt2qsgchCHVBKqf
W3Z0lkzfrcVhXfZDLL/UzDPpHcdQeGc2yeraViwLmm3NThaUI6W7ksZ+R3cGItLmpNUIbXSFItI+
2Ou4JG6dlN2/2Qyn5LnGHkEushWwKnSn+nb6pNh7p9BkCv/bUPyN8btyotkeO94aCsXC3E1wY9ZI
+BeHk9atZRzDydanT9/oW1do0jEyL8/er5AjrOm434ayqyo0L0R/Hd/+8HAkzCp7mxT0zVdUm9jT
CYsCc0tHQi61g/op1bC1iCIddQRd0SGF3cYHxO/EF94EzN6wbOzMpgDj7tzPrzpJ/gBXoEpaaMZD
BLxYUmLb5M5NbgUp2Pplthh4ocnzOtrom7cu1/hy9D7aUq65hpyW/8Kh3g1t13qHzTdTyZ8/0rPd
RGhlDT/m3BiTuFnollfI0xA09hSuM7ZbKSwX/lEBEJOjnm95F3jm53cnKdTHkMH0LTRnMJBMD4QA
rANWO/0Wf1sqgqc+57vgrNNjmGD8CryuuOXrSJONOMHf6iCApBlQg1us3cPI7zI58EgSAnXKyR1/
KvRbfNvQFDOfRxuSHmBM7KKhEzgdyNrEHU9s1H3dKOZvok1Zl7e0pFDMP6Y7VoWguNPKIXkouaej
wTHLYmRnUiqipvYxMciQYNWyHrqyA+qPY1d90kSu++QuF0bId28Ne31NCuQ0jHGLfUFY1SPxwneV
Y4hAbfG5qfxyK9SJlp5B4xudyQS5jP7tzj9wT/us6oh4PF9m7YW1My2OUSb3RNmxibZhZLE3OYsf
7NlAMwG8mCKTPkgA97QfwO+rw00vPtuJ0xcMTk9Ya+tLT/cFGqgHW5tmoBeURUIpQVi/iRluzTqP
6vNW87tSnonWmQRQRMnmpHvYvOX4R7fedhtlTy3B/CkwTr+3N5vr68GEbpoInYuh/5G6QeLbohXP
Sel4FaWl+90ZpzbswiPVH8IZumtyv4J4yA+mI/iUOh8eW2/w8qgCh2t/32c3ul+AjE0YselGKZKl
dwO7k554uCYzgyMTmhshb/DZH5Xa181AhbGJiqBP/dZoW4ELH/EfLNriuToMDfTKj/M1gSjZOZgt
7Y9LeYRUZ+atlk/ntB9HrFscj+Ymy0WSpE1u3jLFLEUerBfvTcQwytpJ/SqiPmoTmk6g+taKZTmQ
pZmJbIucgM2JxeyV1920MaJ/JhISysJuEbz7lngXvFda+++tRMLjJNnlSVrQupY43wXRZQSlVQms
5OJTJz5Ml/BfxoAnm74d8UqjwBHtAXHblbfcjZz0lcbjqHGRIm3Ah97bckSF7m3hXleXApX0bQrL
M6iiF+2K3IZ8jDbrAHZqtBweg520XJebjwu2jlhCAsO8iEiCnCDEbx5z0Y6mCHIQyuVdC5XJ99tn
Aa//tGJsArzHyyLpH2vzacvBwhrD/22oggIJhzMGSuS2ybwadVaYwLtFqOP4FmkG61G5eOwrEGfO
R0lRnmtSAx/J9mdAfOX1MW4/Dqw/sHThhOHQmIq6FBoPI4hu2o2Mjzu5287KCscrj9iVlDOAxBWv
ZCxnhS9j2o7dUzRHZVvM8k+doqHxyskKW9lZMsTRcphPtsI0zUrTVZlcyhf5dlCcpq2WEFWLoYce
QRSRpC2o7+rn/UOjsSrITEFTZz9htPaAMluIfdEouB8WjLG7WBTHKcngqm8mSwNZWxBUKXQ3BozW
F94rnZUmPXd+QtvBdihgRcHSrx5huAXJhUojzWlG0wUgvNz8bi8zCuWspxT6xqgPbvtfMXSLBbW1
jLVJZwhhjeDQck3mx5Jy6fRU/dcEqv4rxyxSSc0A3ap8O7X7Br/G6//gwCYRRSRXk65eLUw1kPUr
aDETtH9sHRgq3UY+cZ8878sIk+4zfwSrEeAflJwcJ88huWPHhl7POihfQBMiAUB9qzKXNvQJuMLd
BEnvGCJ9ch0RnvYxxDqLX9O08P725GnZmWa2o8G4LPoLi1QbtH6mlA6a8/SL3v3t+ovB/fnfibyz
K61FZVreST2XK7VZVb7bts3Ub5n14TDsc7xIuPiimdsI+WbrkVDrYHWMaSfNMHlOC3W5Lohi44i/
TX6jkyW6BwlVqZiqiH5IjF3jAhWA8l6l4vgC3HH0DLBFYYFOrfaNc/B0hCLnA7bo8pAWppLcGi59
9NhK3TIQRr98Dnvjwvt8C4OWbdXOc83XDH5Miuns9g1YhALkB49OPKqYfF+uhp34AQzL0QmBKVFB
fvd3Jega+CMh+mUfS8+esIytE8jFDtN6ZfEJOUCg1wFZakFjymW6aG9AWRiKfawNwo+3Qsf6uXi6
0HYLi6BpbUHEFfSOHZzq5SjXWBPZSLXrUehfRsWtP8O2WOYdA7GMpGzsuUIZ6mZ4TC/5OK43yB+0
FE+qGefHTsLb0QWrx+S9HnBXMrbzVpozA89s5sn/qmgY1g8Ezfvvutdrsu/QTLbtrq7Adn7mFCcv
PlWsXS243x4Rg51CJ/rfs/kiIECjxUOBYcSH4jaQ+hiP5wOk4z1Jxk4DW/Er7P4g3AX2Iz0MsrGe
nkyxgBtynGgvalojXZWD5l88tqcal2EL9feG0YnarmFPFE6cIxaBhyHzfs5LJdw9f0NomZRyXC7A
nC/5ze+oObbkJcmnd/NB8K4oyg2pZ3MA4xEUS+WCtUnPYVx5BhXubXg5xvsL3R6C/7z1cqyohH7y
y9HriiGmDJVI/9cO9vXu8GKlDOiBT4T+7RqwRa6DaNRmU/OQcw+Pk9GPCr05mv9J97hufmYGIPju
t4HJoDnb08HZLpekhFMoWNLZMRU6u1vWqgI0by+W0YvNJ7vIh69lRi8nt25OHx6s675G50yFmzUz
ZysbtI6M7nMz8LK65stNl5fONw4lWH7/t70lUOZ77mH2HvAU0uyIGjKpJb7a6E5SBOcJ9bccDx98
YfEnhQG6eQCqTwwQ+ob800M3Msbh1VCgeSRteBus1RkdHIsJ+wXN/9b5hXLz3/5j90CN5mULKtrT
becXTLcuuD5RGP8TJvT+qpef5q9bBFHHc6eRksbwM7BdjsTwy9e7eMWl5rvDRmY/0jq96Li134df
ecUaN6dLBj586XpgWAjNKFhbzipgQmGviN6HLVVWLlBWBBcbCChg5WoGnscPd3cYJACB2WYgO3fL
NnkWHJkIsy7OqF5L6X3vnk9tQBUpuDvmi6sJT9EPQDli5ERxNZ7D5o0g9eorMQ+7/udR1CCuj3dm
+aKdIXj/NE142gYCi0Z3gZw9NijeKtt1ZB4lDVXiJbIVavRoOutM/6DuOo5yAfRYnIeRIW/Hyfr6
k1Y5hxDqu95c4LGKSQ7jGWzdSp4hRhAbHF62dxQ10gr7mYZGfQ1al5w5Mx/7loMmsIEsdDL+ew5J
ET83N8uZVKQJn8RO49HMycvpHmspmrLIjl46CMsN90yoaSbGcrXOdqQ73Z+EOGuTTn1DjlPy7ALE
54iZ2yxLNovx9F9OLFADkNlVn01nteFsD1S7/PmxHAjZ1hEtSnXkLi00E+D3FI+elaixjgO7axKz
98DrMgzvsb6jRJn6rhg90L4b3oNor0iRjfZFaFmeR2zmL8i0L/gsc/vWl96rj9OnAieTXyaQ70aT
tnVYr/h9YSEIv0h8aixTwMUNPXxniTwL4GSXVuoogDpMv9nT1te7OMkovmL2rRPN9EHBGaaZbvqr
yopM9KSvMLqjjZPA4Vzh/On5h0XnPAbS5fYwc2bK2nRKZE4A7NjveVR2hZS6zVMMLGRnIGdHq7fb
yNQ4wNviyhupvZA/EGO6nscWTDIVP2D94MaXj3HkRxcYOpFX50+Bjar22VdgaSyz2XCpJ7+QT6V0
M9n9p69ui5laxGLtrB/QJ1W00xyUGcF9lwTyUz1d4NVYl4Pnfca85ID5hAAtvahOpxTv0WSK+LNX
fCfPPEaE9l0QHALWA5KhVhDqduRMb3HmE+lj31SWGtmmnYWaW9Dng2VBQRTCzg/TxG1o35U55e0o
JzOPYBAiUY4ilWCRHGhnQa3tA92wnRPgzlN0lSVcz7pBeVs27CzXWzuSGUUeh8YErbEU4nWZzs0Y
gUee/b/v2q8jhVXr6E+D1/iYpr6rvD9n1jpzuVLVn2qxocfQrOhnVLcSCR9QiZvGyCTIQ7SZnyGT
XU47cAeJwNnIyUxq4UWctMC3p/tgT2RsaJmIaFFp0TbZCiAwMghQBwlUZVR/hKf5ebsGRLCRPKB5
qnwkxOI8HGuOW1Wg6rlFf4FIfaKD0Lj6mHs+MfwGxfQys/ytgDgrF4d3uFoSUxjadJsDnAqGESG/
Fgn3r8+eP10S+Jj/V8sRtRYVeTHDkJknQ7KULvyyDYvEQwySb2FfRZ2VcNf5jCGKDbwUBK17gk5p
aFwQZGIgEUK2auqN1GmfzN06h5wyhQuWnrNhm28W7IGRDhRQbDe4w0jOEhWx3pOXbYg12jfW6wkH
uC4N6xvQbYchd7wmVg4CvRGDbIARrDamHd+5ebwQ7PkHlCqG4ncY5TFQqGDCyXuAL4KDdWkun0OG
YWgEYrikyA/li654VzrfdSjvFQEOubrm4tzBua1PgsGdlwbqyqVxp3hE7V7fn2jxvnuxpvmVHkQQ
+xVyDTt/MWCYbof57SJQq7lfWV8g9rKGxx8w56S0i5/r/Oy7lKWqF4Dp8/Msmr2rIzZS5hJn40E5
fWDGsUQzOlGj3zmys0G43d4rP26qOmp6tlc7kZ2XvFewEcY39bvF+BUCb7P5Z05+AZ+gdOm1FDqv
FzLWzLqlv0ppMSPtXEdoCzJdF+erK1t9KEYWQRhN0ICeKO5vgMFmms74KmkDyO9ob4Zupu/wgypQ
KVZMY/2AVA0bdOE0Tg1+OekwougbSh5gUGtMLnXm5Cnzx/yOZJSwDMq5jVZVYz7XaSo9sDuLm5FW
huRJFoJXP7NB0zSjpC51Xz0AwjJ0vLWKHIG1H7wceQViJXaJgHUHx6URQ8TggKFd5vP6kuGYTVus
TyOkR+w32Naaq8ddBS1W52mL8mHy3AYv4CgLxxF25zKGNZUvRPESWPEwc2xnfGw3X+7YfvWyAhvW
yhuUemnAOQqymeuqpovn4ozxNVMxgsJACH7oA0ErtLqCNIrZ1jfzrVD19j573GASDA7/54A9Zq+o
0cUfgaZxXEBOJqvyCxy9JhR0y4MJhQV0KhZhZaEWHiYauynJ/3lTKK4WP6ZNxtKlOuGm3cJ66Y/P
OEYxwl3DhpU4W3VwbKzeVWUenqc2ThQgsqqnYrB9SqRJCqmsunqE8MlY1K1NAfX9lj8UcfyrDz86
PXNC61pqbfRpVDqHpGZ7ge2riDi5uxl/adwSBBoArB30jvs4wygGrbzqiI5Zvwsut86qO7g7K6jv
U3zYF1RFDiOqRL3G4M9V/0K2nDVneWNwR0NY82BKgl7v92ncVhQh645UVqAXE9yL8rY3PSrVcZF0
NjQWUw65+fllW5zf0/ZfjXgdMnNGHrZchZXX1cuunJb+UXQr11inuyQhCFlGHcHV5WCuhFgN73iV
WZAh5Xfpt90PyBGDVuE0SjGJEaDgJSa3OtnnyHgdrkokZsPlLAuZXM9u3f1naTcqDKpz/Ctec2G7
Kagi7agx7JYqPMnuRIv7z52E2xFo0zD2wMnhEdc6HzhenFVw95kTTiiih0Jhwr4miD4TVXRlZzBa
MZJtrvUBhveXFwTUgXZ9DafWEINVUqgZIcTWRhWT3Yw8c4NyG1YRFOdBB2RyDxT7Ek3DOZ9J7qtn
x6AzvsflT3EIMi/LqM+x7zB3fSyKf7TTI+eLG8v7ZAA/LVM0MWE5K052Brn+sKuWQmIjM/bt9GRS
tKdiU1REtnDI6t82vRbcYJSy/drPO2Vl0b2SUgk6GCI+NrgBfzbjYniMw51cG0Azki9q9+aWWhyg
ZVfZ3TEaoxNZNGzOvMdF5DTmfyDOcYzB4TYtN6SDT2qp07GkjDEArqvB0uCLJ/TzWKg4KaoFqHNk
TlAYUh9YoXF6zSu4jCE1qvGajUZ47hIni+GcQ8nvVrUjkWV6l92H2Bnv3iDU+6HEZkkI/hg2jLyk
zlxFDsoupnCAApU45KbsyQPszMnj70SxQCBXdlP6ejiYQnq3WtLCz5K0LHdCgQHtgdU5XpGQJOJd
Wa6VppH0QlG8pY9qm6SSHdyzwk3WqlO1SCbqAxYWWnQKBwjvlkIYGDxb2/jEV3MfCysH+OfgZPjC
oZB1mHngGGD1uYFhCGGVEQIhp7ZW9YHjaTbiQKknlM/BJWfNu10T8gK49+Pn2e6wDf6WEWXdBDRt
ufkhINwX1SlcD5pJwvpcuBWT8DglfRQ9L9ufI0ILFcLoigvXdwvu9vG/4hf7ed2nmfoJZJ3TGfVV
kVcWjPzoKxdGyglyPVD9gF8+ydBZg1w3ZBTMyo8utqya2evyfSQHpKuxQT/OjpY1nyg4oJHrKlJw
7eRPbVN86O60qYnOpAocMDR3f22H5uUzObYuhFJMHVnoaU6FBNQgmbCFH3oHpgSADXkmMiMcljpZ
4MIWh42N4qzj0uivqMKq332AJTW63PECRgipi5jCyuBPBK224Mbb6lttziFl5FWknXvxK0m7WEpF
zivnvQJyoevu4Sf2uLMDboKFyVwk66KdbZ9BNwNzoEZCquGpI4y3L2QHsmaMFYHHipYyi24/1eLI
iV7aZRlQFuOJvZhUWiHv+jF/sqEekdxVb1PzljpyBa7+YzREXOyrbvnAUzo8HJuroGzbBQsrj9Cp
uq0UIGh4cp3/9va6w66dGRZJLyFrxJGdKfX0d/zu0POyJMcpvAI6lIMPArfajl0e2W4WvtfqTR+0
5Qj4ano0I1MfKMGvPinDdzbWOsqDBEU/uDzuhphpcRifCSXSctSnFekGUhpkL0Qgj8Mxgxvf2R6f
D5zcgqxMcEan4pU1pn1QDEPl8p7myvjtbc/8kX9mPl1coydcvlpwcesrciJNY4aNgraO4IAYLrid
h5o/T0KFZDu5VV2PgVteei/Byy5dUFMuWkEaswLWTc4/fdSVDPkPCb2f1bElGD382yw4kLY4OwVW
GWQRDXHIZ5j0TZyo07idpNYtpDk0vSO6Lp1suHMDQikNCW3CL4vy1c5O9wne4V1zadfr3kPc9HTL
TjH11TgetxGg/w3cFpuvlpbcHeUDXV9+S+filHpBj6ZyilaJYP6UBvnhES1hHM8wkYuFmE40QgRc
ohTYSXHZKom4cJFbNZiuuSrycdpOqS9wACzO3vqblBRrlX1suzX+1qTSfFH4mpVMJT/Qye9QALwI
+ZjRfdVm1JPKu6UqkqF5lqDw/p7XCn5QxsbX+/apgFzooDuXwPqi1dLZckvKxM7nHws+YPLa+l6o
jNIIXh2T2dwGupLCLZ2VMk503Rh6LFrHPECkmJVWhSmXtOy3R3WAgunE3hn9tyXPjUHCWEmvXSTW
0GsVwun4hIarauEZGrw1toOYLMcWJ80B+J2ba2IJlB48KS7cBQ5wKD3UV2lnCy24n6X1c50Ra/LV
H+w6S8v6WKXgs3JcFkCQRygTcZKfnpbhlu0HclqGiDsjbJ0KSh6e4bfsYzWlNAaD3PvssZatU1zd
Qf/nd67sMkDr8GTwhQHSy5V8CgFzFNox9voTE9jprlDUvkllOMlcuqIlcEsvEY7BEoxhLn8iLk34
LXT4wrgHugBFFU7oen9EnjfxV8ZfhJgGt+ss9rzmsJv36MGXaaKBSApcyUsurk60cSqpTgT7LX+u
w+tCucgBjzFHN9aDVPYzeHLE03ywgjcuIf64Ne3vnAsZglHDz/A5WbRQqU9ohgrje6fKHp3/y/OC
xEMzKtxCAiYth58gFFSaeoezFOU8YT7zYjrr/FZl4Spmn1epUeknZZBjh4Z30bGv8yfzRPmz0JK1
paFWhtNYzI9dDaSfLTve36c3OtX3JZE4rZlcbCms0+aRcy9PQ1SQQCrVW/FybykD5gPXo/68oK/Q
QofKf2Z81HYgAqvFnTepjOTVoNCzZrjJH30N0bVZETOOoaNDYFsSxtlUvQkvxxtdKoOW7finL8E5
aejw7WSoeTt3FezHLmFZD/C5DBkiXd4li08PJ72Q0EGsOQWt/OTrvBRcYOkhYFQfeAry+6Lzr5YV
KEFILJuGHrfbf6me0BCTxPTIlpPAmv7gdEnygaZb1PlA/KCRqLnheORq+4LbmeWbD7o9z4AuUgHY
BSJ+nG3ltdFGdVLS4gJTgicnnr4qeVKL73zci4ZAAop9LbFpTyQZvx6IsXM/DmxGYErwZiK2l5eV
73aA8y6FwInUBFIgE2DfXs4hKUd4TEdEq/WXuUUbhKS8gH0qIJekuJGUmCtGps8iKX7iayLqLEO6
C/Mg61sJQT9/Ztm8pEVOg/NmNABL0IwZS0EXjnl7TELvh6VcsUFf6eUl54v9E6Rrt0AuGtPWWX8X
ojQP9j+DuIvSPLCBwYcO+kdZLPGQElqX2QTtqHoryzmPYkz62+y8/66/4movRj4JJM6aFUdpMuiy
4M4SFdNGm+cjVI0lcruLM/QRwHD8fmvNXVSLTLQkYw+B22DyfoD6389WHniUTwpyTp5w50Eu8JEI
5gXFZu5EZKjuu6ta+eDdAeW8TYpNXKjbfD78EsLcDP0A/htVpSdkXdxDYGnP5Ipd3/430/TvQfTn
xReaAcevtVMmBuF15nYK5GDSxUtioqnodm9QcYV2vWsupaHILDoZUSFBpnaNrkd0i8nUs9XxG6bC
Efx/YqmQeLzot3Nl6uHhwZuX41kTJrKYH+UiP7l29TJbDQ59beZBW1aeEGTAzU8bbwyB6R5c0fRa
ILHo9hY15poQ5X5QHsZcTE+nDLw1JMe6ZqGx8CSnFyp8coYPFBlmTdrgi6B3iOjIZPW8VWpZp8DM
u6jZq+W5th8D7kc7E6qDiARqSk/ysfclfaoyM4k1dzzUevOi8AfafY108owVH6lWbqXKJYyrYwyQ
qrTUV1TY9IpKSj9uzEAtRall8BOuQLolVRj9jhXJqFYfjBuSS4KAJBk22IzaEfhkQGr9SmttluR4
TjydyQ2IQ75P9LY6/QnSpNuZiGchuDCFCX3yDOVuDzDbkbNZaE9F446sWycs4FgGqHdUU6Nuf54L
HVPwenkeMC2ptkZIMfOrH6Y9OT0U6OWOZ4wYNKYrEuYnvBAXk+ziZCI+4ECMze2OdqeXUmclLf5g
GbbzFE14iCX3Z+DTPHhp8mBLu3bruJSAEv8f0mF+5u1tFZj/CvncikFNMyixELwYJzr6W4PGrYlo
145q0vHewhJFtAO+l8kBGffI7cOfiLTRpgOlAM9axHDkaSPCkRHJyDl+fRlzvxSpdOCOAtUPXQeI
lKyD1qAF99GCdaHvv1ORF7tHmZiRaITJwJWYKVlMW/GDNTLjgWd65Lj/GwQJPIgIhlW9S5drSvSA
25+9E93fOgJaJc/KDzXNNKIcL1pz50XRVlwB2CT7AAS+5FQrE1N8z0SQ4R4IPynKpInt1vA3BR4Q
wD+/dlapukD3mI1TvbE0kapoboGcXZFCaIvhSW1q9Avp9uZIGfpWox5V0+S8fz46mNNxFF3CWXFQ
bI9guIQ64h0FOpAxqGVPyuEhgVXFzsuMen6Ke6/NhMVtSz+Yy+zsKpZOnQ4Z+AcebF95/C6/5CS0
ZA0f+7TodGSh4enWZPiQsaIOX8hsVG6tTaNj0Sn37UCorxz9f1nf192QhuZQYYHQNptuZn7isf4P
byiKCdxzE11F51hd+uqQklzeW4Z43n5RRz/5wsONHVwyfTcFukNT4FDJAzog716LB5g8bOt2nq6v
sLp/bEBY+OFNde2KSE2W1vDRobWrkJEtHgmPjENgAkmgjy9Z3ELP7TKWbFcWpGYd1Ft72RJqC0Oq
v+U/Xp5NU2J7QvmO0B7e+Ldskv/kPNrfwilyuTkCmgpQGTyLBvBJlU7smgn24QdXDYFC6uFBa3JS
THWiZPrATbTexNhKUv+qXSehOjByYCYKhEZefQklYhiN61dM3AxfFfp3/DnbXdRmUOjXKzgvf0Mr
VRch4eiKcx9O/X0vQaXXpX38GKDrgv+/x1YRl8K2wbQ/pX+qJyOgv+yY5G7SFEkkOx2n77FeugoL
cLtNHARoeb7VMoSiNna6rsrPDgeQ8ZQGVZCVGl3FXPfXIIJsiKKhIeCQPdNxWoa8DwaDCYYaXMEl
GxA3fMcgT/lm6xrE4OwUE5HpIyL/FJc6A5WxxQh9W7KBGiUPO8tpXe+PMXGaR4KZay1FtbhjJ8Ve
9PDKfpNb+CplCissWRbB+4ZNdYIfQdBOXXAF7WBlOZ8zD8spSu+CuQc2IDoqnm3DOfeoO41Xo3rx
1gRmjcXA1tsf7YWX/Ln+XSNIG8EEIdl+2YwOU4teOM7QXpOIls3Yco7xmuXtYFHP+UujiwU2sEi+
FjX985QiVUW0i2GpUp6Iysca3BCZLjygakHpFUtf+mlIuSCLRWoyFLLH6tKO+GBBVrz8vmIxye+m
b4GLp7kPzGsN7UsX7P5l7lGAEy931vdPENY/vwjnoiCdAaQzMTiBM6xrNRtybeTFOItB+Ij43v4M
OPW9KjHNgpAsMufCSyYKyIMw1OEHQVEpYHkPEO8Ftdi4Zi3c7yLmP0cCWY99GAPS6bMHbP+iv8ge
V4qccQxt+c3sT/1a5GXpjd1OFkqTW7Uk4qsMbadSFAwPiXXGvWQK0Zfi3SmGe1NevA6emu+z90Mz
4QKo/1cuCq3aSFpB5t7jX9H6s2Ya8Atl3SMfIT8jWzBw2hd0KRudtkmUqC2ETyDmJhdEXyi9VHTP
Il0TnTunvPdRlT9I/sqcjtxQmvCxRjeqT93u44M3JCa0IcAwVTIVJdHHNUusiEAZhQdMctXL+I1V
xDZRAa0XjxZfo9U4wS9hGW/S2bZLKTR/r/aK7r6kRT3qtTeQyJnuB6ifH+wdw8+oq+xT9W3MDOtw
1Fxn7j+wzDnoppqfhdRWXARJfkUcmlEeuNnJONxMW4WjTmALJG4IcArhhOJG73WEDO2vtxcynr6Q
dlf940llXxeVOoicZvniF6DG0z2vLQ3Hu3QGDhyDOOhqKnvVVu6q6iNAZhuH/3Aq/Wmcdam/rO/j
+YIh5xhq7KV9GyLBf2r1EtvUb2W1EX2LkojEVtKxXl6mXfI8ndu9eOH9AHSYtaLuigTQSMbj3mT7
0nAt4Uzc+SaR8BOQnc76Aq5P7plKLCEwTBZsMzMKE5LyyMax1mQSC6dQm9j2D4libj1V+57KtSI+
0bmLLyUT8U/H1MlUt2TghfZHaqV1N8+nNRYLCT/WLvjE7gO/4JThYz1AulrvyBCOV48h/ngBgu74
mCpHUr0LTQpu3xVMzCwQ4rhm3acKzU6pzsXc2yGCSx0B1xIG+HSvx2WhsTEHb40DQlvkH36CaTmU
14vba1IgTJ1atOjxNOmChZnmF76SrNVP0i06T4hp1PtlLfsaUVVBSuq2VHhHxlUft20hEcBGIRyd
PX5PDiTjcfla1f90EEldisjvZR5L+ebWmCz+1pLsfRJJO2YOQi4G9O6iTJCIGPKrhzQn3I9O+QHD
rBdm10vd5oTidAsP/71fB1Ow5EsEkTB25N5ss5meMUG1d0qHQ6pydX3X+c0aZdxJb0HTLVawalaz
jJ+nv7fgK/HR4xoofpm1bytTY0/nujxMitdSAAUTB+brl9mMdE35zo433MIFffCDQjhO77GvY7aQ
z4QISoS57RdRHilCHgjXfiyQKi/efJc6m+kxHscTYzZ3RtbqchG0yXcs9e53m3drTPJVNKK4GVbz
5RVngJSuatboiaCyneHQkFffc2268fOOiYlr4tU8mmjzNJnmm31T1+Dvur1BNXoZSaxocgg3Q8qd
1SQX2ujcVRpIv3ZJZILpK9W/ifSjOyAQ3GrsTrIuBU69xeIEKI7gMQj4N+BhQnOLKQ8275VbD/i1
MNs1Rn6C+5mJL1ePaeOJ9BaVD8pflKns1xom+mO/Y5Fy7eMe9nOokW/WBBTf9g2pVf4ne6QkxQXW
3HTuPvT7prcH8OA9w37VSx4vCFN4jmxNnxz4rIFyeO9HYkZHF+RtxeVHn+fhhf1eGCrl3pMkBcQ4
l6LCtC3Lqv4U+wr5cRTkBmZW+a7wu6S8B6dkyZMwoCf6thq1153XHNSeqB82RD+ng2gIRNWqDNhR
/snni0lE9f4iz7N+VOXB1I0rq8xIQsyvkuXxrtMKiwsmnRdVC8+X36W3Pf1GEzWBQRCwy+3q1UAl
oKASSTzl6naVQC6ganH+C1PFDcnATuV+Ek5JZbZsM5dmD4254letEZu0paP2V+UpNor8reFuCjKZ
iZGmOc8sJQSVd+3hCsXZ5SqVymq5D17luPyYEMkIeM5AoLvSq447ATOBjSjm/hIFBwitOdsuJbx2
a+DLvDHWKP2+ymCzbzxRKDneRHoXCnnCjPxBIG/U98zlWsR5C0565kqvfkffDMsj5Fx8KcB9kvs3
0oJmFsuNKvxDcdUZOdTu8bn+ffuMdEBLGAIL7tJUDkzsrMVo43hEUjm/MNV1FqUdgjeuS2DELmqA
6FWd3nlZTQM1Q5z/wbgJV23Dikr+oMZFeFagbl9WmAgUQ5Ht/0ofz/GB2YBrFI9mfAYmMfWRr8mz
rCx7kvR4wOaIvdkLosr+E3pVW0XCFtSLOAQKSp4XdnYSFDrMn7OeT2ul7497CHCn4fXO4/bL9nFb
nFJGZRaG155eeDPijFqmEPgRVCXyxTxxZ69T7p1QcBL9R20wRuFKyv6bmbI0/qgkU/hrf/PeU8Ge
cTWWMty2DW97lYlj+wwoeEasWDGoCi939HANS9/DrtoM77u/m34uRuGfIdvLWsVccTcYJjfg2sDE
WZxTbeui9W5loZqmzn8Uqnmh0UutCEAF4R+khCzSz2aQiKyTEBrDzyaQwszo5/nFdAfNUAgx/kmi
6nQUtUeI69ePW4dV6uyXKvXFdOaD+UKTRdOsq8scD5MM9grd0NLilKF2sDzQHHLn5W6hHVWHcjim
gRjKoqXBczHnLVI7SzvXsWErYtuj5o3cQi+6wJ8yepmRYpeiCRf3frSMCzcd8e/JZG5pfOzOa8ut
kLSLbNV+//aoBWBLJqhL/ufL+dwww9joZDVYJqK7bXiUh0IL1NB+CSVcDs1NsPl86zZBC8YUwBvW
16/p3e7JMnRWlxrrY0j0G4O/uWDWfwdIrfq53sU476ymZ+BJ6NWjnRRMF2a/x+1+REikkw5nNVq9
OfdOwV7fY86sK6AcROvoq3OojxGFLZ0cY8iq5D9enUvhxPaq2OrlnI1bUsLSeJ9m37pIRTbhE//L
vpZdLVQyYf810Y9oX2PZVzofNXAaW/FiC8sCbB6wO4SmdPoXOs/UNbml7bYUGlmTzsMurhzUefxp
9Bg+jikeAZBsan3bQU9yQSVJAAoTuMKjlaVQqgtwd9p1csQb3rV8k8L0jlJ6wgPjAejxCYssR1l/
iF0Szi5s8F6qpsrLoGGvjyVMkyllNRCxF7cPsjsOlSBW1PNRiMgkZunmU5ZDiXKJOj8KNG4BoqWx
+NhO0AD8wzVS3w2uY9DUpFwlzTv0m0XS1cdOpz0O5ocZRgpq9dvuMqrmOwQnRIETSbSvdR2kCbDX
yG0BKQJ0P2C5t3MSeoyQJFcCFVJCjgIOcrdVBggGBgh/0HMDmlKLRXCC+LwrrbRFW4P5uET28B3R
LHz1lTdhndqELQugW4eD/kdvRwQUrCI3aqfcnBzuqnAAHM8kP70fAtXOLOt8dfMLuSH6asuwjFnd
HjAOauUt2nkfdbJeT+V0Sf72gv0zpCw5WZ2bXQqzxN8G6fWsYefnbZSWsJe34CiYV43PAnPAB3oU
D+7QcoaCuuEcUUeUlCIMf+h/aEAadp+sdYvg3Oia64kD2xtE5XAwm6wfwa4lByys37chF98BSo5j
IHfN3b96I6KRCZboUvLaJyYNl57BVeaKp2sdCCEETOS3f4oPkPPOzv7QGfqVCzJUsjtsBsd63BgO
ociYOzJwz70sOIPV/7bwWWi5aHShuX9RyxZwt1Ysjug1qbSLgsV1TlA+gkdCNAJCfdmHnSnIlPtq
IirH2vv18XX0fL06CCS03+frqvejIWXtX+A+cqoiRgSEyesSTaYBk9Y689JRgltMTnZRB3CGRBA5
nEY+VdBQMe2HVUIeFpaK2KrbphpwZrFXY5sERgCoIq+2YxZe52e/T1SRwM140GOla8Wi1QRN6m4x
6qD/GtJn4ba/HtrkHfC+VsIWEUpx5kPUsC6eVi7k2DR8Xno8wDYvxDwjsBTOVBi77lYg2f+9qP2Q
Wib702Rsyn4Iot7dW1vHB0S/8pwH37qreCEUWJxvjwfRXJo/MutzaoKk7/rJniMBD2KRj4oQ1cg5
CnccHzog52aAAKNxyF+N+/LkBFhGpsHRAXwrVQoWi9l2Wom+wF7dJ3OOhbphWW+Dr1XQTi+ZhP1e
4nqqEC9Hqn29ZdJJCPrpD3AheKdO6ssCbe9lA4ZrKaBolZxdC/wYelL3+tijjyd8rK6sGzMw4MWb
MsRfx49CILYWv86S6Exn5B8aGkJiBuoHIJZVvcW5MGLCuC+OeQjCJ1suNSJ720VAZzJ5ouVSWTQp
wGWAayLlNWpKcVefmZKeFzcjO58H7kZfQfoessycA5UD+Pb8/1dWZMffzlmorPGQNonByWRgQqag
1V0LNUltwHGkMRM8ZtcjDKhXRe72hFrsGsN5L9H1dYhWfShhk0W5gvsft12J7IoFNNfdFdRa1Xai
FbIBBDbRy/auHc3lcUoe3m+xu3o+6squcpZgbPZxAF9cI7sNbwbEAySFDuIdEhlgq8yCMw6LIVVV
CKy5ZKxABq24W+rEW3UqupA2gG61Xw2zYC3Cv3/Whib+DfLDfqyjvzMVhv/mtFQPRmvDOAYvqLCV
oOb7Xco9Lav6USn1wpv+XsZtPza9cgEDy7yPvR+srjE+meJJ7i6FSAG7oHeXiEFkn1f1WeG5lqRI
INBwpql2YF7EysfT6XGnstMet1KWq9rqVk856efoyL/2ziOAfhsd++2thqE2mdXwxekb2wCMiogN
MfM/QdVu2h/kXdIyWiLi6yPhaUMpLzv6lsq5wvNLR7NRbA0sGdUhQA6d3HeKD/WnLCmGs00AaiFZ
15QFLpwAkbIl1vpfov+GbXcNU+ut+JSlfa1k+Oq61BZqLXAbaqkxyeEe1AiXhGblV7GAs1h1SIGd
DJX+regXajbR5+6stUR9WBnjy1UI4uOTV9qQDe9SoSX8kRUDRcVA0H4j95Rw2krS/YaYY0dl5IGH
0KKy6piC5/edg2riPOEaTppPsI2M+3DaU0LKphGfQ5VeUlGboBxOQDUL4Kalx3+RSzlmDljjX4Bb
aSFs+cY++48lzXr9aYwq+Zd1uu5FhycVY2shd8LeNfbXM15NQNQXjSKui6QTlGses110KHCh1WoU
RtUMny+4QpLiAeZ85IVv1fKep7meBhGPDMLtkGKZmU+n4G1wx1ewNDHM9QxMKFap3xg1YZFV8qYf
ytnV0rtdlQy9QJ3K5wdirahjUhoXa5xleGQis6FTa+nF3f6e6jbKHjAESKVsV+DE6DINAnVUsDiZ
DnoEt0WyK8RV6gAe5HTlsTKODx0W3P/7lR/KDydXEwR1wrEj/Yo5QWFJDiE3NZ76HdCG18PY5uxT
JZuakMBuk+p4vkGBVBzP4yBm2mbGgkS+KzknTuWhrzZUHxfYXiCcGoRUszDhiCboC4Oa2E0CfauD
zdXfnHwKK6GFDk20KpfFWKFvyQ7NhKOUNi/cr3wR9pPsj2Z0XoWdq9hK3lRmCCG4GtcIRE9t8f36
ilbIZK6Mk08mtfd/AhjezZA6gaxUedGQgqJUzHWS+OJ6j2TJr9INza2rXMtZCWVG8ExC5vl6cJkz
u2gEyD5mdhl1KwUSgR+UFDwxq0OpqCIUJXtemyaSRURdvO7LNB2iRAxMyjCbj3N8s0d8dEpxajon
hGJLdv2g+3J4kBmBefs57feJXSOpCSasrAYQ4Z5RdU7G3B29ixPTZZzc9NVok9tbfGuLnEWi1F5g
unFh8tNgMz0NNmrNgMu63DLVxF/hnPvgfWwYDoFtuehgHhEDxzbjCLhBoTZh1cVnT0lFP7/dZd/v
Lj+QnHARY6mb0zh1eV7Hf2+kndAQhiZkztMD6yhGONzKGaKwxfuWaZjCULyRo7FqNDCif8TVefxh
N5dvekAShwm/ojzz8LoQ2BpPps7B0nOuwJosul6dTGsjV38SI9fKYnz0vKwcZ+l9pEYtqJcr+/yC
VfMnKUiijSw6QY/h75GrNNOIHZbiJAb7ffir8t6mHMp0XfuqF7/A43znh73TUPQKx9C0kS+s5XK+
W/2e92XabD7cZyfMw762JESU8+/gM+j2ozoxpSsjBI/xhOW2teS5n+3LH8+PF26OZwJ4xtzFkMIy
GRVMfjlqyK6FTC/4RbVp5wkYFeIwHJ6QukTYEonOO9zSpxEqZMa2wUbR7Ag4iqgQd8sux38Li13B
5Utmjb9HSkDXNG5bKXitfEs/Y5krzPM94ubX+8tyE1cJN8IWjRlhSvvAE9QuZTfHrqDn6EuDnBT1
1GFiBDo/jTDJxL0De4TOTvNBej82EGIAYhs1dEcUDEb8HIDjVhtIuD5EwDtmNMXmSfn6/lZdQLb1
8nz7jipHPdA64Zbm65ejQ2xsA2b1o+/S5PkofyqIQ2nvoHzGZjq+6lN4tjIES2VDZxDJvMgHJoG2
ErQ77pmXq0E2kRdxP4XSjz+ECU37Ih4ENEnRkgW0BDkVgmhr0xLr5lQuqr/KgIrIldn1pVS//1E3
0PaONTyGXbENEPIGMK1Ox6kvzbSkiaNAs3xgfdxggnrXFDzCeu/R6w2dAReiUF8VwT32wokxhmOK
PYq5t9oqf53X0VLDukEhEHW4E5cdy4nuEyW7ckFCpNHK0g3hlUf5U47+tyN7AMjGgDoI2dW9UwDR
LtZTksYozF8FuwDFv4s18UVBVNfl/THZgtIZAI40WTKVi6JkxHEhuEpeZsCcjZ4ypprhlBkpTPzX
RbQ74oSKnnvOiTddcfkEgPumFmb7Z2LL36ghKwJWnEV1ypk5ntfRRwPikKCljgaSpQmglgR8PxOR
QX4Z5S2zsqk2i2BqdNBFfuJ6jccj7jmycMgDjrQu7wrSmbpFDlmxVA1/f+UmXAaswbDkGgDm+bRD
i7uOAyKy1m+mlakW0KV5hSPcQI1XrZzX1OiGH0Q6zC0f7w8IewskQ4+RbZ6/BjOZR/+zSFBQLJAt
6L1Po4E2Nl6S1PQA9rlaNjKxSwsct5mzoQRW4xxpYNE6rfdLbAJPBQzlie+UI2fH1OHQsXu9FC9K
OvywaC8Vxn31IAtUJT1B1Els8rjasDlJnSEyEHHeYV3HlczUMSdSNrKMEMRboEOaRy1DINld9OzD
Uj6nSnn/Hz38WJA2DX6aOL+wvSYIISBHX+toruiclBEc1XQtzILz1ZaKfJH4omB4Ff6/td16t9HT
ymnb7tEaDn+ITvHELsa1bx+4NsMBYAQQ7vFhAqc8GqYXMhL0dSHU6vH1NJoBX8mSfWNiBhbfxRn3
mlErV1YQ7k6e6wPSU7+KRF8nO4IHmbqoH12ZfGSORyAUzsP7f4sU2oPBPzPg9Zzsi/jhZJCNxBkU
kGEI1Nn7mOnz8rjUwAfucz7ID2HciSze4C5kC935tbse1vbvdVF4HcZlZ4Zc0tfyHOJgX5R8movO
tjiBqLqijn1wWghqbrucm7W0AMHvTCBII219Bfp2WokRR9/ZVi2S+bcNwlnL2wT5HBsjdOvWa0jG
I9w8Fj9cvrF3717S6MVYNGDF3DpAdnssWmYMWiFaTFIE3oyDZ4fBWdMt4AO54t3p9ybV3WDgSNaR
/L7SaWKavR81iZVRe62MO7/K3OAkrI8lEZ4j02RPbE083Wu5L55iao3SJAYyLxs7uDUbsur+uc9T
ZWDiYfSYKOWpPO+ImWhrmABSqFQYrqAlj+cccpHdMvzCZ21jJT8VK/tLO+u8PNnt5lAa6+ldVVKN
kmBcDVY/0aoJ2yAQ3aAR4qpHw8gldq9OfC88qxzfQH1sT8i234vs+aXypLvud7sZqBEGvow7B5Ai
3gKNLbg4yL3i+yu6/yGg0+AKPQhV+TzoafZBWbK3ZXj1Zm9BPOxcoEmLKcucOc+Dq8smma2OXQQp
PL1X51AHi2ahiyub2sDhLoXNfd3FjioOAErpEHPwaTavh4Yf1pdDb1LqMFG49blTmcKAxdNc6tuA
IL++m4nA3or2/7+l1baZ5RSWIDEAb7YyqJ8tedvlSauY6UOex5vL1AeHMmaeGFzNY+huMtl9BZQG
Z0PmtIAUXsZcJrgddfqAf/8KiZCFmKGGnv1hvCb0Xfe4/Ensa/dMEsNaqM+9QTmapIRfBWjJ/DLr
yfzdAO87nlz/9k1/t3iNwiFBIWijrf2nuPLH+j2UcRzFK3M9e0g1E5zkDNA1uCvnG4MwRu/RhHXc
345v1gzIhNpXtxcUZBNIgvqDokvU545BO386F4v42BTtU0bcuHyUBy5jVdHBLFTB9cwY814zU4Cz
XGuiBu0rFbZEmfh/xETEwQMKdslBotcd6Zi0BSeUsODlP7vAdZUrzdmI2Sn8tkVG4Wl7vTG/NjVX
tKDX/wEmmVrqrArHjFL9U68ApPg8p1QOx93VloRkGI/sZT3HpUQAEzAJxcCcSN7cFWxR9V3g2/DS
PvsokqnYdMpOylFhqqBLWYLH3Nakeh2DZ/b6GWFmmXVw8XpICJcZb2AQahDRimT75EbpE5x1Wvzx
1Avb+SCP0ZDFows8IxrPz3iI3r1KHtq7UVQ/Y5XjWro18NyZmxCI7mlLOCsXtihiZI0/D23PPdhx
EmdfmvSHyfXCBLCipCgdpRs66if8k7db8F6IhFt6D8crZA6itE6QA8BeIncojkQvp6Fyti58K4LH
wA7SZTkv4X2VGjk2BTWTU1pLnFJTOXmYWubxPLeXkmWiFLl/BRz1YxdJiwXMNYoRnZGm1XdolwPD
z+GeQWWBjO9uu5f7uCnxesg6zzgYFgQVeLsVDfKUGpdTccnAd8oqsOSYav794rSUFalfVUPdSoFR
8SzyrIAR+XzL8pm+cLPOGnHU5jJgso90Tp3u0dNEbcvxHJb3CBDVeXlt++ioG2G+LnqDllq54Fud
kzvFEUZzgA9GHtdru0szYYe+1zQWxZMbiYBrG48AWzW3sXH/A8Y8Hu5yIfRHh9J605WIKkXjvFDu
2tAScgHMkE+bJueyN/N2VcwCkQGaB4TRzUiKgD0aT1SPSvVVrVUy33Amta9Y6jKgTNU3dfhxp7b2
5y3ePL00cWLaKRAp0mZd3M6Nr1NM15aBgwm+LqI+8YP/s6oqt8jqP8TAI/IgbGH3OILJa4XqMiRS
BuMLr7bbaUIHczrk24D8gdpT/DE9tPtQ9e4ZX4zAjYUyQngqPZ2qY3/A58tWN467Uyi/MTbleotN
FwBSjGgmMV/VlIsZy2O41yvM/+oa9tnO31X5puYKREsc/xX9zuqoM7qtYN1W8bFrELdvwdhuo18q
mhkPOJZgUb85d4zAIzJOZXGK+unrEkfW/zdDHQYzo1kCiq5vXGOT4nCGBl1MD2uDdGFV7REkQOKP
eGPS1BygaBTaxLRvellM8+d27tjYk1Ii/emEP3eiiYLk3ENz+8vImURVFf+DiNcmUbcwNSb/svTm
BZ2pBY3HbMac6l4o+2KPV4gKDqMnk/Jrzs/qsz1yodb+izZ1OU8yZMq1gggi6jMBZm8IJnA5qDqL
hhUPZyjJbC9q1sheNNSQd6ZOmKG/2Xfso/jxBwa5KbnS4XBb9HPMXfRdbtwua7FC2WQYqZSrvxA6
2amszKmEoINVpUoxDe+LMgYQLEl6iOee1Jqd4miVReeLPLpUtskVB6aMUDqgdHsXkHlgpn7GbfMG
7rnR5TKXJLf07Lv9dSN/3yICdA7DaFu2aSaqDsAyHjWfKDDFesg3U2z+BCjTjFjscjnid/8Jfkxb
O+5fLSbw4kdrEuDgWwk4/UQPd+oTNomAoCjKmcCs64efUPLi1AX8nkrD+cciLXjCezbU+zAC8xZe
PBG6BaV5GRNlWei1NakKCvpPaR5SnZkNmCWttVkb7CvJGXhzwSs5mHAcIShWybnjpFwYsWVbtvlF
zDoKkLO1SzO75tl7/G8G3s6J6VQE9Zlp1Y0KOz5Qp34SDOJtfbVLKby2tAkNRxywVucwjARh4LfX
Sba8M8TlZ7oqN3/Qul2pOlt39zsTQCy2UJxKcPXyYVZRvHoVAxckMENAadxWL2zGJES78O43oiEp
BqQAK3E7ZQt+YR9rKfFBIicMywoexGolrS0TzcAj3wd+t28tYJfyIocB/C1W4O6+30JFSMdZMNwY
og2s5JDCiYZJ13b62SvP299rL7laW8q1VE+hLZRGjl17eMA2e+GRAEbKfkuoM8KU4XLF5/SNI0ht
649MCbEg8hfmiAfBzfZXWDPYZGhlQfbEmyaDZCuR4G8tzCnTxamidt1ji0DigfI4w+4kITJGaGD0
j4NiQ6WKeWNcLp9X8zPJelLL6IoX2Z9zf8WWUBa5C34SocAursJ8+ay3PMX4UsJrQt/FJvkLdRgH
dqBFOz/2oUI0R6BOtxt2JeKC/Xo0Id2fdBMC8OyOKnaW3BKntUGHQhRRsN+0XB6E6NRLbLc1XE7s
fjpsZQVCtgK23qEkcM5kg0NM4Q1FoTRKcoNt8timsRWhcn9crQjn9bJej9lQw8FE5zq+zcEwgIra
YuSQJssArHqrW6UyD5a3DYc8yRXjFEqDbUvwcSU337I+42zF9bVBc8o0FQ+VzivMVVb3kbzBgRxy
EJXH8uJwGenwNYBONkuQEAqi5Ipz2PaqHXqENrvcwrFgO0nN8J23waYG3dHjdcQt9sKvdK7IDlBl
ZOpFmEb0QN8nb+Cge/N6HVnEUFyvicXt93rwt0nCqm5Ekv97c/a593SXatCokUhKmInRb0nmDMzk
vLSWfpiYhIjWhfNSkhX6xM55Lhj/1ZE3rRg8rWgz/8+f5o/WeA/+6OvFrrYWAC6WOCqk3b9ptrGk
mPE7aQPZh8rMpDKr3KN7lvHqJ9v+OAWOc+ZdhwG36L8PEeZ3fE/e2ot3r7AOUXXgbyTI1XTntJ8b
KJP1hwOR7gWbvRqZZ4Eh1nc+m6F6b4lkK+LjYcWooR6vu/uGkHwVJGIHt17pX0uIxZ9wjQewe6d+
/IuyOgEcd3+tgg+a9YFkSlRElsQcvSCWowsIELG1cBWjkXh0i7Wb/AyO1T1RfHU/6b1sD+hRW3ih
qGy9IEeykwTttwqAG8HXFbpKFSn4Foz6jHV9nwtUmugWcMJ1LDwU/FpAdSii8CLH459W1MB0S2/K
ptsEUf026UuS312VYDXKuhRom86V0W4bpWzA1+uQZ2TqIyrDRwNK6MnhUCEjBdxtWux4TU3zZTci
UH1Ef+ME1zcg8T/eNMR/rKD/z8DIEu6wldIsX01ZMvlJH3PFBYNNad0m+165OHYZTEfrRqoNUxi0
GooAWTrVz96oUGGNQFU7IoPbJjU2YBW38XUmHH3iTvKia9tvWHRUXhBSiVo2AsPpUeXjzSDozSh8
jdXIskgIjsLoJs0Vly9giHHQFPrAvrJvOEw9FZ116O+dgO013MhdiKnY7VCwnRoBBXLl5OQOy1dl
9Qz28HA7E9gjM9Y0UebfMb9ouOl0MQkGlQSnMuQfm0jJ9KIuwe3msKNGZfRuCC9A8SgpR5SIodws
6XyNlNICTjhdScYPn6U6qL7fc9M0g4GyhrVh5w3TPVwrA6xmHBJVQebprt03xrdZIbnx8/Tm1qoD
gXGpzHaZsgHRPuBMRVpsUCbQSB/oBdWUapT3jYLntUZ3Lvhu/rk2E8DbGZwjyRnl60QaRY14THO3
Gc1kmdSMY5y5LUuIeIVuJ1IP0XzJ1YQQjAZ1uePnQMk/tS2bkSrnMAy9tvHPfbU1ZIPZCyREMLm7
Jjl4s/Y6oMT0dKZpGPjbrhCsb/nc8uCkn4wZqtuMwGs/THJbh9ya+w1t53nPkRdblRfGL4QLd6Gu
Yhj42n4S5JPLnuWJzm2PbmuCt87W+BwEDrjrPuFcMJXE0mAdOb5cXy/479UOTqclbeOdc6CUk3CP
mNyLxw8+1bBuDsEM6i/jHA2rZ0qJLg58dHrpSpRPUQBZuVRZVzgT4XmAZiL2GOaDsNaERDi5ZrXO
qtY5y7on/TCrc25N7Xmv+YH2rl9peFCa/FI9dF/E19p31AR6FgWvcFG7e3LsQ7aF/mpZEn2ZBw2z
QkbsslS5g6wyl0aSnxMcpU1Hjkf/6pdxPknA8NxoPGqppWiLvu/4bani75hjht/FabDoAVQinjJG
cMvHKj2axM8orKSfBIlOU/Nq5xmaWP+p+IYKgGc2oIixKH6zna1iIKkxnSSTwMrPVR7KL2NMq9eU
KVYghRcSZCObVgK0oV1RLlqok4k8f0ACfW+veyvgG6CcYZKxguuKeVGH10/tJjxBPf+IbeLeV73X
2QiuHHeBLop6EbnIT0LoNLyjMPpMjcKn3keB++8oI3ZQ3OApYTo1ZTPbMtQdr8EG3Vt8qO/Zu2d6
tDk7eR1Xk9emHYSRir0q3DyMHgdxzGq2u6/iDu7E00fx2eZigteo5QmYnpBXq56fByI+tAH6nZaa
Z/OtZU3iotFiCcX0lEbjjxG7FJRs1P64us+y4i1G1pcHHP9hXGC8ngXFhD+gOsCUEAs1EUvdAGt5
qyTcLn5kwwkNOodNzQuls5HhrtKvQxwC4NmF8TEx65KRiEOmnGlho9XVlIKhozMc5UZ/yWRGioEA
B/IOKtsicVAIkJftLbwHwtLDgd4NgxwX4DuOmnDAd6qsa9Q22QzF2HHdpC3qgpB/D+FXrpTSUMUV
SgnWMdmo5GDV4KMoYBn5XbGwzhm9BNl1O3bl5UQ5jy4mUBBbaLd5t+G7568gEh/q93xARB2THG+n
3Zmy7IV/A3WGVE0b56tCXDOEefpsAa2hiiynW1Ljl5lkrHlYURHXA4CMDpCom+rVLEE789I04A4R
zw5HMX593y74lZN3w0wIi65pjm84A41C1mD5nicoGY82TDpVf2oP1bpVRk1BzxuvQhjZ9fNTqnTr
sOlmLrxBz6TSGCrF1yk+odbkvn8PEAMqQ09XaNsP8HS3ycSIKuMEWNbTKeWVmMKt3ygxFTaUsdS9
Nxq2WChEGEPh+nDF3yodc3/Opb+wu7LPATQZBSjwvggBRTrZK1nWdh9fBzDVXgU3Ch97VHibd8RG
adrBgr5Je7z+2NX6YzcNu271de29X22n+MoDDC2B2z2cCIB5rInD2EsmkTMh5aIz1l+b6HZGlpko
mZkciHNnIsHl6SR1t8PKPwJ+NKyw3+T87xfg9jWF5S00b0lZVc3mK4Ynek0lMy+JkV8S5KjQmM/K
h8JVBWcSqW8OyhhtrYiGFaQ6+7iUL0hIOp4NefWSq1ZTys87CyNCMYcQh6FQbiNEPDBizA3ugEqd
FInU3kh2UzsN6QFWvDKheEVzpJw/w9NwNs2QRZnazeLIFP/8XDUrJqO70fX7N5yUFjxG2MwWtSKo
lGucFFFTb7pM7wTGpa2YKnhT+l3A+23gvIuTI7eL1PXLzmKdkB81b2C/ywC2aMk4zLcqwYE1DB5J
J6KSidiHNMrL5GonnlUvZRcevr2W4b6nOtMFZCFEpN7cDTSma27AZjlu1lmQSuWTJDC+3yIj3fhM
KQvW7ygx9Knht2aefY00WbSXBiqyDXN1lwr3+jwz+X+zP5hhEJcdcsz0sms7OC16WTApPBnwszmK
FkpFq2VbWNtGveOTSTVmoMLerjSOcnYn5bySjFx3QA5fkNo1lXwzUXG9etLMmAX1lrW1ChK4xpP9
pZUcFmvn/2/HANRpngJENF8UKPMzGIKXz/UcHEyd385vmZhZLh+05RwvfxorKZUCno41NboG7pyB
a92nIHrWQDROdqdn0aNHnGRYCoPFNkGpW5kStmzMHrzOrWOHFtejLZG0AR28myMP6Gmb2AsTTsbr
w2QQic3uhs1ShU+uFxDqDvxr18NUvqsdxRkzOQiBZ7p/5c9HxBiVWArLKsAV6Hj3jLpbUnsE9Tsi
SrZEIhASImVXyozu/A2JLA9zOFOo5Z/4mdINgfqYxX+h5L+Bc+9qizvsPlg9YwW6aw9X5GqonZGx
XpL3OBDHNhW9aisrSTe1E/rGaj1IhVp2N4LMypDMzO4nGBA6EhaRXR3kqzH77febQF3OlRDkTUD2
A4bWefEu1lLoXbJUCR1yBxKyAS6LxXyxX4RcwauC5Kox7GVazYPyMzUAzV8zgrP8QusYHROtik1y
RnRpYiuedd230KWxyYY5mpCTfOVZtqfDBdvUcdH00tnnylUPu3tfzJWAKLS0dIbClg0zcvsrnWi9
HqGVkI/ifmSlIumbsJeDsnYXlWnaQqR2jPlgPxrsQjLDDu4wqgl0ErNBK6uXt7Sx9F89De7yEsro
w5BhZqW13/E2RZpEt1+kVUhopEy83wZrkkeu6lo+/cvAmaC/ttew3yT5ltu6+sdKQjSigXH8HpVb
dt5Dgn0zqL1qmtJWw9sl80P5MNWXysG01IdVFbbybkepqbaiTv1P1RSWT+PKoYWNXoj/4LNr0N11
IJnFhi/7F82uEbnf1XSK8b8ZAuoRYgvHEnR7BGZpVOe/dlhuMEtFXv9YY/1roQ4ANByKpby1xPgR
uU5qtNSQHLLzV9ROHBVcEhPXZV7a2X7BY65LcvDCIwOHTAHCfEsZmsskiCtWY7K9yEZrFRoO43av
rQ7SdbC7CJXM30vyNB+g1h6mGxRoYZhiWAXql0S9eoFcAFua2UgiaoTJU5RQnbtZq0lxCFX6LWdc
Hy4swF57/TQoDyBXtoHJeYlVlkTksBEPWjWbi4bnqTqX8LjT4yW7EyB1PRmWhfQJ5SGiqnnb+mp0
jUIdyUm+4BgpsGHXkeal/FSlW7PsK0DdpiDzQrXzgzyU1Iou+nwFDOlq2i/55D8+5ttH+87HpCaY
raCPQ3R3Bsg0vYtNQG8ixgo89UQcFdzIE37FYbG/Iz40y0jJXpDwWG3uq2AsNKCFC8insUAxc1hg
g7JwnFdPEPy6GDuwOA1MRNofOpm8X9lGDhm0baNcqxczAsViKLRK8L2ZoklztjxoXrIdK3eZNPA8
mNqM4dpbmg/zkpcvmPEwoF4B4RpBZFbNdKVi/QtxakockjZ6lMtonU3zI4GGmJUFTPQJlvx6pxxr
e0apdtOxfBsakxv+6Mrd/b2T6IDHc9oZT4Sg+o6AgDJ5rBSD1F/dzjIKL7g4PojW+NgQdhEiAoCZ
iIqu2hgXq9lNcboSaoFBmApj4boyEHiCpWRya0F5WyYPFWRgdhweTN/DllBivVDT+lt/NUVhYT7r
JKXfZzwA9N6q/+2ARTZLp3dZsBJnf6zocEDv9dp2KXOFpi5XTLgaAX/+KsSR4yaxeS9IWZQ+Iaku
MRLkBFJjHZp/P9fRkkMhqXcWGchyzoKwvQwpeo0JqbMX8XMSR0sO/gYtz5BD153iCYoAwdfjYm+L
/saeDxLPzS0secbWp6DdBNxRCscM4vn+GgLmIRQ46QVu5VK4+OndF2jEZhjKnQTcg3hbPWd+TRAQ
hkkkmI7/VCWvR/IlmmKA+OXN9L/QBmB4h2lU9BUav64hbTgVeYJCL5X/RV10O8d9kPMbkjxANyBr
FUa8txx78hERUrgkjh9+fhV7ER1JM1wsq6fZ2fDX45a9ZuW4nyG8iT0YJaBtCULx+x2aAUo4A9tQ
tboqhY2NqBKVOZyI8gRGm78vgIce65O19HvRehq1zfhKqqjdCMUnj63S6o7ZwJp6dcg6Ba+gM5JE
mjekPQmQI1Hx6eyI1l3WtJLsvO8B5speBfnwwBGbcnwfmCXZhZhQktKocy0497gWEaCnR2K5FXQ4
tt+u0Swg83m+rHotmaiC8bD0NdjwQXv8dJM6q42mBTNP/oykhAAzI2vCcFfkTXK6YoixSch058YY
QPeprGiHHLhw1oiBRbV+XLPXZPriYsGYxB6RIV3MX/+sztDnzpM5jk6EFDGheM4sUaymuJFDF6Js
gkQguPF+Wjn29zAu/cQN39PEVGwl3B4Sd875CT6HrKKsqea0zlF7BDbLLFmp28sJjXBqsWMBmAa3
iQxjX6XH/VGjhap6P2y89S5oaIiLW12Nj4Bx4Gzkzv6Bie+rFLUoJSMXLY0rvKcAldGdzzcWlOWx
OtNVIGcIdETHDgpZyx4M8/aSrOT/BdNcpSScjk/RVM1fuby43pkVqIRjCdSxMd8AjLDoYDhtx1Ic
XBf8s8PxREOE0amtxpgOhlxpFAJqPJuQq9kGIIwlT5Yk2bIC0pNOGhSAeUyUf+bSva0p07VemLee
k4ReomE/L/f1ktnLhVrRqY7zGWTtn7z7EniyuFSuWa37N8q0EsoqlZmJvqwTf5g5JcJvRUK5Bfk/
RlFu/kmdPcfa5vNbS+MFwYIMKpFDGW0gOjJdNKhlY9oRGiDcDhGRHtgt32IERg5sPRix4db28WGv
moTkAQI4IXhdm4wZkp5Te3YKggY0iqnUQ9fKvJIDRSFQ+hD0zwAV6CamiTwCgzIuaY9kNAYsWmcz
1UmPgbhegTgt4zelvlb2QW3/5h9AlGvsHMM9qMwgHaoIomtnVQhqwd1VUcSTDGPP0PLbwiGF9Wjf
hRfzAX5BuFvRkL9ieIcPPtr45/zwvvLL56M80Jt3LDLtB024SWhSnAhJnAZRoZOY0iZOyThnah52
dUIUgjEoEQqMtvbIvbQPVZqxi2qjcbErK3p3O89LoF6zZKxb2GupYVAZFyTIat7+lYe4z3+Uddit
Zr1G3iT1yw7EDsQFhG8a7WrHMqTeVREbP2pbW0Sqs6QH7a4sUU+1VASp9zYZOCZyu3oTXj9zIoPq
S32/hxxY1LVyvIZbzIMeHE0DnA16tlXToQD37zv9/kzDICvN9mVS0SKBDhT+C8Pkq7XcVERDjJ+k
KnSBbiT09Dfen1iGkmoTbDksdD6ACcrmyod7JSEgNpBTzvRP0xJssE5DUFELWaAjQwztqanPjfcs
kuuyF0gGT2zoFC/2/KtHptSIBsV02jf3wsxdMprFYY149xrMmUR9Up+76SSMhcX/V172QgfsOlLX
fIQgBUjCCDzalCYMBxVEsHZ4mehTJVMFqpR1CkbPiGh8aixBfveWTdh0S7E4yWdGTQFryWkGupaC
PigYvO4eXFvVg1pKN/Exa/WUXEX4N9Vv2whnPVBORk54CDjJMEknbrpcLGNroY1OG7KR+/WNnts7
ucwUl1giwX83ei+RF1CFUrmRkBkmwdDOVAH5LlnxyT/RSmuNDoXicbRZFz3/KMyVSAkGYgkQVmWM
1b4Jyrxr4JG/b+I85WsTpgkTAfhnOSthlT8CZ8YrkdyD3UtsEHrYSn4YfZu4Z4NoXd9gYhlgSWk4
VCAu9CnpUhaHRfZluuW7E/C0z6eeltFQ1tdIOwePcOfAJR1873n5CoTEmahrOgjnUfWICwdySc9z
pyLJMCG2KyDq6/ZSHaCptTCSmo16RCcN1mW4p3JkaCFPl+nCNy3FTKpU/K2Jbs4zuG+Qezty5QAd
7FOQ0l+RqjUjoWYXBXw1w6cgPPqzUH/IM8Y9aO5mkkc76RM8vY0sI6Z3UhhguBDqfOAza/AQD2VT
Y+9I8eMlQxcpnB7wP5uxJfktRQiPXIAFzbWFCsuj34POTAxiZnDDNuI5+qLqUjfP19ylTb0++yd/
wGpLWVEZq9aLku3s8rG7lE7+hVdoQJJOYcun4rvHaLSJKw+ZHt+nYp1/YrbwM6AKx5QEZBLXnIkX
A5f6Wct5LA0N5dHbIHXaWcgOZxnDrIJ5RL6AjWCDWwcBPvFpDEXfkxA4ViI2kuAbtzZKlrnc6Wt1
gMmCVyeR4a4eUSjgseL2qtpiab+MoCKxeAq7o4q0N5HRFQuD/fKhztbt24bAwFuzsAvFRnolBMVq
VQ7ELvsKs1rbGs/J1zfZmM4Om7y6oG2GLPtKOAw7GsGmYvGQTqkMsESCO7UhY4lHR5XBV/22VYRb
utPvgbAFk89a9UOebl6Ts86V9InN+h6JMd1iVGcXGv5qQu4BNpNS5GCtGVNpuNaaPPfl1EMtbjf3
ZVZpmH78iIB61tBGkHBEZ3CLaO0mbsChRu2qHsoWvI4q+6MSxpvYnUDOCR69ka7+dTbSrbt5Uwit
c7zF+B85kTeStT1K6c2l18ISjnkBBYtYmBFrgUHnlBn2PJocRgHHWZttVauwr8WC3jxZQ/uOec3M
U8EO5t3wMjzkocpRlQhAKHIqyGubGShiqOu9/iSOAHYs7/6OB6raqwS61SeWmn1tKQeHuxXbem1J
HHhRMe01fH1t1c/zAjabBebK7/BWHUnG0hK9qdBSzyd0DdR3WL19f/snYLLFXhYDu/lqMnrTQRPC
wAIdQsQWBIsgun2kPSnDMsq2xT+ayTUvxh0Fyt6moSb162Q9ocwLG7BiMVx8y5lUS6nzC+PW9dle
RNqEOlYuappNi+rsDqCyJK7kpbiDILbe/c9qatvuLScnz0BqlHJZLPAQ8CFUXH+5OV9CCkJWs7fr
9RWKV0CcU/GM0+hU6KGksCFbU9h8hVcp93HXKq512hE/TwsLWKKZdeAtgXTTLmSPmk2VjMTNPlpF
Q8mkJagIc65TI3hHZVavslSB/HpZYwAo1lzrISK0OOk8NrA4uE0EwntsEl/mdHqpvByG/JLrd3tD
X8e5FI3GPels5C3cEQJBTg8zZ1+qB8c8TcRXLP08shySlvR4z/9YIB99GxeZV1+DAAVQzhfGd/wO
alha7jj53VW29OHf4jq1OgZj5OEDN2EgKBPjlt3HW/MpNy3h08j04XEeyNXQ1C5QKEDIqqHRAxvC
fqSOf9JSI7XV9fy455vVb55Wxiu1pvlu6d6h506xKJBezKcKX3dMbkoS5gtUBPbFSMhMpOcUaI57
xqU2RTmRdq6fDRjS02Xtk6K58BcWmn4cAp8aXcLJgIK1ReZo6x5r85YZNfO5PznfUExkLs3JbjEM
Nu/AQ73Tkbspid61xx/qdQRveHmuI/6FFakyHg6mZC91I2zmtZTM7AzLpeM/LeKnxUtiPoptzqoD
3BfUrzPo1/5+wZgq2jlJwZiHh1QnCrmty2t/MKJ5hNz2GkKWJgwj6JkzAzFOPRyAjFPprV/9Bs4h
cSMp18XQj9XN+jmE0qzQct6BhVxvQwutDuMNdlgSUxX35koRjws7GzvfOTLANpNd4rcgkPUK38G2
ZnkzAI0Zc42sXZXuJWjyBxAVzt+xW2HzqrtTvzFZzisZ3CoCDTfdGJpMMW2tOkoyL/X84imCEVEP
yh+bIvHHNvPWWTLbdz73XoLyqejDZ9ttuZzPGOdQhxgrTbS3GiqwZXsyoKrOQ9sgE7sC2Rj75eML
ontQkxckoy5CIBxiB2WblqieTDlaWynTXcL5YvuEDCrierFw9AFr63RgS5eLVWVUNP9rWJlZr++u
ZRhZ9GZ9WTCUxErMpusohwz/vPOa2tQg80+fRPVu+TMxfrzTmNOQVgU8Np2yjHpoqsSOLQ2FiW3X
4R1G8e1DMeVNnmxq+bvfAWwgM60NhB65v5F5X9cGAz2HsaMMKPxz0BeOgUmbhGCZaU6xIhAsxyi4
ZxF9etqLH+YONMunBdkjwSKdrVuSLuvFKGeGiQOuKUu32R7gw79mIlJYFkpV/Z6db+UJs1Z1y/oi
j/EITV+NOQSrV/D0RgL3YIZjHv8qHpDSVsp/Ur0dQF/xWOs2gqu4Z8KqJbQor5jHq7iCq40NE6V0
iE/7RPjLiKs5zqMJISowXcPDgYBIG/QuQ213drdtBijrDus2juAG3+dADKivpCHcm6S8mQiHiUKI
grnzhLCl9KUIXAY2i/FhRfhzMUdSnD8LGQeeNDHq5gqWc1StIHflnhJEl8SzXFPqPkl21CMZxajF
SXtcmU765aH6Og1Pj0BFdVEu+XZZoaN/HKo83UBmXthD9hJ8xT+Bc4fon15Xbb/uSWufFVoQoktl
GAAkawHgz6wOPje5xUx7O/pcLBLwX8+UJVhqVPDKXByhZAP7kDolMbPp+m0DXVCjbaZjeGZrSV70
U8xKQFa4XPUPohxR2ZdiogEOV98K1tnjYmqK+c7MQeaL2YkNusA1wabIjTbGOBCvF4STmNaVUQde
6qJcHqrwdTK+nbUk77yV6J2Id47mwLuxiTu3jymhKfPcpfolhKwKKNPaDEnkAvzyykPosULkocs8
huQTGZMTypV1826bwD5fKLYky3RvPK130ipU4n1P002m/V+/Zv4jmZAydAyUHLboCdisq5xxqO3o
BVr2ORONVnY9vkkkDzdT2WYYKqtdpTAwD6wIhxF0yqSGSFGYfoBRs5inwi6k+BaiFXAM6DkJVcr3
wZxTixgYQmpQIM1TAmiK+aT2rPhdU8VULLrgnNYPdpVXXHd0v+8hxS87GXbRzh+pYuJzQqZci99o
vk1OcFYxykIzfxUfaqz+BAu+rxc/ZZMK7+ESG8/+bxjZVaYaZInB3vXZe2rwL3pPi9kCc9XiUHdU
15zotTU5Hfbe/06SrROiZafTPIxWEsm65oNEDzg4XqgvhrF+/ve7GkTnoLJmjO1oVZfjyFm4j2mC
ucfobGVph8CeEwY5pIHMBiOGDh35WYj9JpLWU3ONjLfDeiQoJvrT7anr1Cg9+csM/BEuCDLI/tX7
mQqWtAERABE8l7OynIX7QcPIaF/cYGnmpx76nzf/5n+mBYuspJxW1cBpQReBDVwbUYVQGZVowINf
v27uT0sOdfSQPQG518qPcLM9WTIU13iKJT3pTNzCRYV4XlowYk3+2CM7iSknxriX52I1PHlOtpux
bXXZZtge9cv6LNDetorWh0wZpQkHuTULbJ9Jt2jecCfR35d/gIDVS68ZonPjxXgYmVNeK7yx4zNV
ap/8EPrJ0GtPPlMpu8YI6ixwlplmEZnqQR/v1mQqG0dB+bRdXh1cGwlYYBvCdkrgBgx4I0KVpfOq
gEI1+iYtbB/rBLgTVMLYdk+EojosaWIGW8YUDdeDANY5HsSJT0mPr2i1hAUippMsCXQn7zk7BCMN
sEyHiLa9ah9khok6zdqKeYTIf1VB41i9pFP7lFQuKegUwGNaemI5w/djSYrQYSsXT2KBeBfzhiER
qlXbZRkBOF1XXV1+T25iQ7D8ZiKTNMnyxehe5/kv6qtAfAeIEqx73zNzVTLo57sRpSY7Kq+7gn67
aaHTAJfGw6xBZNsm+iRIJNQ3INNblbag/V9cpj7NcsodA2tYmzaGueYKar3O6mbkUCahOqu+GB4F
dTkubjxEqZz1XprqabdayYqdEwVSN/UNUDxEpB6IkjhLWn4Iiy97NGKke/zSvtnYRef89cJgR1ls
48dVa6zmv5Z0ZDMoOdFe0vtav8NuZnKfeJ2b7cNz54Gg2+Ki+toH7dgJKWiHYuV13iA3Ue6NYqzF
x/6i1K9cbpqGTrGqFSQ3NGit2k+OoqRj/3h++2A+r5l7+esVeKrzEgb6r6nNdH2NsHoY6RjJp+xI
wtnn6Jzyz1/0V6VxyldnYflJbc6nQeYnPZTambIFriHZPkBfs4BF6mQOIdoCSAA09tM2wVzqwoY9
DyJ0bABC9nA0NNLI2kYCoiIYNfOxLgR46k2+kkQnBbOA60TeXeuAzJM//M8xWcFSM8d828vBz+x7
jwZuGdIKfmXiRFb5S324TtESlTlfCNtQX94m6fggd2pvMonmdby8ea+nLW01XligFxuXHkHix1jv
guN1FZ57VvBbHQiIza1jG5SJPD/+JRrg1fEUS3hJu/WGNIi6vhOLV44S0ZA4pdQvuww8eeE7Z1kY
1diOdTSSFrSjbHv/QmbvemrD/PzPr7c3yPlPtMZOp/xHZ048UJnbv8JL0MpslGowAK0gPoe2+TWV
n9aJWykqtfWj4rZFh84PHbUwhHdXRH1L+CVfE+Ps09sytORibF4kA1d++mc3Wqf6KGCFDCBsz3hY
iiCE6nMVFFdofFsGHM9HdMltmAxqv0wXkPkJpR4FuJ54kM7cuqfRf4yCa0Xqa6bJ1UcFcd9W6gss
D4NKwlbWdqZDMPACEqgQOWv8LFaCpheEDsLZO/Ykp7zu+gmYJZ4d/avFahE5MgeUq9QOjw2AXF1H
FcvEV9PaPjaGkhxfiFLQ9jllWbxNCn81cccfHkPjDuihmXEJACBAQGP72jmmWmi8q2G7p8FRMe68
gtQ7Zlb5+yrAoJW2PjD5HcAcA+FaTmPQs9uSC6hC3PF6qGUJ3w+7A8XwcMcQ3qnN+IWIwpi9PDvI
kZ6jOVSSKh3Izjfev6vpGV+6QYWndM3rNNDPr2UikGaAX+xb3DwxmztKp5KLTM+gIRaDRQQbHlG2
IfIV5gZ8qj+hDXj/uQZnyjsw79XhSscKomAERTGpSHC8O8TjK63Uotw+llQ8k+BcDLSLijdOH1ab
d8CvfsMxdN8SJNvxg6Nptx+yu3cZChGI7Y4gQYKnqJODnZ1YD70ueI9984TB/yJHZs8KXFHV4c61
JR0vkMUAtP+kY4ocWaHQHbz2azYT5lPjTTTO5KFnII9OxdMNmuckxcFOnFZByIJ+D0G0w3lO9PJr
aV2gpBV2fpBC5bMyxXiUfgoqA/kJRUCj1o0BqUaQL+ecUCtC1TesGpUgAWorgHuNUeT5tXuj0Htj
76UfBaU3GtIt6dsw5WurNYJHLRJaEfOzrk+GtCu8JiPT282MF7+3MkVDm0q+oi/qfmEe7if+fuKA
JxLPSJ4FA1Z1o0cYYbqUgIwFciC+wxYoNW5l6CkB6X568esmVS0aUyr6h/KkX/fO6JH6tPOaUC6i
8oIRZlosR55eXbzGRbXvOBrDHBjzCHKyRKkfBRxrWbqM0NwHaD4LGqLRxZ9LThnwGlOAa+32Fqbi
8Vdc9sWHfF3hcUZCTOoVgJtkFjynZxBt3WEc26DlwK6701JbmW7eTvS/lwyZ1LtDaNH68XFzDTP5
++Bg6jYQJUvqXO2Fn8BlrcdZSKw6APiRQ6Q3xSryyulm6mF6nYsW2OoIUfYl343XCkqW8+e2DD+P
u61Gdn3mPZTlrkLbEYT7Gvm7DCJj4CXFE2H+WcD/2MWIAkyUQQ87FJJBg8d3dLq/25bWISfCGzaU
Dd7eS7zQMFYCPFMmZSoCp4/U/nQ1peTQ+Gpipl2CKPCrtusa5Xt4yIS02idZlQKh9XWhR75Cjm6+
ujhE28sMtzKpFSuISnfFmA8aXphiCxaAQVwBoM9BDBURTvjjvLUD/R3LN2nRCg8FY58rPVCS1b0Z
eihK0C4EOoFyHzBzDytDgAv/4M9envm+8NZFxU9WG1jxQ2kxMGwYaPly4UF0e8xp6fzXcSeTEFhL
Q5xtf4ZpPCVP+eUtymjOa7uQoeMyi69WM7Nzdr10DGbIbTLwgdK4eafqBuNK1i0r0FZpwJtVtx6h
VGY0bfA/IOW3TGo9CTKTkkrc/XWR3PgcKbZ9m1/9lKnUP9jeL7KiEIZ7S6RhnOvpW/vl3K1TnfbI
e4mYi2X6eYK/hOACdQkIGuQYRlho/AgzWMwC2hcDNNvvZz6A8bB1N/WvmjHaAciFfmMuRPSUG9DY
Y8fGvQV0luhD9KhStSbX3wEgZczqZP3WGYJE3ey2U20U9/mQHByiMXL4ovlzSKJf6V+YvqMiAV1K
LbEAbc/IUdAbi+k6P5RDCWe7lBQtutqd4yi6JGN+MKkt+PMHHEIPPQxfJ+DJv7qn8qoF3B++pEGT
1XQXscKKbc+qaKkR2eycBz8WsOq5CdrAZlRQX2DGK188MpgM4E/rw9Z+7U0Gw/I/zc71RC0pXfE7
gZ/v1btvFoQEcNYALnlomUgzleQ2Gzsbzh5EWxUtQKR5q7gHFQjBLEcAHHuSK56KRpJ8SM5TNZvm
j6U0aDyUpdjfobzWDflAmNJWFRsQDQ688BLlc7CCLQTpgCStcipNqLhloHD6i33fznlMPBnvz6lC
mLAaUkwBRKc5D42mEJ7l9EO8QvZNL35ygeUk9yAnN3AnNHC31fhpk7s0qeiLFeh0v8S2e4FHsgm6
C5PX79qOck6r1MX4mkwDBOhF0xx4wVbzZrVycR2wWnD1KaJ/ticDinEdiMgRCaj5Kp/ksc8Mohm2
T5Ne8AGO/pn12XzmNbVhZ0cJ/TePQO+TsifLlz7jRiP6aOJy3mzSiaQQMnqj0FH/COipdqJlPZGY
X9E2ZylZeY+knQRB3bCeF6ORUVQFI39Vp7ZcOkxBxMLjndRAubDZdZ+feww52TQEDlhM1T6h8EaR
Pmi8sE1IGfS5WQvbnCABQgSK5ZZEpYHDZrjtHnXaXGYRvyjgS8YTDhdsmYlPCJW6qeMVT7tN1Ub0
g0VaxwJCJ6WtUBXXInaEXW6Mg7KjvibDNGn62l5GUQWUtOCJD4c42niHMEc55GxfRL6WV4wvkuO8
uQGCcw+0Zim1uBfricCvD1/EOKWaHYBCvg3k2RceqTXihHXrO9voIIfwAmPe2G6grdYOBruYLmFU
jRM4CTH8qShiw1pUa+F5E3iKZmLfA+ZwlJacpeRHEInb+VG/chIQvBa+ESrzk11Bx6ifX/drjrq1
LszzE2kbLDG6lpxcJSoYfk989a1+lon7hg5zk+f9zzWWAry4SAjr7zY3bdSu4+N9vITbGODBw02U
thUZ52Ijnb1V3kO07bgctgbca1j28kXPi1Z7HzGfD9AYVVXPGqTFV9YsOj1O+qDtdtv9O4vXQZH0
gdohg/KLX8pQEW1LK4B2sFYn64Th7D8eXcCOPrS1UEFKUzccmRHD5Cl0Eh6A07bAvDmeI+VN4pTr
fKUlnThbPCchy9jeFqhIVPkbnwkhDZHo4YYsiFfphy65kQLi3tezsbW3e5dxCmQmyYi9jZNNM/pr
fFz0qdGaRI5P/YgfwaedOMyIBprrmsl5SPdDR3Voh0YH29GIZ02RV+AYfVe0U964fnXDmdIKkXJC
dbEnmY1g85drmDfrfiVSJiKbHVBOiUWTrMe4vo9/87os0FvVkNStjRR5qIupjV4P+sxA1aB3ce/r
5+pS/8xXcksSz6UljpoAmhfHeABR0vxDaZZaPlFgaNL2ryH4NcZAdm3k7dl4EgzFJ1lBQO7kJLb8
VMbj1f2O58dVKb0xPyz5PIIiaptx+ZKW6NEfhmPOwsWSPXEudxFwi/36HjzdTe2+c7l4UafRFQz8
Fu/j5GDeh0EwNPFI0t+6EzKBhWibNQcJa+5UCLSlFMqzPBMDwwVfZVTekSTAFDGSJn7DcbCneeEd
RCHXLSHDrv+b26EBPigD6nXEM+dXJU+Ef+8hMqoy4bxSWzgL6g2S4Ma/yaURh6gZScGnIt8pP52L
Q4S0BxIsBn4E8L253xJBs1iBsTQTEYOQg+vTN4aPPZ5iJ452o8uSaeF/asbI2kXEy3/g3nk0XFQP
DWEDvP8LKlzBM1nVsbF6nBbD8ypU4g8CtaMow8y29y5fyRZeyfgfSSS07DlPys3cwdqmcT18sZC7
78L9xSr6pnfbHSRIXUFis+ICcNdVflU8G5FRMZymAb1XYUJQcr8ZGIkDteArrnLGxUIi9lj4oPSm
rq2ropqQUw7hiUpUlNFcA5kqgrjrxxfKv7oijunzHP0irv0bvbkbMSQkNx9PhRGHPMH8n6DS1v4V
ufQoGxSwz5dXrRkMKebAJosQ510IKhAS1vVh4DWqbaYD5KiBIXU8ANU81fvd6ftHjmWwfBRahNZK
EzAvHhraabGcFOFt82bx2YpzgnoHT+lKGqnyokoDv0XTXk+cBXy7bunLRWXGvhlFQ2QrTL6EsEtf
XQsjnOcOuiBCofcDcPDUOrtYYlHHncjCC1QKnjc9V07grJIX2NU4Ujq0Qrls0jECdnsg5eHMRtWG
+/wzL8bWToPE6Jj+sO9xwPC36Ajkw89n6DghzzBNgzAbXLD2ta9Nq6dbYvwQtEADaAUQjCmkvMZi
TWz0Lry79EUL0wwMWa8cpl/ITgvZqKcJ/EAUz2nmhsQc+wb8BpP4YMf0RVGe7C5m85qB8shMvoQR
lHGcbU6nm3fVzRNr4oJPcs6vHiN+oVJOPq54v+UVk9thwmFcEyiEo8vlGaxaRmISYZDF2AuE8iqC
QSeAEXH12PhBuh8JI/M435HCjXl3i+ihPI3gxKhrXhd/HtLUa9w3Ips0S5RW6nJNAm4uCl4SnlR/
z8QvargQdwz0+3KMZ/oChwZm0FjYNJxzK74CHPH6uW/L4bJ1qHx6XsQhI/zEViQdvoEZF6U0fZ08
CddRwYNcwdzZxolhHJMER7UQmYu+0nLddDfcgPceguhCbNqrDRqx9HkLUgWL0LfGQUFpNj0vAmdy
k2xsM/IUewKOD1SNxy4LNIprzXC4qvcNS2SeU89Luwb6wHjrJz0e/IVnKGvlHqDRRbtWA0GsZKUQ
PJl6i+yIY3k7Nb3IZBA7AefP5+krBzYOGcoP2phBuB3CaSe/f+Ps15xIAkDeRJWGYgVQBqjrCtNP
5L3w1C2UriuWAT4xnt48cNoHnkQIn0nWP+VlMItcCdTuLw7o4isNJZoVLulMtMyWa2xcJG8UL6ed
EUsyZ+oVzx6Phlgrd5a5Zu0JVjz6eRGQxoYvu0E4DRW8Nq0lszzyCGHFP4RKyDvu1mIYZ+9Pt23z
kshxZLdaTxXLAJj4bKXRWggArAF2tEZU69ST+EN48Qvtg7uM2Sy1tBBiClunD+MOLH85mIZe/Db2
EIsIBY12LkhagjVXonhFiDACs9NsJGJxiGU1UmTSuthpclmRyJebCqKcyk+NHxD0tzToCxUdJslw
Wams2ft93ewVITH+Kt5QhIV8VSrB8ITHGtNydp1nZxRJ051XxJKsod8et/6K0qp5itq50a66ld9t
g2ErKFLyHDE7guS2RYxpmPPcDONIhuYJgHUMAclZ3Q8pEpLrv1pHh0JDFRDvDnpTn4mvTzQOESO/
CDzPGsdtLwgvHMRYoQctY/UHwr5k4dh1YjCpAQkbzSJKgYl+aVtHYdISf6GQrIIsryPA7xBKC7Ah
OTnrPMY5cixMdvi0q4fQFvKznZqLGt51eRhusTiOh8C6G5t7gOYDFwV9HH4LPeZB8bnuS7JU2lYX
/lV4txuwxmHaZ9ZKk6lBrECHqzmUSx6awBYd5Ao4YpmRKxeCZx2DRbPHVj96BHaMAHndBacqpQVn
xOOsE0Olp1kBSUpMhjWzLmYXXhdZAZApUHXduoRcOEl42Jg+09BudfYkMe+hQ2P4RGyXFegWz4cN
L7xOhG6X5JHECW1dvbqof6hzc9/JEvebKNdpI3nMGNZ/Eb58J6jPruNcMpuEf+3YOIBpw7jCzKGX
bfCyXTq+sc4hZrDTrmJVGf2H8T/CGjTuNnWq4LOu4RrdM4KpNDmarGyPYJi7OJKoKZZRsyAoEt90
WqWTYbhWwwczvAnAv+cHnL9vzNSHIbpFJY52BxjJJg1FlntHOXkEPFKiasayXODhdHOkVC2asJ8f
0ZaGtycCNG2hrr4MPq2Dia6Ht8xIGh+zfE+1QWaUCyVyYyL3av/JOmokiabC4XxLPFQvxwNkL9R7
tfyk9oIjdF6Zuom83/DfbbWe5eF0vomGu/Ydwkoz8xrawpZ0c4D1066h2DgWemy8RzgcxfHGkC48
STbz+Cp1ScP3NEWPvGt28w1zAO/74xvjeKkP58Z0CdNpiRjxbyZFp4vm54VjmnzKj3IaHq52jMur
/Tmio6beSd4FxrWTGiORSj1qxZvpmUhWEjB9lz6nYzqgKUYhbeWbia6syYS9uKnLs0kxfo8gfzZr
WaxBG6MvJ0XtbeMnNyV933ncp0QiYy30oNpP1E3tNtGRthMbo7U5B3Pqe5iJhikvS7cqzZM8BNpW
WDf2iiGGO94tXQCBw+KewwsLd0LgzXG1sbFYRrOkeUm5iYtkUqE6nZ9G3DinlpjrLz/8uCjS2MAv
3AClyxh1AriQMUCGBhnesSeuD9Qc42vN1/jfSuLYyJPg4MuAwXBVDMtM86zVdLMgR3P0+HCCDlZj
PmwHU75aINHh3ie8hHD1xcy0AoIU0Mmyfo81o1UHriMEhJcVPLKEnpMdgwP+wZq/B/daEtwx5cAa
hdQFjXwK6OIu0ku55u6alTloK8YWV9cMIpysOv92pvspvjiIjS9Blmx74egAHxMw3BFxV5X+ptIi
5hzlkq6UzIFgBid+JiIKETTzu7uOPYSAGCC4UGVrVjiWX3tFTTdVPmd850zmt4o7kXGUzD1bEM1n
xijGRguFgBcP2fx+I6DVZqSZICTPfSNnrq9qMrMrzphFerg0YzzDcPmPt7aYjhE2Ebh1A2UN9Den
o0i3XYHViiuN86ZTh5+EaUo9ilJAE9DuG1MdXcgnPgIw8FXJ4QvAKSRU8VhDgQDrBjBlCuKpYcVi
MLcRYa6UPstrJQSD0QK4B+2Y/ASLZHhk813o5XkyGwCJzpF8msQsU5VhtH1oEDejaIpLq0VTVLvl
h2epynEPVHrIKBj15vk59/wh6aSg822tFEYdvFMcPf1roNXE3JvbY+tHnfXo0r3c+YnngPcJSWFN
NYeNgbP0iWXs7NIJRjEyYVC8PtJyS2IP0559jvUGiIdw6FQYeM0SgILWiuzBhxKjiHpSRoqx0WnW
w381VALhfsOdE1KCoPiNUuL+UnLeUCAJfNsl4GZnH5OpwvjjSIVnKpVVhCFk4Jlo9xg/3Lo55yra
30WBcCJIyjsCRjqZiCTZWfNkFK7QYMYKC1c6vvm8eAVr17QODaDpFAJY8m8Xf3JTwfyh3ysiql6Q
AVmwzDDWkNVZiUtzipgFH1I9Wq011/wpyl/RLQUMOSuOrXcT5aCpVgpGSOMjVJybSBpgy+fovTrG
3dvPnzbkCGNg+sPQFqx1f0Fn38gNsClx/ITgcZWUmcm3P9TO6HFpYPPvpP0+T/tg4xM4JXravJnC
vo+GS37PALE98chPiYzOCxNALY68Du9v8o9jiLoRQ57TSLkwzlfzkE4DLHoJpPrJ6XHVL1vari4s
A/XsKyFDYs90DrjV+BmHBZUMlg7wb6eSERK6/fZd8O1ACvTFP2U5PPCvdMfwJoTkTKrIWvHRUcDB
qfFvlGUU6EGPPUvdOPRBnHAD5Rq0xpq4VPaULUeyPzM4nPRxdn4BkRX5+J8k39V32e+O2tjpw7O5
6z7aY62nATUDm4pSPkzBdhFH0O0tntJLAvNtRftDl+K7k4yqLhZykwHHJBs2znt4But6XHUIqw/6
RfIWyf2W0b9UMMVUvYVlyTSszFc5u9DXgqCsKnfbGcmPUZue2uIxZmczJDcuDU7cAmDOvAp2orXq
E3JdXCONkHHPFWdFx5nj0ZRC53ScMzB5eA8x6pCklycwAmlWjqll1JYYPH04ZEY3LWbqIB9HXClM
htFLaQefok+179mxpFMncSGSHWyznayZoD3SuzAAoxPgN6BT+3ULXi/67PEyhaQIaHeTXHgPyxSC
YfNsddnxBXBJt06EPqH1pPocHRmvH0wXv+jaV+qS5pgMbsdt3gBHxWHs8SRZm7lSVtdDGXioR9ZE
Xmfzyyt5XhplVppdExXp2TljoXK2WjFaue644dRuA3AKjfDoX5RW97wYPs3WAv4uf94Pe3WcrCWB
/okU1jB0a5Z7TPNpz7RWmpLnnRSSVtbYEUAJwFx6SYN6JYLAn5AR2sABquuuhWKTg5lvu02TM5mK
Xm7C1/77FcG9w2FkPzEtzhVHiI0oHBV3fW2eo6gU8eclggfVTSBNv1+CCdQHv6MnC53RoiPe1bOZ
iw/9j6HuG5ZZn4jIAPAKBK7zc5KxK/rD4HuWI2zmubla1kb13fv7a2dHSMBWCI8MOigZog17Iw8o
39Ed82Ekbbqx3zXFjyU2L5exW0QNTFier87suyHsoKKHJcXsXSDTVZs8RfbiUXs4SShGzHSU20Fj
RIEuRPBSxKFBxWYyF/ZbomkaJQ8cij2nHnaUtl8nc6wMt0uBiHmfMVoJ8O8vA6uofBlNruOmXTOB
JzX49baETrERbcVQEvi5oa1diTRz2MkpK3/bZ7+syBCVLb0u1Mseq0Ivatg8/F27wb+ckJrgOJlx
6UxaSlCfPoxbj4LCxNDs5rWLDScEi3eryp4+xcEAvZULJmXrNkxYXCsXq6mKdl/WlNx24UaG+DWR
5MtkAWCcdunTFoLlCkJ71gcI2hA1Fw1cobWM1Mn4fQAo0CCfRPkEaDrMYUZH1tVmcUKuG0kiYeCk
qkwLz3rsUjK4vUyPbm35Du69REcQCPO9YIMbbBYT7hv4jyWsQ9ReAxugddPEZuwMHAsbo3zTtML2
rQBY3s5032b0r/fgGzVXwdqrauC5ZZ+GfKbZveREyhvpaOGnIX/sUBbtAbbPdSjh5KB1dtPebBd6
3lWNwBzYYP1EAj2my8Hmh1bpfkZB+tBYEfdcdWtf1ucAVXdUxoRNHRxYjB/Cs5/Diy2r4tphSKdy
uQMh8lAXmCc3GAgBqcDPIcecSg8CecsDMJDHRan3W2uSLrQu9OAiE0LOUN60zrd3IoS7JJtq7HIF
LTEg2dcijhTyh15QSGtUkXBzgbtl1NftdkHlQWDT44X4zCP4wJB8y0UlEGKV51cZ92nc4YE3mzMH
P0aAuuxuSXNFcCKQZfjp4frPpfHG4aZL8lqVD02FxncAUZP+yHicr/dGsuQONlDHMjBaH49+z11g
+DoPMmfHylkbGVdGCQAjzX6jDTASHNiKTNNKp63WOTFQH08GAbHSEYpAmqID/aozJgF+DfmL2MoY
G4y32OOT415ui/G2r914xlBTzAU9awhedZsc7Wjssyc5p8Mxyke5BAol+IpFXUMj/jjexAjZICgm
zs6vRG6FepM9Y/JxZgbJaMsvTTWCO6lkzA5LYyXxX7lJyfTBbPSWW/kKbAEuPwwdYCuZ+/rRSQc0
E723+O9UGOtblD+W18Irhs5oDf7czzFoggBzcYLXKj+BkFPewdmusNZOf01DYT/DdXhFxmGA3pjm
QnBK/Ferz+GNY8KM/F4jlFQOs0RyFYwMXCX7M4O+h8nQ/ukoap92TmlnO8DEwxJT238btAl1K1vj
ZPOU1wIuaXOaJiF5/IcEMcDXoCIe3v2iLJEVIVOBSEOetx5EAnWFilCJxQPzZZ/fPINu0CEy4x6A
JDpJb/CB21kmSEx/vfj7ERhsUvbo+q78KBa3HqoyoKRZTUSt4ELQRZnP9VALmCGeTqzK+K3b1b9Y
2QELILjDBhr+ciPjf6z6UKSGA+lEJxOplTcrhooYhpjXU4fqPjwNRgvy4W4wVukax1TrYDzZEDcK
B01mYEXPnOF6IVQb1klEJCQDhHFgcJfjaYTWXq4/GGJwoVSGqbJ5unU6qQpC32hkQ0OJnb3OwECG
syhV0J0mhLLZ+BjguS1GwXM3BdEDqbKPCXEwjcLwU5YWJaqo2lqDYxGLAc8zyV87dun4/1jEj0Fh
0BzAVBWGzT0DX3CCzWu8XKmJvDyd/yUn7TTb0YpnjfYv5BkqU2V8j7XQF30ELRzr0SVy8Ztp00ad
djQv7FphPzigDqcb8ztmtuBB9txbCuh+QrnX7PJ7uDMC5jiIEhpSkC3Mh94OHw3dVM2zTzDDl04f
0KFlt12GrmhN9kGzzDYQxx+jZX/ykILMODBrvpmp0dPovmE9VLpy5HCm+aAqNznNPBVpu/EHsaBk
g3gzPF1BUU1Ds185tn9Wj/Dcer2KzfHyLfk7BJu4GbzlJhOq1x8+J2+QLvz2UwWT3okWT4RO4o3V
gdWDunsIXi7CESQFxyJANJDalYAra5PMF5Re94KlA4CIKYwpFzi9W7Je6NtFBDTut35oV33//eSu
5W6AjPF5eJoe5JNxxZhSokdt99+UbX7SlScSoWg/F1KfzcjvbGYOTliOi9gfFhLrHw+0YANQEUt5
ZPaeJD5CCzy5I7jnLgiiUNeGtOGVBoWu3r7nND9w5mh2f2P6yiTjXK8Yd5tHlIFhCJi9s7C6bgzd
M6FDO72B5cQyzK7TYOw2jQSFK8rrObl2XDN/XI5Ajy1BGZBQ1oT076LlanT6jvZ5Pel4DCjeMmAE
La3nPK6bTvv7zmImkxpa+wuYS3o3Az5Pu38VgzRJJrYCvvvpgdLUDPckTr7SUbKtGnEn/xUSzT90
1FbENP8jjdhqBQPsDB9Pui0d+3D2EvZP/VaAnFesTQQtS2UfpPeyLQEN/Lt+kxRvdexYLMNd+cSu
rfG80HGAvBguQBMo8/0wLs6ZjPItDwPTQxT2V0ug5iaJ5p6nf7ZZqf61qYHhnr5/1LOrZNQC/SxS
DwZEvP/Nq4bduQTBQA8NO3rQQAyHOwHu4DdUFAD3OyUbhttF5AUus8WzvRiE/aOef/zXwS6HZtBS
A2z5/KifouvfIo8YQUgQBfOzp3JACRFopsRGgjYRK8mhtJkr8eLMwBFIx3n90RoBqa3GZo8RyqEz
afdsHiqLf76cHkYhkrDP0mxQAUasmZ752+H6yeMOZZqGZtHGqm1GrO6lslCCr/9X3fhPNdhLgvqv
ZOyEA7dJWngqESXelECSIr/wiAvZ1aznWJqNLGgG27IO0U6gebVpO+95EpONYcXTLeoJRNL0DDXG
k+ctALVYEIuN9LVBT1Y0zSkrSGY8NykBVnqDlfbOy41B6uGdyZfGPA/zpstPhKANrL5NP9dF5P2M
lP6XVvaFTzf1b1htZIAYgspcN5Glniiip5v3cqHM8/UyPrwuArVKVUwevrClNzvgcYpOzMxXZ0Eq
TGvfQQFtiJ6d46CdL3wIAq34sqF0GDTwNjibvCaiSXrBWjkeN6v+UEOX0KhJboEl/y4oGtBLiW7j
MpCdllgR9j395ZbWmAlRQDgphl4OFle+mU+blTtXG3d3JvLEkj1Fu+8OLovHp9XgOtz5Ahy0mPTd
ihxk826EvqgGtoKMJFIKYFl6dJn4SM2dq2cIBgh8X5f8hMhECkTOn+Ng7evt2QGsBbUHM+BiJOgW
GY5ogId/V2kV+CAd1qYcpd5CFuJ8MNCgNdxKzpbG2H2wbC9pzlnsiwnSC9+/s0p11PzwBCZTSjbG
wUUdyyQKnuDLIARospC4T4QOLRA0Smp5NHClukjZ2XPAwWYWhDJf00LZe8zx+0Aeet6jdm/TkNzI
cWNCYik264I/CjfL4jrbjLJOYRPTSwGjz5H1hbxiVppC4dF1N1Z3Nwsn2qImacjdo/LBe2/pXBzY
nifrUy/nvPveT1CWpLBzCeHKFIAmb+9K+cdLZKFoNzVxg6/BU1gc/m2dMG9MKYOPWN+af2+IE+MJ
eh/rBdPfW2NJ7ZGCInuW2ih2mvzJALkZj8qFuCRv26Qq4emWtXsRngcJKlrRtPcKf8dPgb6J8Mbn
SpzEKltvucf5jrPukPgpYxlO2rIXE2J4WyrwWz8btN32Ooc6SeLEj6VSBsKif60+RqgHm9lTmzhQ
clZDeEBPmqKto3VSrUS9aDrwdllfuDgsJz56smVsUvEFS45b8gT6hskDoH0jg3gOktsIjcgyP5cZ
vjtxB6qeCUHOluNerL/R/0x3RjCLdHB1FDFh637ZWkPRIJjKupxeH9p2zlOsbgDqsLozkEkOHHHM
cLbeMa71VexIR1B+3+6cVLwJbovBKw3PRgbQYXR6BRqUZTaqwCqgxrWVCPk0zl8nAOGOQ+Uk1Mzm
yN/gNFkOaDIJ19jsqns+b76XWK4IxEmUmH0IcqrtNCbVIbjCJJEDWVtVtv2K/c51DGwKTFvwCNjx
HVc5r5dtXbNKR65qJWdO8eiL39xZvlUXtmaVcZY+Rj+dgqtYSQhbOTSL2vb5qglGYfbOcmKLM7rR
UHWXrO8udf2z+7A3DZMwVhUQHx2lXeaCL62sE7oqQYb0qLBQqWSVCxodOdL4Y2SRwRwW1R3QBv2y
hH+DRyym/ZSEtBsiG2ihjdD5QAmBp2HmsIBmJ48zz1PHS2Aiq49HE1bLJYOJI7KSB0kCkKJfX8f3
4TgfuFRKIaS3eY8Ey+OyxjAI3ycOmSejXT5DvlT/D7IL51r9TcMkUgM2UYR2wjYHMF0hDRwm8QkZ
CQjcNOMw5uFp0WyhyULvaDrNsFKsnh+Zuy6R7LmG9KCynZrz5giAe+22le21BxTTUQXzqcu5El2/
p1Rdzv/+bHfDaAm6LbZVsU49umQt4vODZ6Is+iEvRzCKlQ+fLBDBFSRh08ssjpsvoKKS4EyNaRFV
iBe2jr/cTznRACalOazt5EXCtjn2jMHRTydvk49eVAEhGGPE34sJHaftvNS21ZL3rUBajAqO6MOO
Ot7nQ2ku5wEICnBpHP9M3o+fb0unDd6US7UqHv4NfJHH0BBxh22wwvWJFuH2i6SwH3KIxthlYiVF
TzRd2aU4fNoxonaX1UfIlY6knLZpQMyaWr9CXhi0v1imnfMSM24tW3zLhbTwQsIDMtqOOplIHT1O
EC3noPRmHPjz7839ZE95VtXinpBiz3UeIhYm//NPK653W53A5K2v9Ace0xEGU9MoeTyzNWeFCgS6
iBuK9f2pUnFI/5uiHtx3YbpmM/1PPo/tjyMvRc6c2bO2jKem+FQG5/e/X7lk35Q/7EdOlsBmPhtg
UxpQyavGYKfmJ7WuyQDOEpZ0MJeqeZU6ei3Di2R1ZQ2A1I/smjdzS39n7MUxabvVN7Q8ehxlv5Cx
QQUGtUr+f5JYF0cxsJ9Ixj1x4/1qqfYiUM43lGX88QNIvnh+xNwVo/ofTNBFZ/QCDNaEjMqMDBd/
xhJaGQhCm6sQe3FbDZB0HioRt+9AGHKiajEuisWbbQT+ge9VXNqOFI8Ty57V+oblOk1U7O80ii00
5FhfyrK4xwc+cnn4f6TjfuCpGK2Q2Gr5VFTvIf2/VFid9mxKEa3HipZuQsgplsq0ETqHCaVGz/OR
UE1movqIWyu1KbBYpYheL7dn8XQUu1MmaMjFmC5jmQNvP/BFnndR54j7RfDsVeiaDqsdfrkfRIZv
C7xup5Lneg+lbkMMVAbDVIWPWKmTCtZbSXvnZ/PpwI3Vp44ihXgLqFyKRAuEtda3UirWnpj87GuG
N6EE5beufMksVGq//MuE/kvkquVkOHiePtfLF7ZOEjuXuc/Wisw/ywH1n+AKam33z0rLAB5CBB3n
1cHvuRK++EMiBtpq7RnsEYeJE0EEzuvDrwp5sA4a47tCAArOYR05qGYdxCYwJ2N1dGrvLet+/uiL
OPQET9zIO9fAjMkEnrdHtcP7sAKyzkbg0ZG2HpvtZSubvadrGqZsvT3541sP7Fd8SK+Mo0SLxg38
YJpgV49dG2OPI00otMIwx5f0iNVLEto3FauH/3+1twq4TwicbxDWGjnq/WZc2Xh/WYgDkO3ViNO/
qIOx9dVQzo6BdJanMXtViHozjfGba3PqP5PHXTk9GWuVwQQOKIZ6IIs1eKoNS1UiUllg2eLXnEx5
y30ILhLxLXNxI6JL/oyRNB/1ZYrpkPfb/g/bWQU7JJqI7ETZ/nmAhDfQJe+KX7ToJ4tna+BjJdpL
aHPnZdhiibQd8W3m+KbeC6o71H3ElnS8cMFhwsW0SGwTYE/fG8jP1jQi3BaD/DBjzzykFgss3GvW
Jz9RCnakO0NigmMpmIStq53GvWxqo2mEd0fxWmeHiyyMz56TonJrt+FLoS9I99rXh7fcSBQVjcE2
49MP6Y/cRKaCU9YL+R04sknqVK+qEgWI9FG+cg7TuKdldYTXR2CXE2jUnWcV8KJSrqkxxScw2NU5
IFpul0QX5j6kXHc1jPMs8KnlM1AJZaZEH886tcVYPbGOoN5Mk7Mdxe14khNPGoHIp+AnkDBZ7wu1
TI9R/qV40QdMIR71Dy1kXeJOvYX0vm35g745lqOrLMOjtSv1KJhviPoLaX7XXDmIre9vRYUKqbIm
IE6E7gMTVWpft0ybfHAPswrZuY1UjC9WyVKLMTKgNUgnmAoPfwqHjcSA/KcWv4eq/HYlLKe2UIOS
/fS/3gTh9P23S9wXAhifKZzwvfUBxf4x0YLEr8ylW2Ho8Y+kLCJwI20qGTaKNLHtlGXhu1DiZ+8v
AMnw596nsFLVCHKuLqjFu3vQ+YMU3jyu2l8tTlPGlKk/Zfb4Yxlly1yDoFxHuQKxrjkNjWmTn7pc
RJyDQPB7+S7Mp8hhIcHY3YeS94HFGjFQM9gwP9kffWoWyr6SOw5yKnzMG4cWpZx0mFZpioRA93u2
vXAEarcvoG9GZLv3ICOFK9PJs4ep330yDdcCUZgDbex4CpMFI+vw7RqIuqmmfxXVAKkdpWmJcg+O
I+jzmTPk4SAztJ/W6coOBYvAn+3BcqYnip8/+9RKXFQ0SyYLiyiIznSeuF9Cgpptppvg3yBILDdF
YZcGGPP25zIOh2NOwGD0WlfXBGe3SU47SCyR7QqLrpyHoXq3/Y4B0pcy4II/1F0c24Ad25BpfUxP
Xf4+jM5opf4mFkSW/mPJxK2uajntsMUI+IsxQLdUG4xdPPhuKTDHZzQUAM5yM7HfK9uhw7fncg4b
g097Duw6j71h8UkQ5OXkXcV+VSqV/Lzei9aARcRME2xtE5ceB35wSUKR+Yu6NqPu+dfgceZrIWSg
cyCdTzg3ZNS8VmgSMQSq649hwqdPbPPhtl2mxkJBjSRqYraGbG/c12TDg7W4vBZfFu53/HV66LtI
ez7pbqzvreBTOtrn2wlOTblfJzek4j35BrzLkBEyStYi3aQIU1qQ1DW2UsctGpm1LMYq/6Pn4ts7
xpYQfXVm/mi8+zDDv5dFGlkT+aMkmqyJprxYnO4ExL+yzVTS3ay0p1aO/9A+woFkANu9nzRYz0Ae
FTi5HcFRbke8124kpr3hQddAGgdS7BM+o9qvN6uZI4FvtjIrX7GfxIdZSlyQ1ypmDX0XF4QreIwZ
5d3rmOTHaERerp5f/SobM4105tOrjJ6MuG5iFT6+KE+wzy1S8iiHkdQPjTH0dBNeWVzvBI8tAj9S
BAxOg2AHLWjJMLQw5iokOZsrgJP2cCBZf4SqFtONnxb1+ViC8wkUzN5BsAEEwO8VAYvM3cdi6/kN
IjbTVgOqGRad+k6jsCJFjhfbGAEevkVXv4te0Htl/CFtodx2kiq8Lrc4oUJkkkTBsI5xOoOFF1uV
x7FHsd4WuPXV8kyPhsNutzzgcqK4hwxYZzD2SsGeW1DHGAV6aLcu174VCy0VjfDkCHeUY6lQRA12
587vnsungG3Lxtk2jBoaO87UEUEwapIkVMLulsg0pMxfO53j82l6erjegeoZlOSEdvd6c820He7j
/gbXZRHlsEQDp94gY9qOEDiOKk1selbyurW8izrEgmJpfhL/mVOOX+1MdcIodR+w8j0+rYYvZKD/
nVpqI1X8ZI6KwzdmpT0/o+M7VaT8nh1DWnlVF7M92FfMepa+1k9j6xW1ScYabHRb4X1Bh7+LnBnO
LLNhhNwZHA6rL2QQPvWUl65f99fyr6k8GljrGfTGayZMCWXeMhgsfOOyBqfPXYG3K8R1sUQB6ELC
cPjs7pzF3DZMsZ1Kteha7Uk5iwCL0nv0F0vwi8z2TbMIw5e72I58amztQf8PUSX9rU4jveSCIlHp
TWIVk5sAjudxJaBSKFi5agl+PuZTORCdTosEmogYSbDwXN84Wyvil8PTU9keH+CD2bQJFjIwBE1a
HKjuNv2vuSviR+aaAme3s6dA8/lrJvp7VY9ZqUFehUHj6GU8X6pwEAbKW3GGmxSLRnmDOeDXF/CL
KoYUQiH4AOPx/8fhkpTWtayH/KVwGGyGfgAItl8IEiGAX3x6cDd7KQRWfbFY/P0BYHZh0kGPFfyM
rtsBmS4GhrUIJuZGtLW6jTEDaoaOQhsn2YeAtkSts+LSH94UEJJke3+hShCfrm9qmSh9sbCtaY5c
eTQGKFQPtlVb0D4uaCSoT9GbBjXm9Rt9hMcMfzrwFKoBGYDVffenM/GUJcAvxFYtx4becFlBLjX4
3kKrHcCrgIzJYsrQ99tU4ADlAW/XZRwmWjTQbnMlVIrUGkyoQKZV6fhQbLLXJ5mZWN0QD2R1lPT5
hXWOzhPPiE2h6HVRRt6mUP+1ZKzac9SkcCVqPR2Ib0FJVYG9eaneiou7cDjLTRGfI/LRN9VI/26s
DRSenGqg5+CpIZvYY/Eogxv7yy+0gKu6E75v0qxS9TDMUc3RYnzpThfAItpgMBPwqw49G70Zqg49
yhYJ3zOIlEvdu3hAItWM+ch5Nv2gkuArHckMI8DFz+FYVasEBpwlI20eP8ia6n4CIKrU/399+LUw
W5O82wOjZL5LZ1ROpz8I3wuheftVKsNlCOpV2pLVaw+aTqc9q6u5d8UGCn0p/W0msUCHYA3D61SL
Lp4H4Hrd94ZSfedqk9YBACV53rNp89elW8Ctf33vwGrDLYNrcIjSwFro5J9NQGvdJNwiAzphaR8u
mW/Qw8VP4aMlg5nqWP9wQBvfVHMclUg2frUy2p0it9hFPxNk7EWBkjbkJVLH6rusM36gFlfGVKQp
SXbgBt6xm0eDPjmDKL32HG7Xbr8oifIEeqaO3E0dC26SY/MbGitpnC7taVZkJ0HNDSM7xlT+Hq+k
MrucrkK9ociU3voLLZDEUAkDyWMRH3xqdm0gtEVdHseadUgieaLYzLl8FJOBoHvSQ/f5wsMMyTSL
tXAhPf2GGBvl99kYPR1QXEUMIx2JmOwiJbZKxk3Z9HhNH0kpiAv1YK3HYdCD5sOmO+/EqwLXcw/E
ohoKipv5UJH+l0MOrGPEY8fVD/TXhHspq6sCtwRdKwraPdVIw3lhPll4/aA5r5rQd45xVJm2Wfbi
pD88t76Y4dEhPcoghDhySUNzpFOv7O1Gw35spq47ELjvQXsFx/7jvprYj+Rcx8kiujv/Sbmrxoo6
MSRYxFFrMm+4N5nKWGC7FQ/DeUYSX7dHxjB/AEQ9NTyLO2+McyCXnCnmUiaryBKJR1sHN1vJ/agc
A5xx4YXcxgj4Int2APPtJO/OBx17rJJCZakEoVLc8cS95HfdbmnYiVUSip0wGx0fXf0r1Bf+yJO2
+akv/GcnTwcKpOlhdAHzze7zPdmvZT1i3R0NqRmdiv/6MT3Qysc8KkAWjYpVRVWu506HA9PngWAV
duPwfgZESrf1zmQkuLjqc3WJyAT4IwpvfbE4l4rpw9VDww/fngFYxTevHNK4c9oM3QtlagavAaXs
V2Knnff4ZarCRkNhFPhEWcVgstNC0tR0QYRA0bTqiortkttAIslSfzUyMADWtCEsbUZu9IvfNq8C
1aMoARuwd11+3qVjCUGCVeaMbPgFOrpfa8HJZeyMVXeB6PXlhCYvejfFurXpaAne4rYO9T+V8My/
xiq01RmY8vz2j5eAFjb+4C7/y01kciltdj7A8ZkjE4UqHhezORe+ZjeLcbMeWzWu+JyQLoOrl9Jj
eMxC4RRLECyMyDzmx/XoJaaGUflqPPqvM8Jz0tGLg4hKl/ObAgYpUqJxsClxLLELF4gZr0IAIVJ2
kJadePWubSgVFngQhpQuRJNSxqcQGmQ9VVCkmlRHEpNO96JkXTFtjDvQLzC6xF6gDAyb4HXotA1m
vTqrOcMM/WwMpZLfkuTYhyM4Kb73O17zS4pFNuNkNMRXQEXaYYx4xYE5J8vHJu+jbMLa45RmDrZx
FueD5zQqQQGVRYMCnKhEXBIUTY59n7j7BHgM6kmXI44OKIJffWFLtSWhIscRYeFY4Hq4Ps7V0fA5
B2Q8vORBBMKXBmNTdO/PdBOZFhKUTgHsgzUvhC+5N9i6Q1TWCgQHmPAUGxjwrVQLzK8p9YLSiLsq
CaO5WMxw/mJcFqzwzbR9BioUd4rBF8bbK85TYO4u6AXvKgg+cU78rF2Zxjp0jXL1K6oYJ2TrC3/J
2YLC85IKCz+JToKF1bU9X4mwgddpbXKaQeby4I9moEsRu9lkqxNoKwZDZTlKs5L1PC+SnRN0Ow0Y
xZw22IySPNIpNqpgLC4lGEOvo2qnmnXlDD+EMaQzD0hFna77vLolPHr0O2418JzpsHSzQVIFLG7n
5a/OXy88InBklHze9q5nIGGQhIm6O76Bgz+DEe5j9qwaL9AtwUfTNMjOb4i2tLVW2GzQjZeDdL1H
+ECWKbtNFu8rU/7qwiNPfQI077Rpu0MudZI3kHzkfmhS+Jb1Q3QRQrDK/UbsGQabAe6h8Rf+dPaJ
xoFf/1vRCKl2WKy0thyTaVGxq9TKmxcOsThuUgP2Ly5GdnXlcnbTS47chsGvOXusN3NAS+1ZzlHr
a+XqsQfb8tC4nFFmvJM3SAwnif3ESMuesxf43mHIcjJGBcLy+hYoVW+WNBOPeF/62gIZrMdJbwwj
3OYQAyx4WFaBoSLPgaTamtqhoAxey8+/2wa1tWwAsu/cUrFStUTN8/N8fZ1FqKhQdrnTvCFml/MY
XgODweS4nhDZbu/ZDkSzccC59b5wQtp5Y9rsj6XYfmDP6vMu9XR6vsV/7Z1KGUBv5zi9sHcnj/YL
KaWdczgorN69vpDN4MLghHMrlpq3kzdzC2BWK5/s6REJRk4AUpq0ZaUpfIMSl6xMlRj/VXwe335c
l9jAzb6kB2bdDfHoxveiQZAPYJpG/RWDSFGBb/X9a26foRCqS1s9h5xmh4A49J/3HOSHmSrSMd/k
0h81XHj6Gg/RRf72tm2sSPqUWe8S0aUtNIK0f7aNmdXrMP04t3CYAna0OodcY49/Ve7tL87Tmzrd
NxSrfj+N0zfQhaek5v1FQWpUIpZOulYJ4btgHUR6ZnixlQbYr+LkOMY2fOZKFYoqSCOYBKvyAEAV
18Z3gX8fE59q1mAcyduTW7Mgf54qsvrB8nYmyA9Z1JxGXm68jpju4dhgR3qS6dcs+jaGwz2TIybn
lQGkWwRIMzECN8GejyO8Htn+wl0UHjYMI6SrJnA8UbhSsKG5pOssLuG2dyBa0jTopnrAm7zi/ZLw
zLy4g4zET2bUHZ5/hb+q1R15pPzKv1+K/pf4d0rzdTXiSlnk3t3xIQw2PKOSQfMRFSFossGNq4KY
mCvM48GFlCFsI2fzykTmX84xE/cSft7L1ZkVxVNiz8mPZUVa7nvKEevag56OTxzg+1L1SAruzAN5
fdE4y3YMMjrB7s2YGlJMP9oxiYM1dTYPc5nZAaSuQPN+j/9ximP0Slep6Yzu0Uzo3zCM8sd97JGp
2cFpZSP8eNSIbySHDdU+znFicoJtRwL63YEC/CMVvfZT0WfIC33GaEdjOW+CrGA/TJ4et5j2b6xf
B6UhkdWbmlYRGqNH/89WfmsehPPwLPrCmWw+2L973kobIZXeMJlR0kjgbK7tk/IkYoEmW2pLLPBZ
Jyo51icejlCL5hvfQm61bbWHOSp+B34TmoJEP1fxspJu5dUKKapaPZ8gmdmy2GI7voDz58SgbIcd
QcUA5YK9FzusEUP6ExdEzDxOG2AbkTWpmvrPh9EW12S5Hagi/8+Rz6cUba42u74IVOZyJokNlawr
wDpoK5L012ukN+0yEyWuyGpNyWSUWyyiPku16U02cvJjKzDD9ZsmeBGhFKllOmltOUVPXeYBwNE1
ICBJZ/DcUx4JXKDTZmLUUx4WbYtQOsoXK2RJf/pLEcN0OjetFZbT3jyCNfcxpArihq8QIq3Tgm4b
FQ6vDAQiraDievavx+nbvII0tqw2m9uqF3qzlqfIlDlbWogRnmY7bSdv55CKt3aQJo2KQvleBVgS
0IghF+QTFCtriRrT3y6Lok7mdFxewkeGqbPB++8b0eKQnG1zo8Hx5WE9FdTcF4dBFTlsbpqyZZKb
u0hY43XSMEOmoapjv76Yj06229dyKZKJVr0pW+TtBFgGCDBakD6qLFk9kOHL+clXPIgSoxq7RhZi
RgUHRSIbxbNd/XManGaWlCiuhzgani9jYKyn7ucNQ3kJ6/i3EjVsEApln7/3wcXSVqHj7ZNE+6+n
XuWYX/Sd+C4rPz/TEkd5lqRhJm09y2KHDFeea8/hDtxmh3HV7f4VaYI/znOwQu4/7rS58DyKUwWi
tdBGbkYqE4j4bId838KuxP4hx2OWO52rwomtYfduNE0vfYWbCGzb+T5iz1tCXVQv9bF82mzCR32W
WLZQ9CVhWNrIBsBYL3cZZs6NQMNJmswFbTIrDtxIOnoAmzJaHkMLkzxjaoVK8DtM3RK8ilxJ5BxD
KeNINbEjzsy57J1RfNE4bH6kVFHhzugMptjxY5PGq2RDzWkQTGOUkf3mXv4HcM2DBPtjG+735Mbl
bA+QfqbqOzB3c3hppKhN3ArY0pmkeZtz99Tvh2t526lvgv2NVJg4zJRgMPXByWoC30haSEcg40Ms
EGqxIT8ECLdRSOpqZ1wBs2lJ+wk/k1E0vnOveaZmlZWuzXaDIilWM3iLec32xZvLFDZVAqb1aCPg
rXQRZzW8a98oSUdNknlU7d6qPAmgQcSnoOKqHgJsKdIWv8+C+ruS9Cdyd3CAnJtp5SVKRRm57BRW
vCbRUxk9yGaPBYw2oREppJT3WYv4tCMhizGDQLazEIywkqc/J12/v91n8TkAajbUVlspY6wweuUv
Lmi1q7NPDHIvKq5Xkfz71qgNUiwwuXUYPhEWRtNjcrKD+xkG5izL0oPYczcNqZT2l1LZ7JGVuGkl
EWL3jVKpScOhnAsjG61FmOxbD8375ZuACEWbaR3MeuDHfyFZ8MBuW54zFU1Q3mJGHbenX6chywne
izRod03EaK5iMdmAb3rngjEIZZ2VXz1Y4Bd3Jum8CjY5/QJ1Bt1SE2G5EKMzeynjRx3nyUZUH7Gl
jhxWIz3wTDbALZ8IQXzBhbdRD6SoSNCSlgwfmaX45OBFZp0Xoje+KEQ2v+KoZ07fdKcrz3Ptwjp6
TWJ5Mo5d21PeouAF5kzd1GXl1GUX3Z4wxP98LpD5OFvDiN1qAyvgpccgb9TU1M8guu3gqTmy5GIV
54O41LGkU++Eb3a4Syh6vUguMYvF8kGv9Muj+OANGXrPjWDfVlUzYvRF1yLiLp8SPd2BdlTxAY9y
T6Sk0jlTZrzUpX5L6coVMLx5eC5LpP8ChV7o5Ry7eQ5awM7yxP5elzyDiqlfxdYhpn1gfDtvlS4E
TBxONN4eP02LS/lSW1ICh1EGVw9JUrPZWbUfFWp+0rDJWpIeumJvgYcoq5ncmJ71LOK1syPf/mT6
c1O97BVPziN5Z0HpAfT/1G9yrngrXR7/FjwqYHi/ZdMdnfx4O12F0qFGpCwAOiz97XoVgnVkW2xA
0renRdDuvdWSxipdBTELjFOsCkMSySOUCPMGs0LgQQeErJMuNKrWhjKNduqFVKlKUYgDJB/z6Y2Z
ZZQiSG4HtP8RgdaIyv0B81g8RHtrF4T9kBdLiMZcv1bBJ5kq9hi/uUhFMaAq4hvDyBxqsZo4swvG
3Mz4fcTJewj6kOdiLscbhBX7cFFF/HiHQkDQxiL97/FMgolSYrEqnVGk0lZDYIz14COvSkuHeyfA
B7253+6iNJ4FRpcZRig2GnlteW05Z9I5I2QNIaEGsWT58BFsZTfafJdx426oCN/iKll5t+tAjq4r
OSGhs9uTz51xuq2Dy/mm8SI52kJ9g9o1YhAvGJZ6VD5xFGgOkQR2w46ZHe0KOBqIKxTFMZSJZdg0
JQk306qDET28SVYqrWF5U/5I117XTmXQ9qGs+8OmiX0VATu8AJVlSeKHOqUlSfwwfWtjkwN5T1HN
9I8W4edTqgS0y6bjD0jhtkI028hUqumhPX7/AzqNMI76+NDUVeOHmWHsJEM+enAWoIFSG4sAZg9Z
gQOq9+xc0RqwK7h/nieh+jwilidvEw1uYr2BfVVA8rXQ/Mm57aKXKdmdl7j0IvYSXo4K2+CHILDm
+XdQj1DtrAt+eAefwddBIyF6aKp5YgxVyYREViBHvu/0iGk8C3bDGRRuvo2sFhJZfU1Vw+aIASC6
832sDLD1i8++NEnTtK0MvZl4X5Lek1P1dJh4zuBPs7JGVgGq4OKuWpHcRw6i/8rOp1YUUD1M7QEg
+NB9L5JfpAXCuf9XTU9lnyQrEjis+ZUNPkW2E9izYakkby1FaXe6e7rCH62p8xVQzlmfCEqu4QRG
RQi9Vssxszqps37aUUrCuQeRzOL2ll1syHfdk2KfsT1J0ZPK42YqQ5NR3HmfrKIFOK+K4Sh9uTZY
XD8oxbirNmsMklNNToTWxSLMcgsHep9bhse0UHd/J9nrCWnRkw4kGgx6GA+mWxIVjjTMmqsuvw1x
FJvxzqNTlBZFHjoMFqMNg7GpyADhJNU+0DRsisAetaSvcB6eRwhaJp/mQpdpDX4ZYtFPfahlYNH1
0Y1z3Rbosr/6B5dKpzgLOf9NyDGf4O9tJfUws0p1Ofjg3ugCjCYf69lzY2c1L9NEarhZURRdZzG1
aGxm/Zj7E/JGGD9xZHlJOW0eKV1RjRryGp7pH/D52JZV94uiv2P1Lvfc/Q5xz5G0uy6ouXT3Diob
+7U9fOlmxCdsWM7pKJBNqjOjvwY8fbpQqu0FCEpMN2k1agzQrHtRA5rPy00jcQ/GWu5WaLJLb2Vw
VznXqx+pCYmxyAeeEln3fKlMWgMUzANFZ/X7mpcdkH0+w6VsXV/CJP4L4asQU7u9fRK5EbL5NbKE
qkt82auo0nb9ItynR9Q6RKV5ZVWGvRqTyx3tGc/zxg6jBcRdYzf3yqsX6eF8Y8ma9z5+6PrlDXMt
kS55+z6HuTlTgttl2NxzJCpohoxbFcFR2n2stHdR1cusPjC3GHkvUki7NUW7Xw/0Fwjiq8frhF80
wkiXOjcN1BSd13R4N5EMM+QV4GxNVsX/kpdR33x6E2cPvkoAkI5X+WuGl94vqm8xoYkUU2gvFj3i
NZ0cGmGQdduIG1uqTTojhTA5tCY5L1PUrb1ZEfZbE2QYo/RGZAszLIumdc0BhVKXHnDfOJtgMZRN
h6jni2y/Y9unbowv5quFcRVKMuSAL/k/e5ni6AiDlI2isqPXXLzcGiJnRsmxihhG5YkTGR/3/lOg
bDgehgpZWLAklHKPON8aA6WzFV+bb7a3qBjR6LuQqVYyDxvEUzJ9WLixXxTFmctqQ2FDeMSWx5cv
czbLv+UXy/tyVI/yvL011ZbBc/xZvH+0MhgTN85z2ABCsWumA/iCLCunITdD5LWqpN6LIDFRo5z5
Ia+SE7cBYx51KBO+XnPY0q3XhSB6VI5HZXrjj9qo3rFDhfy9ZtG6Q6I301JYbsWCYRWd8QP1DxoT
omg3lzqqNZxC9yN4wJa6PrvKqgrvbNf06cBO8InrlIzYBNFIajGUZCBtOsaPbLgz/AtdOup+SUro
ly393jMEZjkf6d7iGrQIrIq9OCbypjMHJF0HOq8eaHOAU2O/1FL03Gi0O7PEADCrQLOPluud3u9D
hGT4TV6LJdUwx7e0/ZR0KLjeYNlVgLxts17UebcaFt+GaQb9J92l81pbDCNCua0Oe2W34ACfcM+f
vpCh2RgPkKhhPq8zb+vHIK6bEJC05/WFdnx/7PBYvqQkyfEA3TxW53nofGPQPxYXXJkX2hZiy5mI
yVsLCZY0x58nuwhXa3Q79lteEzYxwtMfDAYiSWgV7k19oA15Qhc2jtW5ANW/WHKjM+hilh+MNQhC
6BiCUoq4EpHaVq124Z+K0/kHew0sRPoVIJ4cRUInBEfUdUKL8VTMxR+A4T/MxhZAS5jkkHNZdflr
tC5OfgJ7EvsPOObNfA01mXYZ6olgR9FM120wCSMb9gS9FB6s1LvLP4P9OkClAPab/6/kX0W+eiOQ
IKoBk+rksXCM50bkbw+YyT/v0jERTRk18SX4pKemJomhNCmijbAujtMhOeqExz6emvt/N/858nwO
UAwDWVZYKkM0Gu7cTDBkRVAjqH3OxDiQg0UKfPHXJ4QagxWWseHpYuT7Ww8elV4FegIbWoqle3ir
umpTWEsavCMAyNOq31gFFBq2VLMchUnjdpJSAAelNr5C3tCkAUPR4OOZBffoQKtdRGwpPrsRSiyz
4N1wQvRRduOCpOXhThwKVeaanXKVyg0FG+BiMKYAvGe03ZLQ00xdE1qRtkWseZ7uHeXH6nx2x2KV
Btfn/+GUeuExwDNXq9FsCutD3KS1xYIkRyJ7COT8yeXqu/DgzNWk0w6hZr7vqHz5joBHQkdsMFXS
nV68ZRxy3BYXLChLtQagfCpfZvWPtlKmuWUMHXjZ2083Ia2mjRRRxwjTVJ3j5rYpVQ+OSNVbub2d
C6z9o+hezBFS5bRM14FyiUnLL5Sb7D+X6AOq6A4ugVHsBCS6u4DZRHs65xov7s7BOdNkLm4yWf+k
7zcy5ThLTBLd7PzEAmpsGITa5HEqmQ6usBG9vRdA59MoLythRkwdusTre2WOVM2turpwYw4X49No
1T4B5a2tUoSlxEnwrFPsG8ipRD8l4Ag5QWt3LMyBbiXH71muiqNEUmoSfTWButyN0GYoIQ1wOXln
btL25uWRHHBwO1keeVmcIp+D+QVZxquDETITg+Y3tMKzYqehmRRm22LefoPoxNWqMhBMTj0LPohE
V+nOCS+xl/jIKemTHMhKn6U3j8LuAnk5MDZDic6R7YIE8npAI4zXjgvyw/GuPYzjR/O3CmxpEHVO
0jnwiqUdNLLvy6wagJxc6MJ4Euk9vCLtqwcaA4cB0dfDZ82XOMX6mSmZBPD+Uxgv61wOrJfYWVpP
+yfHtfJ7g9xPtIt8gtY+UmK8QuHha/M3DYl4YGMfBBYUn2nYKJeathq6D2gFfGrzvIlLTkH4rqPK
muATUsjpG7cK++dgSaVdcYwEt3LHYe1N/DxXst3wMRImlt0I0XH7fdo38Ov3BG4eo+Tva1kV3Bzw
qtedb1NxBPoMeJQaNKwPoGQGicogNGZRsnXLhoGZfPMnZomJJcpzBWfdu9q2YiZBlCJQpgMCsC6S
KxT0TrNA6+WqRD0tST3Eu1mcvzxbWgLNzmGzhIvLy0b1a9m7worht7Kc029i7zgk7yjiXiPmtdcl
SFqIjnP/EIa0sbcejBKvrQ4QIpnf87+NQdRiSkDBMBydy++gA8IFhxDOn+Ay808YZVCNnCGA4Il7
iSboZR4WqhjvYXwXLqw8nDKj7h/n1dqkbKfZxQghaPCxSZsb1DS16NjzZUZM3k6ZIoNgF+fgQ5ZA
m2HX0vGN7Ao7i+BpjKcXm+vuUm6yS0AhM6vLy8LUAngb/E+TP5xDptp2cg6pxU+cZjgrYJYITVU9
MyLHqBYBhj5M34tSOXVFHpwjy9zCEadYKpnMopOuiXQrQLmGiYRIW5kflExY0kPccQou6OblRyb6
9CQxbVwKrRa+BBJceBOtucND5We7qRTGufV5+Ih3rOEoSra2usPRlOxp73l2QP9iWb8gC5T0Zk6O
bUw5oxPpd5NXqMdZNKdZO32ZERyKjd3rZTs5oi3cc327e1/xfENYJ+Ql9HwplcOy5y6tJlufF4JU
cc5eqnjwSi9v9obhVFfb3JTNvETQjagrRuJbm6slE8zmHL31cYpdkC1wIFh/YMWjLplx3IjtQuov
hgKgYFxJjFBolQA72WXZ4OrD2Grb6/t52XtFglje49WYGqnfMEPaJNZ8yCIdUHa6iG1CRzMYK5L3
jEGspT6/Xd5dKIcS5PJgUsc3KNUDDjn3cFiAY+49T2wnECxoJJGVenqtoC3sA/DwT2NTH/X7trR1
+nI1nPbjkVr1mH6TWOZxzFp9vdyEzGBxRuxuDMt7v1MRCSfIM2aQGOzTa19EJgQFzzTwVkf/YsQr
RRS5nw5esTXGKhCV/4PLj+ZcDIrvm4IdhZcwBQ9D3CbASyygIwBASK+07Ez2ktawlyU6JwZWzJ9W
kAL/y728p7PDkAAuTq7tKmnU2OJug3busdVrXtgyaqsq09fiqWytkUvTU5dqeoSfRhhg2aMdNpOr
GF3Tt4eIKiCOWRwxfOsPfqdUw8oZ0f8+tU5R/ax1RQXe7oHdA0oiEyCgkGhmlZQMHPZ3TNmDgOGp
ziUr/ZqYluuxrVqXfQCvSyA5YztBWPrmBsI6TfVPdXkMQak1USFaGjwGWCovm1XWShcQIkTkICc2
/Q+i7ozbkXOdBgcXS+3lPsGs31cAWVwpPg3SHeZibY5QI8qpQgxc0iWZbT4Jist8njGyQPcdvzp3
OMZWvtVToCmjEVrTQy6Runc59g+GHPOU8HS2qcBDvpldVipbDCp5QsSa/0nZfTRFjh9aPN+EXZlP
C6IEulEn8WUXw41NJ6vSpYAH0bpGijXQj3OG4WVOemqUAY2Sw/PmCH35fNXyeWT4UHeP1v9f0H9j
j1OrzqJgS8epy5gy/9wY4HJmVs0HpGuahfpYnmgKcg5u+B+RjlkdiJACJwNH2ejO+boILTA+MWHc
IONyDBGsX2OgOdX+wMRHlvAtoMmhvECfREg11rGH4k6vA7EFIZd8EaXqL35jpGpWogEPhvc1Atn4
fsvg/SOCAZhhc4YbeKtujFunMlESevxBSqC7saXW/lvSudzYl/s5GBKDU0Z+vRqa3fYnLrP0M3Ce
c8i5v93SdrJUDOSJzfWkYp22FAhQW8jZyaNfaSLoA7RFEK8wfMyj6EVUxUADSLVMlG71o07Ho0CB
NA3V+hWpUBvk8XEJ19vSGFiFh98+r4RMZ1vSw5i78hejT7TPsOaHXES6J1vIXORBKQDXDh9OoxP/
J0cXqVfodtqVN7ona3g/3KP+DQj/BRrlA8cZ2crFRsFNmf8b9V+c2+fTlXCtyamzgUJv3q+tOhWI
ZjyabNOhHtSbIyBvujkQ22xgwTbwryVy5qne6Iv09Qotc+Y1Koh6jEc/t66ptT0kn88iShSV3UkF
xjdwo+Pa5YOlvi634LpdpBsIGztQ7etOBoYthjWpBuODIBbfQO9zco1mWMlFSRy/ZCD6u2VmUkr5
2muhO7NBP1wwXrm7ZoSuAUTXPzuRh8k93AXrOTlqmrsMH19QhFW7+vxmscDU6F/8YbEyggfnLh6o
EJOmMYWxpCwMqQrwmAf6VHU8hsm3BiRSAun1FdJwPl1SdlbkZp1kD9T0Yp2y4Iu8JejiZtLwOE7R
YmDDHkkr+btqeqexCdPR6Mx43DA9szr+HYwUmo9sLbUMTwTVBh0LViFOUdcArl/S833sQN/cQUpa
cw9nDcjtQnslIHGTucdjl2+bx1TP1scwJWGhuwNrRbt8cXRxti8tnADZq+qUoUGqqjvWzI7nbvHC
2z8wnepSUIG/mwvoVo27WyE9e5Xf1XntzSxM1/TcJArVfPSLqnsmGF24CriAW8YhCdwWcFZJzl93
ulq9TKg1nUtEqO0Atbyb6nGpW5CI8MaO1pJISfcPobQBKSDhHlrnJG1/yRzk8FTeMJgTjO4MQx7q
UmWMIWpBXpq4BDmsh9q33Hlc/mUQ/rmAhC8dq6SyQZqSWefHdY1Ha1muAikyzc/n6CpN2Jc9iuce
u9mM3z3u5jMmkXK8cIPsdjIDBlYh+ckJG3RrDpkfjZl1mDPRclt5e2aI9iP/73KD7KCC+Um8n+sL
3mFd3nAJciuVKvDAJQfTdulphRtQqRxjamw62UkV0PA7DjqRH2d3nEo7sOgWQ6Nl14s32qNU7ooS
2388LU9C2bEw6J50FbRCRwvhk9tiN5VYHtnWRd7wjjl9eNsLD/M+XNSI7P2M4bZNZKl7kjY8Qa98
4QG+Lxl1/o7QyQMzyHLf8jgSHZ+MmyHpUqlKN55LqGiS6M+41XmSzYMhW4H7j/EjwAn6JLJp7X4V
FXeac7PE9pvyEF8PKP9kL7yhvaU82PWiRbjesGR9ivFjkKEjRgrQ4WoOp43Em2ajVKF7rxMlzyaC
JUH+A404ZMmP4LuKTn/P08CjfH44//NYiG1nNpixyZX/j8/BON0HIkcYS1IgwPASdoG+f2585Zs8
I2bi2TTxiUd4I9Ir3QwNH7JGYdFtLeq0IxRh02gtW0KRBPJw6y6Q+4vwz1U6tAoCFCDKOLU1euOF
cCK39fPTU26X6qyLbFKYnK/BMl4yziq+I2mw4W5dDPYpjyI+TB0dF4mI48RyajkkuZQzEzy1FysY
xcMDOJM9yQVkaRNxEWTLDUsmKMToxfmjn9TNquvyFAa5dvkKWNhYlyK0S7MLVDm2BBjOxkjbKOXV
CQ/XYNTaQTsEz4NnW4nvnxP4GjtazShgM/RV4Uqjx8DonqTLgBPTDARqdxG0fGrVQ9BrG1OoRQzR
P0/oqcMJjD3k6efKgI4hFsdA7vgLMjPGOurT/vOgkVGS2zYxttStJcqjL4E5ThhPFnYoZslCvY5Q
ZoECT4hFQ4yzj27F9iECV/RdhmHbsSJJNu743Yq/RCAsNyN/1WlHQ6EfXJiJB6k5K5+7zwV/eqif
t4eXfxaHP5En+eDbX+Su7gGNdeB7mPdvfurcP62DaLYuO/MI7USLsnpTAo+P0ZpX2jTox5wFyr+d
/GYsfuGZZgvMmnXCuTP9lj70ci6XED0VFUOD55UVRfJtUCUZZzYUI2IRQpZjgdpa4K4YNJ8EHoBZ
2pWwwdQ6bsgiMaoFdMSkPzmBGZfcKtlX9xwNPoefSZP88Q+pHJPeeJKa9KD3BKQKsl31CAvo0sSl
4YJ6mnDjAZrYpxcicnynfoFN29JqVZxjTD1KPtEQTuzoECWJUIrKFUpvJLOhRUJ0iEdgTFjVfqJb
cQ60Tb/B8oE0sbi7wWCWynnDRD6MXaTLoOgLY4xoHOjie6oGAujCgFLU5ntAxttyWTBZWLf4e7Pw
U7tCErGxgWk9LMcHv1ptGRLithNL9es5O3GfPe/zbeYWLIuJctcj6OKPhAH5yQ38k6f+QEnh45c+
azwKwNcHVp9Qa75kYh6c1bxjxbTqBeAKouP5eXLHNme+lq+ndmhV5rPViZK+dqDTnpfaN5ZMt/2o
rEHTKdAzOySdBrke0Cnh81udvOy0SNrmnLkXXKmwAHtXE5Z3ABZYblA9DazLJTvI9qiepoMSB1Z7
PbfhD8DHcFa+Wwirj1ioHcxYAKa6Gsh9myfOt8nkOnnuWCbSAPyi3Z058gAUzuT2S19bjR/ghwMC
a/p4NvGARlt8/LGV7N2o4ufFMqDM7wVkZKnkXXXjszxCmAMXUQwgTOxaekvrPwQ2Vf8P+mvtTcFn
JSPy/NczUSYaR4LDRrDuo4RY/Wd4Nwxh3v77XxPAj1LVUGhOsblfmsyETTno5VEA2rkr2Loc9p2N
FiOm96TC4x72W0zAzDrpGk8mIwaMsUrikvdQLcr0sg0cXR/ET9myB7L7k0MwIy/oDmSmIFj7O1+d
AVOmONUsU+dVXPUJG4KbKUhVCUJbCocGYflsHaEnfCmaarZGKNIi+9vMSNiXy8J+algb6mMBxWC3
VQ25g5v7CKj7z5HRvrH8QlddKqMWOSKavMDQshZZNfamjkEUru0UHGT5CuHfxLyxImi/OPd4hYB+
CFPNz+3IXz9wD8HZ7Im2YddGwcqYEgUbaiz5AOgdjtQSq4TeCGLmU30Bo5xulOnOv91ZEejz2qTW
EtqqkMlHnwg7wybsvKz++8T6XSO9hNopzjLT3JfoyPJjvWuJOJaFTl9w31L+aKa2r3yEoN3GVSoP
68aXuOj+Erv/eh519JA4Ahn1qyO44nRtJpyrhiPNd3vgXPHwrNFoBKK14Q8MVWckbWghggjTnyBM
H854Kdqlh4lRpNPXYt69fckunhNdyk9DeTntdkYprA5nndT6zh3AeRKUEL5rOdqSmlQVCl7sysAA
ip18Gm/jk7k4xNI3qpS32ufF0t3/abedr5J3r7yiAgzCHaC27hWfOiF24q+7njHjfdcH5M34C831
ttVsEkM0jngRYOXyR99fRNzauICoJ+OMP+0YhO6cZMREkiGYLHBdaBIQVh0Hp3uXFQNPeXODu0Eu
qU01TBjR1t7IICYixVHqQ/yc/527cIF5UNK19NrD9ElUFmS5tKGcmmcu22i6mFdLCCAAVkbEXO9M
tr7ixZoTMvPeLf4RMqNWSZMr3AeObPJkjW6JjhyN9lUtuK9dd5CU2CYHt04OuZhjmYGR4LBYX6Q0
mQX/fa5JslChm+MY0SUXQiN+hsIhEuSzi2qyLjEiY6jfgI8//OSPFRRZiq26h6FTnVh/tvhNS53+
BEcTedFTxC3iaRzyqGlEdOTCwmZQexJTpZ6VV8WhA2DOVHSyo/roZCJIEVGIYwu5ztF64LDVZa6j
+S/0gR8pgL20JDcTC7V+NlSTdGxq0NhYdPrRwn5SB4WVZ7ZM/RQ73PHYwSXLthNVtRrjuoSessY5
1Cf9/cMhzaMRntLT3ngsBBdti03uWMAba1RKOJFV2HbHkMwr97pE3U3U+1izyXyrKjypSVb44VH0
wIsVvFdskpZN76K092uVBVzswwRxI5Om4f9zvjFB+4zCixSVp6toIuHAdhHiW1ft2B6sSxB9sS24
UTZItI2gkbi835h1asb3u7nQuuAQScg03KM+wY4J22VH4osNHkQtpPb/CSzsrwEoT97k2l6HZAQP
pkYqiqEM7o2qB5n0C6sblO/QFNvPNbpSK6SF/X/dx+phzJ0r8ZigSzGjRN4HMYhLorRAnZB9qvav
VT3nX/DQFybmVQkUiKiPSodSJPQmVo9TG8PZrTWJk/7foQqedLuOvu56Ncza4YEZqHnyq4LDcrRE
FQXpxEk1zeI4t6uAKoASukKW0ERo+L/vJOgiTDBvPUUcu47koc8BbCXLMxNY66d3UtLiUWFuxSMT
tIIp63HW7PX8s5/QOFCN8R6Knc/o9ZCLmHaWucsFUTtuM8OZRmiHu2TD6J4ZpF4X+3zaoTqlKsQX
1RgAB8emb/lQSqWNru+oKyn5QBnbjNZi6ahMXo71wIDZIukbjw2j9R3MBX1ekiH9WC9n7TqIvRLm
KHH45h03rlgi7nx/QlAh8djY3Hi0nl2fiOs8u6IzxnDbRaavzUIRYRT2GwhnZNyyW+hwy6R8rr2E
ZV1aAZAygtSa6tIZxWQAyqy2y3cQFx08LpixTXC7kWigdYNfGU7Ht9NuoG6GahmoE3ou5PbPKwj2
Aom/UdlOPHgN4l9eVD1KWzxu19z89acmNVBeJz4xMBDb+eDLysGPdJLc0FWS/O5qA4Mt8fpYHht/
FTzwfGqZUUvCSEhjKqS0i3sdNNNC6OuouKHrFs4MDElWlcCmUq8Bm3e1RWkTrqzrvWGfNhrn+NJ3
+Phc9sWjHaLZpo6NhAf6MOG7EW1ht/OQRSLgsODD8epk3JcYxrFXhNPiaaaYZlgi8my3MXEOxli2
Pbxk90whPIjPbgyxNWV1FANXw5ckVB96kMp9tTZe9eThDxYc/GzQJ6A9DfvEcB8slFm1/h+Q/zlx
ri6xasXZgCwKtq9fFAAAbk+t2DJvq++/mXzAr8Ch3gFI79+Jvw2saYj/ADotlHmCEQTMkkZPYPP8
mGjs56Sr8bCDgYl3ClVQjXql1Ry7EwAkgqsu9weUKtTQXV8KgAa0g/7K7D9YKBmV+s82zwcK0EnK
88sKpX4607yII15EKCsZeMtbUmsYOFbGIE5OY7CUx3tfUEa8Z4nnG8UYnhgduddIFOTuYFcrvkiH
ZUqUvjCYOk6WMcZasQIgWH1LLe6rBUF/U+g1s1aFKg0kZn9JvjZpMUS8Rfg/uiHH5iRVR1kuJw9S
mzVSDpEq5sGZHJp05a/CxAvK6xBZhe7nWWCzrD4jCTMYYYQ3YMB0UVVUW21HSj3hx+cpd5hadZ17
mCjID0Pm28+zOtLwaRAE8v0xfeDzMMsQW6WVWtnNZdwkYdRirKs+va4/7tDsG8fdDlXLjDEF9ECb
e89usZW6XZC8Up9xUkUPK3SO+2e3auRIOyX+tmuUXiejkSTqaXpyyIHB4cKckQw96UNSkz1ysjVD
y+NVuGLP8k6x9PC5Uk0TnzEOg9cxYTGLCSAuAX0/gId09GDUeGLVWE8laH4blhHy23IDRvhKBaC1
1x/2i7RIr3wEJQibLQKhWVjuEbE52wV2i0I+17mjpmcLGLHauvCUqRqbqLS2MGWkr6IcvYR/C287
hs09byqM2k0/JrcvNaHGEmjokuqS/S6qzr+2tcm565E5t9+b17WXnc1Cl+JydwW93wxdgaQgPRdQ
t9AtPhK5w4WL2II5OrHDB0yknsKaOKiLAe7wrb1VyPmuiUoc3vkSMbO6ucvQICvPdQagoWY6s2i4
+NjS9on0ye/kYGJGeJS+lbYf81+1AeuldAlea+kz837FFZmpiKTZQIIdhTTbvuHmImej64W3sGs3
LlYIB2rW4fPgy5p+Z9BtozURTziSL1HAyg2XLvjZ4wOTwcZrXDNwvfeHRN93WulI0pHYGWOaz1Xq
HQ8JEWjycdYEklm/Dn3iwnrIqlQgfAPc1bODx3r8Ya8vx3G89eEjUjP7UHTcYhdLhouwKabH5dPm
Fj0e1SX3dJ5d9AhlriTEzv9DnVcE0zXdavVVJEdDVVvfQnUvhv5oGckVv3amN0fgCSGfFJZu5N4I
09Ip7qL3tAKeMXQeL3SywuTJBZdA7CmYhYz6XuuEsTeinEMoGbCmnxi8216NA4D6Tj/413WfjeGX
Q5WXY5NUx9PIZZikLR+0uOOFg4PYUseGPjMLlD6tTOwfUuTzcasxYhieJxeyTMBRWlhSF4z/tQK5
gcj9P/kZT26kU2fEBj/9Dx+Y+aHfcc6SNJb7W64lTtMbfpWoq8bb/YEdFbnfyqvIyeJ71s1xbfQp
Qq/d71RbtC8mDl1K30lYOStiNdl16yxaJ3CpMdWBAxTuGojfwuYE879BqlcSL9E8cpsAFKFXYKOF
5MaBrcNQSmhpENwCMOIeW/SSXJuf9vzXtd0Vg6I48NLeFGzwqoXaHZ96Uv7+t2Yj17vZgysNXsxn
79AZ0bmoIYrkx5htwkQIxB35V08ZYIKoLNl0j6VbaoVlDhs5Dw3C816MtKZ4aLxsR91r2tjeXtYJ
8jU/rdg1XejGKYmWlSpLgq9uVvHJPfmUBzj41VjohGd9eJAHfixL6Lw2he+RZi0TXbXGOCg6CxY4
hI7Sn3tlZMmQPAdMZal+9DHLfOUMQUb/UUkVrgO4eQ5Qe38L+WSt3I5nk0p0h/BJfurv9pHi5nsQ
fOYv4tEGCuzB1O8aVkg45eECG90J3eF0Q4chxa0elgNjgGVTwVgZIGA6CZmWb5mZ0eAKO2nUoqkW
N/cgtGtxJ3IW/DcBIIw95SmDFQGwJmnTA9lrHVfbLCwN/gi3/p5X+nqXRzB7orp/m5NA05olZ3pr
t8AaSwwnYhH6FUSMAD3DiORmUDd4spRTwX/nZq8+MlH94guCKMdWShUeXIMIKZKktebkmJjfgHTi
qyVmyMNmOF8IjSRXJC4SuKIPSxAupD5uYpnG+0EpIVpdKWvbqdj3Lx1E7DMm9G4tLIW2INwQC+wO
JNi0SYv3IRYFFbzqoOaHvYwJ1Jh20/mOnzde3xgk5TEzYVK7rG9UeOpC6Uyfs0/1EmAM+VhBdAeU
3sNdRTY41Q2jexfZ8vl99GGcn0hLDYGn8xXcLrfqpQ3PuVM9lZEqpJ7XuPUQ2dIcFSsX5AwjhPNi
VzCA78duWDqILk9Wgqbkr71ux9NO/6cMEDswNQs6HD9DAattaxnHM07rZfIIhResEA9zNRXBom0u
tm30Uq3UBhF6eiwvSRq1kvr567N1hdojzM9xazCzUB9UQXhIP24hgWRkGvJJQXRQ4qqDwPnlP+H+
vZ8u1HiKSWU1hAcl75pf1QScXg2xYPFsFYZcCeexGFPIb4mEshh/E01E8ngBMnglYiu08+dK/1Au
rHkrS6N3rRTaz03RYtNJtIP0bN+1t5NyIef+dJC05tGsV1aNZTSrGzN8TY5ret1wFFJQdKMoUwAE
V+twcbDu9ALP7gRz9Gdq+evyzlr6aHdUxD6e71YPPRGxiY0cXXgf6djhXWO/uCCTgBcGIEazh51t
LjYfqa0uF98ESIGsYIIXZdG9kkgIjfL5bB7xNyHJK5GtiOs5n5j4qdeEi/ibzpQ4mAYU5+4vnJbt
8UPRGhEjEBq/l18upek1fSWczCci+bX/e1S4V5uElSDfISozwedAC1/KQM4KO2aZk6kLFfERExwr
1vyh+7IOtYYsqcJ0ysccxvjhUfUPmR/ADcefDjbJsPNDdEjna3wCZqDbQg4dquyfj6Rz4b2SDJ2C
eTbfJJuyAodNVBG+YNJCuQIL44es4dbIwsgpqFgdqSHZtqB3xwK3P5+r8Lk485rkCrmnOCIx7lJO
DSLBOsNZycBYgL7Plskz92hxxOO06wyIHF9yAqb7Aks4PPS5W3JB4kcJg5FIHkAT5B4y1X42EHR9
KP/X8j0n7OWiBgQZnk79yL0IpGphjPELW3Otf7ZTzn59gznjqmEIorZwlXOC62YFdjSbn7zmK6oc
0MHGp4uaszpv6l6uKCzBKdxZ8qyEAB1WqNpAt4pIdkHXh5xX8xxT+8L9bvOwRMeZmEktomep5Inh
8/dMiEum0yFtP6aq3xCefzVFR3G3fucFCtlH1lMyhMkbSeXcGnZ+VY7TS+IPxQMk5+y+FWbUiZ3z
u6LZL9YWu2bnukoaCtOTuWSY2zKkRX1+/6/CYb3yNYwcBhEM8AfIcMaB2ErvZFHYbsGVRS2n+ufJ
3A6+K8tBL+DG3CIIhKgyNOT3GOfkxn0eaWiLrKEK2dRJCmR8qkkwppPSJOcNiZT2gzWOo6fh7cOy
6/60ms4sTMdhfbv1HX1kx+4ypgOPniNitvOcILzBnmTfYUCXMUpkKh4RaWauMa8zQSh3HYXwBVU2
/JQ/ZdESiWbDxe9XBpzhKlxlxWSlIp0VncvC59eK5QW4QJSS8kLzzeOLw/0ANZCR9HgCIhtWhRlk
ilQpHuhCs7NKoyNyBBu3hpnGwntvw4f0RJvVyKHXKseHWofE1XC4+E0W/hCPmnG9mW/Ist9YwJ3i
zH9uP+xk1Jkos0KMA1SeOPIRgASMthnrSPV6ktglkdWM1FsiCugqLByghiBldICdNK4OzMhUjhnC
nQdMFMiTQCuR3zFqG+N4v4LXWNcW07fIuJIDRZ32zkdG+Tz2Bbyk+7BtPLhMtwmmK8QlNRZmVmBP
MRg43ZIyt3GIWggRrZ6TwjHetxDXOqrbq060evBjXFNQP6x7HOo04S37XyvfedXmwkU3IrY5b0Kd
e2E47FLGVery6DlKPqWGzzKsNbWWk0Ja0hEGF8PfvP3btvDJbKOQo9z3fROmnMcWFMJpz8QzqwhZ
8pjf+X/HNs6T5jqJhNCJm5jUpGQkj+xnWadbLg5BTTHolgy/6iGNFG1Lj8u/tN3gQaiDFHwE6+Gn
cEwhr0tK2QGLh4QvFknkOvn2gTc14h7GxrZTAo1I8IfAoJDM9lggTN4lc7p+zUKybxcCM9lcsAFQ
JwCNMoL0ZcPC8VbDdIrfdaNGsqynK7FzfqBBKMO1QggIJ9H6u601ROEUAc2luweq3VVHrGAMtVNW
WqDx5+p/0DD9Y5T6YzMuwP6hOYyfUWp9L8oGD9fSydCPUDSYzbpOjkFvwi5oKjOD/3YMI/CC1RhQ
/72Safjn5dUbPTywdl7u0Kc7lRHCwXLgkGC+kGS9UgJGTdsZHkj0MPavecbNns6704f7qKcYM/PP
fXpwMMetklPmgsaFmq3pjQDqC+rwb7ybL97MM3L0/lCHmYMNWz/lJUPJUPEalUbE9AAfdehuWJla
SjW/uDCAnHde64o3yX73Il1upK8P2mpQvJKNORtBe2s3MFmLgMHSjzryCeZdByEC7acFQ2crPLSq
fH0TnDUabr3ZOl5myOjT/Gu0hXGQzI2SMNSZTUQRjBIxiHvcwLftY5/AI4ldHD+wxpWAJA1+/jql
LpeVszxgwgPo4RN36tTFRU3Lh34GG+Y6CTklVvNlvdpQKcQ57crZIAF+Cl/UKuJmb23yUkZ4p42o
lZ0zqQEiCSsJMW3zPEa7rE9PV8KzFRF1cUNlOs7HigiuC3Nt0ccb+vGsyGqnRUysGz7dOz9219O/
oHB6421ThgFEyLct6Ol96r98d3SFUkYgTY24zWbMBYjteKEzKlPkxXSMtg/Ds5bfE9kwAjmVg1MJ
3iFbSIrzXrdXrKPgo+dwWAEPDNtOwtHEw/quldf/mRYrBiSNXJCmEXCO7DSh1uIldltUkmPRgHSU
2TmQDzF6JNCemIcadEyuRLnv7wizO2IDkw9YAMA4/TG2DwmfEIVkClrqSmAxj9nOq10fSC7W72Qw
H1yUBt0Sv6NqfP2RyJ8+mLgCOgtnz1j3OOxAPCVII/5xQB5EwKEul2hIH8heBfFmc9+3pUJygcC+
6DQeXkPbs4h1/zGpbFVS99vNj1nuPWhnvOfgumleL2++ZxjW+lSNxQCiNHHwDJ048YPNGMo7rHwO
AuaejeOlEzDELj9rdqHAnJNU1gVD4Rjq0fS7u0LUkL80Vx0GZ0NkCZElarg99d9Lz+KMA45FWSkI
XlVYTjXHrHfRtfbqvwI3hQTKf2biXWPuoyy5N3KRgBENxr9Wz2ZQ2DJrNdY9L+9ahk1fRszZjDgR
5AY0i+VzwR9pvSEFH2odnvP8EWDjSSUv/p8KZ7Wb4HSwpW0D9ganpIUvuBdVGqGOGySO6KvPsdmY
TBKPnc+EgMLpeFcDM2fKbcwvsLP/YgX5E4iYk+hr+Xms2XTrGKFnrG0MQjNJwpQ5DqrzMzi86vFg
S1TmhmA79+iVHS6G59CD7h4pTcOHvVUpVh0sMREIAUxYAh+VdLfhcEZOgGlolP9D3V5Kh9r/TjOB
uOsHbTYpg1cRWJiPWPd4ZwhSq6H7Qsir+GHA6D0QzH8afQaV392fK6UuUqwvYxLmaBB55DEg+FNc
2a/HGpbPsUGnnGQkBi8mUw9se0J2rv/P2HRpBC1368cZ6u2Y/i0GoWp+sVFOQ1Wp0aNW21UQmktB
coq07MoxF+emGsbW4sjm9XZqmA8no4LKRpsS9OwmFhSWLtiv9ytucqkwRmYcBtzgXYhxxApoNRjV
iiX3PnoRdFy40FIbCLobAXuYFUzIVZycLeeLdoqsv6n8l+429jIVihGCp5N5n9xcZFbGOjKpQkBy
KFendQBQT1JcQsut51BOfZK6ibPD8ibw1B44TsE2t/XtYEpO8BWKGTGOj1lU3H0wgP6A6plz995e
d3stv+AnS8FK69JZPekf+iVVOcReUq00WUSqKeQPuxLEkY4Yi876DrTtoaz0KXx9Gld1VWLQmwdA
+sh3ZOGkxSTWYMrDNQZrL+m/ruRKGXIwwqF2+/2wZ7XnavCsaBpZBJEJcXB9elQgc2MNf/EFQW+Y
CZtkS1jzdzZ3O+kLlHiFO9c/3bjtSztrRnkKVV12FRMlceyv2A1plqIr+z9DDX5RuZ+bfre7OGrC
FzLDLcIjvLvdtRu8lU2NwgWeGb4tjGTjElM4ak7jspN6zK5qb+gECwP4XvBte9vdkDP0H4MIBZh8
miIx6XOqI27nzglJrlGJfraDeFlijLJrTh80HP4ckbtXzstLrigWnPe44jEdTMslTnRPaIzKTiCX
JMUoJqs1zJBAXF9gLpzunT0HQKRGHNE2q3AujheknAc7SJtv7aryw7/0cMxngNx9cfwInwXaOoRr
gkJf1r2dPwvK1vbNqhagRfqDCaJzHf3rRatf4UTQFOPGw/cQh22iqGaeTgNAikl5yjz4nz9wlBRo
ebX3sSjeHu/fMTSTDPH0vGR1Yu1QkogZ2xrmZSr8I4mvI5JkanmR5WFXIPvcStdRdQbHe8/qe+L7
AgDLXeDTsAEd8NTzM0mCheKnt/cWgyyiKHa3MoKaeHtjkSGZrfhoTmL9Bbjq5xrKjZa7J5qeO5rR
0qhWqeAzweqtvsDTzXRvzecy2AHyk4EAjl9l0qXglYcN7Vt8NiYleBANsG+eNY1/oAatSGw86M/U
eezuExz286Q+UDwnGsMJiQLdpxSNM9wP/mi96oSjb/hDS+92v9iUsOosy95a1dk8LqARdDAdvfsz
L6cdNbOBNsyZGtOXbBiBrycCNw6nuIp2kOauDMaYww3w/r8nPT8Bf0d2caQXhby9l9Sal2QeayV/
A61qYzI35SJvCDbwjDu649juSQD6RnXauwSPFsNlzOb0bDhk6y/WscJRGtwgQfkLrFeiPwv67mDs
JfdnOrS787b4Xef9npf2GL719l8qaZoFOD8VfnSXWXXxhJcGs6zIPRDoyQU5g3Zg0Y9h07GfvcqM
Kh4UbJk4hnct1+ttkaFsmL7MaxvdrdhRcxIpi4Q+H4vWbBpyTOCzwVW5jaKYxArU50zfxOqe8l0x
Hp4pkLgk5ghezuVScZCOzh11Tz72cD1i+Xawmex2BZ3ahNJO20McswyZQrhMyc8jVzmGwcxFWWTJ
PEmXBybCditW3mfhg+tsyB+joYLfNwjyvW0dzeQBnlDLlsqfuaosbXKnEqwFtXmOTFpg9qi6Wl8T
Ihoaqf20FGhB7ho8NVHpVDGcB4+2GE6e3Es/0dusKuhlvoJdTQzgNaeQO7WfdiBclCndQhcWuUIs
zxydD+17mQygPmgcc31yGHkbq8agmNaiOrLaVAgDhLgqwFOtASv5ezUbaiTs/0t60ei7ndGyAGE6
hf4arNx5riERLHuSyV9dYP25jGZeMA9J6MiNhgzMIXS5EVSnksoOb76uNws/5etzP3f0uyH4MHcP
pVTNx/wRJ9+lIJYpKIx6jfCfr5xqsBCpItvFr2PUHoG95qJ/JwQPY0WnGf2BkPKPYkf3ULuGv7DU
Q8RXyy4pC5cVqkkPgIimP3Iut27lvK03RYubB+1T6lJ86GChfp8fSpvCaruUD/cyt+gVQHzmel/t
voxlq+zNTHMNbEAiDuw1WtY6yt4W6CWAX9ieOl7amnlkN0A9/f1t75xloESEMGYmLgmBStH0otvn
BMZL1vv6C/bf3eu0iC+iiBgWf/3vxVuRLe7IIkOMYiMyzcZW8t/Lrk+K5WZU1iyu6EZXSKfj29Ki
wzBG3LC5VlG/gAwRL7SbPaUHNqxVua0zYWsecjb7Ef2wD6/d5fm7+hFRb69ebf4Iq1PRnSxRzcK2
l/L5c6VrMgaWv+9bsMB2zXwCheyFtz7c/XwwoA+8Vy0oaUzX6e/7M1NLLrRGtMmO99I47GPtKwoe
cC3WWNnCZ+D083Pj2ldUTPUCez6j80dGQZSheO9Lc7rTxXwtRkZuSihkt5Kpt/7ybg2DVtRvDxML
H1/snKpPHVJR7NOgkpB9JrOQBPX8OpBQcAD/qTi1iQPxIApRzBRDAbhGVJVw9OUAtEPhZxk8Xi7u
jGxreWaGJWAPIeXzrfskMcDeKrB87+HVrj2oy9D4Ee0X1TaEIUdd9YaSP+PGABhwaCaqM9+USyJ5
1WgxIu1GzB+xGvCpsfiKpmngTY6C6YO4ydvYCqTOGemRWML6Xq5qNxCMhyjNq7ydGHT/ofJvAr2r
fPqOkng0/y3MowFZfbQlkzViCzlJHWBdaIO0WHWYjco/22THew/oZdHdOllrLTiZ8RXRX1PVsWjL
cVWRCupVnEPnOeKS60440eJmnpEtPMOEEY8LYIpBiNe6UQ09GeltUjcs82xdly0NNyarinLZ3cN8
uC9meme84Yy/po4He9xmuS40agRFeScys9YR/GCBojalA6cN3SEmFjeI6vaCJeNoJGJs6S7GOPXm
as0MLYC5KLBqrk1Gtv5bM9D/WZLifBptRsuYH3auKzDqMAweSlyH9d/IkDc4Fd3bhwfGRRqYUwN/
m/zVYFPO5Ux/P28aZw7trLfP+IAEyrfRrQl+wf9C8PUvgxXq/tb79jOvpM/jtfulcEMxvN3BXubM
bu8HWI+RVNysJ8CMGLieaeakA3xolUr38QJGeDj35R+bKpvWwIMWm+4Qj/tReGq/cc2DdkSU9DDH
ZaShyEtyzHVZ2v2ynDJZmr0zq3f6s96wYDoOarm5YuAF7LeLIohCsosO4cdmHtH4QpfKvN1nP2u8
Yr6zs7gcsPH8Oak4wM5Q82O/KguMm/gypgIxO8noN+EPgM1xKrSTWwsV1oM5ZG/Jf98Y2k5LoC5+
+38PNxZnJUJbgEV6mAiNd/FGMyQGFZJb7aXDrivoLqhwvx4unaVS+qcVHyN1NGdCuX8yakNIhms3
R6M6OetsaqTqMqDFOBcq1oV1EdjUmBp23wqhhmMMswOnNUWwroB9VNgfDePzfyHkJ3LgW+s6/AqP
RxC904UUmoiLl8kaWTKlVKH1q8Er2ci7JZUtq+pN6nCMeO0n8b5nAN9M2BZrKTwDe8oPILYDPXXI
9lFUy4G2mgEMvyw/YDW3oW+UDACjS0DlfnzNl1BA+UvuqFSD6/8y8rsSR7LiDVN/BTOkr5gu444f
fUVYF9ZKl1NA+7YdmOGOlOyQ79koOdzjPy46CIEqzyJKxpvNGflbraI9H6SC44E545TqVOV4QAqb
2HxXSxw+oZl27a+uJS5HduG4+eGilPfZgBFGa1KCr5J4xc+diB9QVHYFB0oZuQPL0OmiYnYj5amX
wAnDltEz1F/PNrw+ouK1b49ZICyPPyy8GRvAQTSjKy0dI/1dKdtkwbmZz9r1Va8DZBC4oX9ytxwX
DXRDdCM1c2y1bYvrEOTMNmk5gkyEI4HDlb8kU6OSjcwqzMHf5OOIbC1rVMUm/Ep80Aumr7YtVfzh
SIXKwY8JX9+x96TFUXqljG2YXNn48Jg9gUkkFCEI2j675NO23knGs47HHIP44/Exqzy3qVACDTyR
sMYOXwxXBQ4RdZFrIGTTfbsEzIKwAMFKYY4lV5XpcS7NTtl8VTxODGZ4iBZO7hmEhawV2yUaCU92
hDgTcX+wJwa1Pg9rh4iCk9YInMuVXlsKKSpCwV4tBicLK6J4xf+NbJlErrKWpeudrVdzPvmhtxku
2VymGC50pWfvUTmx0EmxjSd70CTQWm8Qt5UuuNySKZlvkjwTzLZklOuoagQnnzL+wuYnbWJM3eoq
cgrFInAEhlk57dCIUojMBAXcjg2Q1KdcDJKzigmKKNSRO3QJcOLNvHJuI7C5YA43o888RIUP6pAK
EysZKzHCEP+3w6nXXIdHnxvKt5atFckI9X8lY+FHxmkWtYm13f+fFi0Yr3DhCqKq/2Fvw1FAgP5I
cV4/TmQOg+dhXPBFwK8XvAMecgxRYZe4NZgg7iOJqpfmNd8GlQNuF6CZqLcfX/+FfDRf8SarCXrJ
xEHTBlNXm+oHyvqsRX088rpCr2/SKhv8uLizJDiiULSvyk39tgVvdtc9Q+DBkRHVD51+dzlo2Wki
l71eL83AnZ2nKVO3yMIX9dYILR+ko3aUjH31DiwO9AdL6vyvTBFeEYxAFex5zMdpvqRe3xiwsE9P
MNrqH4REj043Sy837yL2eB5zkG4CwYpRZ2mtpAGrBVRNn/qt5vqBWFFu83nhJJZ96Ac0VKQlPgNR
yZcPvCn6afkVgkRQDiiGrR/KIBCoBcM1IHsmFh3nuuFNaVAZOvM/J0teE+D7OxIK1p9qJpg0ahH0
tL5ym4vMADWIIMdYtFPpFgwYXWIBZa7sYzfFFVKoIoV/9aTEKm0w0p0X8Z0mzDnX/ohTuBShvKzK
efSabaGZP4Z5HMbtL85elwvRF62TsSbie1E9vStxqiEz25pjSsP/UKRAqEOpaBwhv/P5p19kLAG9
z5qpnVfGpm7J2Mfb83N1wWFpKRfXawDaOxY+l+W3FguVJeT6PbdGAmbR1aXILfvAGUa/1WMdC9qx
awvf8pQDzU/W21+FZayCaoEbtEyUMldcHpB/WEqFSYs9X/B3gG9SGpGF0SzSY7rfWzcSesyQHBN6
i94VrcU8WjRTE9fMalso7h9aZ7o5L9hPAcZQa68Txix6lTRqFdELpAjbOhiZvCL1kh5WktCErPly
5aIW6c1ZaQ4pfdreizqaAhbG7/wN+xuVxfQRJUsNsqifCK2f+wvnwXlHfItPg5YGl3aUusMnhpNt
btmwjOqKnd3rmLKp+Ti2q1ea54x+eyXIuuxu/A48UYDBWuijFmShtR7lkMte8cAL+k3JFfVMuQnd
+hKmBRYiPtUc06aTVN3FB2Xy0jbCccq8xpkt1znA2XNuVrTWI8Fd86/DTYOycq2qtpBhDX/l5o8Y
Z7lqQXlGUqoyQ7bAnRYPRjQhPZbtiSMR3nk+/pF2FQCmAn2fGau1xpsfi5PgoVMITndO15Dg05m7
oSJRLTlZYJssLxN5l/EWjv65asZ7ha5s7suldDLqVUpAlviDm3cgCkfxtMam7KTV+f0qL/o37QXR
1y/TqQWwRM/HJ/TBsUFUHM5NVMCTo8mwDhTqoNLDpwBKQ71mGsG+ua789HqLdVuhjqtYIccplVYy
v3UxbvjGwtFczAktJpqzUsxLE/tHUahCnkQtwVw3umzuoEft7KzbvGwIz1Jw8CSjJd/QJDvs6Kib
+pCZGEQM9uk2Ks+R9syUeoZwsvtomz3NkHeZLHO450+CgUlPOruBdRI3VCu5oNIu0dAcp66SVaZL
k30RLnEeATuNytmRYF0ghJZBm3WDe1hhpliuxXhvEO5mPptoePTur402WBErnaLY7zslTuym3Kwo
Dgb2TDS+KI/8DutvbRdoyB/k9Fo06H5SM9yorW90V93fU1jfietJtZ3cf0CIH1DS4M7C0nb1u8jf
G77uf13zwvkncDeC/sd073nlbZrpTJKSH+Aq0ozEPuMs/s5CkSuh7eFqgPtWkEZVcZCkNiuqjLR7
V+aHKmPM4XFEfY3Iqty68V82jeZvZAt1jmvf2e5Jl+OunJt0pxWJEaICFA+5e5vNHtUb7Hk6rsQp
J0tDx1w8BqfQsFlFyT62RXis8kl+x9dKsvqqYVDQJAATgcoduRA+vHD9cCrQpZlyIJWlgAL3aHix
aICQEAaidcdUEr1w0VyGrNCKYQHWjOozPjT6NPzzVwMsYXgakYW2pzbu2uCT3c1+CUjYSSFmENxr
4UZQlvlPWmhkrAV0mFzOwrpCMexDX1P0kG38pRJ12T5XbkeYxWzyaPRL1eb3WbooJ4av2NVmx4+7
rdmVdB0PcQKXhv90Zdd88jgYc2dcCHn6a3+rN1ukgd033NBLrygc3D0l0mJaP0S7oLTnCrxEfdMw
vl9ZLjW+HqTR/mpVnr9iMem9pXMyMRubYGpua1AjduWys0uNMaT9kJkCWP6dxZnAZfoKadfMSOJ2
QaZOhfa4BwmmHxC3zOyIuM4RxlkaL7xLewmo+cH/bv/j6rtOmq2kFbOaSJ+VpMmSBCuww13H43XY
d3rJCm9tkpMlsjdN8wirDK/lceODTRxssHeb+fUPAY2qlZpaafenG6YfjB/spmBjCYt1dZMIxHJG
x3fAMKB6G7ikimHEpyJbBSFjNYhpvcx39LjAeQ2BaB72EkVrY+PB48h3Knb8ffHa1f6/ALN26rEd
JY7XoJpY8z8EidhZ/P5V5SbDspyCnbOKEsFy+BX/8HE5wqoym74rkII3UZ/iLBd0VYWEq+ruZmh6
HtnfNAh6XFq8Tlqq/aJh44296ls6i95qS/9NHQ7clgMWT9pbZJEBh7pfDMErPvFjwyupVIw4+gZO
5rx2td2o0RCb42GWlEmaVlOJrT7ZnLHW07cBDBGde0L+NvdWra/KcahUNpsC4WVqslQfy+mJ7xgd
xeJ3vtHAeHsMI/qWQWmD/yC8rW1Q1tSzEU2QctY5s9lc43pIqLQWUMT8HSUjgEBK70VRQwruY3kG
qTljgAcL77oSDb3ixmt10BbDY6BriwEcTVx/uc6NcEbzFR+XjR/lkrX/kfgKn/L0ji6rS1rJDa9d
cz7yCz1qJbRHH+oS/hHEJ3qZgWptHdvoUlZz1e1DMSq+EjGIJa3PjzmxwbqKKKLfC4Q157r8VtCY
/PJLSHgnSQkaMsZndruXkchqma9+aV3ygfj7ou9M6fYSnHBIgXP80r7rGvzoQ1NjBQQuXtOHgv+L
8YXxTvKKihyXWZ2pFM24SfMQ5G9Ng866AcAgy7auACFhHSUyGA1B6KB+aBZ7Jc2cS873czF4JIHM
wJrUjz6GWTKHx6QLhnRXoKq3Q/60Rarphjw2S7cGsSI7DgsGPLapHSDldnbXqiGNTGw0vWMD8a14
jJd9YzMIghBCPMf5+0FdSlEW+bCnHTPa3eIbjnt/03aSgp8N5l/pXrFzthH9OuGY7Js0G+HNABTt
oUCeehK6NKB/3Ij5AbwffUzVkhNEki3BB6CUcYavlrW40TRIF8C2KEnWxbpxR1DezaDQa6cOdCDx
ss1PyzpQkkrIYO49DYtgnW2b14DO9tjKHMw5/evVjRx8wcb2MyEQBgIno1N01sWcwhQzDDNFuJav
G6HmmrPHeihyQpFQZzMfLleDme3fqDTAMmb077zqf5nTFR8rDrzORVL5YfipF0Xqo89QoQsnRXQ6
XHf1FyeFEvBMFWpaB4RsS6yZAYjZh8vzjcYnlsHXEuaeaJ63Vt0i8QCCP5ME4eoTc4tTuKhtbvib
PXV4YoYiJ/IfCF8CsR7c5sIbV/So5+gq9oIAn5c359u7Ir65EIcfHHmejy45/Mbgni6bmQRuqCml
68CSMZDaCKbYdBMd9e3Ueie3pQHdo24DwI2cPUTwJEWOW9JGJN66F5RATka9M/2Ah/y5cwI0sci5
EK8/kNd6REeDkZ2qx+/uRoOhxLrM706QU7r8qqy0RSbpQcV2wGAQHRH52asC6oUC3muZw4zJwRMP
MO7FCdPHjch8V673SbUeb8QpKgX8kpcaC1AW2b+J2Sh4DzqhywMNA6numYRxkLB+V1j4hMuREm5p
9h6hvtIsrP5Wm57Sd1BBU7YurcWby+QyW5yBgeOCXXZkvyC/VluyUTB/wJe1Xi0HKLiNrYRSRj2D
YffbB6wW52KSiuBhu1Qr+uvozWmyN40jt+v5Oe4rZKoK9SRVonplv2weSYiqByEbETtJI720F92o
Y/ZKEm8sJVkbCu4ZaeAr8tqVviQd06eD7YPqFCPAOEOPQ1fWnY3aYv8jnI2pjJhvmxj0IIYYvnCS
LmN3YDywsPnJpo51xltPAgJIIJoa1BPdd9oVM6J6slqsVv4ipTI2iU4gf61eYw6IIami/n5+hK3u
u5S2mG+mibETEauiCuWpT3QMWfrliKTyPxxbaj/jm+tiYqzuLOJDFQU7VAKtpTbyNv4hxosVxHM7
iDid9vK3Xs6+K6J33bxoV8AeUWhFhJ1OxiCRwUHgQv/U/GDeT6VlzONTG2mWVQiiMH2q0LvOAYiU
rZ+hInv211EpGO3KST+6tjCr+csv2lRNOJITsyCnVstxtpDM8VoEKq1BVSo8ZVmeqU8pc9lV97e8
jswFwHx8F97ppNueO9AQrwwTN9xTJ3hL38noONJ4XObQVAqUotIwDQzxLNc4XPuIjIkKI9Egvb3W
Slh9YyAjNErdtPK3gqog+0NjNXotOlf2dOe9iLC+72nWnqKNF1mGkB1Dub9wbMaNFoCFzds+YVlb
G8IhX0drGKxOmicCFOyozaIpvNMJMPJT1baxsWNWSNKYUHqtNYTqatOtsA2VLweLK0HePyYJngUf
LaZEuMDOtLs2vQ75LQoTs6vrJ7iIX4TS1CwCAWgTfWsK1+IctfLCxTl2b25IDJP2lwAqUiAlghFW
3rmLAemqiYIAmKHZieG+FYAKriz1LC8M50lYDMsmE6rpLM2vsBh1nkOUmRa4HP8ncFoGNvu6CKjF
o6P1pB/f5sRzQRWGFV1dtIoyNXTwjRkmZh1AfXsRw1vzSioZnpwSkBRnh8geRJVVIoFH3HolfmKz
kglOLdBWM/9oSRXi5/CS8vp+80+GW0THwTvDGrNhI+PBwpJenboqImgX71jooe4Z3cw5xzEbNNCS
FGLdvBMi82nOOovx8BZqtckf520Ib0dhummpQnGpne4dJbzppIWyzitnMdezu24bLBaLmJZJy8IW
anKWbtOKVlblLjBEx4FLiG8P3F8ZVBDMdUF6rVOzWacKfBL8naKJFAaKWAK+aPfbt7379TvcLxHu
8OWahuN1aCqM/1BhqlemJkflB+P+SQ0u9nFohLsNR+kXt2u2LaQ04lS1V0GCJbH9f27jgoVZTzc/
I3YPvssRJg7F93Np6nYoL5PjMUE4GdE9QKoWN0ittCyUtA6zqTfyhdlE57H07Wuzal6euKZGbKwk
fRpB56L77TCnRUDPB2OUFVA8uxiv5lHlQTM3rE8ZOUiCMtiv7JSi0uf5Ga1DA1bLQgmoDxRDiTUq
G9qFrNntz63MoqzZJe1Sw0vK21Lwki3C9imZsaoHeUy/NheUdAhQ66NfeAtXm2T9uo726l1h+VE9
dkGRQ2mlva7Cs393BsHM13FFLaWR87llMP06PprqvzNjWKGyfqMS2pRKIpvOGFstrTdsLG4h8DA3
fCkgCHN+It0aAGU2CpauzyOaB1woGb5ySRGwFLZ00LJ48tIDfL52MqPtVC3ZM7Uj0PDIfkWdWvXF
4JjGoeEEUuAKnHFKY0bmauBnZUWfi6EwDheD2FJbsumuri674SslqvXSo62EnPK2P5nwGRda6tAc
0BLJNJeW8YAxoYZyTElPq5v66olAJZdoSrrfznypZqLdU+dMiFLsuUdDjoH1SR1YGSUvcF17J5L8
DcLctetwmq1QiBq+OmqaZ0bB5glVwuGHsWiqthKVZuLY7vxdO3lXlRn0WVTeBz/IItRlDJHwL4Id
TeW2BCDETuF9Sp08qHqoKTrDjNq21VFt4dpi2mtCio2j7TuySv/7ltYIPTeWVnWqn6t55EFSHkgN
ZQ0nO0jDIl0VRov7ayjwrO4DkF7iH85yfjLDqgEePlaTkV9lM9McZvhivREJf9z0RfU9KRXytm2H
eUgoFWRoBONTGnyuWV9E7+a4zDxEkZd9GVfXO3POLl1wzX3PQNEGumBgMOEaTStQwTgCoiq7XOlC
BG3Sr8WAzhn6pdAOfFEkmQzvJKtNHR6TZEGWZMVNmAs2IayFb0soZNDk2mWezj8dqRzdSkZUJ659
sQhzokBditkee4gZF6tYN/Rq6ANTH4inHKlnhgdFEwbqq4EccaKykmOqf9ZdStIiOp74rG8nbB3A
IVWzmii2/XBqx8XXxluykWq7JnEv583GLblA3ydGQhBKMuHTTPpI+mw8mGd3z9Jk2tGRrlIPP4P2
QOIJUh+fhJv3kR4eHE+8F0a2z2h8BUddMiQlsPYViroowG3JpvESFPxIzS1VmAhhfO04yXL/mkrs
QTP3nxHqgz38SQ66+XlGujZMhy/6M1XHf2px9U3FbKRtQZQsZdgKZMyJJQuhcsgEin4n6UcqDMpM
laaom1eypXy1k0XzhOJk2CfK+WOZlgfjGoIcFJe1wHNwebvR6LphHZZb194JT4aolheXbkqyYCMz
AbBq7the9hGoU010KerYeW7Podd+tOYPRHTnli4BudCs3mnjN63qwT6G15wU2iQ6t8AIlLpySyR7
bJ4hFQGXYp3mx4nt1O1bd8rrA5mE9QT/6AT21S/AOaim38d/05PQt05ssc5WRfZvGo5WPINKPMBH
+cYeAfxIVYZLM+jSDP04D9b/Xk7sGDKeQtgGWnS2m8YZbSulIyUaiCnis2+HTCeqLrFO9JaXmUUh
oigJ4SRkvIvYsJCAYCU/JSuNmkvcNNl54xb5mn23mk3pxUnlZ8jw4Z8R0vjWo+uC6Vm26yJ/q3Aj
d94/MCF5IyjeprtEWTsq0EBUFRMBZATNIRJLyXIrq9LtDCr3JNTtZsLuNe6z4MtkfKPGSnybgF6Q
UR07QRnFN+ji5OWw4kepNuQKJULGEjs3EOidDdgotylxg98c5GgNouxl+LQ9Ild+eHnyJTTdN4zE
sDpxVpBNzYwJLw8YWE0Bfe6AAhQWsJ0ISz1zXksU/zru1tnlrDLQ3p3F8o9xtHp3RU42nVcch7TB
dSne1loNLfBdR2FuD8SKkC/9ZmVIAZz9kxbQwJ1KKGwMWbq/GWF+ja6qNSdsPsjSpsccRtt+PyDp
kMAGEHf/CDnBjQeAt+86kiwfxSQQwj9Sm6Z9RnmsZSuMJd5OKjNhf31jJLvqyrD8eHMnNJxbZQV5
mwmMrGuHC+zNHS/IB+CE3ExCQszlrLt8vDeloNzIG5cG3rRVeC7BgQjGP0g0M73kL4N6ktqfscSz
20gUxeIZw/VNvN4HpXyqTimFvW13fev7KlCk25Bf86ZYZGCL9BgEFIByHOGwM6r55VdEHv4aD7CL
TMvqLQpE6xtKRp82QVTTbe0PIyf/apWm18nlQm1oiVmVzs9vPc8SwVSK6C2P+SxrsH8//LGP8f1/
qLo39XwMMTT1U/qrPbt8IIeFgf4EeRCH68VWK7y69QsL/oX5wcfyiDXPsfPla9Yiu9tCpNzmELyW
0nuOseBFbVcdtoph36TLyoKNenraK+W1B26lAnO0UWsyQnO7iqTaJDJixYimoLCV3riyZcXrn8QI
PQI/tp8lvG8KfJqUMsjlHgd7B4/Nz15ssdxzbQ3Hith1FYeljyjdnXd78upxL5on3i+KXeYlXnX+
G7VKrzuWjXaZecdLN9ExXV12C2uub4N5A2+bRqBlBgf2YCC5QcljQl+rBWEbqhc/ESB4TCfaBFgu
L5Zl5wfJ5flRxyjkjwL9ASPsvQiYOIkm1EfkahnmVvUbixXUYpHCW2PipxQUjr/Jyt3MHMFQRLRK
fAOKg8NHYo/sr9kF7NBb62xacLuVX3SPC2Tr91Wkm4U+YvT4/5kAA8Rh+zSxuFqFaGPEX+KYtyX/
2rJTry57hdoNOkOW//zfI93+dTk5iZv7Cq5kqK+q7/DmVO0mBKNGnCtTcczZuW8cOGv9ViwAVmNH
OzAV70mz8OPIy6NNw6W1xztaMxyAT6fy7DjYWsUwy7Fiyl1IZ3VUtFZ33boBJ6uDotjnbPM8Y9Hp
/ho7FNuNw5YIWSucOJ5O6nj0c27/nx4z1ZwQXTbSDfZ8+v7Grgq7CYZKB09eTv0y8tyPz/jLU799
dm9o4QnTQ+BRJx+GKDWX0Yu16DiwOAisiGl0L3erIdU0jVSwVpR2+MK7rG4+TEixw3hHUa90793+
Q3Qnk+MS+DlLJgYyla8LvrHwp+Nd3DX7Pn3ldG5ua45C6otV/Q3ZIO4xNkTfbwM6Km3BEUYIUwwk
g8MwDOO+9ukiIvzlNb3NsDB7P8mpw/WJCYqnqtSCLS/LVtWt15mCfRhmlYm53wy8AyncohXYdjpv
/RfjopxqSqdugNIBfEbUJQJRQoPUX0JAXpy+rk8AU4jxnfJvxCOgigIUEm9GILqIMyPA6ZfoHeCM
QvmQi1LoqBmOstzAUl8C0e+5ywJp9e1Rw9El180nAtfog9XuHjDYemdTkgtYRGSuPPG9JJiF9SeM
Idhm8Sv+Qnf+Yl1gGrrJi4XDvVDu6OXWCaEO2QLYqq0DStr6y2ZGeYCPA1i223ctGNEo9rtUUOcu
j/SYBTcL/JcrdLfTJTUYsBGk6+0Xa2MT+4JuQmQv1WaBy+clBQVvynXE5s7q4xoy1yIEdzHnFhtn
l3doQn0Dz1++nW+v7EFdN3TE2U0h/mKteDJx5I848LDt31/sXE2KUkeCNOHej1kMEnyA/fW3nU01
L+uuEPsTm/VT9mhfVruEPIMRubtcUc35nCeFhbJl9Wn6wIzChzmzIlOQU125LO+7bG1aY/oaKZXg
l8P2r1qo6gYXfhgcKoiRAbpwBcbeAVdB2uYkfTrV0QHs0j6BUeBzRlX5Q3QmsSgzxCEp+OLxpzwe
pJ8SUmfDYzA/Ahm6DVHp3M2cHDXh7WJ0byjsrnj/oJkgISHbv1DYcNhToNEifmRhqkxdFiwMEBM7
80s6MZ5+LKRmE0tU6zma4/mbYej2QyICHpXZ/xRJcrPhANp+YzVaai0T34vUIZKbsiay3P2QI1Rg
i5ThUItkAgWwcPXmsTVyw8SqaGtK1+SgkX3KY+BnHki+yM88LA+7uv1xxCogPfaDBQLjzAtMuJUG
fyIVzw4pULVjlU+GzqKQOk7vu115bMDGajtJc7VscHqihJVTCj5W7P61p2z0Fy1Uye3OQ7YcHWE5
f/w/pndjHRpXHLc6ZFKhnsW+tC7Wi3IrL8JoIFrdmZSsDyMhEwAOGBhnGGBOeYacm2OpOilugluT
VaENm9LjQhynxbQzQ7DcLdZQCpSdfxTBUKO9SX4Eeyw1q+ovnIPbezYNNWeYbfoETXzquZvmtcOg
mZ9YL0P1gdrXMP7U+5VqS4ZkOTeMLvDg/vrzzI5NdVDR0KjLGl8kxApaRgogd47ZEqYCR/143+xY
CcZ1KHT1fL49IfkcN2/pKUwOBG4wEmClcDQllqBPaMmv+iA2itPnuz1eId7Eky2ppV73czefsKEO
+6Z4451LNrb3f3jTIHRG7WNs45BYxSwOHtMhAVph/zJyyvwgcd6aKdsXpRPaAXfenSe2BYp1wf10
Gxj1miblyfHavZTFkTqjPgTw9VxpvCuozzPNDj9vzOyZWQFYrhxAaLtxrTM0ahNx8mEyGY/SILou
mdxedqFWB09mpAMR48QLaOHvj5QzjljOUpQM2j1So/3ebrgJM5u/zRKu70J7JrbjWhTMnh9hSZuo
zGeR/Ox3M6WB5LEL0g6XVjv9cQ2hH5GfyP4toFw1o7KmTDqLFJrsqVDXYmvaMz9bVmCBU+8kiz9V
P3R6vAj7efRoiDFvhqD+TJa/qCxo36j/8VtffUfC7zBPFOWJT2z98FkCresN7tR6zlCZyatEI2tM
REsbPPe4HYHkmgyGBLhMjmoF15JGMeHz3C7PZ/Ydlr6twOHK8yc00G1dVjuIBTMKw62bZluC3qVp
NNWNeFL8ysRKWjnbusfcRA7+cBnE8Pjyg/ith1YVRIKxDsxtWUhBtKx8H5hQ+UcdDtLia9eK62DI
dQPkiPFO4Uls/4DNcJOORVOt2HMlnKyiXuxqXbpWm/pof9ENDXyTo0+GbyQ5FDXG3OJejDfEaLD4
7bOQo0WK7f+97YMPJPCvvG2jpzYyUVnFR98wz/KW9++nJozXIjH17KfxGr+2bu6Mabw4VNoLfsOg
G86j9zkdSoQZO7W5MAUDKZfdMSW2VFIAz3qZ5D5zgyl0OQSd11KGebsCabvBndiO/inizk+l2heQ
PJOaJPdDBqXq3uF8hYg8ozXd74mg83zGRVCn0xcYd5Oufikn0Z8JiPukbLhcZveiYufxr1ZUPY81
vxV30XbtYyPrSwIQ6K67lBl2QTk8BuZku1CCssLICuThiA32V5+o7BK9WBoxHSOtRYcQNhVzm8Yt
J9a93wE86VTt6cL+CQ5G0ekDHVKhZ4GBuyLOcWslqJ1RLu9mwMcKUOfxqLtRN0Did18x1fAJP+5D
rXdeU8h9OlGTIRFCD1VHRLMDJtel6rc85SLwBxPJHuU8RkhEh/ViWB3KJsndi4kyl9znSDnCkp1Q
G8zw9W0Ph9M6X6Y/THF1yv+1Ux2GE+0UzL5qf/qnS/W1WdzNYhDo4Sc1hUCPYKrv8RdUqLcdU5PZ
+sfo6XHaU5GJKXIt9NHUxMTyGxPJoZ6hD4xULLCeDu4vwyfvJp4kZZF9AQucMYwyxmI1L9csBaHH
IerJ4bA8EnSQmC84gMOuOG+QXR9JJpmgmglvm7dVnJY6X1V+p/NT5Dax7DOz5ImFu075/0rqKwv3
nXNjHqTmbxd6dJUUszTsB/Xa9V3ZyG8QjqlBDpqBWis1m8x7GYCdeWpmd6SD/zbFvyBBKA1kq3NU
3q7yfafhNQpmWLiDK8cpzzBpXijlbrYo7BuYX79sk//oAWhsl2mUru0BHikwKv8zuVPQFnKEzpqV
8vvmZg2nFFOnwl8cWZO6+A0zcxmN9ORYFLLBxjnmVz6id2fNEjD4OKud0HlBYb0vnHyKBURsdq45
4xdk7Pcbo+7DhCbM9U3JKBwXVMoDsxu+oKEdh6MHKXHbp6P0+dSOe3tYpb16mV74Cm2UC2TSzjW9
ZWq8JhIpf/xeZPxoq3XglG5f0+NyK1xEeLbiH/E6TOiA8ZOAG13yl1aY5eWLXGNAbiaunWGgOXRf
LOy6PLdkxIg+PtfCAVZ4LB8uW/HU15s1jr7cEfFNdFJjPhC8UNcxgEmo5fzUnutwgsE7L4Cbgtgy
5/hY2m7KSSTpEJDDit3XZBzdftxZR59Z1gj33pV1Ht7eCi2sBfuOj3CAM+j6HeSijhmof/EIAi70
eBUB6DT9RuxrwXAoB5rr2k9aZsKXsaa/4hurAHdICZfs8iyjOYnvjl9pw7nP0Uix9JVi5DWxu5gk
dsliM71NMAs9iiaifzSgDsJZICaiWjr3c3d1G6lv211lR2FXuckLilh4Q6kaNpGyH5vLyhZ6ni3S
YPNw01UqGxfS6CRWJieMS0Fr4/AKniaebNvQM8O7VbvlABGc9/8WWPTppwmWZOLXhAuHZTef406m
RIx27YXKz80QtN764NWL4EjkjfCDLH1I+Rf7SvqORfzU5UCWHahl8Zisfy0XzRau671azaljbwpy
I1WdihM9Ii3T8d0EMFCdz2QQCeJPpqWGQH6Ni2LloFGVkB+QFx3PTfdS7ky/Yoi+Jit0wmbc5PeX
PH/PW2ODNU0RubsQyX8RVq4QgtP+XreEsId27hFTGmmDmwOsHtUJ28WTnNlW3PJoF4lr7lXGjXYk
MSYTHt2vYQYqb/EJeLrWcStae62fWtSH7h3uPcFpAN04vnD4dahajyulJ0JkUzFFTIDwP4kbjgLt
zHlOgSvSdfyUnxM6E8Bilz1gSakwDq4aL8wrX4jawNm/mHioVd76X+o+XVnmzhx/UJNHOtop5f87
/mX2XiCE54JBaeNTIFlihkaSWMhbjwgk40xD1EBMZq/xLklpPGn6VxPomTNQq84aT0BOHjGyRlym
14Mb84FzSohTdV0D4O0Z2y1IU0XnAwWrMAi1Ou9Ojx7ewdNfrx0EB+ytqoLai+APtNWrgwcXambn
Db5oOAJ4pjyH4LSsD4zdpULu/2KjuwfFFEIpOh6Qs2aoEHKk1En/B0dRJAu/M1K3XK66SQrH5z+Q
Ba1ce0B4+yVsJYv1PMRI3+knJ66JM6i/4Q5zLXMy+kUy+LQJt5O4WaBuIQDpXcCYVSmu8ELGF+Dl
AWOQVPRy6eIGmPcM7oHCkiy+N+8vGmbzRVB8q4BA8RY5qJ0y8EpAmssbboDYz3ExSmm89QagDNwH
5RtYknp5iVZL9Ce9QglVtC60yTz+49VqRoFUS0CkkDlgHQ4JKpdBlnvCHXM/fH4FzKAESrQPx7lD
55VwcPaUe3DCKpQDwGn3XOww1l9bCEnMu0f1kPx/4gDcxo99QWSt+oCGcIGnlOEWT8hRyNeYMbcZ
owQFKHdWOjceSwjWqdbAqi9jDPfJLWA4j/Nz2lEgoJkTlOMrpH41apoT08fGV2XvQiT2/0xmedcn
lnVJvm3yreRFlDLs+T3erDtdzduhKIVLrU/gT0c9lXPbMBLwwD+GfPNDRz8ojjodLeF4FXG0vVp4
F6I4p+6jz100cc1C4ic6JAhU0xeiH8WHmVAvhskQ1nq5Ki2vsMGGZgc+4eR+bA41r951dhUzWGyQ
VtqC/KvG3eJ6SoS1mLbIUWGX02cra5tkCosLj4lfxK+A9EVFjuN112ZT458R1J/PieeFMSoq1Eo/
J7KNpdao4PgxyRXoBgw2wYMXfzOU0fNEkyjRe0FzD4IVIil53yAAs0u/XBmYQ7BCPx8ne07mohuF
ROySOJPDW/IoIvX7RmlSS02fLqrEtQjh8HOYv8YX5Q9RBfJ/nZjDOKHsd/mOH090Qad/D3BgNiYS
sGoI3rOeLPi49JCrsK+f4yxc5Mx/RIW52i4Lxq6oSTeGp+TB9K8gj7pReXHaCX9d1Y1ovw9tEb7/
izcKxhJYx186sAbB1qlLE+TMEFBVnKjlZa0AXP6L3oG+zSOKRiwyluQn5PpJlOQ85BW5J8bDSpSp
xPqemC3GW2dGINn1von0Qt7nzf1QeSxo9xuE0CccwSN4ShpQeV0aIsLmSYAVfGjSV56gMS1Noes2
B+0BTD+0X0MImj8BM+VjLWs3R4F1qcjeM2i32alwOEQUceH2194wPijfWJYWui8ziAP4KEH1QRYW
ZTAC6PDtJyjmz8ZTr0z6cd0QuZby5hv79cYnV34HoDWqvTVEPyKt35JrIYInQz3MoAurC61xo6pD
5ptWe7odJEksDv7bYGFYO4oTfCahv3S2OVy4vWBXGoYbT+upbyKBSiwUdJQvE36dnI2S7MzlLMUU
74XX3BHNaJOhNFGKMyNDDVaHcTPS6AGrjkGyK0Q5U0BsBdItmecybmaAl4b+fyjJU16gY6EMR2g6
izIsvHY2I83zXbxwq5KP/MYV2dmFoNOT6Uuo2z95pfu/QucB4BzvcQ6sUfqLrkbImrUDhkb4hstD
5Vu/eOYL0Thm1nMGX8JSLBAaQTEzO1VzhxPayOOO0W0oJNhP+MZoC4f/6mchP9JJUJdnmE9LyWBB
6hAH0u79F1X4m3Uik8weaEHD3Tda0xcIerCKozYZ1ndOZJe5NF1epuPB1uPoDAWVP11EtsaSUO8K
hJ4+UDKmv17K6A3DuygllBtraSolILHYyDg7w2o2lRZ84n7nn9yZ75IqpkX2sF5e7J0Oc9bYgVdF
BhLlGnW+iFRRGYIqTEd1PJXL4cSoEGC5e54I3PJLFE8ya4YSTfDCAOOVPKy1gnNm4RegOw/mSsZC
zpqjRg/pnIF/ouwKF2YS8lU1szvZlo1RHFs3S5omOgzxG969QkLOIzVI4APDNduz422ZvMFXgVRU
F9p4N+ShOZ7RxaBwHG2TWoB+Chlt4cxFFNS7femqsm3sbppnd/Swhk+WoF85Dy+MNPcmtOUh1lLF
4e4pCxpSwE9uaO3bcvhZNWecWQ8zspNioc1Sjd9HHtvr+DrhwqEzxwuzmvSqir0qsMw+NZLtaFND
k6IJzwmbq+wPkfZhPYTDlrYqgqjNx1b+AGbZZ8HqwiW+0F+w9nhmwhEiimLkBbGVC0I6MgoZaZtX
bjtA1dUxZLrUa536B/pkU/LwM2xuX0W3lX2Q7fsmog529V+VepJ51rwTLm7B4COWeZro0XiVkxv/
va363F2HnbxP7m1sQKSZLQRkV0eD6obpmyXx2sfODpdZjfR4q0J0QVWAb4m2KWiKBR0Em0+SyXJK
6H59DBc/4AhYxnF6EJwnQTLgUVVjj9zPRJehUG5AF2DHBRWr7HSQgtxHf4VSNmhk4RpBZKTwg/eg
k/I4HCUyX6KYxWGTnUeqous2jlnM1NfXDmx4KX6okASnW0tSj53Ke3vuzAwjT7H8tLdejmn9AvAU
a4+aWn1NPsj8CMAuqh0riuZgCAvZOsKpWJFqNF6fX2AaqzL9gF1h7NsCT28NBrl+GnCEqJ0cGerx
Cg4o5TBL3VwIqiRHaz2ME8/Eoc2dvxHHryvBLy7F0OTRWlqKSz00ib1YbwEaVTui9eeZcF/nbNCh
6BKP+kRu7f3yZyO/+WLX9x/uxkpc779cxZpdVea9rFy5i2hnhlGGKqgWHaVZCqjIItmw7ed3+JRh
85XvvlIJrE+N0cayIcOl5fEj6fONQPuHi7Be6nrpgwpYQ/JeBNtFgrczibhO6JZrJwAbJt9T9/dJ
ZAtrSbkxVNni+BFWbV2m29gxippFC/Gy7fXR8hpZ/WELlOQHqF3dVXIP2CBk8xSbPrO8Bcz90B9u
fwa5kijnC8wFdpQd/U5j7Wf3N3TBDEQG/zB8sQ+zrtNc51aLaWQQAyXCTUtnf7Wtd+hd5s+Jz29l
a3MDdcf3YT+14B5jVUQRQPv97bSKNtvGMOAoXqi+9LhD0A9X12eAA6sW1jA1nk/CKHa0terq3PPw
x1PN0WIh8tSdU4/1C6TbAV/odEfiUYgeJATK7K/ZjNqYrB6SVGkdo3v1NGr2hqpx2Jixz2+MdIvT
0K6CkSL500ZCXUsRu1oTPEJGiKEKSh0xjrmM11rkHSHoFYLhOQJmuWSnIVggPxgHglcUHTkkNkY3
U0yL/nGrA/tSiAGODTG5EF/WeZofrfV4itCOrVgHHuoPEpaVU8yPtVjiDOy26JEZk07WNtxGfKUl
gBfwzxJok0hjy+jx3J18gCZpvBr0gOodnhFLtqmrAANnMY7M+HpcM+UexlxNJHREenGZWWGM3Wig
MSM0SDgznceojqC6qqfqUIDo9ajQyj0H3rrbnqs6vDQbPHMqdJWendpnD3mnXBQoFlyTZ9nozdZE
1XVwPCtEam7vHaSixEw+W2Fah815Rw/kVMq3YVWJwE+Mq5Km/OlO9YO18TAHS4EsL3OYOWTL4nD0
qsoEX5ZQOGoaVDvcwQyfDPoK2TS+dimW0VobNXKGh4rVULWsWPjThW8TI6Z2Tmmt4qiCIML5w/Ml
COFhROhXXFB3i+D6DUllf1WjursVhNlRKwO3/w11RsxL6jleSD4CP3QpDjsxRNmXOC0qSLiBoz1u
Fma1VnAt35BhjAW/fBlGi7l18gS62UEk4pmDDzztXEid6ieNMTgwF7cYBFPCeVIwPObW3R6rnrVK
bELrNZ8RE0GLFssvUOZDqb19qV36BL4w6D8a8WMNZ6aoIoCjpI4BAGgJAH921BHMKhOwJQxLAobB
x34IEcRXFKmUUd6xCQFq5bhOvQ+2doWa4MZQwaidS7ODKmY+nOJ+b1bCDpz9SlDTOT1KDeOG2aAU
ohGbsfJZ08HlqjPbL/0mYXdKobpXFtq/2aI95QWSXIfjmSz8bAj9YJw9eB8c8PokV7dNWNjyFeIZ
Fmz9U4GLzjcKSBhOrMbnYybYkCqagOFXRGPi3l83eiaWPr/il0yMFKORCRIqvQLg+DtVC7VaTq3n
GBzKxAgtTIvXpMTUWTHgulHe3WM2Wf+wECCwKiI+lU8Qb+DauChpNFxZy2mNKg+LkG1q7nk7E7kd
z/KnHKNBoOtusOJJgWJddTyrShnrsqOoDQrl8fRbiP2ni/61YvIPje8RLbeK42+RZ3YioYAN4bQ8
fyZYFcvFjzFYaz3Wia4Nrb0Wpaiv326a/T3cQQzYP922slEPPQkeVyPbb/CxsYhClz/Kjd/Lfgdp
8Nn+TuvW50IVXszn/F3KB6m5dpHUxcvpfXN/SdOWgZm4ekUsVoHKxBy6TtofS1JVZbLb8Jg1IAdV
w89IchiJtekha5f0CHXFXDoNJ6vOJWt2m1gWveXmBCPdvw9Cx4C8pvuL8diRJYoQ9k1HXC8fr/Je
AXImn9YUgcOC7s4Cmqz0NVE/SqBm/S/2KB2lOxObkEnA5H6EhvaIIj7F9o2Zk4YhDq/QS/i5/yAe
dIyb1u2YFn+ejjC+UUPde+Wq06kqArQzdS/ygqZwWwvEEJkbaK0sdplZslJrvq/Eu2dv4SgWyhmV
YqKcD3oMrHR+fc/kWq2HG2ccpenkku0T8Bw7pjsJglgEy8IK1hRcBhx23pVfnL+6y9SAGHulIvMh
DnD/TUdVEHG/BuuFYP2u1uo4U7myJ70eX3Jc1effqVdwAGIoFdOhF6msUbGBVNzfyQV2kraPXDpq
MxXqGvSPJjvi7lnyXTM2vCOeDSqk5oh3TSgbQr3UHiFixI8nlj+HZWNT6BH66nLYKw2K2WeqMITa
Rj4XWKAAK6xJV8PgA+EFnmrx+gmN8em7NgFvmcTvxu1PyEiyG1PWrM1dmfNh+tZx+HVmVFkK2LMS
3UHPu/sh5BRYWA2XF6knk6Qr4OkT7YOms5kuC1YwzQPusgK1IANqivSZl9gL8R519+mSof/7/Wbr
ymPjzk8KUX+nSzIAP3/i0n1w0eA61snxc9SmWbl297GDiRXX/4LKugminknRDeYwBhWVk9M0VLZx
1+elS9fBKYTwUeCVIIpzmLy1sSyNGtVewI8sEzX0dRehUMz0L7C/R83OqWpOMXk8jHa5MNaXtWzl
0nUf6VOQaHHxAQ9BhTDXRAeEp+hYm4lxxD8azaGWpu0wtMzMBCDZanPjcIjwirN2+J7Ekrecysja
Xvzg9Im2JHoqnFgUiqvoTMAr+Ppo/WrmMDnBBuAO64qd2qkUrDrZzvwJaqljUm+nwixGHA+4SbHD
e5NvzI+IGYtAwyaL05K9+4vKz6eVho0kBidHzdQgQvCYBrRUPyvZ/oq+bH24bu0u9YBJEd45/tGh
z9JZYdf3wZKHCKL/rYKTzgPYu+93G9OtjR5RxHoROD8clkFvMxo648oUEEbKtQQFp+S6EdYcPbR6
P3bDHwL3fpUJcfGRqV8nBQC3yiu8G1gogGRO15hMPROkKooZvfC8ZFtYdZPr3DVZeIZGRsq3jCR5
D8WjNiEpJKb5IuD7oZzQZKG4AUdzYYEj26SDgmZy8UrGuu44xr6a+WrrFiDFGBqa+kyKNtzWh7ig
t8sdDL0O77u6QXssFO4UfRK5u0JwD26/kClH7IoPb8++MlzjjoMdUijotrWw0CQ+yOJNqAPO4hy+
e8Y6Gg46sDzincoB7j/tyIftCepg1Ow7oX5vxjFdzCJ/gvEScCtmmJaMRRkQ92UYhy53y2nnHreR
PbyGdD8KCJJR1vvzuIar2dtzH4Ay9FpUX2ujraxNb/Z7JtKl+7lcLQXE1L3osuNI+yW9F8E1obyz
daeenR9tEGZLApzC23KQC6eZIWWwatKxicEzQVO66hnUDXkpKJ/PnR52Ux9z8GKPeGs1sBgyBk47
/dXHBacc5zFXXwaxFKQXNFZDUzd9iGDxpXVJaV40U7DSC+HVonOzJeqUSwyI83QJv9k2eWwUxK/t
lKFaZ/Xr6UcCKQrojEyiMcKPpU//3q6ytDPAOF62zBmxBC6RbWX4PqyElFOINU8mqthAoN+QWbKG
p5NfG5FVrRK/RzH2frwQlRylJtViAMJKKpuKGUBS7LrdX95oD0k3Vy5KUj5EtIPLyTmRoBaPbTJP
quIRZ5AkQUfw8n/axAJ0VaozgO9j0FzlL4sJ7RrQXmfutzDvSwXWsf2csbFUULIzEyABanBBr401
aWhfNdQB0vmr86uHF4LwblPZjUTkaDOeo/JivzNEmaLCNX738JeBlGA9TmI0xT6jgoUoPp3+JuHW
Tae+byXhbJOep1w/s6EG7zsWAbfGDlqA03+1JV3R181d+0kD7L0QZ5gYdX0Aj66nJ5WCsiYAeE7c
L7JgZp2GjpMagQycL+CHOKNBSKWXfDxzHCPAqCjpcyU5YGmM7uQg7eBoilG2KqUMJFcI4fMahbO3
+JkBv8yuSg/Bsu7Mq6n7fDvPegTTEmPa7KjuPrcLveMZXFTQoYEWXp6805b1TeHBcP1sCTlaAgGr
+a2aLLk7wy5uLVGaYTRH5xiDDyYbJmhW34+rQDYVLI3gh1gl++Bt8LLS/i59/7r3CkUdPMw5S4Eu
jLgLZFAcXxXGDZeplbOQdh/t3vwjZu4vXDa0aeYlBm6dE20YF3/HfweC45EJzqNPtuqF10SFhixe
Sh5Gk8mVg8+hgD25DrnxlBjg9fQXGTEO59zBgztFsNkGS/q4gbL73kpfiO91QLBeas0sDiRjFm6s
B28+yPbNqbgR4DldCzCZCaA+/T1VTgzQbPbd+tgtXz2379k3Pta0mmrPRD6cXhjoHuPfKzKVksDH
xJ1JY7ERlhl2ST5W/X4p0XRP9J5293trTPzEbDISghTuu5HqjtlNpNB7quURUWlWN/vnj+U0cxan
PhhcBEPo8FN0NiSJTezDUGo6PcIukzd1p7eFindRIFzNlo+guGPMqTqvsUZK0DfDGo0mcjtsr9h+
+rJUWxBqcHEwQw/sDJukoKbbt/Qg0pQ5OepBZU5Bu3Sjpghs+IeLfj51GI8/VKHbza2eSF9D223T
GLwT0iTAgDO7K7istzGSH1KRqGvFt5JRKJFrgywWn1UeS+o3mQkwQvT8NYsnYjylZHU0I6rKAkyo
mnCrmud/M04A/Gg3gdbd00xh4hol0VCEx7qT+07dTkqawOFPqwb35UZUSgNVzlMvP+0Ehm3WNRSv
M0BwgdzSnsNYmwOcLWtQWrpF0Nl1LKib+EAVeRyROBJHI+TnavNoUykv6Z/JKfVIET8J8laO2JHZ
hSq1S+2JfMrZjJtWYXHySGDWncDtv7c4tSRdrzG6KbjGUicr5SyxrNvqRJ2fTQsTsNbjj93/fDV2
m9Ty0Xa48xGHj5vSytURJhI+6TpBlfo49xzJgViE9RWzX/FMX3J7pTn97Dz326lzDZNpomPqToXW
Qvfh7jtKt8j74TTOiUoBChzxEdqCnlrAYBj6Cs7mKesEwoNC/iSwKMXFr6gNf+6RA6pvz1QZjO78
kJGemDT23J8eUwvRpTmZd+19IN5ltlrRLV/T9ZpT5Iri6u8I684nsyAk+kLW9drmnVx9ZpvpNX0R
QSR6q62I6h3r9F+YvdV5VGo/k0+SCUB6LHrtAOW/H0gf6wGU1zeErsZg+QcdL8lh2ZCYt0jfSN0o
8MiZEbNWziL8Ai6Dv202oglzWgY6XAWlxD5iKH/Pennu33/pNGTGLwRIOVXh1Ff+d9rBruL7BW6T
HxC9il34/QK/AiSJLNoDwM4GZDadxZKl7gXZUYIL/h1+/4HYcsCfhhbHbo/fAX2WAZpjB7f7Z8QR
FW+31YdtOO9NN4/ZWl6n0l1oEmGBfckmPgdVCr+EqAYF2cofODL4uLczLTq61tZpb2cwgF0JGSkV
WI3MsWD3sOtN7EoedulXPPKT7lPnFEPmITlGfzHVug0ApYpTFcpI7V5HUy7vNBRiT334grYEjXD1
Y8B0e2qeYpYCe82kZu26VfFxoMe/lITPhmOx3vfTEBdCrSGo8nJHJbrjISMTLZvgPq2lPMvHtND5
NcBqD7j13NCLelByzNU10wtB9CAsoAQIqgf9wph25MxGtCtVTgr8s3okH7VhvrB4MrkaBcePiIRH
ngprAnCsA8Q9SUqze27DjJqTzeSgMqCGjKSPVLkExvCDYeRE2YqgrhbsFLdVUr33jfrcq2y6u5jC
clToY8VsAUy/DSR80hg7JXhXtVfy9Ve+9t/3PkLpq392CialtVtlO1PMjjdyVq0mXizcIppxHGE7
SatRcgMlKlJYHSHxf0NKHQrTGuhkOeyDYTsuOPJ/cpwQPg9TL0F3/BaGLP98ppf7UZ+OS98RRgmH
7j1FeZhcSr36vCzTt3BwA4KIGTWgFdycwRuIql2bSweWcPV2wUl4Whr3FeP8j3ywQw2aRpaKt2Y/
J3jVZQOMVD0DuSzGw3j3YyQ2e9gZFKnMKkT/kFksY5gx8Cz9iOs5G9P4nh6B+/EPyXxO6W6laqyD
+RUI0HHfEOk2Stixj4ZkGOvLgNr0m7RKaq1BAq9umPd8XLzfPqgLvVPV/Yt5jBR/jxLQEu0x8D1C
c3mYpc4MaIolTnsrdsFEhGBIq99pd0ZqyuD6MKOlK2+HSu/cxzd0YCEJ9fpej19pH9egJNow3lGP
C/c5fi9iBIrP0fUGq3xuVL9wOPa8fYjD6raV5T0O1SRa5kivXdD4qZQzEr9DLl+K9avz15psIiAa
dJfTKRSe1cruJU/9f9sVaQI8zoLy1W3xw3EB/dRQYBcNWkTv58TdC2fL7l1unqr8ECyHfK10QBFd
mEB45NLwW3pNqe7wnC5ax8gtGbBR0jbG5RGUkhgfOoCvtnf6uRWag9N0R4NdATlp03a4ps2npEzh
ORV624IEODxfCoRM4UQ+B6ROhdW4c6WXA53tMSnAzlvCnsNtRW/tizt4+bGA08ZNiGAjpFWYFvd1
GYQ9ZhyJwcVDKdo18fkvvUjwLUFOAo2c743cyZx14M+V+SNlbPjALwseJ9AkflSn49sLot+Bzwvb
Q9OFAF2I9MrRmM6tf4n1Ngj1ae4RrTUpFg9qKCVHyMjgVv8qmrjdaK0+8hf99A/Sg9wWia886KtL
iQKHzqwlejh2JV/yUWQrxB/wZTvJAQlm1iTAgq0Dgy/5aMj8zMM9rnN+Op30vK+UgfCEe1H/U7AP
7KekYe/0G/U53mGL1pWxt56eEi3ISxJpBpjwEqiqhZ9q4P8Rcu+JAkUoksn3znSGGddGRFfih3sy
uE4Gmk6Ovs0mReM6yy8BnmlELGpMqjf9pyYXk7pFKVKaioUSNRqsH4fPkGprRstHyV3XuNCmZnXn
b0cyG0OzPStQdjL3zsYi8SkpeF4qyWMf9nAvHsAViUZyTGVv7OZWYQmPOjQZEwgdJglruBJkC41/
eTyNei5ZT9b7aws7FMd5K/xtSmhEFzqARknPdaaqOe46Zn7cgSJuRZS+CPyywsP4VYQPRCUgHIdm
dIEvkZfcGCFC3eM0Ex+bTYPNrek3NNgfBnWRJ0vdABXkiMM7W/XW/Is/82SkZBYQ1OvEyM80feLg
z8+VMLcFVZZNyUuCB7UxVuNaKk9I6IVlH9oOMN255aciD375wxbexQ1C5PzI4GrpDlqjl7nVz3yn
UytKWeNQlm4B6xTd27YiRWqbbxDv06NIj/b8Fz+7LtlxcbX8ra7HlvzaCehrlneYqstiunDHJQQT
Hmj5n9tCifxdoxqlHtfRlREZISFglyBL7mkI7TNp1clRGP6nB3nBP25S1cP1cDiWY9QtO590ZA3J
O0zYtMlaeij4QqqNfitwt1LA3tG5apXyqD0/8qrdQ0J/XmzTIALlyyS3iE5xoqEm3xJUspWWpLo7
2Km4I2RBw4b7jcTnFCmSMKYup3e+TYptosNA4ELfazxXwitEc2W7jtwBEMFj5IF34KG9vpCoCelK
zOqtiIC/3OhRlYb6dTwGPqppARfdBDWmaD4QTtWKOl3Ka4/6ZOmZCh+BwXJlzCsgHkEnUVHZ61kA
aOBZg24SLpYFOwjRwNG9QGo80Au0aBBF1HnyEvSOScS039Fp3YOQV1tZXXgJjoCcUipIpYR/5QXH
MsXJ4fTLWZF0yu7HjngAlJv3fazIkyp4h070klXm8p/qKvBFEpi5nhfXQF+rmJBVtU9gUNNFw6nD
2EAhZU/kZjCTPDG9+rHuiBjcF4eWtnxITq6v4AH3dY26k75shmU4hARrbnt0ZQ78WM8oxs9fZRd7
r20Vs+Xlbl5gNI2P7KMisjaE+oF+89tPst4X9C4kVkDBfQFxnXuAWuNvlq0OkUS5+jn5JjEoRHwV
MSYEjxdVWL71zOHhvM3N7XtLmVFvtsBDrpVTcJ0dKIyFrvrGeI8X7iww0ls6g6aExHYSbXU77BPS
VTk/3RkJUgUH7mbVPxmToACWSI5ndBsIS1YcgXmglfMsQftNjrX/jDMQGlWRQOFqb6DFIMA2sMvZ
VT0B4SyeZeht5xrc2oGWr7Tq4K8DUFOJ5lZSxQOyletYjhtYAo0dTTtdeg2ktn+8lpM7UQGALxJd
hv1PTNSeku5GLggVIQq0CQ6pOxXw7uduaZic9cN5M2/7LgeDsMvawPI/ok1SQVh+8CSCkkgX699y
W+X8sdVf5Ksu2b1UpMxWvD/G8j+H9n8DNiI4Vxp0H9kIg0XqthJ+sbQFaL1voxdEggWIlzx06VJZ
JCsEc1ywrSeIrPr3plcVWQAVeRPGPPxGe1t+HtYqSUNegq64cGdiUs+vPRfjqEzge/ogV/MWe1hI
9wrVyR5bhKqyB6dZg1S84Mhto+ePrYll+1Q5xDrp2KsGadRLh5Fzi0WWHHo07ibtqAN4tP+yJu9n
zHtxbOQO7pylSiDHvnwy3otuvtQtQVoA6Vn9Zr1Obi7yeMayWb+K6JmdXXox5j99WKxwLfWAPBz0
UZTkJszj5ecYk7tpBiUa/yF30u2SQj7GkOljzn1DiVDk1sHPIoI6/eXaIJZRtkLT5HV17luw873t
h5irjCg42027/j+RLV0kXPm63FJ8g8pqZoP0kvFxXUChTI8kq+Q02JcKL+QDVkXR8J8zeq69NQND
BjR7X2aB8L462LHFAOAYftI+wA+IticqDkwzw3a+Ks9m8RTQ0sRE3WHpSnKCHcHErWAIhuZ/ZOTA
wrffuQWH0lsd0TUZ3vHlquO+YTcb/nJUlhBi6KkviZk3yknetDm4+SlLHrCaw7bCaYdkGO7m91WS
zZF1qaSE940nPdSZJ+enQJyvY+Q1eQhMOCng7t+5x/IHLLmLrotiDe53Fkml4Br7mgF1um0sBNwp
bme5PapAXcyDN+fsuvo3UwbC+TSwtV8kNuIHllPTtucaPZ73Nz7KLJzsgDYxl1laBluf/3I/oqQj
tNAksUjSn7Om22ZY35OcoHF88LUFsx/kI8Grqx4x//UsjjuFEjV4SVdpbaLWva26FbpSgUwYP/7R
0vBSLWZ6t8P6D3/siUoX3hC3WYFVBU7v06Iyjmr3uLknpE00dqZxgu3WVWrqpaOvIpx4+dc638U+
zQYhx+O1e/wIW0hVai2S/cU50UD+PACgHc6w01Vjv4/r+v9Kjdhhq1ytCyg8jx8lw3eDXojVNzD+
/zvWSOw1Oqn3QSFK+rLcBRE1PfeYb70UHGUpSiwwLZpo2tzoHb9iVlJLQyQcL+ZmBHQiffudYX87
CH9fKOOlI6xhDy0Hznro3fCJKfrSJRtNoWRYfUMym2iUcz6hmLxtS7hRIZL1E0mXauAMAP+Xxnmv
pIHn+GTGUzMnVsIchndPKzuaZMqPiRT3bhcJWhGg9Ub7AIPERhYBRfvljWK9FIOpm8WeVIoUw+ek
rGKHxeTkniRysg5NH98vodYFOcCNw/+k9agv3wgLGwAm2fxn8EfCpWybjzS/bk08OmsTWUPFonE8
FOJ1kzlcpnqamfigOy88C1osS+V9vqnpMAmei8Q6VggVH11IXrJ9hQi/4tNz7qFAU/ZyavOKernH
sFTQGNI8E6NxVkP8ut5//3tlRC3HNDqz8FBw0BoR6r8xZ8NBLTftWkYFUO0De9j7m/qXM0AOpiqe
nArPzpdD4rGc2RiOmikX6WuMt2BL81wTKEFsphahLLgPGeOiJ2bpbj4Y6S/7nUWm1pxBv4fpSHw2
RAf+X7pH3LwWvevfo0C0fGqylngVAfbYMIwUmdLyQ/B+X6pOScyEfL/mShVwpCrdl2BccD40fYRW
a94qKUS33v7SAiJV85AkaenC0F311Ack+mDmZVyzL6zSPldHNVLat21gemXEXwxnVYKu+OhUjeqA
9yMbv/s3vhMySHPISU0ZZLfJhohmePsW8CWDMv4q1lzkHlqt5BtHbESzY68t2LwN8Zp/qduqkFF+
c79uyesz/HzZ7SDgysdGptKdHcVgsjzYuxuLhzrbCoO/v0VOX4U35T3npBVpd8MRflRLe7TU/aLD
dy836S6Uh062vnmHUCyJPC8+BEij2CcmWGqQJhkVN8Jwj9gf+lTPRPLA71xwgF/y8UDkMjyHqAGF
vSxPH/pheoKg4laExuHOb0g+dwzY1GswoQ9wTAO09X95L+uJlP+SRDGyYBqp8fM0WlsQQrodZPq8
1y2H3kCZkft06kOh7r5Df3SSwzujwpJDQNL4C9cLaciouRfnUGtlmcuL7FSAIi3ZWfDzvGYg6pJP
HaxrvA+6csw/Y12urO3GykIN+KnOqkIROX9VOiuh45QY4jnvMhuw5d/Tld8M5B5JiXalyKuW4t4R
uiuEFCSpwJs/W4TiaTNUHrVA3BcRjy9bh634CODvpMeVxVGrLEsNCXLPxMzzUp924LrZVtebyQlL
Xhd3mWdDrSA43zNHY9bkRNx7h7Yt3msnK40PRnjkMygeGWRcHSTg139q37SZDZAOAR2QlJi37o0G
kU38e/ONykzHQjvVSqx6X6UvDvXDJlB3d/3jXV0X8Mpm6YgeNikbOv9+v+yDTiBVY4oionO47Lyc
K59ZV/zRk3BhIgvxodHPxCYxTw+gMtIZlOzBNjl5+QKlyYg9pTuAsTdupzvoNBVEpKzCrmG7dnJo
+hJjDytAhTs6wBTUxQ3eYPT+kF2xbruagTuCat2igJT/EL2kS9LhhWoL9PqktmpzTJANvKcwToml
igTtsGg5CTJKOyOeHYTa4GAFPrpuTTk+2HdxT3ZX1hlwvslRK1zxFBBkOkFbc/QVmFKzzo1QoKx6
zxITByvlRS5hl5uJdugcIaKYI1Vf8aQHncHsvRScib0I4Q2TcQ4oFmzSBoyTcSyBaxXpywcQsXRo
jirtJEmeSf592LpuFNMMb3BcGneELsawqqJW8GrIX504ULfad+Zq3bIImBacGhvtpIJWOzaY4TgH
e4LKfi4GFWRTxxtDGufeMbFWPDBEzuTP+2Isz3NDdYZ5pxExEqowz0KhT82vXJleG6m83n8KozhC
kd8QWAJNZOBJjlExG+706gYD7uxavuiD/NwkPx0P/O6oKFrPrrNvXsRcriHrf0dFz5UEhfK8dEIT
uf4rIjEtqxjYJ64T573YyELsBkABhjms3G/qekZOPz8iPOWU6RFEk/XQYIjdjDiajgU8dRafYOna
5ovL9NCLwAZp1X+FZtJ6j4SzwU9mFQYI5ldT1Jo1TMxY4T/LeRaqPKKX5+t9+NsEXVXQe6pimz6n
m1MxjwsHjNfVPqwNFzmCFFg/TMmSBQSLmv92LltaQkdeHn/HvlhFZEgeiBwAqJ8mpCXQNyqaOQPs
x1+rhbkMNFoBaRNTMLe5wxKL3UbNvL//ruYUzGsk0s+iwj8BXlm9G76+jlBMDyqiwwqDbosKGRyT
94KKpXlFUYrwnnsLsw/E0jWGCpcnH9a9ldcKoLM9eqpzpZItqnS/ZYayWe5QxZWaOWrHrMZy71Bl
Vqn7jQ4lYTkmagZO2B8OZjsDtU6d07DJnnoiga7yuoFXUQePUIZ1LjIuWU0gco+ZqmwFm/5BW3Sq
k4/F/QRO2Sn0vjEhPmdKPlmt0VgPKSMqsuuXDNMpT+ES02W7jWoi/vaNJfVjx0fS6pL6hzLMIqQY
eqpmVma+gRl/D+I/R8/irIfG9b5tY9jG9jJhNbgBDso3KByR9WO3uqPqliB8txSiCALw1UdvK2p4
LemBMXxpLYlQuHWb68DYPE7EL1vr74XNiU6obIuD20GU/Jm7gKCCOz6oqrpVOmqpuV5PQ8cjJB1t
y8Zsh4XnrcgMcqnECBfcUetHd+K0mCqer0eBrMPxq65XuZhpDOwBCgK+nsZGZ0RhgItn0qnAH64N
5S8yykQwwrjZKWHx+aVnOE03TYoIBDKoGtrvyfQwNPjDmpxQcvfFJi6Fly74C/BuiMBOJD/n+lFe
Dv9DXobCqyI/Q5lVImFYWiy49nH5Z7Zbmse6K0vWLW+b0NlpaYEe+SL8GnbZmDfrGAKU/WBkK7fF
ZFWvDrc0725e+klD0aD5VG+RmumNRLu/ge1D88DByh8J8QX+EPE+02uTNfz/wwE/6SbaNhutYsRH
0NB52Zl9gcyYArlNP7sCy7fX3/I7bhTz5TAc8X4MH+iO/jOuQ417/8Y7DCTLptQZuAa+sgGQ4LOy
vJyn7OgKty/ufK+pWIMDdGq11kBWGd/sSEKnckN1jtZZcw+KgwIyVb2zUwAjsQZhbAeN98ChzXq9
1Ru3rCgBFty+/MmX6vMUxHGI9S47+yM4JO5Gx2wBWWgsPpUrZcvLm/bG+hkbnHlYy+I7fwTyORai
vXHzVS9KX+xvu8fKJ/H3pfaYbGZNfsa4/1TxZFGOjjoUkf91x10cXGIcpNZ/m0uPwmZGg0M2EP4A
A9rNERJIzYzB/5NycB/hn6Z7EZIn0TdwDC6H0Xtic8SLQjT8Pwn175ubLrmfCa5QQWHzQjIba3hG
RpZXDdaOX2xPYFfa4VpRtMen9Uk+r8Hw3iQnq/unHS/+j5thouJI/0REpVItYCDCkb09rGvPxpYH
gKr4TFiFCcJlkU/4EdRl0HmokddcLqbbqe+iwf+6FDdd73VCldG0cqRhjsh1m5tNSW/3XfNS2bzi
mXq7B05ijic0I4RnuqwMTGNV3rHaU9/iOMcVOI8TtNn3wzh2da9ghNPU9O4xVsVsNMI7xT1ktKRG
54A3IVA2sQh+cSzr2YjJqOoW745RoU7KH0Zrbea/f3A+XP8ytgMhwE0k3gWPPJ4ZZdbu2zFy3qTA
DTfwDQ9Pgm383ViBSfEuTQtYLY1XRNXODJSbM9wrTaN0Q3jJzl/wmd2J+EcAb0gZ9YV6VWONeby3
3U/6ZRBBXsKbrR5/JhACLolNq3rrIWML6wAuNFKeAhrTgei6rdC790dSNk6vBrsdHGab/wbaHjvv
SyD2/F1NHaXoR47Lq3BcqEVn2UnCC2Clhpn4davXnYEgLl3e+2o7oHWf3BM90STHNVu8pVpXCw9n
k5kC9DVrJHrkfHp9xK4JDtz+P1G+/Il9116cEjK0+R7Hf1X1hro5HtAOs3GVUQt8fDykGcu8Pyi1
DdfFDFizuoPFUEpEO0XDZ65V0alNlXy8dgyj2FYpHVsZZJQop6UGpso8sV9iEJENYb29xucsfzhS
lcBRYwOXU4Z3I8V+j8LY7Yh89fBSkCLB+U4ZAI1SPWguSsQCN5hnPI4yQRL+H2/2UKuhmzVuhXI0
bfF+L8FF6zFHl4fpmgeA/5ydGbhzeQq8hpzQvwxq99G9eYbO4Cqn7SbmhRNToNyw6qN3/ZWiNmIy
c9O9eykiEYMrDI52tBBR7mSoFYNAcsQLm6r976mtTZ/ukCb0K7CNh7V2Y67DUKLTSyqbW4WxcgSZ
BE1wIihp9N2qF5qGJsp7tcbwhFK0K5f4ltiVQUJ9U0+3yMhY028CJSVLIxkgxEsmsvEvZoLtk8hh
mO5mf9bJc4Y3MBChkAnSZS2zQF4nlB8bo9GvmV0dE3d0aRZa8Cc9KdOBQoxcxj2Tuv+pIWKzLNSN
gdLZwAhnXx6rxba/Hcl8rVxTvPcFLPi5vr41q48Sk7ytH2uvFcXVwMdapvyyz0g2ptbMdhhMN8Kp
SclgYVV0wjS0HTT1JxtIuewqc7eSIkjOq68layDGXBi6tLjI8i41CmCQoxPxYKHqw2JcHevd2CTs
yX1JPtHtDr1oz1WNPcsrN0azAWfwd8VVJpcEj9dgp9NK8+VyGu2g3WkuXN4rLw0udEBzThhCOV9a
aSihK+hf/YN28X2G4IWMOlZtfy5aQATulV/qk4h5RQY5YKImSyLE5qvgKOgFBnb+TTqBUgZru2nA
p+AbTVbZXoVsFskw9VLPH0LLRDuXYlpZLz4IRT2rZ6HZZP/0JK3RKgI90U8hKO2JWOtmV1ANOegO
TegvvKAB50xnDCfl9ixVOMQ7O0+EhVf/bmHEygntufr/N16i5MvRSiyYQA7l6xKrfa8pp16a+5t2
I4MrDaGvtUtAOA6YiHXDDb5WXEXies9rdjSBGE51zs7SUelPdd3pxGJ3I6+Cpo53D+XHBROQGtxa
sHNWuqc+ECbOMJAgBQW8xgwxqIxbB8SJOzTKtcDkr7EsmIysy4dYPuNBkFliVQCHFTjtrENBvPRb
yjLFJBM6f/68FR11FoQLSBx0d0E7nwjKt/6e3cUXUfhI1AzpumOrd7Nrhm5bZgfRQTwSM2fMVtZs
cnTlOQ+BLt5Vn2e/aSTKeqNIEW3+5hTrMN4EmUBjeDxF6p51C5/sPPjDIxXRBPF64WUyq/k3jqe5
U6Hspg8su2d200OaBPeJu4jFfha5gSzlRXckQ7aMrJIf7YrB6IxcgPgMv2iYxuizGi4hyHEUV6pg
Ee78pPGJiaAlAlP3CORW/9wnQldgBFDzM5VBsDGWYm/0DmCIF8gRYRomDErOPn1N6QPGVWFDWBjP
9bpMlgWtUHxU/cEl4OcQdgL8JwixGdFLjc/LAY09melBuBp0Els3JwvHWvLPzBLrfVOsO1xY7ANR
xUC4r3iZrwPZXiliUI357jUFcFkDCiG3v09oUAQI/ro4p6p//v1nBaB3eJf4f1V5Bg3tU3hsi2MH
569GpzNZ6QSi24ktILe22bUSAjcBb4Rqg12vqyy/kfF0lT4goKKR7X8G7lD2Cn71t/rBT2uU7Ce0
SwSRkAOHg/y8jFqZBQmWFIhb56esm/bh0bbI/fSZ2boB3Ekbxq4A++XcZooG3Mp+eUw9RKhLjsX+
SGxQDcNCGA1iuyRwAVmf5GxvqEOXSFgKiOH8d9Z+EmF1vK/OYk4dqa3lZyvBFJWANvEE0goImIP1
+0EO7FtgdayZLePWCbEudVlwWJr+ufYL9XN8wow2HZMDeqRVua0TL+oqnX8x+n2g2C+47LdkTuFF
Xsh3ePzw/FrEY4ETEPWUXQhbl7vhwdb4ZbDS9ig3O7Xo5eCUFem1ePpScsd8zzrLg3PFnX0RWkXf
7pOhjL1WL2c5Y/500Yw2XofZrwEh3oEEnsIGsmyq1TvAj6IcD2fDyt26htwyCIix9yIEpUbtjWWT
YyskJtIPI4HefljqiyyxHDd12OceVgfuAITxYlKj9dFurVyIPjB39M2jZu2ad4k9rb4+UEkixJGm
OVvtXuv//BJgQVD4nbRU2U0XRCyXtdeBnsOnRaCHqCshb+M+ULhx2muj6pxoZenjuTW+YI5XE8vl
Bmd4/YiZVyYWbXsDNUcaeKC2PjC8q3i2FkxtMXh6Qqp39lVeDOV/pMPLjZfDs3rhkJeg7ipqCqNe
7q+pheFmsL4CQ/ZYtf7hten/sHT7mFeaVkaXF1H7vJ4b8UQG73wLbnKFKX07dfYb2X55Ue1jrwEP
8ePgBqeyzSbC6BTjiVG2sehAGkn2Dy53G7wtAbqp4pLdS7SDwnpq1O4nujsbdlPK8+ZT6Hg3gmeH
NvcYImbhL9rqfNQN3LJzuVFyWqro+ybqMs0VEFoeAyMGKwZhjPPUuHbKyhboBp8wVd6xVDMjRd2V
vDAA1fd226ZaWPykzjuObjOq9IQEeOhhyprgWIOgvwBuYVWKCvoJckMhdc4ynPMYTdLYsLH7eS8V
O3FPhS+IYYP8si4Wy4LMF1AuGLhUS3VnN9IbOVCYlPznqsUbKVFXTz5mjgBrgUo5yQXKxa7zhvkc
6yoSSOsuKpTvkEqZWpE6kZhCXxKOMapqYtHlbogDlx0bbgPO4UUtg8eiCmuBXpQMQRrh7GUrWkiM
63Cep4468c9HCPhGymdVInAxQCdIzJmcCbg/NHhA0ZvekyKJbiyhwFAnNApJSQWO3uOQlrmQ9r1F
8b8X3Hvh/VBCDpzbjG7tD4OrKtS9XGVRLqWdP3siFfnBvs9tTz2k6AZiQt9l3+0b//NKNDm+QGjE
72AOsGQaqNCbwJApoZ9KiP9WwU41tMCd0PymMlcm4Mab81ZUf3qCSXT5kmq0Z2Wu6u55vCdOTOvt
n+XzkK4nEc8QHGH8k/DRibEStBzvVFMbCJ7iyoUeb8Yg0zgFJqoYxvjH05u4aN4p7ZJEwUcFpO07
WojOlP8Gm7HK3QO9+jQWS7CuSTTii5pxD8sydHjtcyeqqXsVMPHwhnE7rGuf32QwdxxqdEfUhTtx
c3r0H9oXmWtDLZEXPk3eSkumiG8oMZusdUySjG9i952aUMoGEzPxfGio+l5U/b4Vtrly8/38zItX
ZafEpDxDyY1YBeFA2j7MWEdd6v7wMwX/UzBnnz4ToqP7e4JZvxSi+2wDhCNxxpFxVGsEKJvMMlTn
eNrz/ywLfOxNVrPOWJNZIM5MSpE9j0zQfjCOr0MHuHNA1KwgoIEXZGs2F3xpyirGfTNKPaNecI9b
WNtCylZLiCuMNZmVan6tLqN9IPZkdkYKg3OqReRhIRdnNTIu45WeLYZKg2mesyVIIPKQTegLOKgu
KuiFisbc1By/tnHXVw3khUzji3gES+4Nc5OGeAsFQh6gcpPvlXumjQvMBtYe3bx9BuItO7EG0Lyn
XRXPghmiOEudenR4AdPNf65+yoN9GF73IwTmk3zgyForAMa3FY8aeX8WlbBcuiTWDKjD0Qdy678l
EKfpbAzERySJG5l2IHhLRduemdtRHUs5M9D5TTSVztJYEaKDJEnfARwAYW+TkwFz/Ff4BOFLznQD
ymS1MRtbDNHdiyo5lbvEoGUbSpI4e7X2U5mqeg4Rgs3pTYP/euTrqEvYLXN5DBOZ0NuvodlteOaO
MRnVo53n+Mq13R/39c0hyhVHwt+fpgdx10QS7npy932dKo+ogpdLSWaXuH6XAi7j1WcV9xGd0eDm
p41mTaEeE4EsdpuERjhpJasdMVhD7QWV3q5EMh+f/OpM0ydT1zIv8r9oOKB/jqpmdfb0fZDOJcmL
rFiQLXIIiZHo64TuhpLH3nUHzkhpEoLCCNEOQ/hLaYFVlaKsFj6QqSAi4GHj5vUPtc8XZ4S60zVx
gf2f5mqL74VrJ8FnQDn2oMw6K+OvkM6IdUFXi79Rc5v5bnW5BvTzoFOguYxzpEns4TYWvRJDxxut
nNyhG0dZsSIpmxyADhaMPMFGgIoEiu07GVo/kevBjHHumtYSkhpFLJJIjXrLq84n5lPZ5BFsMZ88
TxeKa7B0B7uYcmWuv7a3WmVmS0HNEWubIrmZm6H/dLP83TxeNE5yzZneSEXOqNtA5oJ+v1CYy+Mu
QL2MdM905ey5ORNmoDxjJweFrfUMi0PYbe9JirqGp5sw5XidHPETotfm9y/obwy8d9jMwRLzM6CU
87btjuH/8/QAxTXgoQfrxdkOYyqi3525MydvSVN3+oSsq5eRwujeywAzEZe5LzQ/VKiBaDVZBY8f
44RqVARSAKEkKWh+E+n4OXtaIurAjMGn0BOFh2U4r2NCRmF2Xsw2NrWt79T3/2GMXUYkeUyNBEss
jSOG5LTu7qwVao7xXjFQHM928Q/fkH87oNvZfEHZu4PB7Y4hER/Cg4R5QQRyFWOOCuofFN86inPP
kJcFMwo6z16XJj7eD21+36xWO3enNaq3Jj53Azk9dQaW5jCvPXlre+JasV7GL4Rat7IsjPVTkQgi
IW5bPJWABdE4l5+Tglc5W/jP5kEOEdmAL2wI2oIkk2/I1a5l//riOn20veVjrcBXRGk+52XUyLrf
g5W0gnLIBCayK+Az+VrLigdZ139n2VVWQGT/L41Q5Xj2Md2i4qmdOMY3SUQ+2FkazqnUOa3d2QOL
N+A01w0vdZyZ/78bEy/4x8n8KbAUgaypIzmtsoCsSDmFBQYGlLWHvu77vW+h/E2TXkspIYWDtPml
hDlynPg06m4AWzr3JkpwQ8v/zBSX7Vev4EKwg3eHAnZJEsg0ld/UEC5ivD47ABLAU9Dw/s7PRwrs
DZNlqouxbZO3xNS6KSetxrl4rqRKayI459CCnyEoR7vxg9vZf6QHrd6UTIQuX/0XejtfV0yc9ndK
Y2Ln7R2Cu9G8tBOgxL8+NkIs+2MrJlSnD9YPo751UyRsKx99FHZU5T6oUoHp8FEYhW7YUByNIxNl
PUG3zoeTGlLoJ8iqCtzYcZqKD5xOkADHLCS3EF52aQwqPz4cWa7ADSUzJRyT8LjguOUiurdiSy+4
q1LPoGu6/r4MdfJk3yDjxFcBzgua88dF1f/qQywMDto3w1NsvkXsXhEFlm/FElwKzRXuTQoMK5Bn
Bq7MZULTx+WLyVMQzcgmLvoVyIarjRDgjG8d+DNO9xP0xioZrV3QqVKTRwlWJnEKDmqfqAwVZuc+
PJGcDF6VG97q3ouIjAM9D8bG0r7ewvU0lRS3ggyubvusPbzSWDGjcOX8o+FfD0qLT0gQVB/m2eQl
GQhM7DPabHqaalFUelEab42QZoRzmAVCPVTGikqZTcUB1wLTGkPkWmvsaGW7Wt6ktpzsXTJpA++p
OVrMHn4KLUDL8bwOXDEk/cQWqTrnPI5+tMWHkyhEGx8sZivtrXmYc75qvOIcZsDYIsmlzSXjeAvZ
r84NcsLH4CeOh37MUhVMWai0Tpcpnt7Ym/zLc9OX3H3jsYx+R0j6U71tfkUtKaeOjHdk5q7qhXsl
Fup8S9T6whUDjxcK8Gtpcs5u+B9Mv2Z+F7Sg6eLqC3IXEKMPVAJCiidOmx6FWyMrCGhBEz3J77ks
dd1HUkJQGPJ2BAvg2WGvLo9z2ii1DwVKk8ekFIcEuHtSnuFz0cSJo1nbNsHy08tVWcsS9EID4cNf
6Pn4EMNQqe5RCu7NMZNfsdrLipMV25Vz1ZBQh+ABJiDCeDKE7IzRKzF+8V2ryGU7J9wYLUmJsvhj
8sDcihrlN9aoKaEwagUWggVhBSaYhvJvNxo5ILwI99vy5gsbzLTQMR7Vvmuw9YjigVidgLAisIdI
WFghKSQxxHbf1xzlDPVokTSieCeW+X1tgf3FhJx33hPQMxLIvvvA9hrMwQDwSc5Ze6wiKZZErLB4
bCStO1TkyWXDLUQz57Zidio+1M/stGAQ6wwzGM3Gd6/F87PADFSE+zX1Ix7F5T4zXdS6/d4UHvj3
gbsRRp2nv7TxWzqYa1yLH50tpMfq6oSaxrQOW689GbO/zJcdPc3gzhNx7qg26pGKSwLLh6JEt3dz
b4ZIjKWZKyyPEQeHV47M7bVet5x05GjHmN6tEitHIvTZ1nlG5jJYX/94fsgwQLPYMSF6fMaO2CuK
Kje03IfXp/hV2bB0aV+rHEyC0CvaOU4MZQWKPKwLuOR08ddBlBhHM2Q4PELMmUQPu5y2DeZ52CPe
/8za9xwdRTJ2HDqzwy1wRp9zNo/bcq/3EErqoZE+EZ+78SfMALmCHv3286ropiIRD2rpMp0Gke4/
rccaFudFFdjEAeWv0YGNCoYp3h3wTxBf/MNq16x4qiyAaorQQDS+Y6zKspSz8cz3ffz+FcQawcvS
n+RPm7+Cl0mUaBgu3t82jVymClKHInRq1khqWUTIWDPDn3McOyDBYIEdzDW6w68//m7n/pr1fnzs
WjDXhbc5maw4kDLpC8UQ9jDQvgFwBVG0xeRD6tzBn6mZ4+U6rO7nUGADCtEW3zJYT6OhPvWXA5J8
GBlsidIMS4fC1yMHu5kfW9haOKMjT9WX2X4O8kC7f40A270d2MVmcgDiGURc7AoQdMd0wLsa80i+
BSURjq+46wMw4b1Cqr6MIVRHOsXtfS89ytkCcLupAcB1RvcLVqIhF3jN25hPnNsPmrCgshPqiu/1
aYLTOZ3Dp1av7125ZpolzoCG+qC1FBpMwKkSsbb1nhHsEj0w9OotunE/ZVV8KduOh6ccbnhG5zzX
Wi264Oo0sI4PUhFQtuj6H4JdKtRF9mvmoAQc81TcQm9Htz4rHu5d+uSrDQvisyTpP11i4eVPBOaC
QrTG1v5pPc1TQT9z7rzKfjp/4PJ7ij4QugsdNUOlsmEx0X6uzxzZIEweKUL1CRk56qRCd+tG42sb
N9FbrLSeGwe0bhnNmoEDS5KRnNJC8YJSGWbr8CXAIsz4mrO0E8zLISIcLIc8y4zrlkaUQX3Jq7nK
w/eZhWogjc+kEqDuQgj5CSY6aLZXQ3SMhYqPOriJMQuaAH919lgWVJHa0JT3mVYZ1GAh9xOOZ5Yo
F/m7l7j7h2RBX2z8VR0orqpFzjh3Dx4DUxXVE01DIN1q3G45XAfhcZsWcyvbxMSIFkAuEyqSSuIy
cogT3bYjqRjh+ZbX/gJpOTZHd6szOCCVHQuT6x6x0wnQX4+MsSzNbSL481FD5YNgDTlyG6HTSU5i
VGSKPK2hGumuG+DhKMmg/AOL5nnkj66VN8Ri/SvVs+wyYfWlqx2cDnsPGJGqupXdMKEXRyZXFbqL
QZ6hoPYK2nNOx14XrHDl+8qNXv5YQgbMTvzCVQ8QVB+zkzCQBsIvmEcF29akA9fwP2Uzk75jW6Nu
Re9ih+z5pH9QGJn3zUOcdrZaAZL6S1tInbpe+uqcsJk8Wrbi8RN0dlv0btvaFnq0bOPvCTigaZc5
ZdjjPXe7HRi+0J5FGyMjS7hsAlhnOcJAmMmEgON8UuzwJhwz/C4yoVUGDVPK/BS9sRJtTkXD1k6a
jPswQI5sN93ufoZNqganFfhIsnsvYI0iNFu+2dwHd5s5DkHjeFA8wJW+5iCFsUFpjExAUTiQYx/j
AO8pHOX2IZ2SnMjQ1/600d/srJLBQU5Vv8yNI8Cidu3PRgpdzC95+bhY/7sZCowtzrWAQjEwbyQp
TYZ+EZsXOej1KLTH144PyC+p1wEeSshCKWdqMivTxJTilzUShLxhEkGE8aBNJROru+oomWx+95HW
QqMturgKy9NdRO5iO/ikyTXKlTNXi269STe5gZRv8GwWMbAOunjhUOhw4dO2iUBxVLb88BttDYlD
LYRiCRNkQy+gNritzqs4JnEGrkxkLf1exCuoFoSAy+Ml0Y43bqCYITlaSdKqnrVP60BOxQ7Aiefp
elylbEIfV7+YaFbtUO0kaTx7QNi3rVQJGzO2SC1BqUdNcRePbT15wYdAXRqKTddPKhDiFCPi8KZJ
4Rl3YJLu/IzovwtknBuPGJQW7GK82Wj8zLs74To4smKZmOiQJTYULvvADNT/XWyeu2tBJvqsvUeF
tMmYsAixj0naRPlhO5MlfLgLEps65En4fcBEMhP6/OaAIShp7RmxZgKai0t20P1J3lvIsAwly3tP
slFqkzxA2/dvWwRzxD1TJxgUTk96JVeCmJTUqn4oLYRVDZhEgq3nyUw3GeexjhDy0vmMNjOj1pe/
tbEOXHKHMhBX2DnIxsHesm+8MQ36IGSu+yORCfQAe5pfFQWGpjFKJ0gzy1tq1/O5Lpu+4XyCiOUj
9OlOCEU4rcYBGi5BzUiQDewaue6CqPgiO7GRBrIxLUpQLRZBZ/y9lImR2BZy2zDrFXk9jXDiMms3
kJsSgzv/H3QkZMpBY0Sjv0XIvrd3nsgbinH8ZYmp/a7mu7L6fS8r4L/iDGyfS3yBCvO4hfIL2MCG
ZC5kCXyZi93+Sw+yrTrwyEj1GFVP3AhyzApuJjLU7Nni58usGfiCenBVZH2/wCHlwQggAUNffvJ0
Zg8mMfhaNx5sRk1hzMHjkmVio1abscN5oeqLtnqXRoRGcBwCUIvuY2HIedxTfgf2PGba+fxxmNPK
lMQowFy+be3Zskek2Xo5n9cuMH7w1bOr9yAH7wS+9acIwQndiHL3r3pidqA4ONXGUwL+9mmB2LAq
QoKwXi0Hpq6CI6O0WH2/QZD3a16DbP+v2QMTBz3xOqczBn1kkK+hsr0gyQGTuSouFGI+nPwEKpg5
H7q/UAR1lSehg3q2D/C112Gc5m22A7RvTRAbUrE/nKPfTVMGWxjTJIW4oAcVo/rmeE+gBhc6XKle
ru7C/+h6Fwi08L/IkoTBnyz4DKeq5GUjeIMzwWfHuXdB4RP93tEqovV0dfVeOzPgG/l7Ue/OWuoY
YuCA7mtSUvcN1CJ8jU6BoO+kFpB/CElopDqpHh7IJm7mAdH1n28caNmDaRgbxoVD03MzQZHpXBkQ
he2qi6CFZkgmbADmygRFbCM0wOON2pNPFxSGJhYSKcng8Wnpmb/dgtiMgwYqZtoRIN5fDIUkvZNG
LHvuoh6lb2sPmVlCpFwlysaqVnYoR7W04Ne8LbTzFoh6jADSinAyOkd6AvHf9GIfyNOkRu+9PWa7
NL/jjcirIPd3YrcvuDwgETtFSsDxyVtNL0z1+MxJaiyLosDB6YQ5jG/OV4Vdj8ZBjML8+7MrCy6O
71K+SXeMJ/P8zx4TLdGxQgkxhIQb6mCOcKeoZJgoBJv8Chs6WxfBu42DPUeA2bnEHeBlP9kLMb9G
RRA63+h/18/X78lAMRJKwaWA1MnZMmTxrq/+rJdPvwXOJud+L+uPVcaD3poKA9R9Lun6HBRdYoMX
PF/5vnmptsUUtjZH1ENM87LPtQl/606XjQi4vTNOd4HF+58h+3yXVCOB76NxymONH1Ksv/Xh1wsF
izKGi9cAoDHTbMFL9KjuDFB7ZsoDJKzAnzo5qPQu8wNGnguYBL6bT11cdvK52uIdepKFPXeNdpyq
k/r1iBjSESfxuN2PGLo98WUgo+PieMbpSJekHqLOiKc4qEl9TrlP1KlJfL0FVpLBIIL7aklw6WSi
tXRBnJwtKSkOeKJwqhp3R/J7gWqqlNIRLmzLRXhFG/NixX1HRNcNfnev2Nq07tNd5uFtxjU915g8
lorZTzRjTLuIJYurRpGdqJ/gdJI+K5mXLjwtCV2fuEjiUerbh1gSR0dblxfVPuRe+tKexnjHXbNk
pYQTd7UWykbwL+WnwvwREQaqbqjsorHyAECEAqnir0+kHhSHzf8g0zWeddMP7ljkZWBIdEkNbvBk
09qY9Gu9pMRrx98t3A6bW1sC1BTHyQjDR8uhX/8CEMETFQ7XLIKmWcLwJSpZES6RdRF7uaI0G3C9
BUAQxu1qQC7oC4NPiwslBMnFSsHKBQp6D6Ew4XUSUOqa75PUdJj6zTaXKS60V2JLarMK50fS+paF
s4JUh7L3baEQLag6UfZbb6yPswCv/sc8MYSC2lCp3VRsBm3cG30ICjpzlIaFRj60Nk5Y19Nel8MT
r13u+0+uoxK0w5S1mjVNNsyGHPJVzupOxqCO2hD7c3+PX7Q7keQ901SalFNS9w8bAA1HI0wachJ1
qe9Qb7arOu4NU5x1fTl2uL5aw/XFqIdtke9E9i1UG3Elt645GdQewcJ3Mj3yPOdhvnuWWruKy5ey
KSR2rA1VYTkfTn5KpOVw3hLj0jdel3IGIfTUDMRUe48OHWHMNfQypj7xYkgQwJaeChjGxYq6ucTN
DhfCDhtPC5BXQHubxJRb6OpCl8e09eS9S+mnPzAlA4QouUsOUgvKYqy/2ySjNloCZDzNM1XC2UMD
ndXQB+ruEJo+N+U0dhtzQ1ZbUeTRWg0eaEKx1yZGxd6TOYgE89N1NHTLfVcsRHl5UpD/mDxaZ/gf
DkT4URNG1CWCtnVXS6uCDqRjpsWOXzYCsV8+gkJJR6uiYch1eXTQOHYBO4W0bhnnXJsvuWAanp0C
xZMgWI43WNH2H2Vo2nEhs+elTm1/F9pAAts9OhlBgjfNQT+LYv6YMes4ZYsttbu3hsByF0pMrlfA
vDGig9jOq1uFSRSKkUIbWbqeGk73ET+NuXnnMkyHb4mFTpphEkaQhS8c+5fEIvFquXfgWMs7XMOx
T/ytF644YZ1QiJbGS20w49Tb+CPso1rRaFNMujpdJqf3Ar9AIZDt/ljtx2lio/UZQ3PP1G8U/YkA
nRMBBQXY1wd8+tiRjhbYo5cP8/GK94k885s8/2OEKRmhd/FgKjFiNsqOYY37VYmgFJg80l/IzHUF
LmUdkYV8LYiKMSMdFE6LnB9zLCwATHMB9L2MRatazeEIhG68zoRGHAUlV4iNpAITFklQMdKHDzDr
2WpekcJPNzLVtSdcwsZKeBrz2u5+df3USxcpeqMuxnI+50oAZ7DbUF9xWA3kxDPhV9RqbNmPOD6E
ZKJUT/Kzc491v9bDI25/eaPQRKb7BSyn5c24a3/q1nvMmqBuW9I4pFchUJ38LyrGEwuqZrhhuUyK
8Ij1mxUwVPJpNyoVEZN/b+Urxw6ymmWEhpEv7+ooVaXeu1sKXFIbSNMEFgqmPSnBr6jT1oZZwSLj
rrAvVBXvavjWbFcqEnhPtqBUpPk/D/hqU0eLUyUvHN4RxW8ao87MSU+e/ggpE0KSr6v2nbI3ztyW
/qt4c3xHo3jMmacyo8CFT93VKBTZkX9zqrKD0qVgeJmGuTxiuOsghBL+81mXhvGlHPFO/nRXhTf9
IiM9SSHS8W2pm17f4Y5r5I+47o3VatRJbthJXK2qQN+eQYyRCdWQQh13RzlnNlwBnHprsCYyISyx
yv2wrzkm9cRdX0sawogEasMxqpKFWaTuQRcMWZVRHqp8pz+AYA1GB16tpq23N4IsulT21eMkhhui
2LYgCYPZp52/STnxbSLqM4QJH4FIE8vHryZFn+hNST14/C4DlDIYIapq0h4V+9Jxe+SqHMZulQP5
vr86KjWAqDmGZROaZWNkVg0pKIe1Rg9XU+8vGlpqMrBsTIQ7JBQI78kdAFatutjvixvSsTNaHEFk
3FcNGpK26BeueFO1v4CmUqLQ/H4Tv92I2/aqyjADw5fMycRIP2Q5j+4m6tF7klw43FX1vP5Sd2Z3
SqroHRb7Up5UZoLwRe6qEvy5bJC3cGbXTHhdQ9n5I6k4wVToSOv5bRVNGW6qK0IaOACcYlHGGYYX
aG4mOWuoRQFP7be6e7mJjfMXIy9WwNIE5e+kAn+5sl1edTwUjbCSdeCNgN5Pw4BAXjXB/OiYssis
aTmQRTu8FfRWIQGKfZ3afj9RwOiDrFLf4UQcBor/fZ51o9F7scRxXiXjVwUnXaaHrIzncNIWD9J7
iSzhf4v36P991Ed0vPlPx0mxphs+Tr4Xwj+rCD9yM9CsnPlMyS7L4DkioTgVQS/CCR6j0seu6Ltg
pjBMDS92B/32JASpM7LurNgxGORqGGhfXbm42AUSZpAUgGWgFppdrQIuNv8mY8VzflrYwRoduwyF
9uGl82BfOBrUlhrYCw6DltMS/GMiiYAdHrlBQnk22ztLQXNSeXJfG3C6qBJzABU2fjEH+eCc+iZA
Z/e0clES487FzwKya2VqUHklm0GLiM0DfgzFotsKuKsDMUpPJoa4U44G9hM7G+ms+c5lKrbeuUT6
oQijtqVa40pjxou2oXlRN90Nm/6hfQVmGRfsffNWu39IIly3LqDmT1yhd5U2435KS5+KojmI5g1L
Y77csUMz59MbbYHf/7L6sjQ0ybCBJ06VdsTb8Ua7Lc2jrchUxDAL61to7jEvHhjC2iqzHlQ9EKAY
EDefFCjru6Ief4Tg0RUNCkWEesB7BySlKuuuXOacsVcdjv3jtRA/6YqHXxncb0NrS1TpGh18fBnY
EOGlj2mYrjeTQQcc299DOwt7d2yc699fovJnXEK91LLmVcpLKZ74PrRsDcpaMgh/3fms6lQWusk9
b2kIeMdwey8asnaQAV9+LE71wDn6/fNuNpgxw1eRK2Opl2NUkUPfbWktkgzLNMRAeqtfydc8mS+5
CgAUbne/shKf0ueXxqig2/1ACzbZdZSOwblAE+a2Htrb6tl45xGMZ7fjsUHosh/I17WQoBM5mZpU
5tibQtJnxn2k2ikUMfXQgsTt82c4llN8dK79bZk0hxKjPhLcQpcFVbGOxHALQuMepVEpnUQPf1h9
i/bPO70WtdasKn2+F+IcQranVgCwrWEmJeKrZmUihZAmj4TpjduPYVoLL+dbcV8KqxLptD94yS5Q
KK3pMrJkvEPwJ2fR5kEfDMUuagowXGUJtZfBq3APqApkI6/+zFoDXo3qEXIwm/EIAUdknFqz2i67
HkEkMdKx2hDAKtIbJFYzkuAOOzrL5qqU2XPXtW2MfO54aob7pdrMoMjCZHY6OuC8ErIpVFrAFr3i
1VFJUMVyxJ/QDOD9Zu/Adi+Sa9y+aLEUJPcGmB35582nA86pAIxZ6DP/4mbPrMjCO2OxnO20dueK
u6Cg7VObABJirXT7pAvQJLL+gMqm7kvSheiR2APTAMeWu0jMKDVtqMAOQWWnCV/3ZLcgQK0OKklG
DkpFFW/fi1ozFgGsdHasq8NEqXGzGu3kh7/peYFyojNKy22FztkDjZN5Dr5l5qlBpVwjXNvsUqJa
thZKY+VhDKIbofA0gUx/s3dzOb8x2rvDVdNTGu5ugokHniuLBbr9Sb1bRUxFwp4UlN2zydpMS9lX
0Rj89t8kCSbi7zzp5Cfx1rIMFKJ0PYP3Ltzsvgd46DQzL913zdDhiV2qccVStKqUhzoD9wx4jiED
0c7TmGmavVuCZ5fLEneQo166bB/EZl95RHwoF9GTgN8leSDCOMGWT8v3xirJVLQkjyvFR4SJyyHS
uynFmAcfqOX4sJS3RpIAhiYD0Hu6gEKlFFyFS7XX2kCZU05YqwCZKYMjIVIxw3hm9ph7GMlDn+DQ
iWEZxufkrz4yGZBsQhd30Q6+AHkh/Ajwz4rWoy+/cfrXO6DrVkgjOBLMoxShz03DgWTQPLy8IJbC
pDOxp9Sb3pdgNu0cTcdfcxZXR31Kd/kRbm1H+3o6ladjB4hYf59BqHDR1iV+WW6F+m0yDw4vSD63
cJvXYY9WYh1TDptxmATMh9xKEwZ705DpHy9Ti6aX/XAF9kk164OTjZHriIKYER10cfN4M6zBPAQc
t/C0xBBmQ8bXBkfG+kjpk0iyIvw9BzA4I+ofXQ+rdwfwVuvs4kQhl1PzskcRCMRb4BY2WR141Ajr
G0YxpBd9fahbefYeLzvIL+78nWVtofnYiod/TwuBdATP3PYm8KFL4FvaNQkjulIR7qTL2nVywyN1
a2hef0SEJf+qLh7UrpVtb9wqPLpjZymuL07x6STHQogEW1XuxyvDK0j9jrQv5TeStzbPUE4QJ9OC
TsBs5kR0HO4I8ZHLYImsWqhiQpL5/I+cPKb6105ifFRqtoFdhliaEJqwerYYCYvQKINKqvZnQ7+/
ofCfB/cQb1FmApwMPDatpTFVGGali2CRTjPe6WE7WDZNXtHu122FF0XKR6vR44EYffpX2FcfeJnk
K5JNJH0Eq9wKSxwX8lPOaYOVaQFESvkn9DCC6ppBa5xsRNZ6mu5WH1veEz3KlTlChhDOFJ7OvM4L
AP9UCiCh3g12OcVLruxVveKxqTpvCl4A7lpOT2q4kwBtdEriORbDCdgwagG6C3LSOCg+BvZTVcI2
g8vp0b+KvTTLoq+882X2Zmh0K0/DnOPMAe57xzLeoDE/QpdvCpHSG429M6iaIG40Uk6Pr+VQFPNU
I64Z4oSIJgZVoFMBZAY2afmaZ6Fl4vrLOs7QFRHzelAdmUg+tw0B2fMfSkYTLW6097dp0tmIAjFS
GmW5cTQkXoFCJamzg9/wBVl+6Xlrthr5oFi+AUzNqoxLkHOWoKQayfKeITdSVzB6qR2Bxb5zo7Ad
K/aYtrJD/k0ysyEOsVaUdUYSox0t4OW85IDLkFJbR3Vz0ywVjAf3jrL/Lu3QfS+HjVbiCmXqAlNU
zUQVrRUx7adzWulhSJzcW/QhUtzem66GHCZLI/XoR2brpM6rD/0JMuW3S2syZdx28CZ6EfSvkcrR
Q97hPGAu5wnZ529rpgO2m4kDnhJT2BqAkJkqklL1ZQTJnV5rtcZEWKJQuCV2TzJDV++d+RdA0IUz
mtWce/dLfvZtYMQMAOA6LuAHzOrvWiLw9PHDUNKJLOIcyhgAGBUpG98NEdKFqKLSBTUtO9kkrYZI
wCCduMeP/ww7b31caXqJE6o3mf+csT5zI6MdFDNrhYyF9JAOS8ccdWcba38uzygK8XiyKQIiwIM/
dULYJrGVdXRPEbbSSLTHSAgY/KZYb9wQQ97gLHCrFeuWeyzcWreAYS6txsS7xJVqARt0N7FI6jLG
/xW9AskSyP6IYILJNG2kH3hIqDqRqXFhhU9ew9Xtm1c3KdsSuVuIjWp0h6BT7E3ybRhhPNsL2njn
CqA3Z+XZQHTtEpGOx5AbsaCGbzt+fiZ5GtXna3UTwTZy9dr4N96+Ci1PzPO4HLjj30oTLWydioH+
5zMasR9qCxslTcterO5/KsXZ3kG6kY0GTLxwsrjg0UiWckcmTH4Iw8mYHtBUnBX4bik65kaUT196
RNhrsEZ4EiSvLXJl9TGcdWlFr5mIjeegNIkZQEdtCjOoDzIxP+Q172jUX2ChcUzhx+v90tU/bUot
iDA0uokDUluGUNOYDDf9fbWHzEMlYIlcks4plJ92Kj/h56T6rOShSVKsJvAqfJkd/zCyMkwUZh5M
p7/jvaRJO5Q9PhlxjUku2cC56B6pBHbpoTY7dcu4rr5sVjKRB3MyFjuAFvRAWEH9E7HivPQSapJf
QSuMRYy4OcCTep9kLAzqWOOJBJPl+gp3V06IylM3qnMpSf7wGxwTUdn/TIUZHV+uYASAkqt8492m
YD+pbmkKqt3W9evWURnkfiZPTQRrFtCypy5shJKH7L3wIokyUDX55T7nr740dNMKwQEqQIspK/Oz
HxynY4/loIOpB0loHiS1s7GlQ+6bFO7RhI0ZG7rclzrSn0MK0/VCHpj0Jz0m69jCIEYJ4twsw3OC
QpqVtcY6gGf5OIOFS85VgOUuM+nkPLgHK/7+JqGPQjSJdMitrjROtsuvK/ptwsMTx2SGtivQDuPX
adi6cvmKt8pYB1rqH2aseAsoFV1clYMDH8/1olUvHs6CO9oJe4xou8z+7zxhQ07GIu19wEq4vyEk
OQrWRzpSXoquIJ3paHWJWBFno8v1l5vsGSR67/+IiCwyinHJ90NhfMdusRKz8uOOQjZoZTRfq+hh
0i40YGuMQlkUo0gFtG2RgthU4fyKqhO3jNEuyx84rkzOUJN9as/KbkTgtbra6LJy7otKFwkkNGXR
6bAwwv5cSN10Tl/D/L/CMOHVa5FZoWOD+OX6q18IlyfPuH61LIScXaqjEWhkaFCo3yzxA9tjexwd
6u/6CIQ+R2pRNsahaBm7uAGY5Bm9Wb7P4xi53me1dXLomaEyQB+pApben3cPKcvYrUDr3GSLQsa6
YsKAWp5j0y0oE8/8Qa15uxzZWjtbekWuljIiNfLk5zMaBookChxtnhHn0R3flOzPI4nqwdQbe5EJ
dGhE1GVObgkyXAxN6nJ/w+f5B9sJcVv10Hvb+gyyD/8m1IairBEBzAU6O0oYOezQ0m7ksEEVAwyP
lKmz3qBhIOUhMHWpRAmuE9ZdxMBqrVj1zp8SDLJ40kU3nWQsEIO6jct5XZS3D79ahsaabJ6MANZ5
cCnoF+PXJ2GlLY13N55auTvq+n2emgj0Y9L6HhbpelW7JOdFWWQpT1Qnyx4IJ8lbZghH6OA2k2H3
J/8vbhAU2M2QNaMN7VrjXBesh84+d7T2S8W+cbQjbPdwfp2pJ/hXOMjXBJHzIzqF6+xLH+Qdw+LK
ydE5W/r/lRt3dXF0MkdYxYafOiVlOVsdXmWpmS2+tLs8BosyS/XTMFqrSxJRV0FYA9i1HomQKt6B
SzY69E7HFi68/cds7JIMcFPuWmd51DZ6zLQRlUq3XoPIAIBqZ99FDfe/cnNEWRoMPmMg4V+g5Jm5
RpABQMRaMHRIGAVwy7qu/IWV31QxgOeUqrkTVMkSIlriXNv2/zQVKyzkrYbDRne/wHxfA9tFTIm6
WPiCcRw0ED/ds+xHGtbDEWgTzcZNeo5/SPebdcqkacriTCcXRpvcljhmNpahIP2VaOVbG7uR9WC8
vIhLwa8gxOsHzoQHOm+STjGklrVUsIu0rQXCww6U1DkCMpz0hSKXS1MEpUXSE2TdA/0LCQnBAhqS
6CXy/e42btmx4shkqw38WRv1VC8gHXgx1hot2Ch7W9UY1f8om61fm5t2rfRtQQOUQoskAGKZhn34
GF3U0BnWrLh2F5dio8yuK9y9iKcXW5djBW924v6Mp1NWoy9LXTjnRRX9N86nfxvxdbU1ZdK+7IAS
z6B79h0mFGkFYIkPdcIUBb1nnafE8t5xkXebrxms1Yf+WFB54l6k2u1qc046yUP0LwFodGUHe6ai
leC3ZFckQGB7ca2RYLaWxeIl9QgkAQRE8xKwcsJCyVBf1X8tJkmj5S0GfNrR5pRmr3sTxqBYlrxw
4muF1PjWVRyCDxNSCBlW6pooUdYlsbRwVu/Q7WN42JY85arQP5V6Xe7jxQsPTN81LQfbzn/nOdLC
c6llxU7zJ/vDniF03F8XQdGkXjplB+03AqkiSaLspsDWhVTK1UZ2J9ydUGrCfREgwpaMnbPA/Tt5
ioSzwAeXZXCFZyF8yMnj3pZ29gM0uyOIWRAb2LO/0CYoeVK9eWs1RIJJMqWcPdF2+FMTxZwErDW/
yOAn7Sxt57l92uUOmMFS4f60X7R+P84sNmwKh+zcREZE1YGgpqBpkevE/03t5CMxzbM5R5n12Dk4
aNvLMu/vNw/bz5wN++CY762yIZFEEEndm2NBuieEpnLe2DdM5+KnissIYloe9YXm7/Mcwefh/oHP
l29587rRcn4e+Od0S8DOHXkSwVzv99LhGb6OTu5GmWKUyg6lJh3wVz0Z8z2ICxP0s4JjK5kzZqLK
PLFqWpATC6OEiCPBAJTru3qgH7zzcb7A/wrUqke5JKp1z7ak36Kz18HY3jNwg+OBnqdOGPhG9m/Z
O3nlgpJxJQjjTn6haqwPgN1BvS7+5sYj3IjRcDHYXipsbSoxEmcYN0+e5znHYPEWD1UlROguSi+u
O9+YH/9M6acmzaSytZFQaIWBnUR5kbSWkZPs1L6DlOmXHg1fLqOd3kqjEXYWgqfIEaGYUZz0AEbj
b/MJ2BVMR5KAN27YsamnELR9qf+wxw6eJPh7RpTv6mEbtM/GVGQOXr3onM6tV/s241TAE5ImRAit
Ruwk2/s9TqybHyGNnADV9icX8octhenEX8TkJwfC/c2681cAtCjVG2V+M8lEwoRUxIFrR/uYdx5Q
yIzmfygMN0gObOANH3xwzwbU2c5YaB2Z+dDQ3d2O/GPvtworFnlQ1STgRb2f8j2nP6Vwm4FpyKc0
qxQaLbtlPKJhLXPV2+750OHGlPjdm+JYYeVoLjq6JAdLCtiNftl8s2BbiUAxAbkLu0XVxJHGbZJr
t+SLsth3uVgA1HY2rnsb6cS8LGkYayzj4nSpMRH3UwhhDtQquzq9yAR8q7Pj37KY37Bg8euAyiq1
aJOP/Et0tN5j3FHnkAueQON1ewM1rDiqDswc8vO7CJcSvR5ouXqdkmKj9MZKqP6iK5lfcAN5CY4b
PKPvvDle+kJXaBEl+8SPnX4VpHgEh2TQf19eGLCPTxwzVtTi3NgKKlto4hGsOzS0NeMr3ClMadz1
OArgu0IPv+6QlyRgA4qvgrkXAzQbx7a744ZmQJG/GfAGhNEyHpcg6K6C9TW8SdpSKMnxF/K9AcL/
YDdb7iug7HpBPK/iuil0DGz5xmbgT4fInCqTzA+JIAUwP3r25gRe930tlk3TX5wyqDeXPNyjaNmt
XC5zenyX5TWPqUXrPlhucby23GjJ6k/6tU/K8PRWpb0wiBHwMIIVR2RHaWT667DLaii+p0Rwe4/H
zMFIzQfGGIo+3AwyDnJBE0EkzQVdIBnVgrg/Ig63M15ID7pWzo87EdtudqBylTMFEw6HWpZuJ4HI
TtyQBNl/B/2JVHb4iIZha+GFq/H/dP+iwyGvQjh0tvtKURRpdxxg3UmFtCgNLl6wM3XCkhsl0/Ih
UiH5aw/5k6afKjalg1WZnQv+rFSr7APeJB40Zt53oKAM5XYKYy0foypgs3iXQ36r2UPKkSfrXP6M
H0++u8584+EMqPiGu/Uow/w8rBBi3bMiqRuxhVNwIFz8i9ZP2ilAF0CcaTMQ85NCn4kK982o+C17
OL2/KK+tAJQOxsGzHDnIzVv/sE3thKu/k/Tn3fpKJa12DLnumIzcoCswrE77N4duYWV0o/LG83bf
+QEs2cWiXgTYFMxHWwcXfV/JAddGYuGgpkfSo8h56ahCWdigQgAzWgHkevK6pzW6NhOrQd9TOXdH
Hy66WMhjz+1+L6EtqYmnKfvGgDl/TcNh5vTl8vHLGQr1kcNyI/tKerCEo5UNg1sVLWiOwGXDmNG4
5wTdbU48gnsNH3K1A/5uMSKA3wqrGLmKFd/JpvjhAe+PIGsOPVBGtIUjnXrOMnEioDika3TyuxJn
ggmf8T3AMG4lUnEl83DRKHCZlz1jHtDD78oUVK2YwSzoHg3ZScTi5zpPXMSxqSTE1u6zwMlReDxu
gYQHbd/cYvfASaHTxb/KVKpbxv5pOfe3nwrs7XgPfSZeYBfPOR3iXy/FLHluCVR8PxAeIdQ14q5o
2AaH3veIcsqEGU9peAF20bIs3EuhGjkfCpBLPHzcF0NjaQmaA4tK3LOVdVUzY4EJCetSkTuQJEho
/g+P9EoLtkbmptQ+ajjuS481iIuE8jAAy6sBRpmvqRDhFBWElulin+iRyKZhMuXm1Eqhov22kodj
2wZ6jcp2a7f+yzAwX3OC30b/7wg3XaHQ9SOUBRouD+WGMGq8gxYZ62X3/gYqaU0n5thNwZUoNDUp
9NmWBjevfC8wc5IsjYB9dc3Y3ODhf8o4OgH2bg2pWjXUT4dLBsEew6+Df9yKR09sEcRgrtsy/Tu2
LGjccSr3zjDRAnAJ3vYJTPupsX5gWGAzdNLD1YPS8fCFUGidDknE18Zs7WH5dAT51lW0G5itBS9y
PpIy6D3YjOsDXNwmHY3c3yfbar4qDnB12AcqzdXasZwWKly0WvAEblDcS/G3d+LE+iJ7RC6Xb4oZ
BYxRi7cPBsq9GO/pwmbX0MKxHxjB+wuVZKZFltxjIWKYWnRx9zFH72sEPHexfC2HGdy8/Uwj9hqt
wA3C0fiyZogjtXiX0So/qBtEKVpEBwmPswVxZb/cloK8oAplyYoItUsKBZfvlnzq6WP3B0UG+thl
SWsY8Muq4pO2iaWDOT5dW+MKddKl8ICTqw06D5Vl4QpXwXgryMdvY+SsOodZAQW8y09MRMStDCge
CplWLhPlJci9nrFHjrigMy3pOQf0DBRKu4eNkn3TIwuQMNczOkbZNADlcKDl4kJBrTuj57vN+LnP
8JaxgUAN4qoydEGQAtHwHA8PofFbiNRMPv94pnK5yiiGHyZDy8lMnHGJkCvkGO7wr8x22suAXFqL
aQ8MeX9SmXwtexy89bF/A+jl5rlVq4UhykuURIXfMEOhh2bbKFqk4irI85woZM3tcsgiZjK+patD
hxdfB5wAfPamR4UwyI4Hy+TDnKCojpvlXs/aDxgl8B1jS9fAnsUcnCeBHennmilQw3l3lrP9+8mU
uZ5O1EgAW2x7YlzkDNBeZxZaVk1XwKxdo3jcYlXlIsVRjHKtjqJ7Mu+73EVaVx6uVGO6+CA+8DI+
yq2jFVGYMT8lwVVFmjCg+pO4m812I0YTkw5JfF7HsG8LN6/shdAefPIrPCV33+t0am80gxzzK6um
+xJm2z7NNKYd5+FNno1dqpiJY41xxHlRB+vkCPALOtzM+GzGWbvQ2vp3Ly3gxvi0GDDnbOqYyXkv
ettFiTrjfoBqUuX0Rkksl+mrY63jvQlxoMHoR908tfZisd6P0u74oyRYT+i6dhCo7iCzRKF61FEj
x4BsxKVpQ3G3oUmYfukNLno7p3NpPT3RTai/Mkq6mzpLkP3FhuBongDyZd7RJ8sosop/AvlgbZ1g
SLhzi2Ilte1rZYaDki5Z7Mq23tM7MZmytFPE5Bl+J9Jk/cLexlijoq7rse/3g4jPuHHaa5RZij3E
9YwfbWWcm9IaTcvxUep0LGCh1lveenTr0s6i15tbgvMcS8EiHzw9mEvfg7LW+iXjMWL+M+mT2n8s
g4iTBo5sL/ELpRiQqXl3b+2Izo7iFQyXLW5vPtLd+OfArr7ppbyoLCByIyfe8jE+Qllk7F990VfO
QoreYFgsDlu3WooQE+0Y4GcA1EuD8TZj9220pXDPr9FXhs96k3ulv+Dw/6TodetVt/KBA1S6NHEB
xbAyeYjwF/kwhI9Q32m7YAkEwby7YVmyX1RQLlobkuxho92Ldbt834BQY+uI7zny7pzgMeHfnC2S
Zz4qJQ3rKSKVkLXzUul6I/KDHbygsPiMOB54Mta8WD3EaHG2hojD3zTTzU4wltDSa+1/1ybnb+cZ
EvDwVdnP1w9Tz61WI2jUiaAgdxsyZupUpjuSsJpoLejfPsaBGDfxNz76UKQiz8AOTA6BNlZB8HQW
Ceth5QWXscUIwV5cf/P1+fpiWwR8vwjOHG+SyL5NGgeiR+jL1WaLVkcfKichudqkDbphnq7mhOAM
/yzw8u9HtifvOSmcgw9ql1e1Az6cveK0QKqO0vkulLVdOADOL9OymapSqk60CzKmxyLSs5w2A58T
LGHXJGitQuDH/y4rTNmjSnDKTu1WodV4s4IZK8BuvF8zOAbpR5JCcUZg/qArZPnFck1bWS9JQw7t
7lKE4CtYonp9HpSJYaPbrTaxaDNeU/O9cVsNYlp3cU9YrD2ZaoV5tx9lxCfbF4ZnCJg28F5KfbwR
maAIHI4i+dphg6bqoQZf5K2a3O3hYeduRBWKRl5MGhCMB6o2rdetKt+X2XcxqlPYe61XHj61wNsK
FaHcKMm8nNHwUsC3qbaNF9ebmWu+WZ5r+JUUYbQJf6VL+3P31y0QafkdY5mGFCJFnBKyD/nvJgbD
m8iJ6s2Yx74a7FYrTTlhDn7sbCmXeKXkFNa3AiX4px4VBziPiSNewuUaBOkD/2GRpZuRtDsDiiiq
b192Xrh+NAThWLKMVaDOalnD2GTH1odFEItxOXZdUJNeTq/GoO/roNYc1D9OWBQSPzWrYqPY3GYR
yhvRYuXuD41BWLOLTWs7pJAS/EoO1AgfDMqWkpVY4flSad9sOzTTT2gHmkz4nZpiZsgK4xYLMaYy
vvxQIUr3R+h4JVxf1X8CfnSWcTDtCmRcHpakY6k+3DQNQbVseQn1whhqTHd9PCTqAj+bUhxC0jlf
puMuMxA4XF9yqRCsBocTGeBUaxN5r5mk3AjjzgjstBC91xXAOK8fVQIPurJacLIeU0eFKZJNYGUp
ADiZ/84jsWxopEMaNiHuGD+dECQpxrMv3qfQkHahO6e54xh5zlLXJIrcDVbag/O3gijUahtMEJv6
WnzkJk42vf69kgaKautTLJNfOgmD6ZWcmG2ntTS6SXQALkx5wx8tzrNafff5bZvjLoJGS6nIgKuq
DO6yvj9Wr8Aq3/HTnT8GGc2H5h8wF4hSFnWU0w4XQ18oOIPdiPV9KZa6QnzX8Mnj6t/gbO+iuhm9
NYNBKG3EP6cY97Cw9bcX66BlmvGfmM0CbhVuDxUhTxkCFFopA1Hp8kTgJnvyBEIOEqzLE/sTeuLp
Slv8oHN+yfaBdUVyq6ioM0sMpIvSxZzhL75B8kz3a1o6NpA4uCEvT92FQV2W43w0KZl5gE2Nt1lJ
eovSVVlbqC5R4sCUA/UY7IrlX9PQ6Y7OhU9TkbLjrKh7eyCLuuDG9z+ZJM9A7Ek2CuLBJi/xPThz
NDsfbroXVL0yh2pVXpX60dZ4QnS817Zr4eUNwqCLf4zK5Ni6A25j735gQYgWp27min3XOn9C/0y7
T6xVp4uEmYzg1DNe3sddnUD5z6ttLWwIT7wvpdp0PlCvL4ct4gc0QGOOyDZlt07X8cFoKFWZ6FuQ
GcacuosdIngJQ9F8xXkr0wYUXkU02GhIfwRijOVH70SsI3OZz2zGJ7Fmbq9G6D3x0PHkom/+nywt
3cmxmlz9Iu12N+RhHAbedLFwjKT0AVPthmpz2ZkM8577Oaw5UwfDKlSb1f6yTw4xkVwpyS03JQOy
kzGI3MFAUimuavkLlGKrpD47r7rpS2Nn7B6JnJvWUeTzPRUXExaWkkGmk0mRj3vHzP8ghvZtSAez
5mFwATQe9V3JYFAJCNcgoym4BiWRCGKHIrtexwKisMfAaUeRXOaxtJzPORK8NvQjirxg0hzD6tJH
fTNoEh3AdzleQVKyPAoS/oq8EXJ7DTm7I8zpat+NDuXdvHbSbTt8vzB/uneJIr6WO9UjqBU7T6xA
TcmHOVuqdjKAssxCex+vtLAcc0giTJSG+7nsEPETaIl7k2P8i0npHb24mWN1DV2/KB+mtoxvB8K8
qNC1RtUVLT6AH3rZvaqyiS/bMQDYKBRGI30xIYAc6HoZNBaaqnPmY82Iucf30HkvI0O0kDcYG3dW
dglBT6vocDXSHHqLm3ggxkS+ANZdYKqzrRoOB/VlpVono/QryqwkkueHmYHerP0bA/TYiliy9FZs
xq/j3Q8uR7JGZIaJsZETQAbJCZtIMTGnb/qqTTEZZM4y48q6y1ELS8LEdlByDVOHepDDs7uCyR6w
wB73uCIHa3zljJmaQfGuJdejyyj/bID8pcWqf4hm+Ne0ayOEnnob4YAO05WMbI3I+ALD+rcdLrKw
jYZw01Bgq1JpokSB+4HohUyRYa+Ukt/1XXokN/NSs+YJEAsqGSha6oQdkol97ylp2j9RfAszLoOY
UBF6+GJYHs0Fd8UB9l+wwEuvjMpKA3y5dlNkQlmyS711pcyW/2qKt9XAKKhE3JTKLZfrqjA7B8+N
V9QLljZTQNNZ5neKpXAsSOkNmHmUH0swAooH0dZelMr8V4xOMdwDWkbad0zetyMwswjsmHT2KrMO
Lp/mbKIdJaZRiwt5Fy2EZRA+P/ZrHZmdNEe73GigTSAkYns2eknOFQlIL2ETIBkSiT92m5g5wrVx
6T22WKuk2IiJitcG+uov8xQt9xLKkuzBFBP6eXZt5V3z56+hEcs71nosrGhQGpjuOQTWCAoxvu2Q
PufuLpYCSMKPFncjtMDzcD60scp8UIwOF49eiAywkeb+1Z0PyPYo25kB/evudlWdboCgKxpGU2b7
eA1WHcC6eGZOZ3RHqLpJnPtp/5mEVuLKuc3PO6x8JtJJZPyrcyc3/Vp7e8de6ahH8ouRY4DzYviJ
0t4s8dxQv1oP/3V39imML6o4bhO07xK1hyXmL34yVmfx+L24EGLHnsuAwR9Q8qvm0jrAS1H2IM6Z
34503IeeHuO5eSfjqyJjaaz4Rue3mTxwk4zCaa+4WvmamHLv/aD/IL3G4zWAgcxAgkdD6QWeba4+
mHw0SQrpqXslV+RyZRFkP6TtCeQG7Gu1eZIcXqyikeQhvjcvIUu3NXK56qep0C9E/YStWW7AugLX
6sdAySSbU0pIU4EKocVZxYWp6mLN73QtPs8YUEMMS4Wn3OdljdLGYATAhYIodQPggzb6+Fdgy6P2
q/DbXZ0/SRMmftETb6WPKSKnhw6bbPxVwF9DgBfAhK9u0JmdlegFtQFFYB7uIbopfBnXICEXWczx
a1vY2Km8+S0A4e6FbXR9Z3tHoF1hzPkViwZEuFU7aOqybsWrSdaGPX+Gt9rD3pcVIhxT4f8bAZvG
Xy4ED0rAtbkBBw0MuV9AedxdAuDIGOQqrzZ4yISKm4d921E30lyfnMRLZsO3NMh3rSdXawGUqCTF
ot/nSEcOEvOV6QO8YTyxv6Pc9LKAlJDt5D+OswkxqV0Sk5cXiMiAASt3h2zAk4Phkwroz+XDu3TC
e3ZnKW7bhMjUmEQii1gBhkK4LDSlnBwxzfuwucviUQMfgNhtUTXzV7a0ZC1fuSHxBGiMhmi7YEXl
JOHerW08cmuSac2Uwz0asBk9LzQrbx6YFt6WUPjtvv9EB5DY4PRSnPUDU3+TJFor6CuPax92PNHN
n0E7YAnFPOPKXvWSSXB63YENc2LQdAltJa0tO4+zm0+Hg9VL0/erge3IP/qKKhXArmF70zFQR0K4
MCkztk1FGtcEeMkRvQMnfz/lke/4kUbaFqkeXPpafQk/i2eaQpsGWPtGbxx57FtVkHzATgrp5W/E
hUTbNza+3NgJZ1ZoF0LuRkPxibl5I1LHQupfvuqp6MAvsvZtrkfc1ODO4HFodTjJp2ylI2DH8hJR
EXUmecMeBFHwi2lFQIN+d3AccM49yxhhHqgbGyTtSHz14zkJHo0kqZ6p7E+xLBxhSNHOWom3UL9+
eg6ZQvsHMD695zcViwXDU5FQPKbivTRuB1q6rXyTD0Y5fJZ/vTXilUP0ACNP9SE9yC5TUDWmUW0Z
5sZJzcqQ4vKPCNJe+hTTzCa/GVhwRAFgECWUTPAEmSRcnTxgBs80z04oPLs33KvEC5F/+GbCFEFs
LZSD/Y40PRDb/EMj8BPmGMe0lMt/nuZlYehNWDyX3DPx1Ea/VfvGuPxXMV4zytO9zRNdmImTbi8S
hW7AaxPeLfmoWJwF3kAeMoQVG8BukLiF4353ySICPb0BBpSj5fQUZLdnRX4uYyib434UEL8DYEQ4
c4ima2V0JETQbFAohm0d0+43H1JES3q/4J2KNIdiaoE5/rMQ48wYmx2ig/YnjhpA78Q+UoCipPcA
tKtCKVIZDNcwuKj6fTHlHabhqBgOtaN6sqnfeYiyLb9JSjf4VHSz0NnPLVEGpdsdItvdKWdttare
+CR1fDvxweejZvajWAoSZ6L4wA4s9SuKwn2oQw+DnKPQtYfeMUiDvMzWyXUTGOTmQm5JX3At/91U
wkbEGSF+UtDnlPGToFo6TldPr8NOq+nIjSIrUMTqGCYvs8lzjWCyL9ScrnNXofdRo9tpJoz/oPOC
nVq1Ibhwy2AgwM45qVg+VaFZkdrF5nOpDMJqkZM7sTCCJARkTfqyTL0U9MBGGf0cH6x3ikHkeu9d
a9Q+jQ/DtFB77LWnvtxIShPsfYCQwRUrm0s8y8rGj7N03+c/xvmJRlE46QA4klhb0FM7N5dfKQBV
KNzLiIrLc0J1houhPJbknPS0CMEu+aZyLMAGR1DKODVxeTURNWMYqMZeuPIlmIQCUO6P0cyv9rN0
uonaBz5Kw/rd/7p7WTOuiMTHppsrENDBlWUM8FsBqJMu35aCmL0Hr4b/Ruh5JXCpPpZQks370N+Z
AeGgXtTo4SM3FYRe5eonC7rwHkclbtw7PbITQaxMDOEcvv3b3Mju3k2GRcgVBkIuTqv0kFtGR0jb
Bpu4xBD9sp8cQy/+fuK+tNxHDHKDvRVRU1AOsFDDoacb+TPkUmGY3c2Nw7Ad5W6xrEW38mkHsqkf
v1EflNzmiZTPIWcwweUoWmqIk9DTkrDXUL6NExV0Huw/3r5ymwPn6M+b5Ng558nDP5w7VtBg2WLT
F4MSxEq5XPN/YGdvL0gMhsi20Lc8vfvA9dKtVeSm2d4OlUD4I7YGQqT1ILQpY+Mtniv5ptsWor/F
hWGtPwEJ0zOUSIiKm2gPpXvZ1D/AvTTnwiTu1CymdxZgB5C+VaxSwffMf8pEGrPxnzOOpAmtdf10
3ESN4nLEDLJ050rZahi7G9ia6NoLf5x7fBlAzLCw7z59C5QjwZpTZnfpGBqeT5RUgMmX4MzJqUCC
nsWd/3YVIl3hgO6Jw5uVFe2d+U8K3iDBvgMH+d5yfDSw5wxox3gLAWVCw3gF3NZiCXNkT/vvR0am
NsxsuEllBbYIDjX8xj7pozqpn5BmHoskRtKEOkW0o6V9sd4cyN0cmd0Yesm6wm+qEgTnxwaWBX0u
bXS/d2h5FpzbvVRxXscLs6HwE8se04v7uhU4r6R2k8wRGyPnF1eiO+8UqQZae/IRsOfHndtzbi7z
jI4Zcu2MQCTXua7UnMTeMteeYzedHXfggYTFWyuEqzwgoZI9Gx2L/WYvwNSHDMAb4Us9YW8x8ai0
cOhZRvIw/Y6ppZQK/fFpY0cQjE91dyt1nKpMv+dnsr85Lm7knZdeDnjrxqhCo+5bLbUdA6Yt/gq6
eJvGCYze6j7+DDEuD2/BnJT7JY+MHB3IA42XmqFI5aIYLlK+j1PWiQ2KDlGmiKuGuoKKuENJ1d+W
uf774UH2J35HYk7onEox8cg+ZhIrX+zh4Ix899Z+FdgPc3YFkJDzDvjNo9hlMLbvBmiYD5+7ry9b
j4dJEz/ucxgpkGNv91Y/CR0SnMQWAlPigETSAtvhnCovBjNszx5vPSIE9tZMhqNThJa7HdJrYx0G
W9lFHya9inZA9TLqkwC3XzrDUHqV4Pi3w74JqI5bCx/8vzSQGo600unEdvzr0rQNbQeU+hF/a1QL
YIvHcjgKU/6lXi2sUBOFkKp4mZ5sNzYnsXn6+e0z2Yh6DvXIsFE+23IFO2yHtBrXaP8dd8fmMFSO
yCp2+fF3gSk5G6D9urDHc5MT591wMgBSzYZeGMVTyOXpZDMyEfpXkVLEGNL+hnNsx5r/k6wH2qma
gHxyKSqBPZMUNKKmmy1U2rkpgWNNw6rrBazHBIVhR3RVG+pRqio2yyXVeYgMukI6Jdd6A0mIipOP
YFFmts5q6/UlB1Q1Wze0hl00ghYYH6KBj5hYcOg+hatHKi9OJIKAhzPRfimjdDI4Sps7m3SbpUwS
p16iD6LIRZoCT2HH20u1CB1Wu6oMFKJRipcTI3NEeYOXSpIGK4KwXGEGKi27HnwKZnR5P+CVpmoY
E9SFSR/Fm0Qqey7FNhhf8r0zoICKDZi1Xgs4lPY0V9X0U54qn/drtNGZxIBhllMY07AVNnoM3IU6
/D0NdBZfF5TwnyfUROnDWUFynbjOaWijPYvAik+hi3cU01WoOPDQJuARCXVOgdLcZ4V/oXoxhdDy
n0vzLCxbG06T47jMK6mAqI6G/yG8v2UGyrNJslbxamNKd+CHhFXjRypWMpI+trB0TLd1C4+wdUq9
NX0LTWy+X9xuKTR/n0v99l20Fsrucai8x2Gp+6lIVGzxz+OafVvJ1aOEWDAIAFXLknx7l0Jd2L6R
sZLApKlT5GnXWSEs/V/NQ72on+KsCICS2rY4KeQZnL16URdQcDKvfy1axbyBN9Rej0lntsNMOdRd
cOFR2Sup0ssxwSbQ2Ik61cxONOcHK066isS+Z7BdKhjmZwmU3zPhWuZKY+/MDzBYqpraA1BSlSH8
gjNx5XWgkgeT9LG5rsQhzkbnIsrP/pScXpua20mqjndRioKS02/goUx6grXqjcQmYRqejEOFmnm5
DsQcEB/rrG5lPtsfv8MOhobbHoY1YRQqfFhcWuIIfJtURU2feDOYhXnmMm1prUNeCOgPDKqHWzf0
6O4fO1avqzZ550LfSA3HOLYizgn1vlt8grLEjiIUBt/S1heJyvDyCpvNQfRGqdO6FuKaLrrcQ1IG
EYmAs4E/YJOVrmiO4X37NGjE2vZrL2pZVwcu3yyAeNc4QNl+aoWAmpY/+tFt2szHDmtke+ovGNsP
Y+8Mz9ilWnANFrQHeQAzf4rPTXEsfqy1t4/hLnrX8yK5UYGZf6NTxXBXcr+G4Kxw/ACJqVxpfmLb
Eq7zM0htrIl/8DcGT2idEt+U/WbsIimnO3QPEJCs4p0sMoUwwk2lvXZIf2e1orDXkJk1V5SS0L7K
cZx5eQPSIuYWVlMcgjOy1/Frk+1rrrAWIOZ1NYNB7xAXlwcr8znr22/u6UtX9OZ3uczpLGPBaVOz
0X18sVR+AMalzAEIMAcn0vxGBuHsdRFyleQulLfbXE4FMprJkmGfulgIQRXk4oK9g6V05SRdfm4e
Ru2UI5/BgYURaWByRDOi8YjatJfH9o2SaYP6JZwan+rF0pr0vZ/bYWH5HEAPTXJelkQwY2mC15n1
md7bRs9a1bmB8Ml9rEj9Yt1P8NkzJla+q/e71aW9FnqTLuad0XqG53PyrHe3SFoVgTIuinaksn+i
mfSWY+eyHla8xT0XLzuM4DdNGvVMACkEuN81rxFVbZLZFZpf9ximk+D471WEIYE5NPYSLj+hwsdl
wiwJEGSe+mubmOmVEOmJzxtNW16dyDaibtmJ79pgB7jjDuiG8kyaY5SYuuUSRTAs1piF2URtrkUc
VSZ12RQSjUaEh4tH1z+0DwgDS+3TbVTmw5pSgblefhHxi6kuQIXcxQmkJM0azG+ymm6ZSDfxAzYn
yQqjf6TDfiQduQK7CO+Czo83Wz61qG/4JLsVlwUt/zL2Sgv9YCtiotsfmmkvls3pHmX6EAwMqcko
1NBdpWYlGP+kN2XieIyBg6q0JPSzjrNpAPELfU8pv37oJDjxaMSClizFlj4X3TrTJrhP4gXKtAA4
lQICVhWMTqQednkWxQjSNMq1ajvey/s0Syv3W2xlWcp7sVMsINvHaorZZfW4j3hB4KQqfpRxiYQx
YqFdMlapSeQdW/C1NlN0C7vprNs/KRdbZCYNqIAmBZj1cKqU+lmgGL2QfZT/dtABSzVcYpVVHvYH
9dk7Xtr3eoBQr26oKZqOcUV/OtclPnC4hznhqHwKwFx8HebYphbEdrlnKEdrgmIbn408uiuBPwTq
utEra+nxkxE3IGcSMoc5o/+mgUdqClYfkHF0jDstCJD6vBcWjtKyzmUeApMlvTPxijZ/voQQ8n9T
N5aruZaW57ykGEnCWNJbAHHPnrfbglOVjzEcBwMrDfEOmdzuqsQOq/7htJdwit74PjHcrxgaGPEz
5Aein7LM0u82dkcsjnRk/hM/pKbiGvlbfVSO9IALV/tAY9LTgydTcG1WvySDhcQ+LT3q2OzlBVQt
mNWMxqcnh6DvezBTe2EAUFRP+CSJIFrnySCCjZIEXdRiQQCsD8mJ1E6F0kmC+i19qMbVCnHTlFk6
BA6VNodYz6LtyGtu+3M/S3cTSnoGH7ODozwOGzJQ+3ouA2eww+YSnb30VQgLdKZnQ1VzSrZz/Xv8
7t+EZUWcp/6FrYEkQLF0HWqbyi3Ovn/Yyl7XwfuNrKxI3x2TTM28NDIjndQHqqB+OUWhC9VFoeWV
JGoYafsMx27XVBLijDVoruOmN5P+EM+NIPrv9FaCwvQXd41a/yvHE/ux74+IO4Lsn17qVgxT5duK
jPJcmvY17TDSX/f8nVPyUHJj/MJkibfozTKVp+2MUTxTVD03Bo/ZM+OYIIrgcw538pcNxnoRBBs4
ZJHh6N8Xl4TWZIS5N3ZdgULZ8toytNfKwrub9L9gUcGqKx30gXNgzsy05qmDPamT+kt53PgrZ4ma
X0nJpbGVkmJsFpA61om0Y0HkoayeBYwUHfaLgEwHv5y4OV084nRnhCe9T5yOVEoF0DAiluzzRJgp
/swsYkOjQleniw6bAwSN7FbhLC2kStfYdXtldD3SSCguxxZ0KqBDYg6jgigFJ924kJcxTVUvWAS8
c9hcR0ryJts3LhEHQtcAT+OzOgnHgxaadQm0Kw3deA0QRiNV2HUddGe4YTj7/hBo/WIi1gm204Bb
52OFu3794jyS8Fd5CUy2S9Uxui4FRki5YFN9dTVBVAaFf+mz2fcU6+6Z4YYKLyZb+rcxr/gkTM2Q
P5fchSq42432kBxR7gG7nHZCL1EjXvODEw40XJMrAY7KEvJsCTY9SBNnHP17DM0llVO+kLhzmrNZ
+Kaq8El1vwSGKEYQyyxL+4JFXnQ8BzSXZD2yh/8ZFSCt7rEPmO5u5XFaEP/MszZXMhlqcXErRTIO
EVsIJLyccL+mRsAaTdLImCSGTCohk1IoN+xuZxuNmQq6AJRo5QRwqOTxIkAyda6l4BB3KFXqVjdJ
rWDNDXOMQzBu28xqZml27wHczdu0sg+QKKiST7nfXN/IgzrK5/xU/6nLSFbzqhPvprawXLgxYsSR
1FubEKnOGAJmsu0TnJZAgTGvm2vAHfRR7X5QqvTJFV2fJUBG/Moo2BKh4ln+wLyyIkN4sWeSnf4t
9qiInBcRZUSsnI81+9/ITrR6sED998aByKb4NIxUi/r1+ZtJnLAFnuMXvR/gEQdSna4f+3yEO7ws
P/VdVEjad7bAsTE9M2kS4yZdIZFSXQ5mUWIbzxNPRz4MgL/CxFEs4vRZndjOSrMltWLzRl+AZhmY
G8HtJDs/0QYhm1x/u2uMpDyjzvtFk1TZNQeEUGk80b5b/cYoDasAPQQDQKrYe0c/6+KVuK+A+9fI
mFGNWLdhYiTbw2BDzi9pz/bJb4KKOrHia989g6Ce9tEeQJeF0/kfZqj3zz7PR7eXdm1AvEeNgSnJ
6OJ757RRIDZN0AVSsjxxYEfYB1Iim7tuzQz0jIiRbr2rTsTYk4XGhOVKegwkWDsDxJfw+N3ygCF8
r4QozWKGP/I5do4Ns9nm7Oqx43lDuRs/djqV49MzUEYO3iP2xpqm6TUL1i8Jt8g000pIhUxv9qWe
rGsKsN85sX3BlK4oIsQFoP4/ANCJhONlqavXpNhSPoDJqLe4JN/jDrBgEdw/uAiGz5Je0T9uF+g2
uV7EOtaJ16iTGoq1J3AGKruU/GbacgFKvb8/rjwz1Ton68TKaQKYFICufsG59ThexAemcMqIa6qF
6aVa3Q58zWf/02R856dJ6clntbsUx7rHUvanACUhWrnKu+UbclaBZ5oOOcAZ6mwRa3pXEx4FDnqP
XDnzQfnEXQYUAFrj4bNTgrQ7d+b2rRwL8G8DAbmVkws0auEfuPCfjGljsTicpHJngkBpkKsp5VqH
GyFIt6GtPz1/Lh9k/OWeHOvtHoUeK0hg/o5kkTj7nvjg7YTbkJE3ebcR2AsrbAQ0yWNum+w5nUn5
z3EKToq5ARtAsvUtXPh7sPvdfUpEcTDaGPtQDaWd409EeZXDBeyT76UCITjtApdqUw/71avarszY
VDzgxWZiF5zPPD7IQTLFhhjNsaI7n3zbsoTK/JlF9o/0piQtWb15l25rYbQ83GNFEfu2uHyXzACP
ZtlQYBUt3YlDYWl1bPI03JRazm0xnGjrw7MNx/M/UhrYLPjGg7v7QMXaxe12j71+tCF3hKkP5RIB
NKnAC02c8UvCIZ/3khJ8rOzvDKat1rPHrt5T77lVUoIrC7+lKqqeJkYwWsFQhoQyY8WJu6qappyQ
cTY1Xvm5LY1notQopM7Xd1svCptc3NntXzeR51hS9KpSLeQnpEaUriPBkLw+iG7hDFz+EBSWySf7
Rg0Pk7kFVMUSUqQJMb3qzS6T8ke0E6VdQ7Yem4UY+fHD37Xwy/EQFBn9SK8WwaNPSTpwUWniXHcw
Gy0XpYfounZkoQOIkHeBErEXY0Wu5X3oO50sCxAAITK3N0JINoZ6Q3tyrqUxCNrfJjzGUKmIqNla
ldLNnm8PxWunzD9r9JjVz3AVMbAv95No+IDSx01FRy+7T+ey2ewgrM6mGKUqYX4PgXztJdAVhmWl
1GL/IjmIFsIfLV03zIuu1fAY2BZGag1LgChwLBUbTbGH94dELsQ2Dq5vhSV0rXjm/NuXy/OEZnoM
7XSKWVWR6qh3Ie6GHw3OppGpKFdBmAXpQlutTYaAY0pIjiwNNKtLDeQVUReRGTDgkHRL9gQLdE+G
N/HpdAIjLhNW4+X5vcwfom9y6HuuG6DcHC730f1y2ykLMEBuiqNjeP5lHmWgv6voK7tmkz1pfoJd
kzWzRTEQFzQW0I5nXhsD8HH4vBlRSJYwvWefKQMVVJQlgJiXPliRyPvdzJFMo4JsCtBoziQhwrxm
GwNH9DG0UxpnXyLyQnSuT99YtN8tHxSk3snJ38GS294AWUwFH9riv3/EAKAQWoR+MQNb6Sq6EQER
we+k/MXq4+kWS3GNcJCBPVCs8yQRh7Q2MygGIvhEJu8pFmxfT1BpNJ5wWyOF/++kjCJSbvT/qkUu
VUgfRwCFgdMJTYJvGCC1FP5xKYx6ifbei4QRn0Q8JQd6lihbsKREscYGnhSPwEKigdcUnd3WhxQ5
x/B/DNjcHjeHvNtFn235PfDsDl1M86KTNXdGhlvLu4Gy0XAy9kQzVddr8NdutQ51PXl+g0NCUhjO
MUEwpG99jgKFPW2X+8kY2jMThAVXrn0sDguNHdjSd7f2D9cgNs45lTP6SxcZmEz/i5U6LYqKhISC
W6B9MsKi8O2jComx+rhREWHWvvwbjVaMJAL1RQzzO4hLH74oxwCAq3oOKuYgcYxkEOJg8brV2eYu
BYQGKIiTgQO6Q5DgwyBSwVDFGxecIPyzENMJI+8rf5Ot6imD8dWoGuFNVN5iXGkU6BtDkWSJyITV
nql4ZO0+YP0NRFgkhIO+7enB9mZ4zMQU0ewvEozxE4XO+zAOCoujpeqOT+bsG8YtFNO8zfQATFM2
aUmMyCx2DpMQ+Sjdi3YhRf9Qlmsu5pvyEo163IpAESqoIOVqs29NOQqN+Yq+5vW4R5fpI8Y7tRy/
HN+qkrT33UvzBeFzo3Oy05xpfXRbCXiBlGZO8EPHheWZW8cyji75GZ2dbl1LCbu7WhT/aeV/Mhjd
RjVMGA9rgNnkOwwDKru1FojJjrEry8qXtLLr04Ku6XxGU7R24L1NGmVrNe18iWZNnjTczulnXD88
wvVLLRkWxhYzjbZf7p9hcWG26g5j0WK/AT2wqhRnRyIc9RMmzGnQdtYbO0zQ+6QEuSd+Rz4092Zb
O7k6LljPvJi0XDHuLMHic5Sgw//I+HnhoAxBjehs1/TtXqvV1tHsqD9O344GO8kzu8sFSdzoVFeH
nQtGrdJfIBZavpK8r6IuyuUpc3cSIKr7RDdaMeii/3EUB9BauDP2haim2nmRDqh3t9kr6eXyR+e9
Uhm6y1qpVTZ5cUnmN8k2DLfLWaizUZRlUooT8iOTSSVCMyqZEfixFdmuReCcZvnQT9hgFkNctjSo
tzdNCDLssd+RTy5okTuovio0XtxkI8BiWWObgTff/xusREToXnqFEKp4D5y6puqg1adf5cDN7pZd
HC7xGPTHmiOGxx8DVijop/hEw14I8m61fE0rpGIr1ECe1bFif44eKHvrxMbq2/CgMuZo47+HwJcn
zwQONKrrykPCr8JwNWX8LprRCuTXfqFdHKO1mEkjK8GJq+zzRVvYa1DR5hLzwasTllSLxf77X57J
+4vgtQBdsX5nQqNIBcNbFBN+RXaCIQxPwI+5YmWNOrdK73IWsKjLG/0Sr15nh8lDtmNMTDofIh+z
tZzrmjuAK6S/C+UgEepMGvTuoOJVTmbcUPgZT1/AFJOt4AO+1VKRFa+mi+Nes6S4ESImIlJkEgL2
pPvd+kJbSfbsu3WMeylhdYJb385jxNss4EV89IybeBSG43LW8v/wnDMZdzGy3sJp9Q/J8jbj8+Pv
pGMLznKv8xN47Xbp0e3z1Npkm81Tk64XR9veSTXd5zM7OOGXLG8L2K1hK3n03Qh02wYjcVKdZ0l4
YERiFcopL7b9r9uxDis7ZHYHF51ZqGPpSACX5UdOLpqL3mMVMcT4+AlL1Zt1zXg34Q+Owp0x0WmO
83EUZebj/l1BX8B1rjdf1SGTf9n0G31mW6FiRnxc0etPmrY/OVDqRZdWHYrCAXDz009bsx9guvSG
n3DkeL4XAc8m0uSa2R3uk445i/gqvwwjQTntvhF/h9yclHur6bj0hzogeh1jJpqHpfqukUutFkRD
X6BoW0jRIfM1DQBl5+dvlvDVQQy7X5Ni46zDXWA45ElRnB0oNMX6qPt6ryBxuL4EbEOxJHyIaIkl
Zc2cbnJFsAaXURDuY636vDU4UClw0WijQK387pBU6HPl180n3TqEgMg00kQFrvS4ce1DPhexEYVb
C6sFVr4ChfF+zwqXALkHGrpRQ3GmV3FSJirCnv/Y2PBqtpMmeC8If/f+4PCRRx5YUX1dH0awEXzw
qtptjuK57MOCF2aA+QdLwQJgdBRmHcoFzdREpW+UFmQk+ig+aZCCuMRvzUTRivw44BYvuaHmIEMP
AvtlhtPBLQKrlWgR58RPiWGNC5iOgf/cBpLs1HcWmDIEkRrGaRVoIy4lEboQLAOztLEb18agXii9
VMmBlL/ty6jcRYVWrzr82QaqOMKXvNWpAMBGwYfIxugJA9TRsIpzZiLbRDrxjgiGsUk3krcnvs9x
bH6aMAYCV4mrkuAuFTXtp9vGnaP3Zi+1rLUP+O1MVGNnLjx8+ckxWkIOPvkZFPdvQ9DI7pnjDIyd
kC5C3Yy6pqsTsG8Gkmpzoobe1UTemgsgzPB5X4mrJMvo9XbRuewmfW+iHmxH+bMtnHeAXcVyEYSh
Fkt5ni3UIdBy+gej8lJ5CZ6Obj4UNe62KiDPTaUkfm63Hl2MQpLShJDDUHtC8t/RLdN+3UZ1MRFs
GRQgQ5ihIuanlmO8BIHufHwQzRhWWsJdtnYZpnxhaYWsuHXHemBIHPcre5DfAdVXm8gfRQNWFo/s
VDBZLC/ra8weMMPZ2lxZxNslYbr2MIwr35M8wPzYnNJX0I9T8uXI8xrm+oBv4hzsXiB04HbroRHd
pznJY2VRh8iMSVZeHP2fD9IsHAHx5XWf1EcByEjaGZVvNEP9HGoAc1muDVOSSDo3jY92o48+pTkW
jisSF9pAp9eRXbZzmYJnab4YPlqDiNRPDJiUXMkoYjVBtykH1cKT2XzZf3IBydnF1YhtdP4hosSK
NHxic/etIgpdQeDABlFe2ZKRpOCIc3Rwkv1EP15pAm/OeNBam+JYcu23EibwgbIom7azo0FNbuqc
lSTnmrTSGPHR5LeHvdeE3Aj+LOkCMsDuYjuZK9lsU/ClOkEc4HZPKz7buseDt3wrryokFv3nq3EF
CmeECnj3Kmx/5miMT3wjUzClW6nWcK8g/isyo+T2m5VUecQcbZXa/baWmiyCEnvgTZoY6Wt6KJKu
YjFcsOCe5X7jvpzJWoGO1MjKgyvP6ubRY/Z+k4gtWrEmbGYlaBH06fHR7BXc3+4YTu5+YvNEFWIF
rbRRYeJQOQohCP8sO2E8b+0R5sHnf+vHPNwjTt3aMkksKMBPqIiSv6H3TXkYcH/Y/j2AMZJ+XAcL
OJdm2l6EtYztHKsYe0tOtmymjHpgFOIRDGwqBmzeyk3tjsQZFG9fhiKJsBeRx8IbZ/j3/8L4Bqur
5I+WnNPO1kAXgz+tnPx81khYbYaklimRIFe+NVv9v7FHbpVTG9Zj3Q0gEsUSC3PlMf5K/TwY70TE
cT//0x9/MGChaQ3udqvLl3r8GM7BfU7JWnJVLmYiCJBuBKJ9Rn3dw91EZadp4mHENF7nk5eDSyf8
Ps1iaw/07XlTRAah7b+HlMqOOJoRo+qduXM4DD3u9fUZDl8ln8jhWs1r88BdYX/bpsos0jFN3Nt9
B6WPNsigeLUfQpH/BQUF49MV0U40C1Jo7MG/mRIjGGLdu/BpZWDvqFlIKTc3rXB0PiZ6Y3Bt5/MZ
kAaohgdhZKnGygS958ZHKkdZHK+aoldwCyUd2+0AtliRDHECCJwmB2tTi8qpfQmzXvU/g9LoGsId
SXxHfUjg5yhQnjifey3OAhXSLJmNjQl1xHt479NX+UhSRvjBB5ppcY//KztpY/vB2a0W/lG4ofTS
2Dr9Dv1l88zqwArhN2AlBfvuAP+DcDlAhx9zWauGonzvGnRiN49ayC+2N8qSJzvN61mWjZmZeicV
5BDFKXKrskXaECkZfFvOi7LRkA9cnkx8E2iMj92J4JX3raLML1mLvVoQ+WBKX5owQv/hVOom4UYo
L1MGIN7umi/KgrcD/oGfxf7JntmmKn5mFYGT+T70TTK+gjxo/dxI8aZdTekzkIM5EcKvDKTSYVL5
Jck0qION+qRglUzr9pT38vl0hMYUCYw+hgkRRNXv0tjr6+1+/dTxCh3mnt9mJJ4sQ3NlwFotcGba
4SLdgAnuJoqtUCyTYnteV6okzS/ysq7kyu1D9FwP7JGv+aV2pJEvIEVzFxv7E6wPwTbUFvSHytsv
r4ZyQJiiqoECEmISWfRow8rfkfVhfZbbEsbk8WVkVRkiRbGWhehU8ndoHUKCnUjHtI7kpcK9Pahv
oD04UEvLaSoV18cn8tS2m9oDJ6uxb3tpawzNNao/WJGT5hTqncg5KeVjPQT0gGOnc9Ke+9UkCWaH
oGiYSymxzRvlvoEplwqA976CRvAtkNiIo5hHShUKkhTLPrX7RckW9Rd3RbEfWNwliNfpkwW1gNSJ
K9+PgmxlBBzLBmj20oiMEuEpM0+i8nzpdC3oeukwgXMd69woREglf7rBU4fASB6Gaoe7KAAbcx0N
GyMHRzNvVOOA8hDuEKopuiReUJXj3LHGB4Y6coTBEFge52j6+HmX0uTVlqdD8JaFrx/3CyPjk5eM
LVduaPnTuwCvoJ4t9WbKkKAXJucDOy/GoNZDlsDND/UKoSdTFxLHcqaboi+Nxvt56bGQ+isMPDOR
IFPgxm+W6pSZ8Cv6+PYybwNwwdBWUhj2krSXxqaLPiCrb8nOCN2s9bfOUzxLcqyPZPp+sEosn2KN
MrvL4NnuleGVEyur0JjOMcPqNWdatJLpvwHDa0jrF/0Ahp9joZv7vV4xLxCLE9gJ687wQ2t2x50o
pO9JYYQxEU9mGiJzL//G4G+cFwfwPkdfG2NLEEjiY21ruThVQaTw5X9pXxP31CEfU0E7ZfFK189I
pOuKKenUcohbQwxAa7U9evdIEmDYbYa/7zsI7m8b0CjcYvHQaLZ7+TxvMYIUm1z3YJn3+R/5skzG
F3BlJ1e8+w4Y5lex9ZXE8x4kOiAXcYpFI/Fe7JfOeWN8LL7qswrQRVxqhGcRPcHjYzZAzi1fmG0I
E8UJOB/AnpYbEKRLZ1UoAqw624ZHVAM70/h+gzg3TjaLcKaRUS7Cf9rS+0U4krs9lcKUVwxKSH3i
erfiiUiRzqVXBe8HKVMHwSFvu55KIG5uFMLNuPm9tL7v4jJE6mhxjdIw4+nlsp/FYIltdmcfhPnL
/3dgNF7+lVlgREREtJTNbRhBwGfcrgDReJThlDe+HHMi++offFT6RqD4P6JsxR3K+SO4x4l89LRA
cnShV3vZA34rCAySrCBSFgTOHhogqRfYJP+edjg9iyMCSsnfMnGZmdFWTV1jdVEEkErYSmm2/HRP
oUo5qRaM2t6m31BIncQKsKIsa7YpLqv81DCVUVqBtTsD+OCkU7Mot51JvdxbpfBpXMG/4KO5xFOP
5QyP8yU7f8CCfoGT5kBTMInB8jOkrOSXN6f0w7bEO6lZe0FRQYP+XbZ5ODWCfDmuD7BN40PMczWK
O93P1GeZ1VHVZRmmaGSJmdygZizg5pirVF5/uhrw4YDAyOV4suBO2NF4BJWA4kpJRXX9pyifLiLP
R4SwBssic79pEfqDjpSFs9slUs9qtlOkkesRAzcayMucqwRSaFP4V3XOhdtO22ZCfzvHbdPaxpB2
d/7W+aqsN2uS3fgelDzsiH3rLnGHJ4Hl8b6BxL29zr5H1U5Wn2fhIZcziyB2abEI5r69B3TlPZoP
zt4j+Mn/UvAbEE/lTwnOjZt+dtDTyDlppzmPklsFSKO2y006iw0ZCtTVFCX8zsNKvMPIabiku461
k/bfDL78bTwLwp1iTKLuq2pWDhTnRD/i4xuEUHSoFgCHuBXPqrNHbaKx632IbOnikOZrJIQrnAnK
gt+MFvl8ZCdW7qgbfJTeWFkk+J0qmKfcLs3SBGI43gcj2wqAqNaZCPaDoG4vQ11BRDMzesHsWOQN
UwZLMlU0VsBbGRaaa2jRUN3FAab25P2rhXDTJVG8e01mJ2Nf+1uV6QXT7YCUmSY/aYLADWHjvYhj
blhlAtb0iOJmj6PBy/tC/jjoYH/sVsVN0ZBI+nxDS1cvfFMi1rvv1DUzMku1G5Mw6JCjtCEK3Vw/
5DYqw78X+gY+9o7jc+ijoeTpwQZ/Mr4T/LEMoQfh5CS1wJea2AKciMFgY0EswCiZmvcRTjUgRkNY
GGf+DQJSgdwxldvsdE8yLT2fTGywXpp7hJifLMqnc/egUG6NJsXWTjXMIBUpQSGXRsgGnfSU8esG
tbn5VQXeQ0DEwdwU2f+hexkvLwWpg84R6uZbXp/vFQDS6HeWdaOBm/cfHmHesk6ooOB2yf2LNTUY
OphdcTFEF8AlXVqS7KEl/cnhagmutP6dvIlNvYUqHcct3uLShp+1jvK9Gk8XDtQH8biMJGI2dYcb
+inIGVXEjG0ULErvZbTASnrTihJ7pjsXZyoijfNNRE9TZREonvQxAKG+4gomVnyMGSmsziQJzfsT
FYytRnXAKzz2JftWYhn0lZaU+C5MPZxWFfWca0RzuzbJvKe+vAhHgHs+VKmpCHb5hTqKazlevexL
guHbUExOu04gWb6yvjzTu1qfnyG8MNxhDYM7SkTUMH5La2UHsO+k/jjneAA0A0Dfq4UVTGto9A5Z
PTv2ycCCpy8eYdgt5q37MvTDeaNVG75QY2zVUBNvQ/5SnvDRapb5DRazqmk8SmTs3i9UL/QWS1Hc
PNGCeicfaKMQFeEkjiIJp9G5v2XH+LYmZtAJ4MrblLGZyY2P64lwjOGT80OwRARqny/Up8f2EiFu
/oiPIBEAGXHFFSOS/m6wd6SgtgTUSxj/NY9m4VA6t60MFQHdRB5OFN8VVp1zDIDaI3+B1ZKiBO2a
YKKhXOS8n4Ptrfz/TyZOHFJTPqQHMDUhBgyB0PaCXGwE/q8FPlKspS/+RQL5db2rKSnGJfEeCmIL
Ro4nbvv86QxT3uo4zqhn5X8jYUodmNFM4YPGaoGa4J2EdhJnEqWrM49N6LEij80kse6VLuGDNZGo
q0AVMi4EyadojUbUMaBLzG6paRiZacniLj+YPG0HKa9HlIAYCBCnCf2mRMmgqFb6AR1qN9YFzXUo
AA9BKG6PjxhJvjH7z+M2nNl2CeFay6gEGy51J7rfdTVR+cZx3JM4mxwUnI6GikFfm6qu7txdQv/J
ASvkh8iPgZ76DFhp6Y25myjnsbixzJz11ZRHzdPBky6gJa4XJa7JEuwHeV3U5pHfUDSXWJABgCD0
Nvdk7dj61Tqh1iZ/0UaVaZ0c0sMmWDXgeOiyEcDwdBH6nBQ2ynZrG+c+szeWYgtGEz4OfnJyf6hy
E/cTwepEdxh+6bbAHYGl1evrzfbC+6bUJ3XQ3rFgXaMcmFo716ncu494BfHhxaNeuVUEAqePzAsb
XYMAnhaIxi/VMkvCjpnKj/BO0FssxUDv30cWOBFJfjUC1QRf/mOm2Vj7xCmNudpvsBf5dAjhzBSS
GCRCYFH0qw3BI/KVrJbZEhAPn3vbROkmHDJSTFmKKdaXf9eK3vGFCX/O8BXJdrssUp+ArCiU46Kl
OEPntDUqKrCh5o+3wD2eVxltuOLvQ2GgwuuxAhNX25+Dc4UWTxa/OAm/W+4zz8U+z1xcDyj5MPyw
sYlcE7DU+e29sNGKWwyYYJxFD4Pf7fbAbQNC07tSvIK+fAxHmjw4601Hw8M6dGMMC/MuvW28k039
PEh8fkKgjU/+LXnT6nvV3CEvLqGeqEbniHJNDKPqyl7ts+DVzTB+oetT+ll4StdkdhlSmWEVzf8Y
q9OcBKda7lz1qVvmTKb0Dotvg/PrITcK90AFPCi3ZQJzbKPpEsv84xWfxOKmNIn4mqqzB+R8g0YM
gxfMZG5gVccjwM08EtQEFsI9aLY2cbPbcsFxLAnLz4B1a+4OydfPNaaPwzBNTv/uK4vplrmDbi7u
dq9/c/m+h+KDtAHXL6plXuBGt1sb80teD921muUqm6pNyUlbvWMVaDDTwVyyBYX0GQXW+9d1VAt5
Ks+Ht+TRW/nG2yElr+cx6Krm0Z9dFBNmEwp0Wv8zw7GfS9oq41YB4BEpSgub1ybcFACO1shOW/T4
drf8/L6GS/V6mZEFGa2VsfwNRCKpBtK6G883KjIGV2MuPrvw1xHZ5EkM4NP0MObwRbomV9oU5sYt
feqTUbd5MO7Uo2tqtt/c3Ua2f8i7Yl3+jdcDIEwQl2KojzBB4DWAsNiUmpShNplnT3fXZmMoKtxH
0ulWat5GLBPOmcYa7cc/Ymg4lcoU1AkYoEDnlVhgsWJlAaL+qFqBZQIEW0NcC+8EeG8/HU/MrXWb
kF1zYbK0WuCPdlxhzsv9KEYnCZCi9bBFwMMYi/b8n3Y7o79AgfJt0asg/xJrzJwV6dnrq/nLJCnV
zG72zhWukO4idVhE6DQSbBRpH1gU/KSgOKJjwkFy5j0Y4X49JKKuCDASHjlgdvpDh/bafM1/rseU
KDoCpBpMIQUPzP5PpqZoSBP54p6XLiP5bn9dRzOB+QhMKTiokk1mc+9p5sk0PAVd4tNv3i2VgpJG
HAD+gW+UPUn/567D0CdVLyN9rlWTAlhTE+bkNh3redvb0AiK8TPy7Av8FIpZhFIYO0vrn3v+ioaf
WOx2Ho+T/RNvOIk1aeDiIJLax9k6UGovm0HllxLPfQy69C92baapXVScGtSzx0wphiS+tcLIrKiX
qCBvZVBxkQ9ScE9EEvWLn8iwIrpKDurAOdoO/v75rTZBymXy8HIWjrhuaH+4fXyS6j5j+Ug3B76z
0EJyHPmE2xBfBZRcW2eoMqbEhcTHBUKhRhTNxSaQw5QN959G072wCfu8PjoiZfluRRbqCmNQuGAH
JZzGCpgPagiSAQRI0L+5RKGZUqbzH/GT6u0fHW77p6MuEKY9gpjZ/Qrcz2RFKRO3MBpxjlrMylhb
yKFdJbnMt9DRhLklnyINQqDKKBw/0HZsyTrrsMkMOVFJveHWVpXTK+eo/zx+G2KPUN3+wsQjpTWV
npOjdT53p452NCAJy/V7blmYXFxx4Gw5p0//TJV77stCmrgxPgBjWyhAUjnqZEWQ9sn587Kuncl6
R0z2KK2p+4kp0uDz1KG4pfCY4S4xghOhR3Tu06ifNk53wBh0niN3j6Zs5gDhNgHjt6Vwa7Wbj/nw
bsXKXHe4e98HF2WNu84IsWafDy9c3GlTbFXlxy7AynWPnqumrTYx+C695/229rH/62T1EoULK8iM
+OSNNHieIWz5lPFqp9/9n2zdzzQWoIFHid/aDFcyCV/r8mCpGBKFYs4mPaFj52x98UQxJqm3pmAr
PcrbmDVE4L4LNoteOx1zLjFF0a7JGPephtLHdWT8nhyNwI9eV/EQqLqq8h52K9dCmjEUjsZuj1gk
ldSt010rpkxXmKOa+Rv4NNvhufTNp8irKAUa0qWlK7A+2l8pYKkTximItL94aNQ+HAD5J29iRKZr
2YoJgXmzvtBsrKuvvUSXZFJaLNY2i5C7CSKDoca+rsWJGkbVrzHrJ/EGrTF9RvDwRqmdgjEMeHnZ
Wflb+3pAG+dwF+BhfgGBvjLcjOdCLzo015MwSFGPH5BmP6T1vVM0ZEVZeq/rERfIpItEht8HL24A
fijgVPF8Y5gx8iOoNshofMWCGHj6RtE9mbX/pTsPKaWBX4fyMpCqy1jy27qJgKlDBe25SnHXml+p
KSge1tlLb3pajehr3dnrUchM8jPm092bOmzdDTc19VRc2JKT+FDp9jBprYoBIF2X7zs1rUActV2r
6mw8Uq6zY7LpgvOYKPzr56NYyoSdDxo71nf05D+LcAtcdeTxX2CzXJrW+W3uncvG/2pR5BxkLCYS
BGnFKweA4ShmxeDrkKGaOtJPumvV+qkweVUeDa2KvMtQ23WbStAV+IoDoz9eZHW+hJDSrOgrDy7D
i13xIDm1gunGVlcsOuYbnPGmqkI+39J2F3vbFNQ0fHnVePOmeRKSCU/e3kIBKx4DkAbaFPxSdG2E
OgXy4TNfnl68rukCQCElN5UX4oGDmAVJtKm3W2Y4bKgFBH/TvUt/oCXtwb1+7TDPQuK2paI2r4jo
kdh3NeHVcnyzRy7U5sfspBZYinjPi1llQ8/OQ2S7xy3pZVzGr16yZBBAXy0GsWMHuDmRENV8Tf09
AOYEy3n8D2vNt4/MVaK+YrxcyfVOMpTjdRSSvz5lmFfDKluE5AwWg9lUlgXdO5+pzwbqAMfYP2DA
vJOb8vKqZGbZBEgr3Fd7egbk1hkgqgfY83q/HzoYckFasgBi85T3Ai8nPUullKmYrJ5Q2oIn/n/5
5DoPzQ9Wcg6vjFJhCpjOMclS54E1TgAH39khAIrq35hYHhqZ8ucP3EXOqSOhxQ7MNq1BN7OykfbO
BNrHZONvzh/h4vZJSnNoF51XA00H6GSu2G2Rwhoeo5RR+pddtx2ZBFglH9gbEfMGt6tQC3QFXIGA
LFddeSvTNGHJ6wMebhdTkQMBcTEg+J7KHf+UPvMaT9030BycAvr/zEXgf3a1sbrz0ID3lsNXMj8c
2EhDaAGgSN2fye7YuM99F2FysEpdo3YbTgIKYB9p13Dj+rHNHV8B6KiIGT/CwUeqdwUyfRGfpS0K
X2CfKAizaWfHjWA+27oDkaGGFHA0lSjaSU6n20PmjQH/i64CmXZoZcP3xiAPl3RcMxa6cYWIK/VH
x/HlQejxh/MVa61FArDs7LLbYJ3dywuWZrJuxii4YgKSb0yeLwxrK/zuU72tFhFGz91lItfTFU2t
fnBPvtx01mrhdS6TTKd5ydV1ceDkMmo6J9Z47uRcwd25RyJxhidr/9KC1+TMXy03GlEqwcWR5vEc
XweY/97pkjFSirbFNSxtc80UCh7e6PNQi5ontwvqPbVfkHfq+/+W0Y5msvH3j1F5Ye6fFC2f5082
wcsIlCD4qY2JRTJ+s9u+ErWMPVhs4NwStDM/saeoWvfqwmh1Ht5PuqkPEHFuF1BmjFwW/Ii36kuW
miwCgSadEpNMiLhIZznwt02LMiU9klJBrT2szmw2AXZTUNlblp+fJA+UBe+HLUMjZn7ICYvmSgpH
39j37IgERWbln1ZZpLTVvT3okj/fcMWkqtPCUvCIfxso4NATJ3+Vx9FHZRc8MvUor25sQ+dujbs4
Uq3C7ZOCK0iptLsx//EoRevR1UJAHQbI2SFk6E4iSgfyHOxa27VlcA+geoXbAArboKvsnSva1uVy
+Kx0WHAvxBipkFg1gAd25tN85WUVuE+XLp916y1eVPDU/scQlwksVifVyp/QiIGExyDO+Xbg7QO9
R71gLQCcp+Hil5l1iQ7WglISVAx2emZbMIhNLvvSBwv/TWbNyPAGNKe4VTNmWNYo+YfdpYycnNq9
voGu1xKREaKtJcdbglAl3cllwjfnD99HRaKOdtiYrkFcP3lDjjrOdIYnGPO/iYRb9HQ2yI/uG3e0
9ulcMD0/S16VqRg7xxcfG6dulA1tU49NJhDiultkYtGU7Rf5JpRcDK74b/AiVTdrH9F1dFM5wWmk
atGN0LEk/Yjy+CvzW2+5jMrAcG1+aj0ttUXmhVfzWGsRhdZ9AFeoMD/t1zRueMeJ15ZG7Ltc+q+i
vrClzTBVwBfyYTVBuRaOAy4WliGXDhWJwZknlvvyhYPUHPv7caqJmdkJYm2q+6GZ0ha4xnLCiRkK
D6TNQBlDykBWToIkZsGxgKWSlA0VshBbWCzrk2qP6Wd7HI+Rgo3Wiwv7ia0jzhnn6PRFNsMfL/3P
MT7Xji43JVLdjAilv+ORicBk1rtNPLhSy5Sj8/i9V5E1tzZGFZ3C6H4gqDmC33MW3FarehCOaagh
XAcfqY5u6Q+k+jk6vCd0i5LkONAuy+8F6gahqkqcwL/6xjs+i66SwvV0QIQyo79dCn/KEcGGLNkL
W2x4x5c=
`protect end_protected

