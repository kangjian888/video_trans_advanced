

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Kv0N+ODrJQAnD45jVEsSEPytnysm3pvAbJ05V2JaqTdEQNJrijqrY29nJXOyqQOIioMFCyAehxdh
SS8dEy2RvQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
wl26nrMFXa6fm7UAkMFkRbwMiWczBO907OqYX8JeRapSfb54ShwQXeaNsbVvqp4GNYQWgD8fiWsc
Rg1ZH/ALNgmzzsXH1hqu9qf40O6LpbgjO9M5gvRZkEo/Tsa2oqZnRuXHxvGdfSUWwgm16QfnXWFD
HONMKYo+TnX1BbyoHuA=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cF9G3LQheZJrMO7arGfYkxyoON6brspPywtxFKpTvNhoNGqsA1QaxZgfesvqKSR6jIrBuWrdpeSm
PoQl517JxEpEF310dys+9f254GuonHdyipWsWNgWjbTCuw6rYLvLG1y7lYwgHlSqKUNrBaGYERTL
bx0Arf8JZijWzxoSQ9FVJxjXj/PfvGzrh6e0n/oHLpafMxMPZcDI+yx5HuAhNXSr705mAXB8bgRf
GS+N50n6SUyWqcyUqw3kHjqQ2U4vJW+j5ZC3mQaQb3xJkZgzHfCaBKMstoXIjqY6XkB5Su6aeqKF
tsdYwq2h1uyBfljsOFo3IsRsUpNIiryBaM1j5w==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fN4hvSzwAQXVTyvBcSPI9qSFGq1b0QWYvne9odu5QkpUwhn44DFKeJSRI90o/blLQLnT5fdJ1IVC
mwqzRlL7DmT25nQgDxB1mM1knf9aPQaDbovHFOWTzAPBPJqGcsU8B7iu5g++kkRlIJA/0D9NUZP/
zdeXDuR/f3RpGDQ9X3WIBcSwde7JdAaZPxu8gycDj+eAg//eJ+Ch+IApwl6KjZF7Lov59CHOoVNR
udrlY4+R4MFUEO48SwDCDlqVGTYZykUVxSqzXifsrNKc0qKvKF4GbqbVHDidoVCoh7f7Jnj0snvM
x3DFGPDnokqNpDBX7xF9L6+GYPELuxQwMV3Yog==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MECPOWJAU4w/UvBGQeSeElgdlWQuUK1on5QTAzUF7zMKC1Dzhpw/yWAmwgERdTOHF4jFwSXDGCYX
dcq7yoSgrYHNe1Z9FD7/4uOTgF7lUDYslV5k/HR/cVW9QWbwl5jLUaoa4U/BsWl+xPk3gCXBhT1o
1qrFxMGkr18FyvER+gYFNuGtJOdwhkp3EWSeT0uUZpww9gD8GQxRUyHQJxyLO7OrJ+p6c8iZL8us
t83ykRj64BZ4A7H8a4gi13wX2JOPHaLBMG6QaY9NxFK4P+cAlJ5tz1UR5CiOSua4Nbo8RZAnEv5U
qSe9Ctk2cb+fZHyT1Jbe89K38c/68dSDrW+q0Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JGQumRp5idVwKA3zzoqht/27epSOGyhvfg4tXP+tPHgo6OfP/FU3H6/X1Nd4Y66ilN9i+iugj0ng
ehLY04ISDe8fLdY/NaZ+qOkmAGDYirT/RxSo79rIeXhylLKnHv9FphaO49Z/wGAPNVJcMj7acDAt
BmSxt3Wb7gOV2zsovZM=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FGXHNsFzSGXjbxp7bvoF47vhF8reHgBm6BrifhO2QcSTwMmIfvC72GA44UQ8v8jHIWHgPlay/nGH
qq6loQoHzagZ/voRdMzWla+HchA2la644cxBm8f8Fq9WGjAfrRKdp+ka7tSEmDbdQiKs1i43XT8z
Q9z55GPf5g5GdS4wXPj3ZM9TkEPcyM6MWas1txHsPj+r/l+N/OJNLRx9g9A23yQcrqoY/ibZoyFW
/7no0S9W9Nh+BPh8OXy4CwqtsvPd0/Zl0/JDLnm5d0hcEAn+3TkTvrZq0NgpjAEEOfrxtp+HqvpD
SE2gPjJVpUBZWou1zkZKYyakXZCQodq+NDtzNw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
NQN5+826PyiSfAsnig7eFyqNf82PxS9dbaGhSI3iDb+4lgwWm9dcpXC10jVERerFbZEeHRjtDGbk
h9rUVMIeySzKGdGq11sDs6m4TsUyuVGDG9JrNGNAjy0Pw7cgeIqKX39FSy8HYj9f48THjGjHEOEh
i5vezlqssCPL+3utI0fKiUHdD1Hz8DwZCKux0lBmSubq+neQMBKPzX4VsbGtkXsX9LCFEyplahNt
AaMV63ORYAxI6PszqwLAmjaWhdBYnhMgj+FLzBFlu3AO0eufhxQanAn6f+fwstW13R7ReEOryGVx
CCkDNipm3dXwPysu2dGxUOWt18MRvlxmjirAS0vfyGhMqBpr39gHmOlj4NT/+tG7l8gAg+BsJ0+y
IlKOw/+hQ8gmPyrQr7ZZcZkKTAdabMMZd7a3tAvwRRIr1I2oWy5gAHXb/jH9i1iPTiKicNWwDifU
CFQWk2J6dApoUC2sAdmH8wyubCKrzmqwgAomhrjFlHk7DnASY0Wq0oyVHIS81bMFogO0n9Y8FjhP
/NX+i7MjU1RqbKMX5w2X73ylOgSvhoVP2VCGKNvqQ1cR9YNXEdJRhu9xah4iSi4sdTQDieA49rKD
Ii4Hx3Cts6zf5Ms19Bwn1S+/bq9KX0l1q+Nka3NBoRq577MIupaP0NtWzJaUTKACdaEjAbK2Wl5b
B1QMC7xUEsrbck0+TKPVubjWQS9kZSzKmFQ8pa23BGPGMB/6/3Nv/obp72XoEImaJv8uCQsmY11m
weUtsfgSW/mqTJp/K2VZxOLK12kWKL690H5GOP0mTEiC/otzCekYyXRrNx+5UxoR5iNK6wVet/c4
OuDj9paCm7TZAhH7/NnuNV3Rb/ripPwVsBP4tGdri5cKBM2UdONjPVdKyk0uKopdj01Qt5ZGZsag
0p1owFNOvZAMY74eaZBel1TIow25rCMqIt9eM8B6c4zriJX4ptohKo/VB6RCR0m/LMrzpGWOUYgj
B7tOYt2nlkgBiyCK3k+XfPMC5NjO9FnLxZtOY3FoZUo6t+oFNHhAeex6ldZa2QoCUKuzipDGGTUR
ccnuTSJs2tlJ9UUpeHwrBC/2OwNu//39T3TCVPAfy42N0ASYf0uzYN5FogIq7vrsiY4O0H3rjAhv
oNVOUFvUtlJ7wA5NnbMwJwm6dZ+w+aF1FWgMNQ6i8gR8Img6TgaQlx+L1wFExBJzn0nixKc6Zdp7
2tzpExF4k86RExN5udUKqTLacnmfPwkoxx3zf/gvVVPk/Rlvq/VVpSIxnWV3Y7Psyg0M2NzCDW4O
Oy7TnypiyTonsXRAIbjOSDZRDJbg1bYy8fPZdV3l6pjYu2Ttp6J603yHNxTdsjf2mtpBdW+RBySs
iQ7BvN1F5iAUWyq+p1RR7e9qULEbMqTOUWMpi58TGC8m0cvFOb6t3rP6jqc/dJmnmFjO05z8jtA1
3sBzdBv1f32ytxh47VUkS74l8ecdaEganj0GCe67yb5eWlElEu3TC+vWN/dXfhCscukIO2cU50Df
ccowa/R5geSwMMP5XHh4UgXcQCxeDW7JEUD87ui2OnCRWtwyS17+50+Nz8j5aPK+D7jg9CSAgLo9
FF1GKFJoLI9i0m1e+tFW8xhQOLIPZKTkoplmSiAmBp8aw+6YYqCS9DIvkxs7kv2fDFAUEPMCkCa6
1T3Cu56g1WuqoGuwPVx0XX9Pc61oGqrQeu1Xk2JT19PKIxgJwGts0Bn2cgAndCJVrwV72yEEwyvz
3lhwrJ/WEzovH9D48gaPf5dQInUhDQgM1PK4DV9leuR+aS6hMRYqtdAnP7H96rENV7KAAMFF3ncx
otAWAZDt+gNv7jZgfIJksmxSpXmV4nujemhfEmLijfUDdf0HXAbik2P3+GdFkGccnULZb4HHt8EI
Nv5J+YEXl9Ug6Gv5h0191af9X75Sfeo3aasyKCxQ4h+APHCyR4VGUAkN/XIlFch7P9qXN6/K/MaB
Gz9HEmPD6XIEWZRqn6Z9aqKM9Kjk9WecNRY8q0Jh5fz0o6y59Pl+iDNOyvvq++XFmIff2oJmgyJs
wwzI3Maqo8TRtVhokxtDj+jJeO6o3YTW+sqEbgUkUdy8lDpbPobReI6E3P6Q6ngSW2HZKaJEh9Rk
FSlPPrhwR5pj+MLfGJwmwT/ZXSo5FCYsM04ZRMO06iZwvAqrVR4QqYe0ZoOaMW4cxbk34TGVA9n8
UoNwSdxWagroUrP9mOXBqmuJLBwvi2aemxhZRiQtpoWJftRO3fc3Lj04k06N/jDzYN+BLeyCcWqj
NJ8Mh7d5/Nf9qxJ2H+A75lB/t9NQufi89r+yRBLdg4zV9znBe0nTPivIGH0CYKkGFww74ntx+id7
KtJz5c35KCISafHJkQM6yfDWjZEszklkCjDgznkhiv/3cSv4MBoVj/OhKMeHQnUOeJoU+WIm9qNY
HEI3IOkjovEhaG0leaO3WKXv6offx+Mqw0+6L5WcvxTtIsMO9eyJMG7GVMvS+pExLZyj9G+O3pZK
oaTCG2PTkU3gCmQBU8sQpuXAJz8t+jpo8FJelmWWub1nwHqSRDpQYc+0CQKmVjAJYRK72URngLJt
ckdwEQEt3YVPi5fuPZkJucxDjcIV/O9FCsb46H3uOVIfyVjhunvYwXBLn6AMXesmyY670yRdb6Gt
s6Qe68iorHW1Y95FAnvRDOxcumSAYxy9KIZ/wl+2cwxKc399S0qGw9NeUIoTG97l8ullYYEbU6yd
HhYukWotFvcicvohmCTtli9KGuKbz2x2SNj5g/ZhmP8czeWmyCESSSXb2SdPkEZdDZq87IMq/H8y
BL60nPcNB1vPWggf6seELLs0uooToSpYCBSXfdBpfnN8EQkV2jQ4QgOfdoEc/7uo42E/tkxhcmKL
i+KNq/MnExelA0lL/2p7j63EqUVcvL004D51eUPXgfStEAZ/oMEnRDEoVv9TdorvokFqRPIJ/AeD
6OknJVZYNdK431i3AVdJYjY6CmbQ1YXGCbGKNGcaImFKUHPzwrdp3HMk71/JDpmXS44kecYAJbhs
Qw+w/2wMewS9ktMq9ypxvQdgAof0NjxU57X5HwZKO2a753NQ5q4WomzQ+8RsFLCnQKKSIYXbRkJl
tk3s/3e3an4isKiauDd2uNMjl35FnlfsoAnMTw3JwW0gnricfRIGLX2eh71eTJ0QGTNfNl/hDDQs
B7j3jJ4f6G4ds9K9VMwLNsLqgBMTHxQDssbj7LRe/x/kCzWGtUhzk4MH1m4vQzWtG96mIeSqbedS
7/4CbtcXm5WaaB2oZ94BGPPk/R0nM+irgzd4z9CDWee37u1agJOHf+h9q7DHmjR1nFKWQ4hM57I1
rqxQseD6kQ4kfo2lwWcPTpujzOCweFgBuuWKJBgK6spqWVSHHKD+ISKH5TPLs+G+VF0f7BpdDQ05
GHOEz0W12JBamY1PxxF/qA52w/yTFjVtCzRTChLYP6XaOmK5+8bC4W7yDKtNGhaW1KX7z12Z6iJE
9XAYpQ9+q0xG2rflPxwrjownQaGPGg8JfsSaCsnX7PeeCZI4Ahcr9XUFK0ZkkEwKTdo5x/vOVWYH
is72z4TkVkcvBHTOA9COE0njB0XShUhjB3fdKpDNilFLjmtf2TA8LX4DfCWAtmV3kKhDmLhOLsuG
yuttM/l2cPvrOQWfAAhnbm2udvAkV2pC/S7vy8FQspQej/zRGTZwU5xBl9c8V4nFmWfYdtWCJil3
ovUZonohuauTP77O5cfbEq+mqOZ/EyWEwRfiMP6+Zo2JtSUOZIFXNa38uApLJw7gwH177RWcxBSA
ABbCwYIoCKy2j7zFBAKjkwLeI5JW2EN6JJEKTTd0f+m/ykHCmjaXmKQ6iL1/WqLsgrq4XuiqtlEN
XBUJFmaV6TjpX5SUUcNtA2GkduK0NKlp1W2idMsnLIx+NzdleguCp9BINpvI22CHk1Ib7gwXRTIQ
nJ39lZXbE1XTD4R4aUBhxHyo2PXM7zzG28WOV+YQavuQ1K8MZzjBTz48eBVk6KQJ2ehD6WTF/LZf
v97PFX1AimB6bJ+M4Pm15wTpm+7J8OW1Bp4B623QCHKWAGc7VIm3fvIhyi/9+mVhNjJb35zyHfoL
4KcreKdf4+LS+rT0n10y8GejIMY54CxtrIrGFeTuzTU1GkZxAaNUjVCIiwdE0mWKv1AGKiIr641P
qucZdS59Qqi3XMcq7u6Od8cdYlz47LjwBvErPKqUtIAPQo8EmxcEeL72k1H9E4p0GhaYtYdCETgX
YgEDeUqjV215SoxdYQkV0o90VKw9GL3cIhXUDOmfGbWZHQXoT4CGl6ZBL+4lJX/JE4hfVQgXpHaN
pw2CtHSHMfbas8cAqbO/8DcAbFa6Q1Rr5/B/b6Vcj0yjM9G+cLU4wjlP0aLXJeQ+uXp7Fy2k0IQV
IrUL0o6j4xY+su0jwUKs3/RbXv+iGyxZGfphF2Rf8dSUnlJTv7h0ls28QUYnvkiT56IiZlxbtg5O
p+Bz+cO6OnmH3pinJ4dihPy9FHdni2HpMo2quvb+zj5FR5jmfqhuHIWvB0KWdzxgCwALKn05+4L8
d9pM27SKTBndZU+LoEar9gJbkYxzqvG7xdnflgtdwpUiyX3CmgU4Fzab1efJUmH1wlb0JF+oruxp
NH42BWr6nhMpRIvtUud3sF70C5ctGhneInWJSlor5jReqCVIyAvaR3fF8f4j+RG4A4Ur8kiWue/N
bKkAfDExM/g79tSMl888WS+s2r78xRMhqNV4EICJ9n8JnwTXE2CGtP+NHOTd9OJ9KiFxlsFY0Hds
UqrLuYUjYFdV4bQ45CQVR9RsSorHTZ1YZst5tF0nfLnyz5E7xJocBv/yOf0nszXvTYjcP6cYM+CF
GY6E593Evb9N0N8NNMWyDZ/odk1jJ3p8FZQj2vRz0ZnPTdm+Is8tcmz0rNr5DhLNjWR3Ejm5BxDG
tADMuLKcFxxikHMpk6bS7o9L2eV0Fq7Tt+St+9Hd7O3tlrMSwQ1cxKl0zJIGw6+DDTmy7eBL5dMI
9qjrwupgJoDHmNi55WbBG5GThzyJpsBOaz4NO4I5Md/KlsTn54I51512KX1hdzZ9VppGFJMp2/oa
SNcFgxdIG3NIPIRCU43nbt8RCbUSdfCkqQ2b2g66134J6di9xQaSV4awJoeIRU81iNAEQ3Dh/C1B
MeAYh3z0VqHg0JPiJsl8H6q85wvBI+6qr0Q8l3xVIU/vp5C6Ekf7cWy4uZF7QuJ4Uq0P0jX1deg2
K/R9JbH4Ub8nrjR4/YaoXIm4JhFkhky2E7BghPWZ6XI3xuzg8oU8w6YwBBZ3YKqnmdZcteUA4Wnv
fvSulghDQrmqlVo8fWTI7N6q+ogBaM1oZPxrxmJoNycbNngwIozXORAW6bp+MZjpfS2jsOnsIRev
pMo9s9V/zTlZN8SJiFuRk6D7zKRAqZrCfHNkgbLq+7MYwMx+NbPWnfA44jz7mVu0s7N2wMxvsYOq
qGwBSkGLWTo/AOYGyIbH1L3LUUsXxeA/vfhAyBXP65BQqQUodA7oF+ZUq0D7SI7oBVFJmWRlQJWJ
ZIwJaQ7NebNhOzbzrbDU9S4QR9Zj+mpQdJo06ipt3cQX2Z5JBlN7AavTKbybLrySzwOulMo2q04p
9TfdoRTSNjbwzFE0LJOySUGmZY1kTaD6t5HfsCtklkZ6350HE3P5dQ5Z0Gx9xqGQT1jRvO0s3Ze1
55uS1P8EJEC8i/hoMmVYynkzi6Phgh87PGXecBT7cR12rV7kNH2IQvoVDP/zfZqAZYINWGZlygtD
D8dTr3KS40K9dE5ahQhPg7zWtX9IYYdRuOSXWJDJp1lpWvW5EGGLxDIKHGr/4gaWyY2IppUdV3tN
+jrhJBuHUBM89NWrcQ7G7bqBbcQ2seCGQ9A+wR4oU5MChN/84koV8BHrBFqNzrVT08GarU3Zitpn
4tyXaenJKTVsbh8ylEUAHsBbsIhtb5mNhcuu7YvNfXcjT9860fmIk1clpj/jToxZgeaTVHo4Abq3
ceivBl69uZXN1Ibs++BYKEY5YeHJgTy0XRQEbYU2GM/OBZn7W0oB+/mw9kCIosnkufwokIo2kkFM
vmiQBQgni32LKRv9Qh8lZtY4icXjKWpcFMy/A2Xyqx/Tj9IteilzJkXo/7u/LjWMRFUdiCFWkEs2
/y7VUyJ6aZkveAoqNco8LWTij1dm5F60vR+SR2jOEdNGTgfODxj+dSdLDBMJ/92DRZ/ZiQ/iP+r5
XNejfwDBSc9EoCuw7qF0/Ml/9AVS+8D+43ROHuqcT4jbZ52bTSDWJswB2ivoUoh4XAhlbXUjg247
hMBZtsd8/GbAcIJL/dNIcFOjKwaL3KsaKfjPaECyXyW7GCrvp0sgIm9zz3Z0xzNQWpKhKEIHitc0
q5ZH0b2DLKnLP0QqbBfIJ8nDFHTgIyu27fJxWbJNMptSm9Bqah3KT7adrGkvDr6/0UgsPdveK9xe
z9buLqVTQkS6W6aiT1m+wAo4MJURfONW8MvDB1HSOhf8GnQuXWC64jZQqreFMhdGDKqAKNYIKbMA
T4VQkFQPfcCs1uD2g0rzx5QstpOGyfwAnU9xoZdm75ks3lKzsSpAbwX8OohB+bKTGD0pTQzmUOE+
ZyKAoc1FL+GWRaylmwGw+ypIAGh9pl48JbhSO0LausgL5jAZ0X7+JyuPSizgZODyMJpLE94m1Rnm
OBUVGj0HbNvWgPg8oDOS92XSLKsRW2qU3riyMlrhNHYszaml+rqRsQDwy84P6kEKRU3f4flRAYUD
Hu2Udk1/Us6NLrjYQ+UDQ2rnisH9ckIL/cGAijTn2Cx8SuAzRTDFDnywxzGO5ZeFJGW8geBDzlur
4LXzppAqZnrwzbvWJ75187yzInOOLfHxCxqPklZn8xQLZJqX0Lh5x35EN/po+hWIPsaWqHGngru4
8JZxeLvUE0N5Mg8wKsMgQkimVmftdhmvxF7ehJ9pSALE4SH+Gm4zRys7hhYafP032JjhdCd80xni
uKo0oZwW0ClTS8v9sLROrl+YKhWhQNUWK0mRSNKXEGPomopNN2xJ+PIrw4JwIMRN7EPiYnakj7dx
sf+JMg9iQajqAr0+nCTuLSK/BsOXwBXmfteI5bNlIC0lDHf4wkG3yVeU+ddHSbSJvUcoLZJB7i/S
bMdTd5u9XqcVVtAYpJsy/TajvgXHHbuOFqKyspC+bULVNgPB/pLUc8KrpMURmmgTBghk5oZwCB0C
vZoTUsyMJjQnSTWAAToKCi3zc92rm55+wR4QobEP/1t8jtyJmjMUvLRESWrMvOPbslFRDTVz7VNb
g3nvqdAvdHaFboyk9RKyPxYbZRxBsjr1mfEgYNwQWZD1UF8yvIs52WnDr7tjGprllqle89qgqsRs
saBPQzUXDMYpMFqoaYUT2WSRwjZWNhLmFf4JwvodUQO7i19tNCHGt9r2wuEF/E4cNHx2vTINvVPU
5PyjRjyJ7Ui5JDV1Rgu57y9Da9D9qvUuTYu9exErtpExxJAHa/wKVKTGd8eqtQkY9l6DAZzP+kUC
qYYjSnYgyjaEywYfpthjXGzqeGi8aTWndOLPA0A818KiN1b6McMPmT8Im1wurAyq/gLipJ8l89BH
3oUZpEoJnH2yEcfqrSwEOVcgrH9OcUtpF/Wht8bKa6c76rrAwipaPU/qdrTFFJ8/YFiZZuhz7zUC
wsYJmF7FzUJmLDrdq1DzRj3QoFPCKkgvj0L1QjhD136EEC3O5VHs4ETV5wIN1HLKdTHXvF5IwyCI
gBUAFwuR1N1k62OBzLrfisVH/ZoYediJfM2w9G5uFTFNVhVv70tjCSHDt+OUic6SOJUeyckMdecu
W7uYu2A/wdrJNFpufnALp4AQqF44/XK+2E3dTDuV3E1Spin6JliwyMaF0swRehTb5f9MJrzT+dDk
ZvUAcpUx3TAP0ryqlWY/AebFhg91saHhdoowEu4wJzCJ7j24Yf6RstO1fX735+qiybYDJTOy/kR2
++jXcJ7QOUtyyfmJ8KN1VTjdDNGyYbo4tTiH6U3oGflEMTGB0tT3JTTlknSZJrrQLTzCMHWswz1s
70r/z7ubmBy/Dba3XDaZNANRP8YEM34gjG4l09caXeyT/Y8lLX53jm2fzzVrr0iqg9ifAWkLMhuu
YYF9X57v5uYSTejsxT2S7MJAgJWNlzDH/hr/MWSp7uRSs2zvsgpSABsRuBu+gAB4saybqmaqUTJl
LL+OwIJneN7lzlQ3bUeDqvbmnLyvpe2Gqtr01G3etuCaeheAHmsKIUh2ghxoy5sXz60ixRyhDQi4
2qHbhx9lxAUwe2yx+FxVe0oIYelaOwONZpb4QlNzBAZtwR3XtJOdScrQ/cEAwcFjR8I13J6xGI66
SZ05c0wMy8mIQyxUh/fi/FjqRkoHGiQDhZxjeMgweiJXXaOCveTc7QkMpSMIGNpA+tNFv7OFNGWE
AFW4fT6ANJvbadhXO9XQYgP84H06i8tNRm4vncaNEqAUEKj3OjtrVJK3jPxPzh4xRnfomOHNHXm7
t1T2rUE6XArAjafJL+fFBBVVELl0sLAA/AGdjIwjTgSCkutouWhkxH+DwiqHKJ4CFtFw3Zmf4ahT
1T7BsO/ifBHRAJIXOy6tZCBcFTPCeOcMiWo/Ec1lCf/9fD7sTDhjtuKk11A+2eM22DGFKWykFShg
EfGqMAvW99J5fcMGRfpGtgrbOiO6XQsNorFNJ+XAAUHdSWxfNtX6ZuiQxxAi8uu9zcHmyTwHHbe6
Jotq6+QkOlsjsVSm2uNSRJ1gq3VhQxqG0KdYJstj4nvEIr4+KAqqEmrn5T2Li+JXj6i3rbysP8J4
yLvx+0umrtROJcYRwPfty69O2qC+h5qhcpM1SLoOrGnpVr2zkIrdAhHFzDsZXsPnpYRKlIQ0jhrE
SA/Oqs805vA6iqoSMbiJyVm/pnPvEe1Nzy884LUR0x6UNTnsnfpw1Ej6ALEuXtGg9moKBxu3DE+p
O5DJ4TrHpxBW/y8mfBEUg3TPl4n2BU/rRKH4Uw1ceu5mXI0+WSyI28TMw+7OS8EwHhS7WsEQcNXf
pUzCOS8GNg9/EPnEHGgxWFPoQTIPW9adaCEE1WfCWexWm1htIDTDEgST+UMZ8cQgKG+a2s8e8CA7
QpdvS7rf7QIDtdtYYMLUUmlyxx1HmfgbiSqNvf61aM2DdqtZW10E6bxD1Sid5pPA0x/wb30LQOgT
I1SqFSmyTIBPiFE8ED8zJ7m+diPH6NI62EBmBo/Lyvj761MUZkdiddD6iw21uUPYf18fJ4jjbJZv
UQIt1Myuv09A7wlsXilw4WpV71wZODcdNg4WakoDoiFkK8B7lPbJMeYZr33cLaTpA00cM3ryQJ9h
BVESK26KcOYiRiSEmaQxaLHbWwq7DZjHFHHacKzaoB+W+wTbM081lSB/uExYEuCVzcpiLOnmRZwK
cfN4xB+O23qWtyIjC5P+FCOOoi6x0jJiPAxPi2JAykuddUdhzri9DL++JURPfGhIujc9fvA44eHa
cryZ5onUhAgvNPCf4cPusjAJOB5DjhGXfl6S9Lx90ne09IbFbSPH8fb121R/hBLui5VJErDUOJyf
C6cozNrAaBWZj1ZXTLUgH7ERAj/KXsS+G32MO7+svkQokVHFCl788PJplhbPdnLASioOx/j5rK5H
6uaL7I8Vjr3sjrUkemjQPKstaFe/4YElzlDkPPylYWeFWKhJ3gFhqgknQ2x1GYRa10P+Wulub8ky
T/A9BhX8xi0Aix34pHLrZoW2yDOivVm+bs7PkfFdhbaDEMCGfcEzZtsKrHPzhWpc67vMyQ2j5vY6
/HIlp6ZegbbG2q3XMJ09bbGMh6H9nkwxbWMNoN/Mxam2OUMyapW8F7r7ScpJYc9lNwMISs2gR/bm
5X4swQW7p+6KX7GbYdzCIZa0gYJPSbf6QNCH9XjlgUI/BUxaUzYLQfdVNIFR9S/uDzmthdOly9XJ
MSQNVNUSJ7y2BN1hfykV5Nlzg8lfLOb7XMJ+zLQfP7/WI7M9+XQqFLnA5VMN/aPfS2o+ee84tMBY
aviqd/fDWphrO7UqEA1eILE/hJIBTqUx8J9JpHc+BbGs493OttIiFWdIPmhV3ZsHsmD3eWMyaysd
XldfezafRGGod4zzVMxgx/JIU6pZmsuSbRwCpSKvgSIi1rdSFLSl8SJ5Pva6IlV4wlG0hFWkkxSn
C/imkYygP4lIuHhm7wHHLaD0DI4hi/n6siA0oHvbU5D1bZQr3kypdYgGHggtyAPqcufgQ/FR0Nei
TNidQenYhYQcy2ZFEsYsakve1smZIWmP29yteMRMJ09egcasLp+m9YGmckERpZQ+7+f97cZavLh7
H1f99RFxP7iqBmOd5Ig93P5D6S8K8gg2ttfGB7/ts/BPgFTV4g9skuP8p8+7M0nfe1yslP/av39k
RvfVRflnNToTM5ZOXpNstOIbnUWGGzu2uLoBESZtRINI2PsLTELGOqx2HWNqLEcFYgEJ9hdbiuhP
j7x47lafPoeKEESciseUP4wfLJZtuSJMyz7W8bHUi15GfojlxNY/HqZk9NzJCUY2vw0Z0jWOUDzU
5aOhZYekIh/iSJSqeIIWu1Dx0RTcO6U/g7m0PlY3hMIhXfrTRO4uSs3ESNpI+ibFRQ2eG5J7/7xs
GgkJPLtrA05EclJAf9gJCiC2ERpMPJ5OgZu6aLVZvyAboJSiZpf0iy/5DCUsR6C+4IULuD4dqGrK
1kSvsKsrrmSdXLX3apGhXxYBz2dWPrZzmosUUHN6lyVQZCZCqUMp8Aw0uDJP9IT3+uOwK4WFyXoE
UYTXCys4oxkt5k++Jg86FQSsnNgOaZSjI1bgSzliMwGlNz8wyXajKlgiGlhDShmd4hXaE28KQx07
Lr3ezh0edQXCigf+rYUPD4DX3/CK2iLkcuZBB1jWUodoJeWgFsTpGGGgqk8Id3X5bjBjkQhT5t43
QdeHRHjKwZ66uMS7lLgxhpBjW96tNPgKzx+XCaKUTi5Q+1ve/xxxd4PGHWj93Yv/1J65eOpipkdC
q7ap3I7Ey9Mu+Y3ezvvm3NHslJ5lHE39ZvVjtvIa4230CQUm89EFlVY02S7tQkeL9aKnpEIFvsc5
cxwCRtNNvsQ51nGEfEYJMSVgVTp0Xz7aQR/I4YC//7S2rJMtGeV9HgDNhW2YOK4w+GbfKfDeJrOB
NjwFiw7WQcwHUCMpUZ/4AWV58hil/AbazYUOQLVHZwxOJ5TTYx5TnUvnpkALtAt3fj72qUNYHFxR
H7x3qhgS5rqJIlEeMRUe2et+dcpoOSd+ZJ7alGRVDS1RBZ1W3tKocGUKhewnZ1WRksoo8CNUX3HK
kQ8c/cyW8j/Jg62vMLKeYsiQgSWZ/deEvbhhhHt6wwR80zb/vQsw0eum8Aim9fsHbzoWTWVwVhgW
oY2Cftr1R8G3vturrfc0HlEMZugnBzXYcT4iMHhHaEvgvswENwKI4+1LabAKZRIwPG6AhflJ4Tsh
K+ohoLt363yHpD8bYBYg9fg+dgeDQ+f9F+uVdLCqeZYYUYY0VAyyoXGDiSd7+pSMpg7yKncXMGEv
AjX8yulP0w+/Zt4crr3XnxKW/ak/dUbwPgOIOAvzXCXtq7F+7IoB6mFTswUlclDL/Otb9Cyn87tw
8YieLjRfFADqlKIT8TFVq7cPTI4Vd8dty/7Fn/cePJoon9U2vptpfEYYwyONpmuLlZVhR4D6Vnml
Izj2bGjAt+Go4Pnd1yZf0TTIgtim6cWBbaLcsLgAizwtxKqeflso4sy76QM/wJsLFUfvZn4VK+fN
rXjGOos2cTK2pkGEREpwNvghPGtEz/CVbsJeE5NKoZ5TyfXoR2vDH94VyylSS0xTIutPm0nUWYYw
atTKbh6TJHUE4/wWPCvNeHl++J63xUShwDmYpxQBjQMvMsyfwWkMFifW7hvRxCkFbhYYL13kZS1D
REvaq53UE9lna2ApFFRyksKxa7XNILW8fXdCEouG0nyns7skJUKE305eddST3K5iQkoh6KwxDR5z
osho2Fy6crvHJyJ6vHbkXmj9yHV+8Xonhqst6OWeadEeiWJWGy52pX0njxDVUqhBehHKWW/6srpX
cWMFAOptIOzjBScGNpLeD9RsZBjxB+tTm2FJULhoBkG/7qdP/tXCYIBwkKwEkA+R5ryZ68QnIiBu
xi6RDqko4h+EgqO7G49M9HCtDZs8PVKUFCJkMU1skxSeDl7EfLfNSpHNljhKBBOsk+AF82I5Hq8N
RHcmU0hcAa+Yk1XaTfAEe7dQ45t85Q3grrIdqwLM4WTN/46DpRKRkqMzg1/00WuKZoZ8KW4vOQEc
LZ364wOhR3EY2KJd3H+/YxXRslHCCXqCrJx0XTDLPTvXqCOlWOpa5Qnx0F0C94/9tRjD/oqEw2u5
QJnH6RPNZX0ptE9GXmqb8R1aIOi9LYdkXyYWQLt+Fle8euYvKcAugziacke3VjmEwQbsgeqhqHYm
o9twDvXu8tC1XlnmwNHZ+oNgLkLXCuMGfscXEB2+XX0Xjt/michNCneBS+J/cmiMSaTWqX0I57fp
4p6JoelD1oqBUz2BfYWV4oKM6rbHy3IGeTYHiDYAXXVE/K51hct56Zi/53RQx0dShlUUNzkS626A
I/a9btgssZixGxmyVcJlvVlJluG6T7o4a6CCM3IdTGbXUA682uboC9+6d5R+30Mc3+PSVTH26uSY
YOkwBP30672sUKdvlbGwxmbHnQmxlqYcJno0vi+1P/aULU0VKbyxobQznR9FA4VxqQcyVhkY7BLM
GMiGby9jXChQg7C214rjN7ucJI0/h8qk+KgPA17UVBaHaRehcBkn0LsaqwjeYn9gguxpHACXneOg
xc8HjKSZliyZFtNlfCLXkZEIIBurxD6K5gOg7/tKtS58KNFaQJR3+8z+y5SQwCwht53WJgMwnJ9C
V9NwmN0DLF3jAk0gwMIS78pRDaySQ+fNGR//uQCP3LegNCT84QPd+yGXLB/1G3wOEuYEHx+8UzBU
LkruwZCGM5hcb53uoxeVlC14W5q1vmoaMV5IVeSwPIxp6H/d2oF1WMe472FHIYB662dcFng+xAMB
8lG4I7StTmllj1E7BqddJqgk5hEeeDpfvIZ8mZFK69ol6PHW24kMpKFME7pofJ7Mvs2BKH9Ggvnv
FAqye6nJr9yIk9x/Ponl4H8DYR65FCxE4FZMojsmIiME6odvaJBh2cmHbScBUOo2aK+JioxwfXSg
Tn6LsDeyfHRhOizqJW6WYoMmVPJRcaJuac6VigN5rzRaz/CpHuXhsjNSY8KeU2LVp46E9bT8Zb9p
FQp0wIOO8rjKkZNgOhPTAJwlfEOSlmJB4xCtiD+KtTp/nMxDxT+5V+BJOhFWbmTX4tQ9Aig7pP4j
j3ueMD/ZjMG2gtjzXvN3nYL95kWLiFCMYEsf19Z0O6WrPHRk2+GdT1hVgN4Eby/qkzKWgm0XLr6u
X6A2p0sYxS3SyDCV71q/QKMcmuMtsvaAAkjmmHfA7n5DdXzem0Yaw+l5fMnntcypy52Ob4FEoW8W
PJkPV17ndff9Zt0J34SvpukdhqsFHAPo724Pujwnub11zIcY6OnUHO+5oL1c/UMNr9EjZJ3or+oV
pFaLdXIiC5GN6/io6CfINisMVpHG+ZWtUJJClmoQ6FDPJAT6ETuK5Hd7E+hJ7I4lP4BlKLk5maZ9
w8OFVH2ahbGCCh8col0gBOB58zSrLmbH+iClJWNw6YxaBGPT7jWa4AaGJzevrxu8Uc/ZAETNgDu9
jla5Vrj551eFMXS9IcHBo0ECst/9q/jNo+9hs5Dgt36cAA5OmNYDWjxXZXWkO0TxBXMaO8fljhgD
G77J02C9qkkbxq4SAL6AgC5aYAk2xhrAKj/6weGPt4qK6QZFyJbqtJB1Ao0MFqoEeZY1Zq3rYmvg
zuA9ORgmKSEJ6RZ8um5sV3geXmmEbjiJUjIe0u1IIBEgtW+fykYk96HhuNXsQ9DpmDYZ5HkR7fCf
Ccdf0JK3jbJ65v/9PnXyvU7m08SmArBI9sHxjEoY+RU69REwQ0BUaFh56DvT3INmdkxUow4VGdzk
RxOPIjTKdRz408QsxI2oT++Oi0i0yYjOraIoUfCN1+D8Q6cHenCm3XlK9MYAAxrYMnrQBeNwoDzX
lehvcPfL/RNVgr/3DmVRYKA9IDiOCbbo8u/ihAtkSbhWh8bx9yDUBfD8kK1cctIm7c0BL4K3VzW5
haAqI6bHIhCKm/5ESykphJ84DGXfUUyl55QYdwir78VLkiO7wOGWlY8B61B9ALy0icT2sBJglpU+
7lyuGW7cbLJC3Izl7uOTJEYWKRGZ4cCSBa2hqXGhRYJDmq4LX/KcfyRhQGY0leU0xStDK3wxD91t
ts5hqLNnyrmpjamVhx/cFPlH8VSv4BK8TzmRqTcHgxbQQ+gkRN1ghhOm3Qg+Sn56FRS7oQcwD3dh
gLLd+4gyLR1vQYUwXvoLr0GZ/37wxCw+BnFZspxSf064hwuSqCp9jdG6nLGn2ZsLqWlAbLoIyp8a
p1vKd1VhdE70XBYYGDRgfjEo6srhCQ9zT7qZuCaKhhCbuSYuGT/z3GHEO/2x1SqMqtsWhV3SxnN9
OPlHTiGKGf4Kd5NWuhDvl31hWekcxPXz7wHlsXHJEd7zL1AALelqctpWPbLTvFPCMQXdhq8buNjJ
NSgb7r0lYpapGFLrKghsgDrgYWi3VR7vTBNMVrEzbqKBkqh4C3IqLsGw5BEIp+6ak3jiCHrJ3JPp
ij3HbO8c4DDZHK6PS/JDMdrtnYQnBDbzBOF54VvbAIZMQ5qLy/oV2uhOSOKdUqEYjX+P6iqEWR8S
3ZQZE1p2KEpikm3R4xX96FtnSHL8KQYMBcy4vf+OTrRObrK0MeOeHnb5vQ8qvzVup45mYe9UqAQ+
Q6xAJEL3VMTCiDb78HmZavjnWFezAuFEsgGDUBQzT9HiUn90mCEqBgHjEk0BVB/h7U/NF3ZS0WNK
2QBO8E4FNYsCtDOUDDkpRXr3DqNZmUk+46o3PQdeHs/mAovFcYlIXqWc5cOcI1FlfxEMXtzjlCac
t94u3L+yTqO+KJNHYtg80XlhDAQf3AYtB1EtjKa2urC7uz4doCZ60wZZVUVMrlCzhVOGTy2IvoRw
ys01jgVpMasT86AnieQM5U6mPqvX6wDKyqziTIz2NwO8sY6+w8fyYbjEUuq1VhQpquzPVQjHa7vn
naK9zd1LG2TtDSo6+YHbxHBu1olRlChjk60ZMSUwoAQiR54t2feejIbjvszKClaSGGNNYZ9bOhgR
5qKzP3Ja+n3XphAD0EKmP6/uZRA9cdEzJ/x3pV4J1uqlNzb0B31dPxZbtQ+Ffw5f3L8NJ0iSJaTd
2T2PzrtM5VIRigUzjuMDiSJv/5rIQSEZSGGlzKEy2qg6Gg7blLjEjCINlJkUdvoJuEoXt0bOuPSE
7io9whLjAFscVZRWybOp/fg11iiR4TFFihreNvjmz9RDPXh0haa3ki2gIFfYVEg01mc3htSz2dL9
wTZIWztGvRcorgDKKNaIgzGZiP4LfeYJfi6SdqAMJqUc/gryBZ5tZPEVaCXId8CFEdJRruK9xvR+
VaO/6Fyt2oUqKfddyQ0FRPskQBxHgPuuolKvaxWi1ciNIQCsrdDAIo3FS8k4l5itKYPHJqz78DrM
iDsWiYqAG1MTM6m/HntOk56lyg8nhW68BHxN0AXeNL6/5uWYtK2LBpAEkS9RxS/2ddCfFPbvHb5r
plBGKvQerX3D5BdDQfHxfMHjfoZXeb1ytGzLPYrw9u1r0YqQPYJgGbsWleS97Th2c1f9GPqROD96
nzQjfoO5Lxb+VZlPmPExLT/+kilyol6UGt0Es8LhsJPqt0UsU0rpOLLX05CavuxnM7T2aty1b/Xh
nRqyHHcXeemeIdU0QhEXyYhQa8KFDjpnFYp+DgMXDD5MNZHZRsOQQpV9XBkLslwLOO9R1qTt7mMo
mhqITvtx7lPa9//I3s6oyfw3yVVMdCdZ+3gy/AFouwKNBF5+Bgp/RTgX2HGmxqKQBZXSDQT7U/fm
Lb9E0hy8Nq/9wKegET6S8uSc1iIjVJN85m7hx2tj67L0uuk6ZnZ6PwlTKKVxrXbdmxYio8gtbJo6
BkkOYHoiOurNzSETm5ceU6ak5au9gsExhIEBqH7Vs/a9U/BU+pC6pNPGFIQqAC7VJmzDFbpDXl8f
OhmT65VA1Q7DCIuAEbU1FH1XRSjgpAW1AubhKuEKmwjrhnoOLTEIkMfgIkubKe1RMpnDfXpXur9V
wrYLju6DUrS8VTG3cdDfE71dtsF5ERMjsFOS0l29n4i+tTqA6PesIbWad5am6UPf0+OP7eLY5tAx
YIarYvaUqBy50KYQIKPSAicaUXC+phhxhaymwF4IgsAPwNYYq76g+yKm9bXvxdWmp4+zoQfwuAZ1
F7pFaNAG1U8jslPbabdHeSpkz4d45gkDNkI1AAEVz97THP5Q4Sq5gpGNAaqmnnLoxGNsxTa8z3VH
0OldgTshNULkGA+tD71aXGZmyZl/00aIVC/GSoNHIeFgxb99GryobvQlE1kC+78MOKCtbjxT8MiK
GiB3SaRUrqD7zmMb3ussV73rtTztzohet1dRLv7dQ4TWrcbVYmx8e9ZmHkCoMxvdPFxOrrcnRBvb
qXzFSQoOVvcwh5tsCJOT4cLmm95+u+bF/Gan/w7Tn1adp0p314Qb3WYqkKtSr1ZMACKPFn9i9q5d
7ZYYsbWk/f6iKa1X087JUnSE8ZxQsBxkWJIVNLGOVIYXAtBXjzVLFlEbk8YvdkfnGI7uvOC9WiZ7
ml5bfsfPShUcanmJsuFMQhalLdBFbXcabCUAVu55agLu61AN6WC/USDkpMSh1LZ20HpneK5txzPA
WTu3vbajpifcXzG52rp9k/ApsAxJqtOTDY8ce0wTNu3ezAk/ffUZsRI+vrW80qOAQdPC1kRfN9Ic
JefCK3G89XUlCGuW917ij8A34JPYCP/Tl8fkY3N0yK87ub09bvOQh2SB0tsU7Sqcbr2LthVtOhz5
2PFIDJ0qEmWe5qSJFfd/JfCW5eIO03sAhQh+Svi4YmRTwu6YPlubkOo2qToxyI9zkLuzmtS+LeoJ
Zu12Aqoz0jvG1/r4OjZVNcQfksKFlCWj+x79RJBIPDVZ28Ipez3/575YAWvkF1lHsygqh8hGBk1z
r36O5Co8LrXMRNa/YdEmNfPlyUUS05ij5HFBmPZChPhWEVsnqBTKcRSGRD683GY/fKkDyDRRd0wP
ICyPHjEkdXAYvkjH0masYjj0yt8nbkZFfg1mIaWEjLGHJO6XFf+ifo6lMaa9uVe+KGUol4XDtk+d
qpdNfQqHFpES0ZMomJklovYuOuy1+UR8ro8apx9qngJ6TGVYdZn+pTadhsHHzs6t+EBi64wBdE2k
SUq6Lx4/pyq/Co94WYYN5+lUoiS+t54XaafX1HRHtLbJmrKewIsWmdrZTP1O/6ATyC8BqynwGoH6
zJetUQty55dGTQY+ht3Irvl9W7zSD7vdZDVlkZzfI3NP28zRjwFVKIEJxP7lt1vuzpJNIemFvLIu
lndmfJi1Sx5XfpjlN3keTX0A/FHk5mi98oI3R8pxHA5ZOzemIsMlN5UNubKCq/Wly+Acsqijuydo
tZSC3kP/TAdgOKig4UKvueNdJra7GhRZr0KuvqNZ+ieHDiUgaGZ0Tgg5RqO1q6Co/dEBZSX928ce
fmOwqQUdFdV5I/9IJF8xSYkNsBl/Kc/MR3LVTOb1v7jeK1YmnzxXaty8YZwuFTDg4doJi0XCWiFo
E3G9Yqi7O0ZKLlLawsf/MrjY5f8hDidOVN4Hs3qmmSaSoMJd26Y9grhYdiDfykY0tNeCrXKbhl+z
/j4fqFFjNrKNt5Wf9Tdp5AVdjH/vypfoTgw93gR6LGsokK6YvBLcNNZHAB0m2d4RkvMM8ohX7bfM
I9/+YRY3jS1nUlRE5nTl1Ujj9TIfR1sQGTjVK6qzt6iEGna6OHD+Bnpvf+Zg7cRfnAF+OoYl1WZU
KihJlSfe799pTk21X/x3pTGD7At0xdC1iDgJyjdMFhr+BrKT/IfmRwth1p/P7djkM+jsu5NeMoWr
a5Fp86hR/IGgYK+vT4lPRjWRK3xbnJfWhzVtmOP6j3XI+I7mEK7hjiLkO4Kaxy+NQPo/GUeIY113
Fyho6CgiSlfDcJzigPAWg/Wj8BSwCrOnU2eoK6RSj0p4Yie1wTZ02N8pT8moqo1oNt3+28G35Qsr
3T1UE/oWMzz/6DCV4ipkRrQ2g0NiTZfPUlphAPNpwnGfEYPx+Ni2bEogp5rFfZvCTuxRnV/g0Bij
m7SRXVS3Rj2GOtxKztK3lyXTR1BDFgVvkOQPhaA1j+XUO/z5zcFunwshFOP8wr7xHGF849V5QmNA
NUnAgGo7ZlNm77qYqdietjGuJNOMDUbl82phVfY71V8H9Vzz2Xegx6DprJgmGgezHoZMblsqE9io
LZ7kBKg94cAfJMF92GfKpov6Np2w7NuzjYInNOogvkuouyON4dZvRHq7+lsXE3Vy4eFFuoQC/oj/
1CE1ZgHwXpsoFZYvbM6owUQnvL5aa/494gMoYfv717ZeRbWAexPFyL7e0rpWA6tAXh7Kkvz7dFVP
DYFrcxh9D6pS+Ge0M+vVGUdiDo0SoVN7sdhilEBvyvMav0uml4Ql1+MUhSHCSa/A5gHVQbytu5ln
zC6hv+zxaLNNdk1rC+6u8Tl14gKgG1/olzkVRCUdHSBtAWt0dFF6AG+7wPRZhRfZvUA5SVQc8yOW
/1idbk7IQH2E1pAucRCfWvdR+UaKq/+w6WfWA/0xB6DMMJNgX6qt64Qu2KQuHZf7Oj1o3DNOrtCZ
7fOv8dBggv2ntfhVCleYhhs2tNqs6nFkpubTTs2yANHdPeeQ/ZMQJBbaENutim+zg/uRUWGdy0vn
W3/Tuvek/Z17KyoxTxDgd1B9+e/VCeLBHKz/7gSpcZvP5Yzpwcbl5Huy+DGRRTmQHaM8PmIc9pOA
11CinrIPlGKpnpIvZ6uAE3flNTGvEorF8z43ToPvfMFQzBEp05N/tEx9LBMaZvXOKRTi3/u/yQTH
q1PZJoLdTw02FGHVeuXix1aOT7h21uMztY5DTXSbvRWxF5iI/PgoBAFPNhRu7C3WJ/1QDtWYbA/2
0kyLXgzbOp8nlXZ0zTV6Nb3b8YRXCsW1TPGgzMyBYPDEGoRz+TP08soEqH7x0FRhTpztbL5CUglH
zH6GW/6LPvHSwxPNDCmzLx5lX8HBUY1OugBrTqsGfnP9/jB0JS9cLY0KsIyjbdE7/cEZeGhDBA/z
8FwxKqx9SnfLt2SrvujxG4Ct+hil1R0eg4N+k7hdI/Rv8AoFogTZbcnVZ3g3olRHaso8kATqUyXU
GlpKdgehbH4QOQM2CSIPbvyNiJhfJc90bp65GSxhl0k0fFm3lZJgcpLrg2hbWaNhWI743ZXjkfWm
zrMALIF0d4oaENvFc7Ct9nxm7g6QfxULczFU7AZVPQ0bg4SgGYbBCVvGUA5dTWI9hv0ybY3ltDMG
vTo3cvS9+Yfy3zsOr9xo+hbhzx74TjH2LnCBgoC/+ZhSZkxeGTZfZTfBDDBhBX0Oh444PL53WOt/
PstQhRF9HEdhwvWvJzftf+A8PVf1R0CS+jxeEQfcZLZF9sYvyB6s8y+7l6Ot9LImQ9ZTEFrU9SBA
KkhZHC1Fu5kB9xKIqkdOTPmuu/cFzXcRcvgbgaKgxuSQTkpoH+JejpzmuMx8qryJilwTueC49GQN
Duv+/JrvBXIR50XqIA68KQCMr4lZVv5jVk5v4yRMnSiburGw8g5WDuQN61shILZRQ2967O4Nz7+a
oroEDFQ+dRHEu6oOx9A6H1em55iUjRGQfLWJTduI1BUCF3hnk4yLF1J0wbiaggkVzyZUaH3sEv9t
OlCVOe0ON5PhmtWp8ikUAQq4sJtC5On4WcYwuhY6EjGXjSSiBGxmJCeF9yWwUUGH78yhbtxudYag
MSppXhnH0KaAA1FnViXIdA6GNPgvH/LEN+m2ijK9Ctavs2NwdPasWN6UgnpOH78frGu02fVN0LAj
A6hJb9HOX3+VAm3Q2vUNssisaO5yaJqLCFCQeaTDY50Fqs9j4FPtXkxD0OIHDMCYwB+Pj7dm+ii7
zq/q6yrMkYFuicAwsmljxQlW8G0pOKq1dvlDNtJxK9NQd0ZD3bbfIJDH+WIdglKY4mUaSF08Hjrm
/q6SXcybFOghOrX2yRJgL5pwkhX9eo6SA+vYcwAtNmsCkOiL+kIWMHMtgnNyRe1sdbwmuHj0UwMS
q4nOkoHM0ZS8cuKa1+uYLIai5oo7uGZoRWmr3wdvQaE7H6L+bqs11RBUkVyAAXuI8b3vErSVwtbr
Brt5Xy3kO3+jERUFx/sLZ6FVrmvl0ljbVJWV6Bbjc393T9VsajPN8gnLaqUZJcrFvShSXwChZZz7
IzEV3cp/Ad8tOKBvt79eNKZoCUI2nwhuIhGHYbO4m1bSFIcL3lQ0659Diq9i+n/Dp2yFx1EJMZEh
vDNLeNLm06jgyRxadchd/eJHXfQH29OooxHxNYHMoEfGDWvd1shskxV/Mx5kl9rbhGrrnnNb62kv
VEljoFEu+FFqtICOEZgf0B/vesXwysDTM9KaK+eTI99WR45FBi9WPy2J01Y51MvBBjzuDQqYm/3P
dmq5PdtnQGkWoMXWY44QnLVw0o9rimxNEUbaWYcBDc0WAmjoXkql1+FzZDTv8ny76x1l5kBHKFJ7
LkK+bohZ0nxC7t/EgaGiexFIBsy6Kgh2VaBjithRN3zIKLJCbaxADao22ONhzrNhsqMLBCGzIRmI
gtQquIGkQHDLkhlGIm/wcuKHD0EsCJ8KA55ExPlcABCILagmw2iLoeKO+LYP0N8VfKM6KS7yhoj/
E5pYj3tFm7HIDcZtSE7lbJZEnTfmCCQzAsaCytjZS5O4yo/3mAtGY8Yw2zaXaDC6NDnIvgL786uK
s5fuZ45aW8RqqEbNbTvWRimedwMRIKU7p5MyWrefWjDpW3VN1utvw7aWoxsLO0BGEJhJ1UAAcE7L
J6u0eiLqdOAUCV9woiWYJr9swTZSQUVqtG/2SACLmTEJ/Hw0Yz+vBNWt1fpJBz7F2xj3dJeosrzc
0E5tUvQcRFgMZML+PeM+EgV2A7UAqNR25lsScXOIARcUGo2YnYWoPhfr959t2GknVkUeMV/WgozY
LMrpzFNlFeQOfkEZBHVAU25DPQpK5q7Oqge8GV9LDkI4am++Zz2ku78aw5kgfemBJNT7rL9eKY0+
CQ934dF42z39u9vjkNRyNtCrnvRBGOcc22lj/nSHo6bWChQOM4na4wR6id7HZCChllLs6B7jGYtd
xEUR/TA8ySKxCKLr8XP2DsI5qeVNXREAU5Ba1syXFWZQIXz0KFsd+y5Zc+8PAvvSCg295sGOpNGL
Utq2zmo6rGYd2UCOzbJZXEzUN7E+w19JVIFeiCgTfEukjpRll6lBNSthOiIwnenQqV9RTdrpyDaT
25ZDUqVmYuzvh3tIx+K0gqlz9unOdEB3yfUsXRmD2oG/sRRkv6z5XM3yafAYYNE122JukFMPkg+m
GtgW9CwwNQhBw3x1mCiJZwOcja2eg/DxY3pJM9x5QHSGf4Mt9/TaBZv8RS/Tt2SNSbrsanxAQHfs
CvxzJzWUFvodxQVs0JwvcK53NMMl/o7fubdzpvfJuF+OsRkgsMKNOenFaHnE3PZyZxEAr1YwzWba
AR2W68XZ+nPiejDQYt2FfhWEt8cdtpMuc8NgxmpvhoHT9H4v5eCMhi6Ing9eUhRD3VYjXkaCCPfm
VbzW3VycdHsOjuL5kJIV4ED2K7DTMPA5nJb3/pYCueFevKrkLNYyLjfvKO+wIiddyyGXIwAVv2zG
/NU4OO7igOMBRSjFma9FVrVEmMSbTcU2/lHbWGmILuU8tr+V/uqj8LzUKivcKhpvTZNZPiWT7d/X
3W546g5Q8pEOPqpAueIhKdFOXKgbw6K64qZSnqU0KdDOOIWtPp3+NvCBZADuu8OfhLJ0/YcDREjl
PkkXa/83kHUywpvbBIpV2ujeaRx5XazbIb4L7eAho6KEE4MB4Z0p1/FBLei9MalbFx7TnP0PL2Ox
588Hydza9+SSbI7kdXT1tMNN7JR/s8dUgPw9Oea+4NYRfF+sAi5qSXara2N9cMj0S6a8kw+JV85d
NftU0NeWnoJRPwQKN1X+DW3ybzKmILL0C4PxQj3p2uBFcQlzcvRDMjfV8tQD/uxoFp17RMKaeIrl
3JQmJx7BRHhTsuKZ3GfN/iY7u9kw2VM3XZPCJwXq/eMIYmztdqXt5ps9XmYXAY8FyokNy31Wmdn8
O6lZcJeA0BjGPU5uun/Z3iRwXx0vdxjQS4ODiBx7JGV4Nb0IVZZlxeMkCodAx8vvLrVNZgMDZC94
DcTtQ5VcQjZjz3ksPPXbKY3xfJKf9geBkImR+coMpSHPh9TDfklUotfQTR1EUl0Qx55DC/9ibUHx
g/IYjVXoV0BR5PRgrNgSCMQdyHzD6k8Mu1l6UXhzezDquKZkDkfMzmu4g/Nm1/8vBTRbn7pByPOb
i+ca4s25clrVkg39ikA6t6o5ZPXUKea75FDLUa8w1wWfd9cO6F1LKbLPKYcqpe8kpCctfJ2dE/2u
Ie+N3xbhS9ys8ysn376iTKfD4DxnD2pDR9R2q+Yzmt5pUwaglqHrLy/mwPpTo4K5H5mLGtXKYwRC
Y4DBKVKVkXEZ7NItkzguOLYI1SSIkRGzJis1v1rv9hvrIgz+y5v1osSdr5DgNWyQnPI6cHXdqQQr
OB5jxiZkkrm6z/sY0iIdkdwemri0iNwUaoqCZY/TJMvSwjSLMZqfipBtPpsRnOfxG6U2IDlH8o6M
FyOxq+Eu78P0xMXSf0OmQrp9vDFxOIYDwRy4roVXOPm7XqxM3AuQhbm/hMfx1CmxZPUEcQKBD3wq
zxb+SpRfzlN1TSCH8V6sajtn201z59BOJJ99KegqDQQCrNneo0CFBH8FUvNt78jcb3JtBwQQUpqa
XYKItEwJK1KlIKBlM8CtrnN64pFeNCGsmZSXgoioT6o9qyuv0EqS3vi5MXa7JErxA7+UyBhpxBjT
tcfzU9aPuPLqWxfE9b/scRlI3gMN03zDuIa+8kaDJcy0gOUecAP8+KMBEYGY9LzlfEhygL+R97AT
xaQQMZju5Ew38I5FBcLspTHRkFtqGwqTyyjhTQBi/qF8GkPFxflRPFk+o1DUWPNm9RwbQP6+1x/H
ZfLez+BmBQCnxWx4jbF5ZNflnld7TQtJ/sft6wJ1pwRQ8hnnTwUvdBfc46kkVSeSBl2ojavoDb/b
GJI/6l6naTsICLlpDj7RoYJsnCXNo/kk8UVuVZlB6S9sdQeLqwnYPDMAYd7vM4ii6blJMRKUl3rE
d0U/L30oVdukbALdH30uMMZ+ly9kHU+UJOjA/Gnlx+rJwoHhJUdfYdFUXbzSErWs/OdL2eRHAn50
VZgcmdixsZytiqhZRK+c4xGM8vCz0DIgX3nHesAHi0ei6T7Hv36SfyqgrY8H33p308CkKl9NzDAu
SIXiOYunLeSNeiWEBFrKHJScEGp/IdxbpU4+WZDmw7tZVloALf+8a0nvyH6D3Hf3jhk65ISd5CL7
4lFKOixnthnXYrk2k5MezBVOYuaUSw/A8yPlIPM0aepGtO7Ud8gCyap9s/3y6jLcXtf+hbRO9+mi
+moJ4C9pn5BhpqtEZaXM1A29Z46ne+0WJCcwCZ0k3gTwnIkBPJglbwQNbxAlgSeHjjGVPRxVMTGJ
jp1gK/yft0kbQyyXuBSvCZyC3iSTw9cXxcImamNCSz59rwQnAoM6qdqFK3q7you8dHG+ekqopgGy
uq+zlHg3XC8SS1QRqprnQ2ad7cpSPs20t8BNbFaUbT7gsI85/NjmegRkXhMcK3CxjoPfTjdXaCFk
JVnK019guJPXgMhTy5eTUNPqskM4emgDhbGYG3b+gwaGKZsMIgZn8aQZ41P4+2pSabB3DUBouHg3
aPQyeEkQTyyeYbffgR+9E/uEJd9tdwwuCu3COc69pms65QQ+OuYIXL94IBJ1TF8bYysQQU1um9WM
MW38Vr75od94y99Ys2a6Jvm++NGuHRrAqA9zAvzEwMbuo2iQJJ7XceVL+aFUCkKbB1ZP6bOs8IgS
yAA2EK2C9v7ToIJZrCeNEV0E6hn1iQpfRsMoDq+nav1KQlXjYmzUtOtCv+d0BRWB6GRhnx4Tc9JH
ZBGxyZghNbllrHfvwJY9pw8PHpHCwaOtZZnDyy0fi427ArMxan+pMZK1nR1rPsNaGmAtXplHe8Gf
S1iSCoivsVDGd2c3hlQnooqPRqMGLQmduvnJclU2j0c80k/8qmu6ov0NzcSOI5gLq/FXb03XLRsE
6T+ov9lVEFHinAfZ+56qLCltQgT2kotp6YxG0nhqLAdX2pA5uiq26VZD6qgVN7wF2k0CPB8CSBEv
ha0UHMHVxUV/9WYt6vupGkbjI+m9+z+yqOS+NjtkrIpYZQRyj/W9supUSvVYA0XIbUkJ1p4NwSA/
CjysT/XLf6peswcUtmXMhneKRAS4YEaJsSglOQermPsAJXbyRSXR63CmonC22uxvvBmcoRyX0svt
25zxf0UD4afske+81vcsW/tv+pluY1YGOyEIs/tTi0ggIdSLMOf2/dBq0b0TZyfB+Ldak+XMGWZ/
BoxH4XaqA99O23ePRQITahvOMDGONXJVkTgfxWIffoZNd3gPrkaeYZP2wcUpqKYjO+6r2Wog+ewW
tnRw54pA0TAs14EuFq0UCB7R/zV4i7BB8JPlzafND+ZmUrcM9YGOUz8r8udsywmu8UV4Nx6JPfMI
HqPGDndKPdzDWl56q/6T5W3YvCfRTbvdVt0mj4RxT8hT2SvMoyyed/FOKvVSdE6nvqYHXqdvbydO
7capF5r5VueS0PDkI15088H/PlGJcPrr37kx20sQRl/gQUwGZEXMpY8Ng4bpRkkQqH74lcWUNkv7
Mme9UpjjqG2BM0+BtVqnadMDUHOf/BrM5PuoRqB2X3q9n71MdtJhDmBm3PT2OSoyGgSuvKd+cecy
yYZ5B4mf/zzupBE4FdkYvy2o9cwksLEpDPAxTPGdL4U2l/kPh2kDuLg+2kKB4lxfIpYQIYBhe5t1
h69gWnCBSINDZ8TRqCR4Gn0GLc0hPeUeMr68rswaV2Xc+78jzZ3lOndrNH3Th68OTrnm8Q18Zy/o
VQdY48efEpdmnKzprhE1YREDIOWsQpAz3kOYahCaN7+u4X1EgxeHB145dJ5DNwCgjOojDAPFS7DE
6RpDLY+MNGJw1GLE7DQXnTPeOP41O4PAMqackC4Syv6NZhQk7rJe7xEfOIzH2s6xTn4a5qqN+sXL
j7gG70H0HjSAYTLabsx+YN2gVnXupGn3feBpNk2pdHz/rXjBm1us/LGjZC0/zsDFTI/OP1GUHQNr
Gr+7kTE4aXznso+2HcCZSWR+J0GJezzU5Isx2+t0yeeyuygxXK8mP07/1BJaUl7ADZc9aYmJ5JBq
Bcn+z5ctGlLJ5roA07offrPLqOTrd/s221PA7PazAbj25i9K7TfwDIYTjYsSq6q7cO3JQtkAgHAW
NvkAezILh8zw1llUOnWb+g++oxU7qkJSxx8/40PJOj/BkRXnGeqhyOLJiLar1oN/W1lMGAw1Ku+q
/80Wa/bV2gvEJrpAn6rTiaQPAAWLSnw5G60qEfATMjyQ+RjQ+ZdNeYwhO2CPqmnQKTQcjRhiyFLf
l1gcD2ZrhoGYw9hTyKaeSR0C5poGy11b3k3r3VVcOqpKSTib3VNzEG6S5XuEPIh/Hau/m387/9ip
CO2AdOqxEi26cLBK1ZOtYUAVbBJO35J+cG6wcBXY0AmehVsDjpBZ+g0bOv+46Ni9WZzstyVkwmOS
P/CZUsUH72GgVsac0WBWCPlMce+lAc74ck9eocsF6Iai3mlnHuOl55/BtunUYQ92HN7JYAUtbIjT
NVye9jePHXSXpzPqAuGQ3NPIpJuDIK8Co8y4kp0gny/25Xos1ScawIh4P/KjhWpNyjEobQqJe+12
9B+RcIS6z5q8nJF4P577HlDNSghM1pPbkkgqWQj5gLFfIVEg9ZyakwEWjwmF3AGb67GQaurvtrZf
lsP5NKdkXZrkniVrKBwYD1yrLCusKhTkm/ssA1LrkqENoUfvoA4o5R1Qk6FhhfIQZPLFH7iTt3Az
mQA+oGCilwKLtoG7NrMCQc/0/IsvBCYJ7v5p/Fg/WT2Oe4dbDDUobWzNED80babkil+XYWfmUtKv
AIGgPc6ANQ9vnK5ZtECVqLi4PPrqiXwT9uEvzFTPqrBeniHs9ueI6uRWUllpsvKXO/g+ZeF5dGbu
lPxVxqs44hjP1499JD+dkb/fRF3F7HRRoaMLRjwODPyJWLrjhAT7VCb4Sb0+R7URK+nG6WpMYUid
wZ0O3+S+G/brAioz89pfsY/meum9SLZ2g0fRiMPBt+wKCl7Zcxl6k6cIVA+hRqa4vBbspiRrnVCC
tlPn8a26bQDep4T7bvnYiGNlzs57guD7MGb98F/vdjMBg40ekb2DjS4UpjkNHyDMwyMcU26VF22W
d2iRcFxACxszfZepZtCZ+0rYM3pVxV7M3LlbRzZyhlUrxayHSvlWVkAoYVnNoAxb2hzim/yB38Ry
czfA5+6t8UFtgmrIPkJ/chuDlkZumeEyXtkvgjX0jZsTONN9wz3tcaIBcefywxdzsT4ZoG0rdRQU
UJkDtDAwLu6QiQxNnDnfeuCJRM8t39uE/fvsrsxY5OZ/r6YTeTWC6EMOZwA0D2UH0sf3nZJAxLpI
TbikwrnFcg==
`protect end_protected

